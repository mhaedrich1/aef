module dtc_split33_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node11;
	wire [16-1:0] node12;
	wire [16-1:0] node13;
	wire [16-1:0] node14;
	wire [16-1:0] node15;
	wire [16-1:0] node20;
	wire [16-1:0] node21;
	wire [16-1:0] node24;
	wire [16-1:0] node25;
	wire [16-1:0] node29;
	wire [16-1:0] node30;
	wire [16-1:0] node32;
	wire [16-1:0] node33;
	wire [16-1:0] node37;
	wire [16-1:0] node40;
	wire [16-1:0] node41;
	wire [16-1:0] node42;
	wire [16-1:0] node43;
	wire [16-1:0] node45;
	wire [16-1:0] node48;
	wire [16-1:0] node49;
	wire [16-1:0] node53;
	wire [16-1:0] node56;
	wire [16-1:0] node57;
	wire [16-1:0] node61;
	wire [16-1:0] node62;
	wire [16-1:0] node63;
	wire [16-1:0] node65;
	wire [16-1:0] node66;
	wire [16-1:0] node70;
	wire [16-1:0] node71;
	wire [16-1:0] node74;
	wire [16-1:0] node76;
	wire [16-1:0] node79;
	wire [16-1:0] node80;
	wire [16-1:0] node81;
	wire [16-1:0] node84;
	wire [16-1:0] node85;
	wire [16-1:0] node89;
	wire [16-1:0] node91;
	wire [16-1:0] node94;
	wire [16-1:0] node95;
	wire [16-1:0] node96;
	wire [16-1:0] node97;
	wire [16-1:0] node98;
	wire [16-1:0] node99;
	wire [16-1:0] node100;
	wire [16-1:0] node104;
	wire [16-1:0] node107;
	wire [16-1:0] node108;
	wire [16-1:0] node112;
	wire [16-1:0] node115;
	wire [16-1:0] node117;
	wire [16-1:0] node118;
	wire [16-1:0] node120;
	wire [16-1:0] node122;
	wire [16-1:0] node126;
	wire [16-1:0] node127;
	wire [16-1:0] node128;
	wire [16-1:0] node129;
	wire [16-1:0] node131;
	wire [16-1:0] node133;
	wire [16-1:0] node136;
	wire [16-1:0] node139;
	wire [16-1:0] node142;
	wire [16-1:0] node143;
	wire [16-1:0] node144;
	wire [16-1:0] node147;
	wire [16-1:0] node150;
	wire [16-1:0] node151;
	wire [16-1:0] node153;
	wire [16-1:0] node156;
	wire [16-1:0] node157;
	wire [16-1:0] node161;
	wire [16-1:0] node162;
	wire [16-1:0] node163;
	wire [16-1:0] node164;
	wire [16-1:0] node165;
	wire [16-1:0] node167;
	wire [16-1:0] node168;
	wire [16-1:0] node171;
	wire [16-1:0] node172;
	wire [16-1:0] node176;
	wire [16-1:0] node177;
	wire [16-1:0] node180;
	wire [16-1:0] node183;
	wire [16-1:0] node184;
	wire [16-1:0] node185;
	wire [16-1:0] node188;
	wire [16-1:0] node191;
	wire [16-1:0] node192;
	wire [16-1:0] node193;
	wire [16-1:0] node195;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node203;
	wire [16-1:0] node204;
	wire [16-1:0] node205;
	wire [16-1:0] node210;
	wire [16-1:0] node211;
	wire [16-1:0] node212;
	wire [16-1:0] node213;
	wire [16-1:0] node216;
	wire [16-1:0] node218;
	wire [16-1:0] node222;
	wire [16-1:0] node223;
	wire [16-1:0] node224;
	wire [16-1:0] node227;
	wire [16-1:0] node228;
	wire [16-1:0] node230;
	wire [16-1:0] node234;
	wire [16-1:0] node235;
	wire [16-1:0] node238;
	wire [16-1:0] node241;
	wire [16-1:0] node242;
	wire [16-1:0] node243;
	wire [16-1:0] node244;
	wire [16-1:0] node247;
	wire [16-1:0] node249;
	wire [16-1:0] node250;
	wire [16-1:0] node253;
	wire [16-1:0] node256;
	wire [16-1:0] node257;
	wire [16-1:0] node259;
	wire [16-1:0] node262;
	wire [16-1:0] node263;
	wire [16-1:0] node267;
	wire [16-1:0] node268;
	wire [16-1:0] node270;
	wire [16-1:0] node271;
	wire [16-1:0] node274;
	wire [16-1:0] node275;
	wire [16-1:0] node279;
	wire [16-1:0] node280;
	wire [16-1:0] node281;
	wire [16-1:0] node282;
	wire [16-1:0] node286;
	wire [16-1:0] node289;
	wire [16-1:0] node292;
	wire [16-1:0] node293;
	wire [16-1:0] node294;
	wire [16-1:0] node295;
	wire [16-1:0] node296;
	wire [16-1:0] node297;
	wire [16-1:0] node298;
	wire [16-1:0] node300;
	wire [16-1:0] node301;
	wire [16-1:0] node305;
	wire [16-1:0] node307;
	wire [16-1:0] node310;
	wire [16-1:0] node311;
	wire [16-1:0] node314;
	wire [16-1:0] node317;
	wire [16-1:0] node319;
	wire [16-1:0] node320;
	wire [16-1:0] node323;
	wire [16-1:0] node326;
	wire [16-1:0] node327;
	wire [16-1:0] node328;
	wire [16-1:0] node329;
	wire [16-1:0] node330;
	wire [16-1:0] node332;
	wire [16-1:0] node336;
	wire [16-1:0] node337;
	wire [16-1:0] node339;
	wire [16-1:0] node343;
	wire [16-1:0] node344;
	wire [16-1:0] node347;
	wire [16-1:0] node350;
	wire [16-1:0] node351;
	wire [16-1:0] node354;
	wire [16-1:0] node355;
	wire [16-1:0] node357;
	wire [16-1:0] node358;
	wire [16-1:0] node362;
	wire [16-1:0] node365;
	wire [16-1:0] node366;
	wire [16-1:0] node367;
	wire [16-1:0] node368;
	wire [16-1:0] node370;
	wire [16-1:0] node373;
	wire [16-1:0] node374;
	wire [16-1:0] node376;
	wire [16-1:0] node377;
	wire [16-1:0] node381;
	wire [16-1:0] node382;
	wire [16-1:0] node386;
	wire [16-1:0] node387;
	wire [16-1:0] node388;
	wire [16-1:0] node389;
	wire [16-1:0] node393;
	wire [16-1:0] node396;
	wire [16-1:0] node397;
	wire [16-1:0] node400;
	wire [16-1:0] node403;
	wire [16-1:0] node404;
	wire [16-1:0] node405;
	wire [16-1:0] node406;
	wire [16-1:0] node407;
	wire [16-1:0] node409;
	wire [16-1:0] node412;
	wire [16-1:0] node415;
	wire [16-1:0] node417;
	wire [16-1:0] node420;
	wire [16-1:0] node421;
	wire [16-1:0] node423;
	wire [16-1:0] node426;
	wire [16-1:0] node428;
	wire [16-1:0] node431;
	wire [16-1:0] node432;
	wire [16-1:0] node433;
	wire [16-1:0] node436;
	wire [16-1:0] node437;
	wire [16-1:0] node441;
	wire [16-1:0] node442;
	wire [16-1:0] node443;
	wire [16-1:0] node447;
	wire [16-1:0] node449;
	wire [16-1:0] node452;
	wire [16-1:0] node453;
	wire [16-1:0] node454;
	wire [16-1:0] node455;
	wire [16-1:0] node456;
	wire [16-1:0] node458;
	wire [16-1:0] node462;
	wire [16-1:0] node464;
	wire [16-1:0] node465;
	wire [16-1:0] node469;
	wire [16-1:0] node470;
	wire [16-1:0] node471;
	wire [16-1:0] node472;
	wire [16-1:0] node476;
	wire [16-1:0] node478;
	wire [16-1:0] node481;
	wire [16-1:0] node483;
	wire [16-1:0] node486;
	wire [16-1:0] node487;
	wire [16-1:0] node488;
	wire [16-1:0] node489;
	wire [16-1:0] node490;
	wire [16-1:0] node491;
	wire [16-1:0] node495;
	wire [16-1:0] node498;
	wire [16-1:0] node499;
	wire [16-1:0] node500;
	wire [16-1:0] node502;
	wire [16-1:0] node506;
	wire [16-1:0] node509;
	wire [16-1:0] node510;
	wire [16-1:0] node514;
	wire [16-1:0] node515;
	wire [16-1:0] node516;
	wire [16-1:0] node517;
	wire [16-1:0] node520;
	wire [16-1:0] node521;
	wire [16-1:0] node525;
	wire [16-1:0] node526;
	wire [16-1:0] node527;
	wire [16-1:0] node532;
	wire [16-1:0] node533;
	wire [16-1:0] node534;
	wire [16-1:0] node537;
	wire [16-1:0] node539;
	wire [16-1:0] node542;
	wire [16-1:0] node543;
	wire [16-1:0] node546;
	wire [16-1:0] node547;
	wire [16-1:0] node549;
	wire [16-1:0] node552;
	wire [16-1:0] node555;
	wire [16-1:0] node556;
	wire [16-1:0] node557;
	wire [16-1:0] node558;
	wire [16-1:0] node559;
	wire [16-1:0] node560;
	wire [16-1:0] node561;
	wire [16-1:0] node562;
	wire [16-1:0] node565;
	wire [16-1:0] node568;
	wire [16-1:0] node570;
	wire [16-1:0] node573;
	wire [16-1:0] node574;
	wire [16-1:0] node575;
	wire [16-1:0] node577;
	wire [16-1:0] node581;
	wire [16-1:0] node582;
	wire [16-1:0] node584;
	wire [16-1:0] node588;
	wire [16-1:0] node589;
	wire [16-1:0] node590;
	wire [16-1:0] node592;
	wire [16-1:0] node593;
	wire [16-1:0] node595;
	wire [16-1:0] node598;
	wire [16-1:0] node600;
	wire [16-1:0] node603;
	wire [16-1:0] node604;
	wire [16-1:0] node605;
	wire [16-1:0] node609;
	wire [16-1:0] node612;
	wire [16-1:0] node614;
	wire [16-1:0] node615;
	wire [16-1:0] node619;
	wire [16-1:0] node620;
	wire [16-1:0] node621;
	wire [16-1:0] node622;
	wire [16-1:0] node623;
	wire [16-1:0] node625;
	wire [16-1:0] node626;
	wire [16-1:0] node631;
	wire [16-1:0] node632;
	wire [16-1:0] node633;
	wire [16-1:0] node637;
	wire [16-1:0] node639;
	wire [16-1:0] node642;
	wire [16-1:0] node643;
	wire [16-1:0] node645;
	wire [16-1:0] node648;
	wire [16-1:0] node650;
	wire [16-1:0] node653;
	wire [16-1:0] node654;
	wire [16-1:0] node655;
	wire [16-1:0] node657;
	wire [16-1:0] node660;
	wire [16-1:0] node661;
	wire [16-1:0] node662;
	wire [16-1:0] node664;
	wire [16-1:0] node668;
	wire [16-1:0] node671;
	wire [16-1:0] node672;
	wire [16-1:0] node674;
	wire [16-1:0] node677;
	wire [16-1:0] node679;
	wire [16-1:0] node681;
	wire [16-1:0] node684;
	wire [16-1:0] node685;
	wire [16-1:0] node686;
	wire [16-1:0] node687;
	wire [16-1:0] node688;
	wire [16-1:0] node689;
	wire [16-1:0] node692;
	wire [16-1:0] node693;
	wire [16-1:0] node696;
	wire [16-1:0] node699;
	wire [16-1:0] node701;
	wire [16-1:0] node703;
	wire [16-1:0] node706;
	wire [16-1:0] node707;
	wire [16-1:0] node709;
	wire [16-1:0] node712;
	wire [16-1:0] node713;
	wire [16-1:0] node716;
	wire [16-1:0] node717;
	wire [16-1:0] node721;
	wire [16-1:0] node722;
	wire [16-1:0] node724;
	wire [16-1:0] node725;
	wire [16-1:0] node726;
	wire [16-1:0] node731;
	wire [16-1:0] node732;
	wire [16-1:0] node733;
	wire [16-1:0] node736;
	wire [16-1:0] node738;
	wire [16-1:0] node741;
	wire [16-1:0] node742;
	wire [16-1:0] node746;
	wire [16-1:0] node747;
	wire [16-1:0] node748;
	wire [16-1:0] node749;
	wire [16-1:0] node750;
	wire [16-1:0] node753;
	wire [16-1:0] node754;
	wire [16-1:0] node756;
	wire [16-1:0] node761;
	wire [16-1:0] node762;
	wire [16-1:0] node764;
	wire [16-1:0] node765;
	wire [16-1:0] node766;
	wire [16-1:0] node769;
	wire [16-1:0] node773;
	wire [16-1:0] node774;
	wire [16-1:0] node776;
	wire [16-1:0] node779;
	wire [16-1:0] node782;
	wire [16-1:0] node783;
	wire [16-1:0] node785;
	wire [16-1:0] node786;
	wire [16-1:0] node790;
	wire [16-1:0] node791;
	wire [16-1:0] node793;
	wire [16-1:0] node796;
	wire [16-1:0] node797;
	wire [16-1:0] node798;
	wire [16-1:0] node803;
	wire [16-1:0] node804;
	wire [16-1:0] node805;
	wire [16-1:0] node806;
	wire [16-1:0] node807;
	wire [16-1:0] node808;
	wire [16-1:0] node809;
	wire [16-1:0] node810;
	wire [16-1:0] node813;
	wire [16-1:0] node816;
	wire [16-1:0] node817;
	wire [16-1:0] node820;
	wire [16-1:0] node824;
	wire [16-1:0] node825;
	wire [16-1:0] node826;
	wire [16-1:0] node828;
	wire [16-1:0] node829;
	wire [16-1:0] node833;
	wire [16-1:0] node836;
	wire [16-1:0] node839;
	wire [16-1:0] node840;
	wire [16-1:0] node841;
	wire [16-1:0] node843;
	wire [16-1:0] node844;
	wire [16-1:0] node848;
	wire [16-1:0] node850;
	wire [16-1:0] node853;
	wire [16-1:0] node854;
	wire [16-1:0] node855;
	wire [16-1:0] node856;
	wire [16-1:0] node860;
	wire [16-1:0] node861;
	wire [16-1:0] node865;
	wire [16-1:0] node867;
	wire [16-1:0] node870;
	wire [16-1:0] node871;
	wire [16-1:0] node872;
	wire [16-1:0] node873;
	wire [16-1:0] node874;
	wire [16-1:0] node878;
	wire [16-1:0] node879;
	wire [16-1:0] node880;
	wire [16-1:0] node885;
	wire [16-1:0] node886;
	wire [16-1:0] node887;
	wire [16-1:0] node888;
	wire [16-1:0] node890;
	wire [16-1:0] node895;
	wire [16-1:0] node896;
	wire [16-1:0] node897;
	wire [16-1:0] node901;
	wire [16-1:0] node904;
	wire [16-1:0] node905;
	wire [16-1:0] node906;
	wire [16-1:0] node908;
	wire [16-1:0] node911;
	wire [16-1:0] node912;
	wire [16-1:0] node915;
	wire [16-1:0] node916;
	wire [16-1:0] node920;
	wire [16-1:0] node921;
	wire [16-1:0] node923;
	wire [16-1:0] node926;
	wire [16-1:0] node927;
	wire [16-1:0] node931;
	wire [16-1:0] node932;
	wire [16-1:0] node933;
	wire [16-1:0] node934;
	wire [16-1:0] node935;
	wire [16-1:0] node938;
	wire [16-1:0] node939;
	wire [16-1:0] node940;
	wire [16-1:0] node944;
	wire [16-1:0] node945;
	wire [16-1:0] node947;
	wire [16-1:0] node951;
	wire [16-1:0] node952;
	wire [16-1:0] node954;
	wire [16-1:0] node957;
	wire [16-1:0] node960;
	wire [16-1:0] node961;
	wire [16-1:0] node962;
	wire [16-1:0] node963;
	wire [16-1:0] node964;
	wire [16-1:0] node966;
	wire [16-1:0] node970;
	wire [16-1:0] node972;
	wire [16-1:0] node975;
	wire [16-1:0] node976;
	wire [16-1:0] node979;
	wire [16-1:0] node982;
	wire [16-1:0] node983;
	wire [16-1:0] node984;
	wire [16-1:0] node985;
	wire [16-1:0] node988;
	wire [16-1:0] node990;
	wire [16-1:0] node993;
	wire [16-1:0] node994;
	wire [16-1:0] node996;
	wire [16-1:0] node999;
	wire [16-1:0] node1001;
	wire [16-1:0] node1004;
	wire [16-1:0] node1005;
	wire [16-1:0] node1008;
	wire [16-1:0] node1011;
	wire [16-1:0] node1012;
	wire [16-1:0] node1013;
	wire [16-1:0] node1014;
	wire [16-1:0] node1015;
	wire [16-1:0] node1018;
	wire [16-1:0] node1019;
	wire [16-1:0] node1021;
	wire [16-1:0] node1024;
	wire [16-1:0] node1025;
	wire [16-1:0] node1029;
	wire [16-1:0] node1032;
	wire [16-1:0] node1033;
	wire [16-1:0] node1034;
	wire [16-1:0] node1037;
	wire [16-1:0] node1038;
	wire [16-1:0] node1042;
	wire [16-1:0] node1044;
	wire [16-1:0] node1047;
	wire [16-1:0] node1048;
	wire [16-1:0] node1049;
	wire [16-1:0] node1050;
	wire [16-1:0] node1054;
	wire [16-1:0] node1056;
	wire [16-1:0] node1058;
	wire [16-1:0] node1060;
	wire [16-1:0] node1063;
	wire [16-1:0] node1064;
	wire [16-1:0] node1066;
	wire [16-1:0] node1067;
	wire [16-1:0] node1071;
	wire [16-1:0] node1073;
	wire [16-1:0] node1075;
	wire [16-1:0] node1077;
	wire [16-1:0] node1080;
	wire [16-1:0] node1081;
	wire [16-1:0] node1082;
	wire [16-1:0] node1083;
	wire [16-1:0] node1084;
	wire [16-1:0] node1085;
	wire [16-1:0] node1086;
	wire [16-1:0] node1087;
	wire [16-1:0] node1088;
	wire [16-1:0] node1089;
	wire [16-1:0] node1093;
	wire [16-1:0] node1096;
	wire [16-1:0] node1097;
	wire [16-1:0] node1099;
	wire [16-1:0] node1102;
	wire [16-1:0] node1104;
	wire [16-1:0] node1107;
	wire [16-1:0] node1108;
	wire [16-1:0] node1109;
	wire [16-1:0] node1112;
	wire [16-1:0] node1115;
	wire [16-1:0] node1117;
	wire [16-1:0] node1120;
	wire [16-1:0] node1121;
	wire [16-1:0] node1122;
	wire [16-1:0] node1123;
	wire [16-1:0] node1126;
	wire [16-1:0] node1129;
	wire [16-1:0] node1130;
	wire [16-1:0] node1131;
	wire [16-1:0] node1135;
	wire [16-1:0] node1136;
	wire [16-1:0] node1138;
	wire [16-1:0] node1142;
	wire [16-1:0] node1143;
	wire [16-1:0] node1145;
	wire [16-1:0] node1146;
	wire [16-1:0] node1147;
	wire [16-1:0] node1150;
	wire [16-1:0] node1154;
	wire [16-1:0] node1155;
	wire [16-1:0] node1159;
	wire [16-1:0] node1160;
	wire [16-1:0] node1161;
	wire [16-1:0] node1162;
	wire [16-1:0] node1163;
	wire [16-1:0] node1164;
	wire [16-1:0] node1168;
	wire [16-1:0] node1169;
	wire [16-1:0] node1171;
	wire [16-1:0] node1175;
	wire [16-1:0] node1178;
	wire [16-1:0] node1179;
	wire [16-1:0] node1180;
	wire [16-1:0] node1181;
	wire [16-1:0] node1183;
	wire [16-1:0] node1188;
	wire [16-1:0] node1189;
	wire [16-1:0] node1192;
	wire [16-1:0] node1194;
	wire [16-1:0] node1197;
	wire [16-1:0] node1198;
	wire [16-1:0] node1199;
	wire [16-1:0] node1200;
	wire [16-1:0] node1203;
	wire [16-1:0] node1204;
	wire [16-1:0] node1206;
	wire [16-1:0] node1210;
	wire [16-1:0] node1211;
	wire [16-1:0] node1214;
	wire [16-1:0] node1217;
	wire [16-1:0] node1218;
	wire [16-1:0] node1219;
	wire [16-1:0] node1222;
	wire [16-1:0] node1225;
	wire [16-1:0] node1228;
	wire [16-1:0] node1229;
	wire [16-1:0] node1230;
	wire [16-1:0] node1231;
	wire [16-1:0] node1232;
	wire [16-1:0] node1233;
	wire [16-1:0] node1235;
	wire [16-1:0] node1236;
	wire [16-1:0] node1241;
	wire [16-1:0] node1242;
	wire [16-1:0] node1246;
	wire [16-1:0] node1247;
	wire [16-1:0] node1249;
	wire [16-1:0] node1252;
	wire [16-1:0] node1255;
	wire [16-1:0] node1256;
	wire [16-1:0] node1257;
	wire [16-1:0] node1259;
	wire [16-1:0] node1260;
	wire [16-1:0] node1264;
	wire [16-1:0] node1266;
	wire [16-1:0] node1269;
	wire [16-1:0] node1271;
	wire [16-1:0] node1274;
	wire [16-1:0] node1275;
	wire [16-1:0] node1276;
	wire [16-1:0] node1277;
	wire [16-1:0] node1278;
	wire [16-1:0] node1281;
	wire [16-1:0] node1283;
	wire [16-1:0] node1286;
	wire [16-1:0] node1287;
	wire [16-1:0] node1291;
	wire [16-1:0] node1292;
	wire [16-1:0] node1294;
	wire [16-1:0] node1296;
	wire [16-1:0] node1299;
	wire [16-1:0] node1300;
	wire [16-1:0] node1304;
	wire [16-1:0] node1305;
	wire [16-1:0] node1306;
	wire [16-1:0] node1307;
	wire [16-1:0] node1308;
	wire [16-1:0] node1312;
	wire [16-1:0] node1315;
	wire [16-1:0] node1316;
	wire [16-1:0] node1318;
	wire [16-1:0] node1319;
	wire [16-1:0] node1324;
	wire [16-1:0] node1325;
	wire [16-1:0] node1326;
	wire [16-1:0] node1327;
	wire [16-1:0] node1329;
	wire [16-1:0] node1333;
	wire [16-1:0] node1336;
	wire [16-1:0] node1337;
	wire [16-1:0] node1338;
	wire [16-1:0] node1342;
	wire [16-1:0] node1344;
	wire [16-1:0] node1347;
	wire [16-1:0] node1348;
	wire [16-1:0] node1349;
	wire [16-1:0] node1350;
	wire [16-1:0] node1351;
	wire [16-1:0] node1353;
	wire [16-1:0] node1354;
	wire [16-1:0] node1357;
	wire [16-1:0] node1360;
	wire [16-1:0] node1362;
	wire [16-1:0] node1363;
	wire [16-1:0] node1367;
	wire [16-1:0] node1368;
	wire [16-1:0] node1370;
	wire [16-1:0] node1372;
	wire [16-1:0] node1373;
	wire [16-1:0] node1377;
	wire [16-1:0] node1378;
	wire [16-1:0] node1379;
	wire [16-1:0] node1380;
	wire [16-1:0] node1381;
	wire [16-1:0] node1385;
	wire [16-1:0] node1386;
	wire [16-1:0] node1391;
	wire [16-1:0] node1392;
	wire [16-1:0] node1393;
	wire [16-1:0] node1398;
	wire [16-1:0] node1399;
	wire [16-1:0] node1400;
	wire [16-1:0] node1401;
	wire [16-1:0] node1402;
	wire [16-1:0] node1403;
	wire [16-1:0] node1404;
	wire [16-1:0] node1410;
	wire [16-1:0] node1413;
	wire [16-1:0] node1414;
	wire [16-1:0] node1416;
	wire [16-1:0] node1418;
	wire [16-1:0] node1421;
	wire [16-1:0] node1422;
	wire [16-1:0] node1426;
	wire [16-1:0] node1427;
	wire [16-1:0] node1428;
	wire [16-1:0] node1429;
	wire [16-1:0] node1432;
	wire [16-1:0] node1433;
	wire [16-1:0] node1435;
	wire [16-1:0] node1438;
	wire [16-1:0] node1441;
	wire [16-1:0] node1442;
	wire [16-1:0] node1444;
	wire [16-1:0] node1448;
	wire [16-1:0] node1450;
	wire [16-1:0] node1453;
	wire [16-1:0] node1454;
	wire [16-1:0] node1455;
	wire [16-1:0] node1456;
	wire [16-1:0] node1457;
	wire [16-1:0] node1458;
	wire [16-1:0] node1459;
	wire [16-1:0] node1461;
	wire [16-1:0] node1465;
	wire [16-1:0] node1466;
	wire [16-1:0] node1468;
	wire [16-1:0] node1472;
	wire [16-1:0] node1474;
	wire [16-1:0] node1475;
	wire [16-1:0] node1478;
	wire [16-1:0] node1479;
	wire [16-1:0] node1483;
	wire [16-1:0] node1485;
	wire [16-1:0] node1487;
	wire [16-1:0] node1490;
	wire [16-1:0] node1491;
	wire [16-1:0] node1492;
	wire [16-1:0] node1493;
	wire [16-1:0] node1495;
	wire [16-1:0] node1496;
	wire [16-1:0] node1501;
	wire [16-1:0] node1502;
	wire [16-1:0] node1505;
	wire [16-1:0] node1507;
	wire [16-1:0] node1510;
	wire [16-1:0] node1511;
	wire [16-1:0] node1512;
	wire [16-1:0] node1513;
	wire [16-1:0] node1517;
	wire [16-1:0] node1519;
	wire [16-1:0] node1522;
	wire [16-1:0] node1523;
	wire [16-1:0] node1526;
	wire [16-1:0] node1528;
	wire [16-1:0] node1531;
	wire [16-1:0] node1532;
	wire [16-1:0] node1533;
	wire [16-1:0] node1534;
	wire [16-1:0] node1535;
	wire [16-1:0] node1539;
	wire [16-1:0] node1540;
	wire [16-1:0] node1541;
	wire [16-1:0] node1545;
	wire [16-1:0] node1548;
	wire [16-1:0] node1549;
	wire [16-1:0] node1550;
	wire [16-1:0] node1553;
	wire [16-1:0] node1556;
	wire [16-1:0] node1557;
	wire [16-1:0] node1560;
	wire [16-1:0] node1561;
	wire [16-1:0] node1563;
	wire [16-1:0] node1567;
	wire [16-1:0] node1568;
	wire [16-1:0] node1569;
	wire [16-1:0] node1570;
	wire [16-1:0] node1572;
	wire [16-1:0] node1575;
	wire [16-1:0] node1578;
	wire [16-1:0] node1579;
	wire [16-1:0] node1582;
	wire [16-1:0] node1585;
	wire [16-1:0] node1586;
	wire [16-1:0] node1587;
	wire [16-1:0] node1589;
	wire [16-1:0] node1591;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1599;
	wire [16-1:0] node1600;
	wire [16-1:0] node1603;
	wire [16-1:0] node1606;
	wire [16-1:0] node1607;
	wire [16-1:0] node1608;
	wire [16-1:0] node1609;
	wire [16-1:0] node1610;
	wire [16-1:0] node1611;
	wire [16-1:0] node1612;
	wire [16-1:0] node1613;
	wire [16-1:0] node1616;
	wire [16-1:0] node1617;
	wire [16-1:0] node1621;
	wire [16-1:0] node1622;
	wire [16-1:0] node1623;
	wire [16-1:0] node1627;
	wire [16-1:0] node1628;
	wire [16-1:0] node1632;
	wire [16-1:0] node1635;
	wire [16-1:0] node1636;
	wire [16-1:0] node1637;
	wire [16-1:0] node1638;
	wire [16-1:0] node1641;
	wire [16-1:0] node1644;
	wire [16-1:0] node1645;
	wire [16-1:0] node1646;
	wire [16-1:0] node1650;
	wire [16-1:0] node1652;
	wire [16-1:0] node1655;
	wire [16-1:0] node1656;
	wire [16-1:0] node1657;
	wire [16-1:0] node1661;
	wire [16-1:0] node1662;
	wire [16-1:0] node1665;
	wire [16-1:0] node1667;
	wire [16-1:0] node1670;
	wire [16-1:0] node1671;
	wire [16-1:0] node1672;
	wire [16-1:0] node1673;
	wire [16-1:0] node1674;
	wire [16-1:0] node1675;
	wire [16-1:0] node1677;
	wire [16-1:0] node1681;
	wire [16-1:0] node1684;
	wire [16-1:0] node1685;
	wire [16-1:0] node1686;
	wire [16-1:0] node1688;
	wire [16-1:0] node1692;
	wire [16-1:0] node1693;
	wire [16-1:0] node1695;
	wire [16-1:0] node1699;
	wire [16-1:0] node1700;
	wire [16-1:0] node1702;
	wire [16-1:0] node1706;
	wire [16-1:0] node1707;
	wire [16-1:0] node1708;
	wire [16-1:0] node1710;
	wire [16-1:0] node1712;
	wire [16-1:0] node1715;
	wire [16-1:0] node1716;
	wire [16-1:0] node1717;
	wire [16-1:0] node1721;
	wire [16-1:0] node1724;
	wire [16-1:0] node1725;
	wire [16-1:0] node1727;
	wire [16-1:0] node1729;
	wire [16-1:0] node1732;
	wire [16-1:0] node1733;
	wire [16-1:0] node1737;
	wire [16-1:0] node1738;
	wire [16-1:0] node1739;
	wire [16-1:0] node1740;
	wire [16-1:0] node1741;
	wire [16-1:0] node1742;
	wire [16-1:0] node1746;
	wire [16-1:0] node1747;
	wire [16-1:0] node1749;
	wire [16-1:0] node1752;
	wire [16-1:0] node1755;
	wire [16-1:0] node1756;
	wire [16-1:0] node1757;
	wire [16-1:0] node1760;
	wire [16-1:0] node1761;
	wire [16-1:0] node1765;
	wire [16-1:0] node1768;
	wire [16-1:0] node1769;
	wire [16-1:0] node1770;
	wire [16-1:0] node1771;
	wire [16-1:0] node1775;
	wire [16-1:0] node1776;
	wire [16-1:0] node1777;
	wire [16-1:0] node1782;
	wire [16-1:0] node1783;
	wire [16-1:0] node1784;
	wire [16-1:0] node1785;
	wire [16-1:0] node1787;
	wire [16-1:0] node1791;
	wire [16-1:0] node1793;
	wire [16-1:0] node1796;
	wire [16-1:0] node1798;
	wire [16-1:0] node1801;
	wire [16-1:0] node1802;
	wire [16-1:0] node1803;
	wire [16-1:0] node1804;
	wire [16-1:0] node1805;
	wire [16-1:0] node1808;
	wire [16-1:0] node1812;
	wire [16-1:0] node1813;
	wire [16-1:0] node1815;
	wire [16-1:0] node1817;
	wire [16-1:0] node1818;
	wire [16-1:0] node1822;
	wire [16-1:0] node1823;
	wire [16-1:0] node1827;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1830;
	wire [16-1:0] node1831;
	wire [16-1:0] node1834;
	wire [16-1:0] node1835;
	wire [16-1:0] node1839;
	wire [16-1:0] node1842;
	wire [16-1:0] node1843;
	wire [16-1:0] node1845;
	wire [16-1:0] node1846;
	wire [16-1:0] node1850;
	wire [16-1:0] node1851;
	wire [16-1:0] node1853;
	wire [16-1:0] node1857;
	wire [16-1:0] node1858;
	wire [16-1:0] node1859;
	wire [16-1:0] node1862;
	wire [16-1:0] node1863;
	wire [16-1:0] node1865;
	wire [16-1:0] node1869;
	wire [16-1:0] node1870;
	wire [16-1:0] node1871;
	wire [16-1:0] node1876;
	wire [16-1:0] node1877;
	wire [16-1:0] node1878;
	wire [16-1:0] node1879;
	wire [16-1:0] node1880;
	wire [16-1:0] node1883;
	wire [16-1:0] node1885;
	wire [16-1:0] node1887;
	wire [16-1:0] node1890;
	wire [16-1:0] node1891;
	wire [16-1:0] node1892;
	wire [16-1:0] node1893;
	wire [16-1:0] node1894;
	wire [16-1:0] node1898;
	wire [16-1:0] node1901;
	wire [16-1:0] node1902;
	wire [16-1:0] node1906;
	wire [16-1:0] node1907;
	wire [16-1:0] node1908;
	wire [16-1:0] node1911;
	wire [16-1:0] node1914;
	wire [16-1:0] node1915;
	wire [16-1:0] node1918;
	wire [16-1:0] node1921;
	wire [16-1:0] node1922;
	wire [16-1:0] node1923;
	wire [16-1:0] node1924;
	wire [16-1:0] node1927;
	wire [16-1:0] node1928;
	wire [16-1:0] node1932;
	wire [16-1:0] node1933;
	wire [16-1:0] node1934;
	wire [16-1:0] node1937;
	wire [16-1:0] node1940;
	wire [16-1:0] node1941;
	wire [16-1:0] node1943;
	wire [16-1:0] node1944;
	wire [16-1:0] node1949;
	wire [16-1:0] node1950;
	wire [16-1:0] node1951;
	wire [16-1:0] node1953;
	wire [16-1:0] node1956;
	wire [16-1:0] node1958;
	wire [16-1:0] node1961;
	wire [16-1:0] node1962;
	wire [16-1:0] node1964;
	wire [16-1:0] node1967;
	wire [16-1:0] node1970;
	wire [16-1:0] node1971;
	wire [16-1:0] node1972;
	wire [16-1:0] node1973;
	wire [16-1:0] node1974;
	wire [16-1:0] node1976;
	wire [16-1:0] node1979;
	wire [16-1:0] node1980;
	wire [16-1:0] node1983;
	wire [16-1:0] node1985;
	wire [16-1:0] node1986;
	wire [16-1:0] node1990;
	wire [16-1:0] node1991;
	wire [16-1:0] node1993;
	wire [16-1:0] node1996;
	wire [16-1:0] node1997;
	wire [16-1:0] node2000;
	wire [16-1:0] node2001;
	wire [16-1:0] node2004;
	wire [16-1:0] node2007;
	wire [16-1:0] node2008;
	wire [16-1:0] node2009;
	wire [16-1:0] node2010;
	wire [16-1:0] node2013;
	wire [16-1:0] node2014;
	wire [16-1:0] node2018;
	wire [16-1:0] node2020;
	wire [16-1:0] node2022;
	wire [16-1:0] node2025;
	wire [16-1:0] node2026;
	wire [16-1:0] node2028;
	wire [16-1:0] node2030;
	wire [16-1:0] node2033;
	wire [16-1:0] node2034;
	wire [16-1:0] node2036;
	wire [16-1:0] node2040;
	wire [16-1:0] node2041;
	wire [16-1:0] node2042;
	wire [16-1:0] node2043;
	wire [16-1:0] node2046;
	wire [16-1:0] node2049;
	wire [16-1:0] node2050;
	wire [16-1:0] node2051;
	wire [16-1:0] node2052;
	wire [16-1:0] node2056;
	wire [16-1:0] node2060;
	wire [16-1:0] node2061;
	wire [16-1:0] node2063;
	wire [16-1:0] node2064;
	wire [16-1:0] node2065;
	wire [16-1:0] node2069;
	wire [16-1:0] node2072;
	wire [16-1:0] node2073;
	wire [16-1:0] node2075;
	wire [16-1:0] node2076;
	wire [16-1:0] node2080;
	wire [16-1:0] node2081;
	wire [16-1:0] node2084;
	wire [16-1:0] node2085;
	wire [16-1:0] node2088;
	wire [16-1:0] node2090;
	wire [16-1:0] node2093;
	wire [16-1:0] node2094;
	wire [16-1:0] node2095;
	wire [16-1:0] node2096;
	wire [16-1:0] node2097;
	wire [16-1:0] node2098;
	wire [16-1:0] node2099;
	wire [16-1:0] node2100;
	wire [16-1:0] node2101;
	wire [16-1:0] node2102;
	wire [16-1:0] node2106;
	wire [16-1:0] node2107;
	wire [16-1:0] node2111;
	wire [16-1:0] node2112;
	wire [16-1:0] node2113;
	wire [16-1:0] node2115;
	wire [16-1:0] node2116;
	wire [16-1:0] node2120;
	wire [16-1:0] node2123;
	wire [16-1:0] node2124;
	wire [16-1:0] node2126;
	wire [16-1:0] node2127;
	wire [16-1:0] node2131;
	wire [16-1:0] node2132;
	wire [16-1:0] node2134;
	wire [16-1:0] node2138;
	wire [16-1:0] node2139;
	wire [16-1:0] node2140;
	wire [16-1:0] node2142;
	wire [16-1:0] node2145;
	wire [16-1:0] node2146;
	wire [16-1:0] node2147;
	wire [16-1:0] node2152;
	wire [16-1:0] node2153;
	wire [16-1:0] node2155;
	wire [16-1:0] node2157;
	wire [16-1:0] node2160;
	wire [16-1:0] node2161;
	wire [16-1:0] node2165;
	wire [16-1:0] node2166;
	wire [16-1:0] node2167;
	wire [16-1:0] node2168;
	wire [16-1:0] node2169;
	wire [16-1:0] node2171;
	wire [16-1:0] node2173;
	wire [16-1:0] node2177;
	wire [16-1:0] node2178;
	wire [16-1:0] node2181;
	wire [16-1:0] node2183;
	wire [16-1:0] node2186;
	wire [16-1:0] node2187;
	wire [16-1:0] node2188;
	wire [16-1:0] node2191;
	wire [16-1:0] node2193;
	wire [16-1:0] node2194;
	wire [16-1:0] node2198;
	wire [16-1:0] node2199;
	wire [16-1:0] node2203;
	wire [16-1:0] node2204;
	wire [16-1:0] node2205;
	wire [16-1:0] node2206;
	wire [16-1:0] node2207;
	wire [16-1:0] node2209;
	wire [16-1:0] node2212;
	wire [16-1:0] node2214;
	wire [16-1:0] node2217;
	wire [16-1:0] node2218;
	wire [16-1:0] node2220;
	wire [16-1:0] node2223;
	wire [16-1:0] node2226;
	wire [16-1:0] node2227;
	wire [16-1:0] node2230;
	wire [16-1:0] node2233;
	wire [16-1:0] node2234;
	wire [16-1:0] node2235;
	wire [16-1:0] node2236;
	wire [16-1:0] node2241;
	wire [16-1:0] node2242;
	wire [16-1:0] node2245;
	wire [16-1:0] node2248;
	wire [16-1:0] node2249;
	wire [16-1:0] node2250;
	wire [16-1:0] node2251;
	wire [16-1:0] node2252;
	wire [16-1:0] node2254;
	wire [16-1:0] node2257;
	wire [16-1:0] node2258;
	wire [16-1:0] node2261;
	wire [16-1:0] node2263;
	wire [16-1:0] node2264;
	wire [16-1:0] node2268;
	wire [16-1:0] node2269;
	wire [16-1:0] node2271;
	wire [16-1:0] node2274;
	wire [16-1:0] node2275;
	wire [16-1:0] node2279;
	wire [16-1:0] node2280;
	wire [16-1:0] node2281;
	wire [16-1:0] node2282;
	wire [16-1:0] node2284;
	wire [16-1:0] node2285;
	wire [16-1:0] node2289;
	wire [16-1:0] node2291;
	wire [16-1:0] node2294;
	wire [16-1:0] node2295;
	wire [16-1:0] node2298;
	wire [16-1:0] node2301;
	wire [16-1:0] node2303;
	wire [16-1:0] node2304;
	wire [16-1:0] node2307;
	wire [16-1:0] node2310;
	wire [16-1:0] node2311;
	wire [16-1:0] node2312;
	wire [16-1:0] node2313;
	wire [16-1:0] node2314;
	wire [16-1:0] node2315;
	wire [16-1:0] node2319;
	wire [16-1:0] node2321;
	wire [16-1:0] node2324;
	wire [16-1:0] node2325;
	wire [16-1:0] node2326;
	wire [16-1:0] node2327;
	wire [16-1:0] node2330;
	wire [16-1:0] node2335;
	wire [16-1:0] node2336;
	wire [16-1:0] node2337;
	wire [16-1:0] node2340;
	wire [16-1:0] node2342;
	wire [16-1:0] node2345;
	wire [16-1:0] node2347;
	wire [16-1:0] node2350;
	wire [16-1:0] node2351;
	wire [16-1:0] node2352;
	wire [16-1:0] node2354;
	wire [16-1:0] node2356;
	wire [16-1:0] node2359;
	wire [16-1:0] node2360;
	wire [16-1:0] node2362;
	wire [16-1:0] node2365;
	wire [16-1:0] node2368;
	wire [16-1:0] node2369;
	wire [16-1:0] node2370;
	wire [16-1:0] node2372;
	wire [16-1:0] node2375;
	wire [16-1:0] node2378;
	wire [16-1:0] node2380;
	wire [16-1:0] node2383;
	wire [16-1:0] node2384;
	wire [16-1:0] node2385;
	wire [16-1:0] node2386;
	wire [16-1:0] node2387;
	wire [16-1:0] node2388;
	wire [16-1:0] node2389;
	wire [16-1:0] node2391;
	wire [16-1:0] node2394;
	wire [16-1:0] node2396;
	wire [16-1:0] node2399;
	wire [16-1:0] node2400;
	wire [16-1:0] node2404;
	wire [16-1:0] node2405;
	wire [16-1:0] node2406;
	wire [16-1:0] node2409;
	wire [16-1:0] node2412;
	wire [16-1:0] node2413;
	wire [16-1:0] node2417;
	wire [16-1:0] node2418;
	wire [16-1:0] node2419;
	wire [16-1:0] node2420;
	wire [16-1:0] node2424;
	wire [16-1:0] node2425;
	wire [16-1:0] node2427;
	wire [16-1:0] node2428;
	wire [16-1:0] node2432;
	wire [16-1:0] node2435;
	wire [16-1:0] node2436;
	wire [16-1:0] node2437;
	wire [16-1:0] node2439;
	wire [16-1:0] node2441;
	wire [16-1:0] node2444;
	wire [16-1:0] node2445;
	wire [16-1:0] node2447;
	wire [16-1:0] node2451;
	wire [16-1:0] node2452;
	wire [16-1:0] node2456;
	wire [16-1:0] node2457;
	wire [16-1:0] node2458;
	wire [16-1:0] node2459;
	wire [16-1:0] node2461;
	wire [16-1:0] node2463;
	wire [16-1:0] node2464;
	wire [16-1:0] node2468;
	wire [16-1:0] node2471;
	wire [16-1:0] node2472;
	wire [16-1:0] node2473;
	wire [16-1:0] node2474;
	wire [16-1:0] node2479;
	wire [16-1:0] node2480;
	wire [16-1:0] node2482;
	wire [16-1:0] node2485;
	wire [16-1:0] node2488;
	wire [16-1:0] node2489;
	wire [16-1:0] node2490;
	wire [16-1:0] node2493;
	wire [16-1:0] node2494;
	wire [16-1:0] node2497;
	wire [16-1:0] node2500;
	wire [16-1:0] node2501;
	wire [16-1:0] node2503;
	wire [16-1:0] node2505;
	wire [16-1:0] node2506;
	wire [16-1:0] node2510;
	wire [16-1:0] node2512;
	wire [16-1:0] node2513;
	wire [16-1:0] node2516;
	wire [16-1:0] node2518;
	wire [16-1:0] node2521;
	wire [16-1:0] node2522;
	wire [16-1:0] node2523;
	wire [16-1:0] node2524;
	wire [16-1:0] node2525;
	wire [16-1:0] node2527;
	wire [16-1:0] node2530;
	wire [16-1:0] node2531;
	wire [16-1:0] node2534;
	wire [16-1:0] node2535;
	wire [16-1:0] node2539;
	wire [16-1:0] node2540;
	wire [16-1:0] node2543;
	wire [16-1:0] node2544;
	wire [16-1:0] node2548;
	wire [16-1:0] node2549;
	wire [16-1:0] node2550;
	wire [16-1:0] node2551;
	wire [16-1:0] node2553;
	wire [16-1:0] node2557;
	wire [16-1:0] node2558;
	wire [16-1:0] node2562;
	wire [16-1:0] node2564;
	wire [16-1:0] node2565;
	wire [16-1:0] node2568;
	wire [16-1:0] node2571;
	wire [16-1:0] node2572;
	wire [16-1:0] node2573;
	wire [16-1:0] node2574;
	wire [16-1:0] node2575;
	wire [16-1:0] node2578;
	wire [16-1:0] node2581;
	wire [16-1:0] node2582;
	wire [16-1:0] node2586;
	wire [16-1:0] node2587;
	wire [16-1:0] node2588;
	wire [16-1:0] node2589;
	wire [16-1:0] node2593;
	wire [16-1:0] node2596;
	wire [16-1:0] node2597;
	wire [16-1:0] node2598;
	wire [16-1:0] node2600;
	wire [16-1:0] node2604;
	wire [16-1:0] node2607;
	wire [16-1:0] node2608;
	wire [16-1:0] node2609;
	wire [16-1:0] node2612;
	wire [16-1:0] node2613;
	wire [16-1:0] node2614;
	wire [16-1:0] node2618;
	wire [16-1:0] node2620;
	wire [16-1:0] node2623;
	wire [16-1:0] node2624;
	wire [16-1:0] node2625;
	wire [16-1:0] node2629;
	wire [16-1:0] node2631;
	wire [16-1:0] node2632;
	wire [16-1:0] node2635;
	wire [16-1:0] node2638;
	wire [16-1:0] node2639;
	wire [16-1:0] node2640;
	wire [16-1:0] node2641;
	wire [16-1:0] node2642;
	wire [16-1:0] node2643;
	wire [16-1:0] node2644;
	wire [16-1:0] node2645;
	wire [16-1:0] node2648;
	wire [16-1:0] node2649;
	wire [16-1:0] node2652;
	wire [16-1:0] node2655;
	wire [16-1:0] node2657;
	wire [16-1:0] node2660;
	wire [16-1:0] node2661;
	wire [16-1:0] node2664;
	wire [16-1:0] node2666;
	wire [16-1:0] node2667;
	wire [16-1:0] node2671;
	wire [16-1:0] node2672;
	wire [16-1:0] node2673;
	wire [16-1:0] node2674;
	wire [16-1:0] node2676;
	wire [16-1:0] node2677;
	wire [16-1:0] node2682;
	wire [16-1:0] node2683;
	wire [16-1:0] node2687;
	wire [16-1:0] node2688;
	wire [16-1:0] node2691;
	wire [16-1:0] node2692;
	wire [16-1:0] node2694;
	wire [16-1:0] node2698;
	wire [16-1:0] node2699;
	wire [16-1:0] node2700;
	wire [16-1:0] node2701;
	wire [16-1:0] node2703;
	wire [16-1:0] node2706;
	wire [16-1:0] node2707;
	wire [16-1:0] node2711;
	wire [16-1:0] node2712;
	wire [16-1:0] node2713;
	wire [16-1:0] node2716;
	wire [16-1:0] node2718;
	wire [16-1:0] node2722;
	wire [16-1:0] node2723;
	wire [16-1:0] node2724;
	wire [16-1:0] node2725;
	wire [16-1:0] node2726;
	wire [16-1:0] node2730;
	wire [16-1:0] node2733;
	wire [16-1:0] node2734;
	wire [16-1:0] node2737;
	wire [16-1:0] node2740;
	wire [16-1:0] node2741;
	wire [16-1:0] node2742;
	wire [16-1:0] node2743;
	wire [16-1:0] node2745;
	wire [16-1:0] node2749;
	wire [16-1:0] node2752;
	wire [16-1:0] node2754;
	wire [16-1:0] node2756;
	wire [16-1:0] node2759;
	wire [16-1:0] node2760;
	wire [16-1:0] node2761;
	wire [16-1:0] node2762;
	wire [16-1:0] node2763;
	wire [16-1:0] node2764;
	wire [16-1:0] node2765;
	wire [16-1:0] node2769;
	wire [16-1:0] node2771;
	wire [16-1:0] node2774;
	wire [16-1:0] node2775;
	wire [16-1:0] node2777;
	wire [16-1:0] node2779;
	wire [16-1:0] node2782;
	wire [16-1:0] node2783;
	wire [16-1:0] node2787;
	wire [16-1:0] node2788;
	wire [16-1:0] node2789;
	wire [16-1:0] node2792;
	wire [16-1:0] node2795;
	wire [16-1:0] node2796;
	wire [16-1:0] node2799;
	wire [16-1:0] node2801;
	wire [16-1:0] node2804;
	wire [16-1:0] node2805;
	wire [16-1:0] node2806;
	wire [16-1:0] node2807;
	wire [16-1:0] node2809;
	wire [16-1:0] node2812;
	wire [16-1:0] node2813;
	wire [16-1:0] node2817;
	wire [16-1:0] node2818;
	wire [16-1:0] node2819;
	wire [16-1:0] node2821;
	wire [16-1:0] node2824;
	wire [16-1:0] node2827;
	wire [16-1:0] node2828;
	wire [16-1:0] node2832;
	wire [16-1:0] node2833;
	wire [16-1:0] node2835;
	wire [16-1:0] node2839;
	wire [16-1:0] node2840;
	wire [16-1:0] node2841;
	wire [16-1:0] node2842;
	wire [16-1:0] node2843;
	wire [16-1:0] node2845;
	wire [16-1:0] node2849;
	wire [16-1:0] node2851;
	wire [16-1:0] node2854;
	wire [16-1:0] node2855;
	wire [16-1:0] node2856;
	wire [16-1:0] node2859;
	wire [16-1:0] node2861;
	wire [16-1:0] node2864;
	wire [16-1:0] node2865;
	wire [16-1:0] node2866;
	wire [16-1:0] node2868;
	wire [16-1:0] node2872;
	wire [16-1:0] node2875;
	wire [16-1:0] node2876;
	wire [16-1:0] node2877;
	wire [16-1:0] node2879;
	wire [16-1:0] node2882;
	wire [16-1:0] node2883;
	wire [16-1:0] node2887;
	wire [16-1:0] node2888;
	wire [16-1:0] node2889;
	wire [16-1:0] node2892;
	wire [16-1:0] node2894;
	wire [16-1:0] node2897;
	wire [16-1:0] node2898;
	wire [16-1:0] node2901;
	wire [16-1:0] node2904;
	wire [16-1:0] node2905;
	wire [16-1:0] node2906;
	wire [16-1:0] node2907;
	wire [16-1:0] node2908;
	wire [16-1:0] node2910;
	wire [16-1:0] node2911;
	wire [16-1:0] node2915;
	wire [16-1:0] node2916;
	wire [16-1:0] node2917;
	wire [16-1:0] node2918;
	wire [16-1:0] node2919;
	wire [16-1:0] node2924;
	wire [16-1:0] node2927;
	wire [16-1:0] node2928;
	wire [16-1:0] node2930;
	wire [16-1:0] node2933;
	wire [16-1:0] node2935;
	wire [16-1:0] node2938;
	wire [16-1:0] node2939;
	wire [16-1:0] node2940;
	wire [16-1:0] node2942;
	wire [16-1:0] node2943;
	wire [16-1:0] node2946;
	wire [16-1:0] node2947;
	wire [16-1:0] node2951;
	wire [16-1:0] node2952;
	wire [16-1:0] node2955;
	wire [16-1:0] node2958;
	wire [16-1:0] node2959;
	wire [16-1:0] node2960;
	wire [16-1:0] node2964;
	wire [16-1:0] node2965;
	wire [16-1:0] node2968;
	wire [16-1:0] node2969;
	wire [16-1:0] node2971;
	wire [16-1:0] node2975;
	wire [16-1:0] node2976;
	wire [16-1:0] node2977;
	wire [16-1:0] node2978;
	wire [16-1:0] node2980;
	wire [16-1:0] node2981;
	wire [16-1:0] node2985;
	wire [16-1:0] node2986;
	wire [16-1:0] node2989;
	wire [16-1:0] node2990;
	wire [16-1:0] node2992;
	wire [16-1:0] node2996;
	wire [16-1:0] node2997;
	wire [16-1:0] node2998;
	wire [16-1:0] node2999;
	wire [16-1:0] node3004;
	wire [16-1:0] node3005;
	wire [16-1:0] node3006;
	wire [16-1:0] node3008;
	wire [16-1:0] node3012;
	wire [16-1:0] node3015;
	wire [16-1:0] node3016;
	wire [16-1:0] node3017;
	wire [16-1:0] node3019;
	wire [16-1:0] node3022;
	wire [16-1:0] node3024;
	wire [16-1:0] node3027;
	wire [16-1:0] node3028;
	wire [16-1:0] node3030;
	wire [16-1:0] node3031;
	wire [16-1:0] node3035;
	wire [16-1:0] node3036;
	wire [16-1:0] node3040;
	wire [16-1:0] node3041;
	wire [16-1:0] node3042;
	wire [16-1:0] node3043;
	wire [16-1:0] node3044;
	wire [16-1:0] node3045;
	wire [16-1:0] node3046;
	wire [16-1:0] node3050;
	wire [16-1:0] node3053;
	wire [16-1:0] node3054;
	wire [16-1:0] node3055;
	wire [16-1:0] node3059;
	wire [16-1:0] node3062;
	wire [16-1:0] node3064;
	wire [16-1:0] node3065;
	wire [16-1:0] node3066;
	wire [16-1:0] node3069;
	wire [16-1:0] node3070;
	wire [16-1:0] node3074;
	wire [16-1:0] node3077;
	wire [16-1:0] node3078;
	wire [16-1:0] node3079;
	wire [16-1:0] node3081;
	wire [16-1:0] node3083;
	wire [16-1:0] node3084;
	wire [16-1:0] node3088;
	wire [16-1:0] node3090;
	wire [16-1:0] node3091;
	wire [16-1:0] node3092;
	wire [16-1:0] node3097;
	wire [16-1:0] node3098;
	wire [16-1:0] node3099;
	wire [16-1:0] node3100;
	wire [16-1:0] node3105;
	wire [16-1:0] node3107;
	wire [16-1:0] node3109;
	wire [16-1:0] node3112;
	wire [16-1:0] node3113;
	wire [16-1:0] node3114;
	wire [16-1:0] node3115;
	wire [16-1:0] node3118;
	wire [16-1:0] node3119;
	wire [16-1:0] node3122;
	wire [16-1:0] node3125;
	wire [16-1:0] node3126;
	wire [16-1:0] node3128;
	wire [16-1:0] node3132;
	wire [16-1:0] node3133;
	wire [16-1:0] node3134;
	wire [16-1:0] node3136;
	wire [16-1:0] node3138;
	wire [16-1:0] node3139;
	wire [16-1:0] node3144;
	wire [16-1:0] node3145;
	wire [16-1:0] node3147;
	wire [16-1:0] node3149;
	wire [16-1:0] node3150;
	wire [16-1:0] node3154;
	wire [16-1:0] node3155;
	wire [16-1:0] node3158;
	wire [16-1:0] node3161;
	wire [16-1:0] node3162;
	wire [16-1:0] node3163;
	wire [16-1:0] node3164;
	wire [16-1:0] node3165;
	wire [16-1:0] node3166;
	wire [16-1:0] node3167;
	wire [16-1:0] node3168;
	wire [16-1:0] node3169;
	wire [16-1:0] node3172;
	wire [16-1:0] node3173;
	wire [16-1:0] node3177;
	wire [16-1:0] node3178;
	wire [16-1:0] node3181;
	wire [16-1:0] node3184;
	wire [16-1:0] node3185;
	wire [16-1:0] node3186;
	wire [16-1:0] node3189;
	wire [16-1:0] node3191;
	wire [16-1:0] node3192;
	wire [16-1:0] node3196;
	wire [16-1:0] node3197;
	wire [16-1:0] node3200;
	wire [16-1:0] node3203;
	wire [16-1:0] node3204;
	wire [16-1:0] node3205;
	wire [16-1:0] node3207;
	wire [16-1:0] node3210;
	wire [16-1:0] node3211;
	wire [16-1:0] node3214;
	wire [16-1:0] node3217;
	wire [16-1:0] node3218;
	wire [16-1:0] node3219;
	wire [16-1:0] node3220;
	wire [16-1:0] node3224;
	wire [16-1:0] node3226;
	wire [16-1:0] node3229;
	wire [16-1:0] node3230;
	wire [16-1:0] node3234;
	wire [16-1:0] node3235;
	wire [16-1:0] node3236;
	wire [16-1:0] node3237;
	wire [16-1:0] node3239;
	wire [16-1:0] node3242;
	wire [16-1:0] node3245;
	wire [16-1:0] node3248;
	wire [16-1:0] node3249;
	wire [16-1:0] node3250;
	wire [16-1:0] node3251;
	wire [16-1:0] node3254;
	wire [16-1:0] node3257;
	wire [16-1:0] node3259;
	wire [16-1:0] node3262;
	wire [16-1:0] node3263;
	wire [16-1:0] node3265;
	wire [16-1:0] node3268;
	wire [16-1:0] node3270;
	wire [16-1:0] node3273;
	wire [16-1:0] node3274;
	wire [16-1:0] node3275;
	wire [16-1:0] node3276;
	wire [16-1:0] node3277;
	wire [16-1:0] node3280;
	wire [16-1:0] node3281;
	wire [16-1:0] node3285;
	wire [16-1:0] node3286;
	wire [16-1:0] node3287;
	wire [16-1:0] node3291;
	wire [16-1:0] node3293;
	wire [16-1:0] node3296;
	wire [16-1:0] node3297;
	wire [16-1:0] node3298;
	wire [16-1:0] node3299;
	wire [16-1:0] node3302;
	wire [16-1:0] node3304;
	wire [16-1:0] node3308;
	wire [16-1:0] node3309;
	wire [16-1:0] node3311;
	wire [16-1:0] node3314;
	wire [16-1:0] node3317;
	wire [16-1:0] node3318;
	wire [16-1:0] node3319;
	wire [16-1:0] node3320;
	wire [16-1:0] node3321;
	wire [16-1:0] node3322;
	wire [16-1:0] node3326;
	wire [16-1:0] node3327;
	wire [16-1:0] node3332;
	wire [16-1:0] node3333;
	wire [16-1:0] node3334;
	wire [16-1:0] node3335;
	wire [16-1:0] node3339;
	wire [16-1:0] node3342;
	wire [16-1:0] node3343;
	wire [16-1:0] node3346;
	wire [16-1:0] node3347;
	wire [16-1:0] node3349;
	wire [16-1:0] node3352;
	wire [16-1:0] node3353;
	wire [16-1:0] node3357;
	wire [16-1:0] node3358;
	wire [16-1:0] node3359;
	wire [16-1:0] node3360;
	wire [16-1:0] node3364;
	wire [16-1:0] node3367;
	wire [16-1:0] node3368;
	wire [16-1:0] node3369;
	wire [16-1:0] node3372;
	wire [16-1:0] node3374;
	wire [16-1:0] node3377;
	wire [16-1:0] node3379;
	wire [16-1:0] node3380;
	wire [16-1:0] node3384;
	wire [16-1:0] node3385;
	wire [16-1:0] node3386;
	wire [16-1:0] node3387;
	wire [16-1:0] node3388;
	wire [16-1:0] node3389;
	wire [16-1:0] node3390;
	wire [16-1:0] node3394;
	wire [16-1:0] node3396;
	wire [16-1:0] node3399;
	wire [16-1:0] node3401;
	wire [16-1:0] node3402;
	wire [16-1:0] node3403;
	wire [16-1:0] node3407;
	wire [16-1:0] node3410;
	wire [16-1:0] node3411;
	wire [16-1:0] node3412;
	wire [16-1:0] node3413;
	wire [16-1:0] node3414;
	wire [16-1:0] node3416;
	wire [16-1:0] node3421;
	wire [16-1:0] node3422;
	wire [16-1:0] node3424;
	wire [16-1:0] node3427;
	wire [16-1:0] node3430;
	wire [16-1:0] node3431;
	wire [16-1:0] node3433;
	wire [16-1:0] node3437;
	wire [16-1:0] node3438;
	wire [16-1:0] node3439;
	wire [16-1:0] node3441;
	wire [16-1:0] node3442;
	wire [16-1:0] node3444;
	wire [16-1:0] node3448;
	wire [16-1:0] node3449;
	wire [16-1:0] node3450;
	wire [16-1:0] node3451;
	wire [16-1:0] node3455;
	wire [16-1:0] node3456;
	wire [16-1:0] node3459;
	wire [16-1:0] node3460;
	wire [16-1:0] node3464;
	wire [16-1:0] node3466;
	wire [16-1:0] node3469;
	wire [16-1:0] node3470;
	wire [16-1:0] node3471;
	wire [16-1:0] node3472;
	wire [16-1:0] node3475;
	wire [16-1:0] node3476;
	wire [16-1:0] node3480;
	wire [16-1:0] node3482;
	wire [16-1:0] node3485;
	wire [16-1:0] node3486;
	wire [16-1:0] node3488;
	wire [16-1:0] node3489;
	wire [16-1:0] node3493;
	wire [16-1:0] node3496;
	wire [16-1:0] node3497;
	wire [16-1:0] node3498;
	wire [16-1:0] node3499;
	wire [16-1:0] node3500;
	wire [16-1:0] node3501;
	wire [16-1:0] node3502;
	wire [16-1:0] node3507;
	wire [16-1:0] node3508;
	wire [16-1:0] node3512;
	wire [16-1:0] node3514;
	wire [16-1:0] node3515;
	wire [16-1:0] node3517;
	wire [16-1:0] node3520;
	wire [16-1:0] node3523;
	wire [16-1:0] node3524;
	wire [16-1:0] node3526;
	wire [16-1:0] node3527;
	wire [16-1:0] node3528;
	wire [16-1:0] node3530;
	wire [16-1:0] node3534;
	wire [16-1:0] node3537;
	wire [16-1:0] node3538;
	wire [16-1:0] node3540;
	wire [16-1:0] node3541;
	wire [16-1:0] node3543;
	wire [16-1:0] node3547;
	wire [16-1:0] node3548;
	wire [16-1:0] node3550;
	wire [16-1:0] node3551;
	wire [16-1:0] node3555;
	wire [16-1:0] node3557;
	wire [16-1:0] node3560;
	wire [16-1:0] node3561;
	wire [16-1:0] node3562;
	wire [16-1:0] node3563;
	wire [16-1:0] node3564;
	wire [16-1:0] node3565;
	wire [16-1:0] node3569;
	wire [16-1:0] node3572;
	wire [16-1:0] node3573;
	wire [16-1:0] node3576;
	wire [16-1:0] node3577;
	wire [16-1:0] node3580;
	wire [16-1:0] node3582;
	wire [16-1:0] node3585;
	wire [16-1:0] node3586;
	wire [16-1:0] node3588;
	wire [16-1:0] node3591;
	wire [16-1:0] node3592;
	wire [16-1:0] node3595;
	wire [16-1:0] node3598;
	wire [16-1:0] node3599;
	wire [16-1:0] node3600;
	wire [16-1:0] node3602;
	wire [16-1:0] node3604;
	wire [16-1:0] node3605;
	wire [16-1:0] node3610;
	wire [16-1:0] node3611;
	wire [16-1:0] node3612;
	wire [16-1:0] node3613;
	wire [16-1:0] node3617;
	wire [16-1:0] node3620;
	wire [16-1:0] node3621;
	wire [16-1:0] node3624;
	wire [16-1:0] node3627;
	wire [16-1:0] node3628;
	wire [16-1:0] node3629;
	wire [16-1:0] node3630;
	wire [16-1:0] node3631;
	wire [16-1:0] node3632;
	wire [16-1:0] node3633;
	wire [16-1:0] node3634;
	wire [16-1:0] node3635;
	wire [16-1:0] node3639;
	wire [16-1:0] node3642;
	wire [16-1:0] node3643;
	wire [16-1:0] node3645;
	wire [16-1:0] node3648;
	wire [16-1:0] node3650;
	wire [16-1:0] node3653;
	wire [16-1:0] node3654;
	wire [16-1:0] node3656;
	wire [16-1:0] node3659;
	wire [16-1:0] node3660;
	wire [16-1:0] node3661;
	wire [16-1:0] node3663;
	wire [16-1:0] node3668;
	wire [16-1:0] node3669;
	wire [16-1:0] node3670;
	wire [16-1:0] node3673;
	wire [16-1:0] node3674;
	wire [16-1:0] node3676;
	wire [16-1:0] node3677;
	wire [16-1:0] node3681;
	wire [16-1:0] node3683;
	wire [16-1:0] node3686;
	wire [16-1:0] node3687;
	wire [16-1:0] node3688;
	wire [16-1:0] node3689;
	wire [16-1:0] node3694;
	wire [16-1:0] node3695;
	wire [16-1:0] node3697;
	wire [16-1:0] node3701;
	wire [16-1:0] node3702;
	wire [16-1:0] node3703;
	wire [16-1:0] node3704;
	wire [16-1:0] node3706;
	wire [16-1:0] node3709;
	wire [16-1:0] node3710;
	wire [16-1:0] node3711;
	wire [16-1:0] node3715;
	wire [16-1:0] node3718;
	wire [16-1:0] node3719;
	wire [16-1:0] node3720;
	wire [16-1:0] node3724;
	wire [16-1:0] node3725;
	wire [16-1:0] node3729;
	wire [16-1:0] node3730;
	wire [16-1:0] node3731;
	wire [16-1:0] node3732;
	wire [16-1:0] node3735;
	wire [16-1:0] node3737;
	wire [16-1:0] node3740;
	wire [16-1:0] node3741;
	wire [16-1:0] node3744;
	wire [16-1:0] node3745;
	wire [16-1:0] node3749;
	wire [16-1:0] node3750;
	wire [16-1:0] node3753;
	wire [16-1:0] node3754;
	wire [16-1:0] node3755;
	wire [16-1:0] node3759;
	wire [16-1:0] node3762;
	wire [16-1:0] node3763;
	wire [16-1:0] node3764;
	wire [16-1:0] node3765;
	wire [16-1:0] node3766;
	wire [16-1:0] node3769;
	wire [16-1:0] node3770;
	wire [16-1:0] node3773;
	wire [16-1:0] node3776;
	wire [16-1:0] node3777;
	wire [16-1:0] node3778;
	wire [16-1:0] node3781;
	wire [16-1:0] node3784;
	wire [16-1:0] node3785;
	wire [16-1:0] node3787;
	wire [16-1:0] node3790;
	wire [16-1:0] node3793;
	wire [16-1:0] node3794;
	wire [16-1:0] node3795;
	wire [16-1:0] node3796;
	wire [16-1:0] node3797;
	wire [16-1:0] node3798;
	wire [16-1:0] node3802;
	wire [16-1:0] node3805;
	wire [16-1:0] node3808;
	wire [16-1:0] node3809;
	wire [16-1:0] node3812;
	wire [16-1:0] node3813;
	wire [16-1:0] node3815;
	wire [16-1:0] node3819;
	wire [16-1:0] node3820;
	wire [16-1:0] node3821;
	wire [16-1:0] node3822;
	wire [16-1:0] node3826;
	wire [16-1:0] node3827;
	wire [16-1:0] node3831;
	wire [16-1:0] node3833;
	wire [16-1:0] node3836;
	wire [16-1:0] node3837;
	wire [16-1:0] node3838;
	wire [16-1:0] node3839;
	wire [16-1:0] node3842;
	wire [16-1:0] node3843;
	wire [16-1:0] node3844;
	wire [16-1:0] node3848;
	wire [16-1:0] node3849;
	wire [16-1:0] node3853;
	wire [16-1:0] node3854;
	wire [16-1:0] node3858;
	wire [16-1:0] node3859;
	wire [16-1:0] node3860;
	wire [16-1:0] node3861;
	wire [16-1:0] node3862;
	wire [16-1:0] node3865;
	wire [16-1:0] node3866;
	wire [16-1:0] node3871;
	wire [16-1:0] node3872;
	wire [16-1:0] node3875;
	wire [16-1:0] node3876;
	wire [16-1:0] node3878;
	wire [16-1:0] node3882;
	wire [16-1:0] node3884;
	wire [16-1:0] node3885;
	wire [16-1:0] node3888;
	wire [16-1:0] node3891;
	wire [16-1:0] node3892;
	wire [16-1:0] node3893;
	wire [16-1:0] node3894;
	wire [16-1:0] node3895;
	wire [16-1:0] node3896;
	wire [16-1:0] node3898;
	wire [16-1:0] node3901;
	wire [16-1:0] node3902;
	wire [16-1:0] node3905;
	wire [16-1:0] node3908;
	wire [16-1:0] node3909;
	wire [16-1:0] node3910;
	wire [16-1:0] node3913;
	wire [16-1:0] node3914;
	wire [16-1:0] node3916;
	wire [16-1:0] node3920;
	wire [16-1:0] node3921;
	wire [16-1:0] node3922;
	wire [16-1:0] node3926;
	wire [16-1:0] node3929;
	wire [16-1:0] node3930;
	wire [16-1:0] node3931;
	wire [16-1:0] node3934;
	wire [16-1:0] node3935;
	wire [16-1:0] node3938;
	wire [16-1:0] node3940;
	wire [16-1:0] node3943;
	wire [16-1:0] node3944;
	wire [16-1:0] node3945;
	wire [16-1:0] node3948;
	wire [16-1:0] node3949;
	wire [16-1:0] node3953;
	wire [16-1:0] node3954;
	wire [16-1:0] node3957;
	wire [16-1:0] node3959;
	wire [16-1:0] node3962;
	wire [16-1:0] node3963;
	wire [16-1:0] node3964;
	wire [16-1:0] node3966;
	wire [16-1:0] node3967;
	wire [16-1:0] node3971;
	wire [16-1:0] node3973;
	wire [16-1:0] node3974;
	wire [16-1:0] node3975;
	wire [16-1:0] node3979;
	wire [16-1:0] node3981;
	wire [16-1:0] node3984;
	wire [16-1:0] node3985;
	wire [16-1:0] node3986;
	wire [16-1:0] node3987;
	wire [16-1:0] node3991;
	wire [16-1:0] node3992;
	wire [16-1:0] node3993;
	wire [16-1:0] node3995;
	wire [16-1:0] node3999;
	wire [16-1:0] node4002;
	wire [16-1:0] node4003;
	wire [16-1:0] node4004;
	wire [16-1:0] node4006;
	wire [16-1:0] node4010;
	wire [16-1:0] node4013;
	wire [16-1:0] node4014;
	wire [16-1:0] node4015;
	wire [16-1:0] node4016;
	wire [16-1:0] node4017;
	wire [16-1:0] node4018;
	wire [16-1:0] node4019;
	wire [16-1:0] node4020;
	wire [16-1:0] node4025;
	wire [16-1:0] node4026;
	wire [16-1:0] node4029;
	wire [16-1:0] node4030;
	wire [16-1:0] node4034;
	wire [16-1:0] node4037;
	wire [16-1:0] node4038;
	wire [16-1:0] node4039;
	wire [16-1:0] node4041;
	wire [16-1:0] node4044;
	wire [16-1:0] node4045;
	wire [16-1:0] node4049;
	wire [16-1:0] node4050;
	wire [16-1:0] node4051;
	wire [16-1:0] node4055;
	wire [16-1:0] node4057;
	wire [16-1:0] node4060;
	wire [16-1:0] node4061;
	wire [16-1:0] node4062;
	wire [16-1:0] node4064;
	wire [16-1:0] node4065;
	wire [16-1:0] node4069;
	wire [16-1:0] node4070;
	wire [16-1:0] node4073;
	wire [16-1:0] node4075;
	wire [16-1:0] node4076;
	wire [16-1:0] node4080;
	wire [16-1:0] node4081;
	wire [16-1:0] node4082;
	wire [16-1:0] node4083;
	wire [16-1:0] node4087;
	wire [16-1:0] node4090;
	wire [16-1:0] node4091;
	wire [16-1:0] node4093;
	wire [16-1:0] node4097;
	wire [16-1:0] node4098;
	wire [16-1:0] node4099;
	wire [16-1:0] node4100;
	wire [16-1:0] node4102;
	wire [16-1:0] node4104;
	wire [16-1:0] node4105;
	wire [16-1:0] node4109;
	wire [16-1:0] node4112;
	wire [16-1:0] node4113;
	wire [16-1:0] node4115;
	wire [16-1:0] node4118;
	wire [16-1:0] node4119;
	wire [16-1:0] node4123;
	wire [16-1:0] node4124;
	wire [16-1:0] node4126;
	wire [16-1:0] node4127;
	wire [16-1:0] node4129;
	wire [16-1:0] node4132;
	wire [16-1:0] node4135;
	wire [16-1:0] node4136;
	wire [16-1:0] node4137;
	wire [16-1:0] node4140;
	wire [16-1:0] node4143;
	wire [16-1:0] node4144;
	wire [16-1:0] node4145;
	wire [16-1:0] node4147;
	wire [16-1:0] node4151;
	wire [16-1:0] node4152;
	wire [16-1:0] node4156;
	wire [16-1:0] node4157;
	wire [16-1:0] node4158;
	wire [16-1:0] node4159;
	wire [16-1:0] node4160;
	wire [16-1:0] node4161;
	wire [16-1:0] node4162;
	wire [16-1:0] node4163;
	wire [16-1:0] node4164;
	wire [16-1:0] node4165;
	wire [16-1:0] node4166;
	wire [16-1:0] node4167;
	wire [16-1:0] node4171;
	wire [16-1:0] node4174;
	wire [16-1:0] node4175;
	wire [16-1:0] node4176;
	wire [16-1:0] node4180;
	wire [16-1:0] node4183;
	wire [16-1:0] node4184;
	wire [16-1:0] node4187;
	wire [16-1:0] node4188;
	wire [16-1:0] node4191;
	wire [16-1:0] node4193;
	wire [16-1:0] node4194;
	wire [16-1:0] node4198;
	wire [16-1:0] node4199;
	wire [16-1:0] node4200;
	wire [16-1:0] node4202;
	wire [16-1:0] node4203;
	wire [16-1:0] node4208;
	wire [16-1:0] node4210;
	wire [16-1:0] node4211;
	wire [16-1:0] node4214;
	wire [16-1:0] node4216;
	wire [16-1:0] node4219;
	wire [16-1:0] node4220;
	wire [16-1:0] node4221;
	wire [16-1:0] node4222;
	wire [16-1:0] node4224;
	wire [16-1:0] node4226;
	wire [16-1:0] node4229;
	wire [16-1:0] node4230;
	wire [16-1:0] node4234;
	wire [16-1:0] node4235;
	wire [16-1:0] node4236;
	wire [16-1:0] node4238;
	wire [16-1:0] node4241;
	wire [16-1:0] node4242;
	wire [16-1:0] node4246;
	wire [16-1:0] node4247;
	wire [16-1:0] node4250;
	wire [16-1:0] node4253;
	wire [16-1:0] node4254;
	wire [16-1:0] node4255;
	wire [16-1:0] node4256;
	wire [16-1:0] node4257;
	wire [16-1:0] node4260;
	wire [16-1:0] node4263;
	wire [16-1:0] node4266;
	wire [16-1:0] node4267;
	wire [16-1:0] node4270;
	wire [16-1:0] node4271;
	wire [16-1:0] node4273;
	wire [16-1:0] node4277;
	wire [16-1:0] node4278;
	wire [16-1:0] node4279;
	wire [16-1:0] node4280;
	wire [16-1:0] node4285;
	wire [16-1:0] node4288;
	wire [16-1:0] node4289;
	wire [16-1:0] node4290;
	wire [16-1:0] node4291;
	wire [16-1:0] node4292;
	wire [16-1:0] node4294;
	wire [16-1:0] node4297;
	wire [16-1:0] node4298;
	wire [16-1:0] node4300;
	wire [16-1:0] node4301;
	wire [16-1:0] node4306;
	wire [16-1:0] node4307;
	wire [16-1:0] node4308;
	wire [16-1:0] node4311;
	wire [16-1:0] node4312;
	wire [16-1:0] node4314;
	wire [16-1:0] node4318;
	wire [16-1:0] node4319;
	wire [16-1:0] node4320;
	wire [16-1:0] node4325;
	wire [16-1:0] node4326;
	wire [16-1:0] node4327;
	wire [16-1:0] node4329;
	wire [16-1:0] node4332;
	wire [16-1:0] node4333;
	wire [16-1:0] node4336;
	wire [16-1:0] node4337;
	wire [16-1:0] node4339;
	wire [16-1:0] node4343;
	wire [16-1:0] node4344;
	wire [16-1:0] node4346;
	wire [16-1:0] node4349;
	wire [16-1:0] node4351;
	wire [16-1:0] node4354;
	wire [16-1:0] node4355;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4359;
	wire [16-1:0] node4361;
	wire [16-1:0] node4362;
	wire [16-1:0] node4366;
	wire [16-1:0] node4367;
	wire [16-1:0] node4368;
	wire [16-1:0] node4372;
	wire [16-1:0] node4373;
	wire [16-1:0] node4377;
	wire [16-1:0] node4379;
	wire [16-1:0] node4380;
	wire [16-1:0] node4381;
	wire [16-1:0] node4383;
	wire [16-1:0] node4388;
	wire [16-1:0] node4389;
	wire [16-1:0] node4390;
	wire [16-1:0] node4391;
	wire [16-1:0] node4392;
	wire [16-1:0] node4394;
	wire [16-1:0] node4398;
	wire [16-1:0] node4401;
	wire [16-1:0] node4402;
	wire [16-1:0] node4406;
	wire [16-1:0] node4407;
	wire [16-1:0] node4408;
	wire [16-1:0] node4412;
	wire [16-1:0] node4413;
	wire [16-1:0] node4414;
	wire [16-1:0] node4416;
	wire [16-1:0] node4420;
	wire [16-1:0] node4423;
	wire [16-1:0] node4424;
	wire [16-1:0] node4425;
	wire [16-1:0] node4426;
	wire [16-1:0] node4427;
	wire [16-1:0] node4428;
	wire [16-1:0] node4429;
	wire [16-1:0] node4431;
	wire [16-1:0] node4434;
	wire [16-1:0] node4435;
	wire [16-1:0] node4438;
	wire [16-1:0] node4439;
	wire [16-1:0] node4443;
	wire [16-1:0] node4444;
	wire [16-1:0] node4446;
	wire [16-1:0] node4449;
	wire [16-1:0] node4450;
	wire [16-1:0] node4451;
	wire [16-1:0] node4456;
	wire [16-1:0] node4457;
	wire [16-1:0] node4458;
	wire [16-1:0] node4461;
	wire [16-1:0] node4463;
	wire [16-1:0] node4466;
	wire [16-1:0] node4468;
	wire [16-1:0] node4470;
	wire [16-1:0] node4473;
	wire [16-1:0] node4474;
	wire [16-1:0] node4475;
	wire [16-1:0] node4476;
	wire [16-1:0] node4477;
	wire [16-1:0] node4483;
	wire [16-1:0] node4484;
	wire [16-1:0] node4485;
	wire [16-1:0] node4490;
	wire [16-1:0] node4491;
	wire [16-1:0] node4492;
	wire [16-1:0] node4493;
	wire [16-1:0] node4494;
	wire [16-1:0] node4497;
	wire [16-1:0] node4500;
	wire [16-1:0] node4501;
	wire [16-1:0] node4505;
	wire [16-1:0] node4506;
	wire [16-1:0] node4507;
	wire [16-1:0] node4510;
	wire [16-1:0] node4512;
	wire [16-1:0] node4515;
	wire [16-1:0] node4516;
	wire [16-1:0] node4517;
	wire [16-1:0] node4519;
	wire [16-1:0] node4523;
	wire [16-1:0] node4525;
	wire [16-1:0] node4528;
	wire [16-1:0] node4529;
	wire [16-1:0] node4530;
	wire [16-1:0] node4531;
	wire [16-1:0] node4532;
	wire [16-1:0] node4536;
	wire [16-1:0] node4540;
	wire [16-1:0] node4541;
	wire [16-1:0] node4542;
	wire [16-1:0] node4544;
	wire [16-1:0] node4545;
	wire [16-1:0] node4550;
	wire [16-1:0] node4551;
	wire [16-1:0] node4555;
	wire [16-1:0] node4556;
	wire [16-1:0] node4557;
	wire [16-1:0] node4558;
	wire [16-1:0] node4559;
	wire [16-1:0] node4560;
	wire [16-1:0] node4563;
	wire [16-1:0] node4567;
	wire [16-1:0] node4568;
	wire [16-1:0] node4569;
	wire [16-1:0] node4572;
	wire [16-1:0] node4575;
	wire [16-1:0] node4576;
	wire [16-1:0] node4579;
	wire [16-1:0] node4582;
	wire [16-1:0] node4583;
	wire [16-1:0] node4584;
	wire [16-1:0] node4586;
	wire [16-1:0] node4588;
	wire [16-1:0] node4591;
	wire [16-1:0] node4592;
	wire [16-1:0] node4594;
	wire [16-1:0] node4597;
	wire [16-1:0] node4599;
	wire [16-1:0] node4602;
	wire [16-1:0] node4603;
	wire [16-1:0] node4604;
	wire [16-1:0] node4607;
	wire [16-1:0] node4609;
	wire [16-1:0] node4612;
	wire [16-1:0] node4613;
	wire [16-1:0] node4616;
	wire [16-1:0] node4619;
	wire [16-1:0] node4620;
	wire [16-1:0] node4621;
	wire [16-1:0] node4622;
	wire [16-1:0] node4623;
	wire [16-1:0] node4626;
	wire [16-1:0] node4629;
	wire [16-1:0] node4630;
	wire [16-1:0] node4631;
	wire [16-1:0] node4636;
	wire [16-1:0] node4638;
	wire [16-1:0] node4640;
	wire [16-1:0] node4642;
	wire [16-1:0] node4645;
	wire [16-1:0] node4646;
	wire [16-1:0] node4647;
	wire [16-1:0] node4649;
	wire [16-1:0] node4652;
	wire [16-1:0] node4654;
	wire [16-1:0] node4655;
	wire [16-1:0] node4656;
	wire [16-1:0] node4661;
	wire [16-1:0] node4662;
	wire [16-1:0] node4663;
	wire [16-1:0] node4665;
	wire [16-1:0] node4668;
	wire [16-1:0] node4670;
	wire [16-1:0] node4671;
	wire [16-1:0] node4675;
	wire [16-1:0] node4677;
	wire [16-1:0] node4679;
	wire [16-1:0] node4680;
	wire [16-1:0] node4684;
	wire [16-1:0] node4685;
	wire [16-1:0] node4686;
	wire [16-1:0] node4687;
	wire [16-1:0] node4688;
	wire [16-1:0] node4689;
	wire [16-1:0] node4690;
	wire [16-1:0] node4691;
	wire [16-1:0] node4692;
	wire [16-1:0] node4697;
	wire [16-1:0] node4698;
	wire [16-1:0] node4702;
	wire [16-1:0] node4703;
	wire [16-1:0] node4704;
	wire [16-1:0] node4708;
	wire [16-1:0] node4709;
	wire [16-1:0] node4711;
	wire [16-1:0] node4715;
	wire [16-1:0] node4716;
	wire [16-1:0] node4717;
	wire [16-1:0] node4718;
	wire [16-1:0] node4719;
	wire [16-1:0] node4723;
	wire [16-1:0] node4724;
	wire [16-1:0] node4725;
	wire [16-1:0] node4728;
	wire [16-1:0] node4732;
	wire [16-1:0] node4733;
	wire [16-1:0] node4735;
	wire [16-1:0] node4736;
	wire [16-1:0] node4740;
	wire [16-1:0] node4742;
	wire [16-1:0] node4745;
	wire [16-1:0] node4746;
	wire [16-1:0] node4748;
	wire [16-1:0] node4752;
	wire [16-1:0] node4753;
	wire [16-1:0] node4754;
	wire [16-1:0] node4755;
	wire [16-1:0] node4756;
	wire [16-1:0] node4758;
	wire [16-1:0] node4761;
	wire [16-1:0] node4762;
	wire [16-1:0] node4765;
	wire [16-1:0] node4766;
	wire [16-1:0] node4770;
	wire [16-1:0] node4772;
	wire [16-1:0] node4774;
	wire [16-1:0] node4777;
	wire [16-1:0] node4778;
	wire [16-1:0] node4779;
	wire [16-1:0] node4783;
	wire [16-1:0] node4785;
	wire [16-1:0] node4786;
	wire [16-1:0] node4790;
	wire [16-1:0] node4791;
	wire [16-1:0] node4792;
	wire [16-1:0] node4793;
	wire [16-1:0] node4796;
	wire [16-1:0] node4799;
	wire [16-1:0] node4801;
	wire [16-1:0] node4803;
	wire [16-1:0] node4806;
	wire [16-1:0] node4807;
	wire [16-1:0] node4809;
	wire [16-1:0] node4810;
	wire [16-1:0] node4814;
	wire [16-1:0] node4816;
	wire [16-1:0] node4819;
	wire [16-1:0] node4820;
	wire [16-1:0] node4821;
	wire [16-1:0] node4822;
	wire [16-1:0] node4823;
	wire [16-1:0] node4826;
	wire [16-1:0] node4827;
	wire [16-1:0] node4830;
	wire [16-1:0] node4832;
	wire [16-1:0] node4833;
	wire [16-1:0] node4837;
	wire [16-1:0] node4839;
	wire [16-1:0] node4840;
	wire [16-1:0] node4844;
	wire [16-1:0] node4845;
	wire [16-1:0] node4846;
	wire [16-1:0] node4847;
	wire [16-1:0] node4850;
	wire [16-1:0] node4852;
	wire [16-1:0] node4853;
	wire [16-1:0] node4857;
	wire [16-1:0] node4858;
	wire [16-1:0] node4862;
	wire [16-1:0] node4863;
	wire [16-1:0] node4864;
	wire [16-1:0] node4868;
	wire [16-1:0] node4870;
	wire [16-1:0] node4873;
	wire [16-1:0] node4874;
	wire [16-1:0] node4875;
	wire [16-1:0] node4876;
	wire [16-1:0] node4877;
	wire [16-1:0] node4878;
	wire [16-1:0] node4882;
	wire [16-1:0] node4885;
	wire [16-1:0] node4886;
	wire [16-1:0] node4889;
	wire [16-1:0] node4890;
	wire [16-1:0] node4892;
	wire [16-1:0] node4896;
	wire [16-1:0] node4897;
	wire [16-1:0] node4898;
	wire [16-1:0] node4901;
	wire [16-1:0] node4902;
	wire [16-1:0] node4904;
	wire [16-1:0] node4907;
	wire [16-1:0] node4908;
	wire [16-1:0] node4912;
	wire [16-1:0] node4913;
	wire [16-1:0] node4916;
	wire [16-1:0] node4917;
	wire [16-1:0] node4921;
	wire [16-1:0] node4922;
	wire [16-1:0] node4923;
	wire [16-1:0] node4926;
	wire [16-1:0] node4928;
	wire [16-1:0] node4929;
	wire [16-1:0] node4931;
	wire [16-1:0] node4935;
	wire [16-1:0] node4936;
	wire [16-1:0] node4937;
	wire [16-1:0] node4941;
	wire [16-1:0] node4942;
	wire [16-1:0] node4945;
	wire [16-1:0] node4947;
	wire [16-1:0] node4950;
	wire [16-1:0] node4951;
	wire [16-1:0] node4952;
	wire [16-1:0] node4953;
	wire [16-1:0] node4954;
	wire [16-1:0] node4955;
	wire [16-1:0] node4957;
	wire [16-1:0] node4958;
	wire [16-1:0] node4959;
	wire [16-1:0] node4965;
	wire [16-1:0] node4966;
	wire [16-1:0] node4967;
	wire [16-1:0] node4970;
	wire [16-1:0] node4972;
	wire [16-1:0] node4975;
	wire [16-1:0] node4976;
	wire [16-1:0] node4978;
	wire [16-1:0] node4981;
	wire [16-1:0] node4984;
	wire [16-1:0] node4985;
	wire [16-1:0] node4986;
	wire [16-1:0] node4989;
	wire [16-1:0] node4990;
	wire [16-1:0] node4992;
	wire [16-1:0] node4993;
	wire [16-1:0] node4998;
	wire [16-1:0] node4999;
	wire [16-1:0] node5000;
	wire [16-1:0] node5001;
	wire [16-1:0] node5005;
	wire [16-1:0] node5006;
	wire [16-1:0] node5011;
	wire [16-1:0] node5012;
	wire [16-1:0] node5013;
	wire [16-1:0] node5014;
	wire [16-1:0] node5017;
	wire [16-1:0] node5018;
	wire [16-1:0] node5022;
	wire [16-1:0] node5023;
	wire [16-1:0] node5024;
	wire [16-1:0] node5025;
	wire [16-1:0] node5030;
	wire [16-1:0] node5031;
	wire [16-1:0] node5033;
	wire [16-1:0] node5036;
	wire [16-1:0] node5037;
	wire [16-1:0] node5038;
	wire [16-1:0] node5043;
	wire [16-1:0] node5044;
	wire [16-1:0] node5045;
	wire [16-1:0] node5046;
	wire [16-1:0] node5049;
	wire [16-1:0] node5051;
	wire [16-1:0] node5052;
	wire [16-1:0] node5056;
	wire [16-1:0] node5057;
	wire [16-1:0] node5058;
	wire [16-1:0] node5061;
	wire [16-1:0] node5062;
	wire [16-1:0] node5066;
	wire [16-1:0] node5067;
	wire [16-1:0] node5069;
	wire [16-1:0] node5073;
	wire [16-1:0] node5074;
	wire [16-1:0] node5075;
	wire [16-1:0] node5077;
	wire [16-1:0] node5078;
	wire [16-1:0] node5082;
	wire [16-1:0] node5085;
	wire [16-1:0] node5087;
	wire [16-1:0] node5088;
	wire [16-1:0] node5089;
	wire [16-1:0] node5094;
	wire [16-1:0] node5095;
	wire [16-1:0] node5096;
	wire [16-1:0] node5097;
	wire [16-1:0] node5098;
	wire [16-1:0] node5099;
	wire [16-1:0] node5100;
	wire [16-1:0] node5102;
	wire [16-1:0] node5106;
	wire [16-1:0] node5109;
	wire [16-1:0] node5110;
	wire [16-1:0] node5111;
	wire [16-1:0] node5115;
	wire [16-1:0] node5118;
	wire [16-1:0] node5119;
	wire [16-1:0] node5123;
	wire [16-1:0] node5124;
	wire [16-1:0] node5125;
	wire [16-1:0] node5126;
	wire [16-1:0] node5127;
	wire [16-1:0] node5131;
	wire [16-1:0] node5135;
	wire [16-1:0] node5136;
	wire [16-1:0] node5137;
	wire [16-1:0] node5140;
	wire [16-1:0] node5142;
	wire [16-1:0] node5145;
	wire [16-1:0] node5146;
	wire [16-1:0] node5147;
	wire [16-1:0] node5149;
	wire [16-1:0] node5153;
	wire [16-1:0] node5155;
	wire [16-1:0] node5158;
	wire [16-1:0] node5159;
	wire [16-1:0] node5160;
	wire [16-1:0] node5161;
	wire [16-1:0] node5163;
	wire [16-1:0] node5164;
	wire [16-1:0] node5166;
	wire [16-1:0] node5169;
	wire [16-1:0] node5172;
	wire [16-1:0] node5174;
	wire [16-1:0] node5177;
	wire [16-1:0] node5178;
	wire [16-1:0] node5181;
	wire [16-1:0] node5183;
	wire [16-1:0] node5186;
	wire [16-1:0] node5187;
	wire [16-1:0] node5188;
	wire [16-1:0] node5191;
	wire [16-1:0] node5193;
	wire [16-1:0] node5196;
	wire [16-1:0] node5197;
	wire [16-1:0] node5198;
	wire [16-1:0] node5202;
	wire [16-1:0] node5203;
	wire [16-1:0] node5205;
	wire [16-1:0] node5209;
	wire [16-1:0] node5210;
	wire [16-1:0] node5211;
	wire [16-1:0] node5212;
	wire [16-1:0] node5213;
	wire [16-1:0] node5214;
	wire [16-1:0] node5215;
	wire [16-1:0] node5216;
	wire [16-1:0] node5217;
	wire [16-1:0] node5218;
	wire [16-1:0] node5220;
	wire [16-1:0] node5224;
	wire [16-1:0] node5225;
	wire [16-1:0] node5229;
	wire [16-1:0] node5231;
	wire [16-1:0] node5233;
	wire [16-1:0] node5234;
	wire [16-1:0] node5238;
	wire [16-1:0] node5239;
	wire [16-1:0] node5240;
	wire [16-1:0] node5242;
	wire [16-1:0] node5245;
	wire [16-1:0] node5246;
	wire [16-1:0] node5247;
	wire [16-1:0] node5252;
	wire [16-1:0] node5253;
	wire [16-1:0] node5254;
	wire [16-1:0] node5256;
	wire [16-1:0] node5260;
	wire [16-1:0] node5262;
	wire [16-1:0] node5265;
	wire [16-1:0] node5266;
	wire [16-1:0] node5267;
	wire [16-1:0] node5268;
	wire [16-1:0] node5271;
	wire [16-1:0] node5273;
	wire [16-1:0] node5274;
	wire [16-1:0] node5278;
	wire [16-1:0] node5279;
	wire [16-1:0] node5283;
	wire [16-1:0] node5285;
	wire [16-1:0] node5287;
	wire [16-1:0] node5290;
	wire [16-1:0] node5291;
	wire [16-1:0] node5292;
	wire [16-1:0] node5293;
	wire [16-1:0] node5294;
	wire [16-1:0] node5296;
	wire [16-1:0] node5297;
	wire [16-1:0] node5302;
	wire [16-1:0] node5303;
	wire [16-1:0] node5304;
	wire [16-1:0] node5306;
	wire [16-1:0] node5310;
	wire [16-1:0] node5313;
	wire [16-1:0] node5314;
	wire [16-1:0] node5315;
	wire [16-1:0] node5319;
	wire [16-1:0] node5320;
	wire [16-1:0] node5324;
	wire [16-1:0] node5325;
	wire [16-1:0] node5326;
	wire [16-1:0] node5327;
	wire [16-1:0] node5329;
	wire [16-1:0] node5332;
	wire [16-1:0] node5333;
	wire [16-1:0] node5337;
	wire [16-1:0] node5338;
	wire [16-1:0] node5339;
	wire [16-1:0] node5343;
	wire [16-1:0] node5346;
	wire [16-1:0] node5347;
	wire [16-1:0] node5348;
	wire [16-1:0] node5350;
	wire [16-1:0] node5352;
	wire [16-1:0] node5355;
	wire [16-1:0] node5358;
	wire [16-1:0] node5359;
	wire [16-1:0] node5361;
	wire [16-1:0] node5364;
	wire [16-1:0] node5365;
	wire [16-1:0] node5369;
	wire [16-1:0] node5370;
	wire [16-1:0] node5371;
	wire [16-1:0] node5372;
	wire [16-1:0] node5373;
	wire [16-1:0] node5374;
	wire [16-1:0] node5378;
	wire [16-1:0] node5379;
	wire [16-1:0] node5383;
	wire [16-1:0] node5385;
	wire [16-1:0] node5388;
	wire [16-1:0] node5389;
	wire [16-1:0] node5390;
	wire [16-1:0] node5391;
	wire [16-1:0] node5392;
	wire [16-1:0] node5396;
	wire [16-1:0] node5397;
	wire [16-1:0] node5399;
	wire [16-1:0] node5403;
	wire [16-1:0] node5404;
	wire [16-1:0] node5405;
	wire [16-1:0] node5407;
	wire [16-1:0] node5411;
	wire [16-1:0] node5414;
	wire [16-1:0] node5416;
	wire [16-1:0] node5417;
	wire [16-1:0] node5419;
	wire [16-1:0] node5422;
	wire [16-1:0] node5424;
	wire [16-1:0] node5427;
	wire [16-1:0] node5428;
	wire [16-1:0] node5429;
	wire [16-1:0] node5431;
	wire [16-1:0] node5432;
	wire [16-1:0] node5434;
	wire [16-1:0] node5438;
	wire [16-1:0] node5439;
	wire [16-1:0] node5440;
	wire [16-1:0] node5441;
	wire [16-1:0] node5445;
	wire [16-1:0] node5448;
	wire [16-1:0] node5449;
	wire [16-1:0] node5452;
	wire [16-1:0] node5453;
	wire [16-1:0] node5457;
	wire [16-1:0] node5458;
	wire [16-1:0] node5459;
	wire [16-1:0] node5461;
	wire [16-1:0] node5464;
	wire [16-1:0] node5465;
	wire [16-1:0] node5468;
	wire [16-1:0] node5471;
	wire [16-1:0] node5473;
	wire [16-1:0] node5474;
	wire [16-1:0] node5477;
	wire [16-1:0] node5479;
	wire [16-1:0] node5482;
	wire [16-1:0] node5483;
	wire [16-1:0] node5484;
	wire [16-1:0] node5485;
	wire [16-1:0] node5486;
	wire [16-1:0] node5487;
	wire [16-1:0] node5488;
	wire [16-1:0] node5490;
	wire [16-1:0] node5491;
	wire [16-1:0] node5496;
	wire [16-1:0] node5497;
	wire [16-1:0] node5498;
	wire [16-1:0] node5500;
	wire [16-1:0] node5504;
	wire [16-1:0] node5506;
	wire [16-1:0] node5509;
	wire [16-1:0] node5510;
	wire [16-1:0] node5511;
	wire [16-1:0] node5513;
	wire [16-1:0] node5514;
	wire [16-1:0] node5518;
	wire [16-1:0] node5519;
	wire [16-1:0] node5521;
	wire [16-1:0] node5525;
	wire [16-1:0] node5526;
	wire [16-1:0] node5527;
	wire [16-1:0] node5529;
	wire [16-1:0] node5532;
	wire [16-1:0] node5534;
	wire [16-1:0] node5537;
	wire [16-1:0] node5538;
	wire [16-1:0] node5540;
	wire [16-1:0] node5544;
	wire [16-1:0] node5545;
	wire [16-1:0] node5547;
	wire [16-1:0] node5548;
	wire [16-1:0] node5549;
	wire [16-1:0] node5553;
	wire [16-1:0] node5556;
	wire [16-1:0] node5557;
	wire [16-1:0] node5558;
	wire [16-1:0] node5561;
	wire [16-1:0] node5563;
	wire [16-1:0] node5566;
	wire [16-1:0] node5569;
	wire [16-1:0] node5570;
	wire [16-1:0] node5571;
	wire [16-1:0] node5572;
	wire [16-1:0] node5573;
	wire [16-1:0] node5575;
	wire [16-1:0] node5576;
	wire [16-1:0] node5580;
	wire [16-1:0] node5583;
	wire [16-1:0] node5584;
	wire [16-1:0] node5588;
	wire [16-1:0] node5589;
	wire [16-1:0] node5591;
	wire [16-1:0] node5594;
	wire [16-1:0] node5595;
	wire [16-1:0] node5598;
	wire [16-1:0] node5601;
	wire [16-1:0] node5602;
	wire [16-1:0] node5603;
	wire [16-1:0] node5607;
	wire [16-1:0] node5608;
	wire [16-1:0] node5610;
	wire [16-1:0] node5612;
	wire [16-1:0] node5613;
	wire [16-1:0] node5617;
	wire [16-1:0] node5619;
	wire [16-1:0] node5620;
	wire [16-1:0] node5624;
	wire [16-1:0] node5625;
	wire [16-1:0] node5626;
	wire [16-1:0] node5627;
	wire [16-1:0] node5629;
	wire [16-1:0] node5630;
	wire [16-1:0] node5632;
	wire [16-1:0] node5635;
	wire [16-1:0] node5638;
	wire [16-1:0] node5639;
	wire [16-1:0] node5641;
	wire [16-1:0] node5643;
	wire [16-1:0] node5646;
	wire [16-1:0] node5647;
	wire [16-1:0] node5650;
	wire [16-1:0] node5652;
	wire [16-1:0] node5655;
	wire [16-1:0] node5656;
	wire [16-1:0] node5657;
	wire [16-1:0] node5658;
	wire [16-1:0] node5661;
	wire [16-1:0] node5664;
	wire [16-1:0] node5665;
	wire [16-1:0] node5667;
	wire [16-1:0] node5668;
	wire [16-1:0] node5673;
	wire [16-1:0] node5674;
	wire [16-1:0] node5677;
	wire [16-1:0] node5678;
	wire [16-1:0] node5682;
	wire [16-1:0] node5683;
	wire [16-1:0] node5684;
	wire [16-1:0] node5685;
	wire [16-1:0] node5687;
	wire [16-1:0] node5690;
	wire [16-1:0] node5691;
	wire [16-1:0] node5694;
	wire [16-1:0] node5697;
	wire [16-1:0] node5698;
	wire [16-1:0] node5700;
	wire [16-1:0] node5703;
	wire [16-1:0] node5704;
	wire [16-1:0] node5708;
	wire [16-1:0] node5709;
	wire [16-1:0] node5710;
	wire [16-1:0] node5711;
	wire [16-1:0] node5714;
	wire [16-1:0] node5716;
	wire [16-1:0] node5719;
	wire [16-1:0] node5720;
	wire [16-1:0] node5723;
	wire [16-1:0] node5724;
	wire [16-1:0] node5727;
	wire [16-1:0] node5728;
	wire [16-1:0] node5732;
	wire [16-1:0] node5733;
	wire [16-1:0] node5735;
	wire [16-1:0] node5738;
	wire [16-1:0] node5740;
	wire [16-1:0] node5743;
	wire [16-1:0] node5744;
	wire [16-1:0] node5745;
	wire [16-1:0] node5746;
	wire [16-1:0] node5747;
	wire [16-1:0] node5748;
	wire [16-1:0] node5749;
	wire [16-1:0] node5750;
	wire [16-1:0] node5753;
	wire [16-1:0] node5754;
	wire [16-1:0] node5756;
	wire [16-1:0] node5761;
	wire [16-1:0] node5762;
	wire [16-1:0] node5765;
	wire [16-1:0] node5766;
	wire [16-1:0] node5770;
	wire [16-1:0] node5771;
	wire [16-1:0] node5772;
	wire [16-1:0] node5773;
	wire [16-1:0] node5775;
	wire [16-1:0] node5776;
	wire [16-1:0] node5780;
	wire [16-1:0] node5781;
	wire [16-1:0] node5782;
	wire [16-1:0] node5786;
	wire [16-1:0] node5789;
	wire [16-1:0] node5790;
	wire [16-1:0] node5794;
	wire [16-1:0] node5795;
	wire [16-1:0] node5796;
	wire [16-1:0] node5799;
	wire [16-1:0] node5800;
	wire [16-1:0] node5802;
	wire [16-1:0] node5806;
	wire [16-1:0] node5807;
	wire [16-1:0] node5810;
	wire [16-1:0] node5812;
	wire [16-1:0] node5815;
	wire [16-1:0] node5816;
	wire [16-1:0] node5817;
	wire [16-1:0] node5818;
	wire [16-1:0] node5820;
	wire [16-1:0] node5823;
	wire [16-1:0] node5825;
	wire [16-1:0] node5826;
	wire [16-1:0] node5830;
	wire [16-1:0] node5831;
	wire [16-1:0] node5834;
	wire [16-1:0] node5835;
	wire [16-1:0] node5839;
	wire [16-1:0] node5840;
	wire [16-1:0] node5841;
	wire [16-1:0] node5843;
	wire [16-1:0] node5844;
	wire [16-1:0] node5848;
	wire [16-1:0] node5850;
	wire [16-1:0] node5853;
	wire [16-1:0] node5855;
	wire [16-1:0] node5856;
	wire [16-1:0] node5857;
	wire [16-1:0] node5861;
	wire [16-1:0] node5864;
	wire [16-1:0] node5865;
	wire [16-1:0] node5866;
	wire [16-1:0] node5867;
	wire [16-1:0] node5868;
	wire [16-1:0] node5869;
	wire [16-1:0] node5872;
	wire [16-1:0] node5875;
	wire [16-1:0] node5877;
	wire [16-1:0] node5879;
	wire [16-1:0] node5882;
	wire [16-1:0] node5883;
	wire [16-1:0] node5885;
	wire [16-1:0] node5888;
	wire [16-1:0] node5889;
	wire [16-1:0] node5893;
	wire [16-1:0] node5894;
	wire [16-1:0] node5895;
	wire [16-1:0] node5896;
	wire [16-1:0] node5899;
	wire [16-1:0] node5902;
	wire [16-1:0] node5903;
	wire [16-1:0] node5904;
	wire [16-1:0] node5906;
	wire [16-1:0] node5909;
	wire [16-1:0] node5910;
	wire [16-1:0] node5913;
	wire [16-1:0] node5917;
	wire [16-1:0] node5918;
	wire [16-1:0] node5919;
	wire [16-1:0] node5923;
	wire [16-1:0] node5924;
	wire [16-1:0] node5925;
	wire [16-1:0] node5928;
	wire [16-1:0] node5929;
	wire [16-1:0] node5933;
	wire [16-1:0] node5935;
	wire [16-1:0] node5938;
	wire [16-1:0] node5939;
	wire [16-1:0] node5940;
	wire [16-1:0] node5941;
	wire [16-1:0] node5942;
	wire [16-1:0] node5943;
	wire [16-1:0] node5947;
	wire [16-1:0] node5949;
	wire [16-1:0] node5952;
	wire [16-1:0] node5953;
	wire [16-1:0] node5956;
	wire [16-1:0] node5959;
	wire [16-1:0] node5960;
	wire [16-1:0] node5961;
	wire [16-1:0] node5964;
	wire [16-1:0] node5966;
	wire [16-1:0] node5967;
	wire [16-1:0] node5971;
	wire [16-1:0] node5972;
	wire [16-1:0] node5974;
	wire [16-1:0] node5978;
	wire [16-1:0] node5979;
	wire [16-1:0] node5980;
	wire [16-1:0] node5981;
	wire [16-1:0] node5983;
	wire [16-1:0] node5985;
	wire [16-1:0] node5988;
	wire [16-1:0] node5989;
	wire [16-1:0] node5991;
	wire [16-1:0] node5995;
	wire [16-1:0] node5996;
	wire [16-1:0] node5997;
	wire [16-1:0] node6002;
	wire [16-1:0] node6003;
	wire [16-1:0] node6004;
	wire [16-1:0] node6006;
	wire [16-1:0] node6009;
	wire [16-1:0] node6011;
	wire [16-1:0] node6014;
	wire [16-1:0] node6015;
	wire [16-1:0] node6017;
	wire [16-1:0] node6020;
	wire [16-1:0] node6022;
	wire [16-1:0] node6025;
	wire [16-1:0] node6026;
	wire [16-1:0] node6027;
	wire [16-1:0] node6028;
	wire [16-1:0] node6029;
	wire [16-1:0] node6031;
	wire [16-1:0] node6034;
	wire [16-1:0] node6036;
	wire [16-1:0] node6037;
	wire [16-1:0] node6039;
	wire [16-1:0] node6043;
	wire [16-1:0] node6044;
	wire [16-1:0] node6045;
	wire [16-1:0] node6046;
	wire [16-1:0] node6050;
	wire [16-1:0] node6052;
	wire [16-1:0] node6055;
	wire [16-1:0] node6056;
	wire [16-1:0] node6057;
	wire [16-1:0] node6059;
	wire [16-1:0] node6063;
	wire [16-1:0] node6064;
	wire [16-1:0] node6065;
	wire [16-1:0] node6066;
	wire [16-1:0] node6069;
	wire [16-1:0] node6074;
	wire [16-1:0] node6075;
	wire [16-1:0] node6076;
	wire [16-1:0] node6077;
	wire [16-1:0] node6079;
	wire [16-1:0] node6082;
	wire [16-1:0] node6083;
	wire [16-1:0] node6084;
	wire [16-1:0] node6088;
	wire [16-1:0] node6091;
	wire [16-1:0] node6094;
	wire [16-1:0] node6095;
	wire [16-1:0] node6096;
	wire [16-1:0] node6097;
	wire [16-1:0] node6099;
	wire [16-1:0] node6102;
	wire [16-1:0] node6105;
	wire [16-1:0] node6106;
	wire [16-1:0] node6107;
	wire [16-1:0] node6111;
	wire [16-1:0] node6112;
	wire [16-1:0] node6116;
	wire [16-1:0] node6117;
	wire [16-1:0] node6119;
	wire [16-1:0] node6122;
	wire [16-1:0] node6123;
	wire [16-1:0] node6126;
	wire [16-1:0] node6129;
	wire [16-1:0] node6130;
	wire [16-1:0] node6131;
	wire [16-1:0] node6132;
	wire [16-1:0] node6133;
	wire [16-1:0] node6134;
	wire [16-1:0] node6137;
	wire [16-1:0] node6138;
	wire [16-1:0] node6140;
	wire [16-1:0] node6144;
	wire [16-1:0] node6145;
	wire [16-1:0] node6146;
	wire [16-1:0] node6148;
	wire [16-1:0] node6152;
	wire [16-1:0] node6155;
	wire [16-1:0] node6156;
	wire [16-1:0] node6157;
	wire [16-1:0] node6158;
	wire [16-1:0] node6160;
	wire [16-1:0] node6164;
	wire [16-1:0] node6165;
	wire [16-1:0] node6169;
	wire [16-1:0] node6170;
	wire [16-1:0] node6172;
	wire [16-1:0] node6175;
	wire [16-1:0] node6177;
	wire [16-1:0] node6178;
	wire [16-1:0] node6181;
	wire [16-1:0] node6184;
	wire [16-1:0] node6185;
	wire [16-1:0] node6186;
	wire [16-1:0] node6188;
	wire [16-1:0] node6191;
	wire [16-1:0] node6192;
	wire [16-1:0] node6196;
	wire [16-1:0] node6197;
	wire [16-1:0] node6198;
	wire [16-1:0] node6200;
	wire [16-1:0] node6203;
	wire [16-1:0] node6206;
	wire [16-1:0] node6208;
	wire [16-1:0] node6211;
	wire [16-1:0] node6212;
	wire [16-1:0] node6213;
	wire [16-1:0] node6214;
	wire [16-1:0] node6215;
	wire [16-1:0] node6218;
	wire [16-1:0] node6219;
	wire [16-1:0] node6220;
	wire [16-1:0] node6225;
	wire [16-1:0] node6226;
	wire [16-1:0] node6229;
	wire [16-1:0] node6231;
	wire [16-1:0] node6234;
	wire [16-1:0] node6235;
	wire [16-1:0] node6237;
	wire [16-1:0] node6239;
	wire [16-1:0] node6240;
	wire [16-1:0] node6244;
	wire [16-1:0] node6245;
	wire [16-1:0] node6248;
	wire [16-1:0] node6250;
	wire [16-1:0] node6253;
	wire [16-1:0] node6254;
	wire [16-1:0] node6255;
	wire [16-1:0] node6257;
	wire [16-1:0] node6258;
	wire [16-1:0] node6260;
	wire [16-1:0] node6265;
	wire [16-1:0] node6266;
	wire [16-1:0] node6268;
	wire [16-1:0] node6269;
	wire [16-1:0] node6273;
	wire [16-1:0] node6274;
	wire [16-1:0] node6275;
	wire [16-1:0] node6277;
	wire [16-1:0] node6282;
	wire [16-1:0] node6283;
	wire [16-1:0] node6284;
	wire [16-1:0] node6285;
	wire [16-1:0] node6286;
	wire [16-1:0] node6287;
	wire [16-1:0] node6288;
	wire [16-1:0] node6289;
	wire [16-1:0] node6290;
	wire [16-1:0] node6291;
	wire [16-1:0] node6292;
	wire [16-1:0] node6297;
	wire [16-1:0] node6298;
	wire [16-1:0] node6301;
	wire [16-1:0] node6304;
	wire [16-1:0] node6305;
	wire [16-1:0] node6306;
	wire [16-1:0] node6310;
	wire [16-1:0] node6311;
	wire [16-1:0] node6313;
	wire [16-1:0] node6315;
	wire [16-1:0] node6319;
	wire [16-1:0] node6320;
	wire [16-1:0] node6323;
	wire [16-1:0] node6324;
	wire [16-1:0] node6325;
	wire [16-1:0] node6329;
	wire [16-1:0] node6330;
	wire [16-1:0] node6333;
	wire [16-1:0] node6336;
	wire [16-1:0] node6337;
	wire [16-1:0] node6338;
	wire [16-1:0] node6339;
	wire [16-1:0] node6340;
	wire [16-1:0] node6341;
	wire [16-1:0] node6346;
	wire [16-1:0] node6347;
	wire [16-1:0] node6349;
	wire [16-1:0] node6352;
	wire [16-1:0] node6354;
	wire [16-1:0] node6355;
	wire [16-1:0] node6359;
	wire [16-1:0] node6360;
	wire [16-1:0] node6364;
	wire [16-1:0] node6365;
	wire [16-1:0] node6366;
	wire [16-1:0] node6368;
	wire [16-1:0] node6371;
	wire [16-1:0] node6372;
	wire [16-1:0] node6376;
	wire [16-1:0] node6377;
	wire [16-1:0] node6378;
	wire [16-1:0] node6379;
	wire [16-1:0] node6381;
	wire [16-1:0] node6384;
	wire [16-1:0] node6385;
	wire [16-1:0] node6389;
	wire [16-1:0] node6392;
	wire [16-1:0] node6395;
	wire [16-1:0] node6396;
	wire [16-1:0] node6397;
	wire [16-1:0] node6398;
	wire [16-1:0] node6399;
	wire [16-1:0] node6400;
	wire [16-1:0] node6401;
	wire [16-1:0] node6404;
	wire [16-1:0] node6408;
	wire [16-1:0] node6409;
	wire [16-1:0] node6411;
	wire [16-1:0] node6415;
	wire [16-1:0] node6416;
	wire [16-1:0] node6417;
	wire [16-1:0] node6418;
	wire [16-1:0] node6422;
	wire [16-1:0] node6425;
	wire [16-1:0] node6426;
	wire [16-1:0] node6429;
	wire [16-1:0] node6432;
	wire [16-1:0] node6433;
	wire [16-1:0] node6434;
	wire [16-1:0] node6435;
	wire [16-1:0] node6436;
	wire [16-1:0] node6441;
	wire [16-1:0] node6442;
	wire [16-1:0] node6443;
	wire [16-1:0] node6447;
	wire [16-1:0] node6450;
	wire [16-1:0] node6452;
	wire [16-1:0] node6453;
	wire [16-1:0] node6456;
	wire [16-1:0] node6459;
	wire [16-1:0] node6460;
	wire [16-1:0] node6461;
	wire [16-1:0] node6462;
	wire [16-1:0] node6463;
	wire [16-1:0] node6466;
	wire [16-1:0] node6470;
	wire [16-1:0] node6471;
	wire [16-1:0] node6474;
	wire [16-1:0] node6475;
	wire [16-1:0] node6477;
	wire [16-1:0] node6481;
	wire [16-1:0] node6482;
	wire [16-1:0] node6483;
	wire [16-1:0] node6485;
	wire [16-1:0] node6488;
	wire [16-1:0] node6489;
	wire [16-1:0] node6492;
	wire [16-1:0] node6495;
	wire [16-1:0] node6496;
	wire [16-1:0] node6497;
	wire [16-1:0] node6501;
	wire [16-1:0] node6503;
	wire [16-1:0] node6505;
	wire [16-1:0] node6508;
	wire [16-1:0] node6509;
	wire [16-1:0] node6510;
	wire [16-1:0] node6511;
	wire [16-1:0] node6512;
	wire [16-1:0] node6513;
	wire [16-1:0] node6514;
	wire [16-1:0] node6517;
	wire [16-1:0] node6519;
	wire [16-1:0] node6520;
	wire [16-1:0] node6524;
	wire [16-1:0] node6525;
	wire [16-1:0] node6526;
	wire [16-1:0] node6530;
	wire [16-1:0] node6533;
	wire [16-1:0] node6534;
	wire [16-1:0] node6535;
	wire [16-1:0] node6537;
	wire [16-1:0] node6540;
	wire [16-1:0] node6543;
	wire [16-1:0] node6545;
	wire [16-1:0] node6548;
	wire [16-1:0] node6549;
	wire [16-1:0] node6551;
	wire [16-1:0] node6552;
	wire [16-1:0] node6554;
	wire [16-1:0] node6555;
	wire [16-1:0] node6559;
	wire [16-1:0] node6562;
	wire [16-1:0] node6563;
	wire [16-1:0] node6564;
	wire [16-1:0] node6567;
	wire [16-1:0] node6569;
	wire [16-1:0] node6572;
	wire [16-1:0] node6573;
	wire [16-1:0] node6574;
	wire [16-1:0] node6577;
	wire [16-1:0] node6578;
	wire [16-1:0] node6582;
	wire [16-1:0] node6585;
	wire [16-1:0] node6586;
	wire [16-1:0] node6587;
	wire [16-1:0] node6588;
	wire [16-1:0] node6590;
	wire [16-1:0] node6591;
	wire [16-1:0] node6592;
	wire [16-1:0] node6595;
	wire [16-1:0] node6599;
	wire [16-1:0] node6601;
	wire [16-1:0] node6602;
	wire [16-1:0] node6606;
	wire [16-1:0] node6608;
	wire [16-1:0] node6609;
	wire [16-1:0] node6610;
	wire [16-1:0] node6614;
	wire [16-1:0] node6617;
	wire [16-1:0] node6618;
	wire [16-1:0] node6619;
	wire [16-1:0] node6620;
	wire [16-1:0] node6625;
	wire [16-1:0] node6626;
	wire [16-1:0] node6627;
	wire [16-1:0] node6632;
	wire [16-1:0] node6633;
	wire [16-1:0] node6634;
	wire [16-1:0] node6635;
	wire [16-1:0] node6636;
	wire [16-1:0] node6637;
	wire [16-1:0] node6641;
	wire [16-1:0] node6642;
	wire [16-1:0] node6646;
	wire [16-1:0] node6647;
	wire [16-1:0] node6648;
	wire [16-1:0] node6649;
	wire [16-1:0] node6651;
	wire [16-1:0] node6655;
	wire [16-1:0] node6656;
	wire [16-1:0] node6657;
	wire [16-1:0] node6660;
	wire [16-1:0] node6663;
	wire [16-1:0] node6664;
	wire [16-1:0] node6668;
	wire [16-1:0] node6669;
	wire [16-1:0] node6673;
	wire [16-1:0] node6674;
	wire [16-1:0] node6675;
	wire [16-1:0] node6678;
	wire [16-1:0] node6679;
	wire [16-1:0] node6681;
	wire [16-1:0] node6684;
	wire [16-1:0] node6687;
	wire [16-1:0] node6688;
	wire [16-1:0] node6689;
	wire [16-1:0] node6692;
	wire [16-1:0] node6693;
	wire [16-1:0] node6697;
	wire [16-1:0] node6698;
	wire [16-1:0] node6701;
	wire [16-1:0] node6704;
	wire [16-1:0] node6705;
	wire [16-1:0] node6706;
	wire [16-1:0] node6707;
	wire [16-1:0] node6709;
	wire [16-1:0] node6712;
	wire [16-1:0] node6713;
	wire [16-1:0] node6717;
	wire [16-1:0] node6720;
	wire [16-1:0] node6721;
	wire [16-1:0] node6722;
	wire [16-1:0] node6724;
	wire [16-1:0] node6726;
	wire [16-1:0] node6729;
	wire [16-1:0] node6730;
	wire [16-1:0] node6733;
	wire [16-1:0] node6735;
	wire [16-1:0] node6738;
	wire [16-1:0] node6739;
	wire [16-1:0] node6740;
	wire [16-1:0] node6741;
	wire [16-1:0] node6745;
	wire [16-1:0] node6749;
	wire [16-1:0] node6750;
	wire [16-1:0] node6751;
	wire [16-1:0] node6752;
	wire [16-1:0] node6753;
	wire [16-1:0] node6754;
	wire [16-1:0] node6755;
	wire [16-1:0] node6756;
	wire [16-1:0] node6758;
	wire [16-1:0] node6761;
	wire [16-1:0] node6762;
	wire [16-1:0] node6763;
	wire [16-1:0] node6768;
	wire [16-1:0] node6769;
	wire [16-1:0] node6770;
	wire [16-1:0] node6774;
	wire [16-1:0] node6777;
	wire [16-1:0] node6778;
	wire [16-1:0] node6780;
	wire [16-1:0] node6783;
	wire [16-1:0] node6784;
	wire [16-1:0] node6787;
	wire [16-1:0] node6790;
	wire [16-1:0] node6791;
	wire [16-1:0] node6792;
	wire [16-1:0] node6793;
	wire [16-1:0] node6796;
	wire [16-1:0] node6798;
	wire [16-1:0] node6799;
	wire [16-1:0] node6803;
	wire [16-1:0] node6804;
	wire [16-1:0] node6807;
	wire [16-1:0] node6810;
	wire [16-1:0] node6811;
	wire [16-1:0] node6812;
	wire [16-1:0] node6813;
	wire [16-1:0] node6818;
	wire [16-1:0] node6819;
	wire [16-1:0] node6822;
	wire [16-1:0] node6825;
	wire [16-1:0] node6826;
	wire [16-1:0] node6827;
	wire [16-1:0] node6828;
	wire [16-1:0] node6830;
	wire [16-1:0] node6831;
	wire [16-1:0] node6832;
	wire [16-1:0] node6837;
	wire [16-1:0] node6838;
	wire [16-1:0] node6841;
	wire [16-1:0] node6844;
	wire [16-1:0] node6846;
	wire [16-1:0] node6847;
	wire [16-1:0] node6848;
	wire [16-1:0] node6853;
	wire [16-1:0] node6854;
	wire [16-1:0] node6855;
	wire [16-1:0] node6858;
	wire [16-1:0] node6859;
	wire [16-1:0] node6861;
	wire [16-1:0] node6862;
	wire [16-1:0] node6866;
	wire [16-1:0] node6868;
	wire [16-1:0] node6871;
	wire [16-1:0] node6872;
	wire [16-1:0] node6874;
	wire [16-1:0] node6878;
	wire [16-1:0] node6879;
	wire [16-1:0] node6880;
	wire [16-1:0] node6881;
	wire [16-1:0] node6882;
	wire [16-1:0] node6883;
	wire [16-1:0] node6887;
	wire [16-1:0] node6888;
	wire [16-1:0] node6891;
	wire [16-1:0] node6894;
	wire [16-1:0] node6895;
	wire [16-1:0] node6896;
	wire [16-1:0] node6899;
	wire [16-1:0] node6900;
	wire [16-1:0] node6902;
	wire [16-1:0] node6905;
	wire [16-1:0] node6906;
	wire [16-1:0] node6910;
	wire [16-1:0] node6911;
	wire [16-1:0] node6914;
	wire [16-1:0] node6917;
	wire [16-1:0] node6918;
	wire [16-1:0] node6919;
	wire [16-1:0] node6920;
	wire [16-1:0] node6922;
	wire [16-1:0] node6923;
	wire [16-1:0] node6927;
	wire [16-1:0] node6930;
	wire [16-1:0] node6931;
	wire [16-1:0] node6934;
	wire [16-1:0] node6936;
	wire [16-1:0] node6937;
	wire [16-1:0] node6941;
	wire [16-1:0] node6942;
	wire [16-1:0] node6943;
	wire [16-1:0] node6948;
	wire [16-1:0] node6949;
	wire [16-1:0] node6950;
	wire [16-1:0] node6951;
	wire [16-1:0] node6952;
	wire [16-1:0] node6955;
	wire [16-1:0] node6957;
	wire [16-1:0] node6960;
	wire [16-1:0] node6961;
	wire [16-1:0] node6963;
	wire [16-1:0] node6964;
	wire [16-1:0] node6968;
	wire [16-1:0] node6970;
	wire [16-1:0] node6973;
	wire [16-1:0] node6974;
	wire [16-1:0] node6976;
	wire [16-1:0] node6977;
	wire [16-1:0] node6982;
	wire [16-1:0] node6983;
	wire [16-1:0] node6984;
	wire [16-1:0] node6985;
	wire [16-1:0] node6986;
	wire [16-1:0] node6991;
	wire [16-1:0] node6992;
	wire [16-1:0] node6994;
	wire [16-1:0] node6998;
	wire [16-1:0] node6999;
	wire [16-1:0] node7000;
	wire [16-1:0] node7002;
	wire [16-1:0] node7003;
	wire [16-1:0] node7007;
	wire [16-1:0] node7009;
	wire [16-1:0] node7010;
	wire [16-1:0] node7014;
	wire [16-1:0] node7016;
	wire [16-1:0] node7019;
	wire [16-1:0] node7020;
	wire [16-1:0] node7021;
	wire [16-1:0] node7022;
	wire [16-1:0] node7023;
	wire [16-1:0] node7024;
	wire [16-1:0] node7025;
	wire [16-1:0] node7027;
	wire [16-1:0] node7028;
	wire [16-1:0] node7032;
	wire [16-1:0] node7034;
	wire [16-1:0] node7037;
	wire [16-1:0] node7039;
	wire [16-1:0] node7042;
	wire [16-1:0] node7043;
	wire [16-1:0] node7046;
	wire [16-1:0] node7047;
	wire [16-1:0] node7048;
	wire [16-1:0] node7051;
	wire [16-1:0] node7052;
	wire [16-1:0] node7056;
	wire [16-1:0] node7059;
	wire [16-1:0] node7060;
	wire [16-1:0] node7061;
	wire [16-1:0] node7063;
	wire [16-1:0] node7064;
	wire [16-1:0] node7068;
	wire [16-1:0] node7069;
	wire [16-1:0] node7071;
	wire [16-1:0] node7072;
	wire [16-1:0] node7076;
	wire [16-1:0] node7079;
	wire [16-1:0] node7081;
	wire [16-1:0] node7082;
	wire [16-1:0] node7083;
	wire [16-1:0] node7086;
	wire [16-1:0] node7090;
	wire [16-1:0] node7091;
	wire [16-1:0] node7092;
	wire [16-1:0] node7094;
	wire [16-1:0] node7096;
	wire [16-1:0] node7099;
	wire [16-1:0] node7100;
	wire [16-1:0] node7101;
	wire [16-1:0] node7103;
	wire [16-1:0] node7104;
	wire [16-1:0] node7109;
	wire [16-1:0] node7110;
	wire [16-1:0] node7113;
	wire [16-1:0] node7114;
	wire [16-1:0] node7118;
	wire [16-1:0] node7119;
	wire [16-1:0] node7120;
	wire [16-1:0] node7121;
	wire [16-1:0] node7122;
	wire [16-1:0] node7124;
	wire [16-1:0] node7128;
	wire [16-1:0] node7131;
	wire [16-1:0] node7133;
	wire [16-1:0] node7134;
	wire [16-1:0] node7135;
	wire [16-1:0] node7139;
	wire [16-1:0] node7140;
	wire [16-1:0] node7144;
	wire [16-1:0] node7145;
	wire [16-1:0] node7147;
	wire [16-1:0] node7149;
	wire [16-1:0] node7150;
	wire [16-1:0] node7154;
	wire [16-1:0] node7156;
	wire [16-1:0] node7158;
	wire [16-1:0] node7161;
	wire [16-1:0] node7162;
	wire [16-1:0] node7163;
	wire [16-1:0] node7164;
	wire [16-1:0] node7165;
	wire [16-1:0] node7166;
	wire [16-1:0] node7168;
	wire [16-1:0] node7170;
	wire [16-1:0] node7173;
	wire [16-1:0] node7174;
	wire [16-1:0] node7176;
	wire [16-1:0] node7180;
	wire [16-1:0] node7181;
	wire [16-1:0] node7184;
	wire [16-1:0] node7187;
	wire [16-1:0] node7188;
	wire [16-1:0] node7189;
	wire [16-1:0] node7194;
	wire [16-1:0] node7195;
	wire [16-1:0] node7196;
	wire [16-1:0] node7197;
	wire [16-1:0] node7199;
	wire [16-1:0] node7202;
	wire [16-1:0] node7204;
	wire [16-1:0] node7207;
	wire [16-1:0] node7210;
	wire [16-1:0] node7211;
	wire [16-1:0] node7213;
	wire [16-1:0] node7214;
	wire [16-1:0] node7218;
	wire [16-1:0] node7220;
	wire [16-1:0] node7222;
	wire [16-1:0] node7223;
	wire [16-1:0] node7227;
	wire [16-1:0] node7228;
	wire [16-1:0] node7229;
	wire [16-1:0] node7230;
	wire [16-1:0] node7232;
	wire [16-1:0] node7235;
	wire [16-1:0] node7238;
	wire [16-1:0] node7239;
	wire [16-1:0] node7241;
	wire [16-1:0] node7244;
	wire [16-1:0] node7246;
	wire [16-1:0] node7249;
	wire [16-1:0] node7250;
	wire [16-1:0] node7251;
	wire [16-1:0] node7252;
	wire [16-1:0] node7254;
	wire [16-1:0] node7256;
	wire [16-1:0] node7260;
	wire [16-1:0] node7263;
	wire [16-1:0] node7264;
	wire [16-1:0] node7267;
	wire [16-1:0] node7268;
	wire [16-1:0] node7270;
	wire [16-1:0] node7272;
	wire [16-1:0] node7275;
	wire [16-1:0] node7276;
	wire [16-1:0] node7278;
	wire [16-1:0] node7282;
	wire [16-1:0] node7283;
	wire [16-1:0] node7284;
	wire [16-1:0] node7285;
	wire [16-1:0] node7286;
	wire [16-1:0] node7287;
	wire [16-1:0] node7288;
	wire [16-1:0] node7289;
	wire [16-1:0] node7290;
	wire [16-1:0] node7291;
	wire [16-1:0] node7293;
	wire [16-1:0] node7298;
	wire [16-1:0] node7301;
	wire [16-1:0] node7302;
	wire [16-1:0] node7305;
	wire [16-1:0] node7306;
	wire [16-1:0] node7309;
	wire [16-1:0] node7312;
	wire [16-1:0] node7313;
	wire [16-1:0] node7314;
	wire [16-1:0] node7315;
	wire [16-1:0] node7318;
	wire [16-1:0] node7320;
	wire [16-1:0] node7323;
	wire [16-1:0] node7324;
	wire [16-1:0] node7327;
	wire [16-1:0] node7330;
	wire [16-1:0] node7331;
	wire [16-1:0] node7333;
	wire [16-1:0] node7337;
	wire [16-1:0] node7338;
	wire [16-1:0] node7339;
	wire [16-1:0] node7340;
	wire [16-1:0] node7341;
	wire [16-1:0] node7344;
	wire [16-1:0] node7345;
	wire [16-1:0] node7347;
	wire [16-1:0] node7351;
	wire [16-1:0] node7353;
	wire [16-1:0] node7356;
	wire [16-1:0] node7357;
	wire [16-1:0] node7358;
	wire [16-1:0] node7360;
	wire [16-1:0] node7362;
	wire [16-1:0] node7365;
	wire [16-1:0] node7366;
	wire [16-1:0] node7371;
	wire [16-1:0] node7372;
	wire [16-1:0] node7373;
	wire [16-1:0] node7374;
	wire [16-1:0] node7377;
	wire [16-1:0] node7380;
	wire [16-1:0] node7381;
	wire [16-1:0] node7384;
	wire [16-1:0] node7387;
	wire [16-1:0] node7388;
	wire [16-1:0] node7390;
	wire [16-1:0] node7393;
	wire [16-1:0] node7396;
	wire [16-1:0] node7397;
	wire [16-1:0] node7398;
	wire [16-1:0] node7399;
	wire [16-1:0] node7400;
	wire [16-1:0] node7402;
	wire [16-1:0] node7405;
	wire [16-1:0] node7406;
	wire [16-1:0] node7408;
	wire [16-1:0] node7412;
	wire [16-1:0] node7413;
	wire [16-1:0] node7414;
	wire [16-1:0] node7416;
	wire [16-1:0] node7417;
	wire [16-1:0] node7421;
	wire [16-1:0] node7424;
	wire [16-1:0] node7425;
	wire [16-1:0] node7427;
	wire [16-1:0] node7430;
	wire [16-1:0] node7433;
	wire [16-1:0] node7434;
	wire [16-1:0] node7435;
	wire [16-1:0] node7436;
	wire [16-1:0] node7439;
	wire [16-1:0] node7442;
	wire [16-1:0] node7443;
	wire [16-1:0] node7445;
	wire [16-1:0] node7446;
	wire [16-1:0] node7449;
	wire [16-1:0] node7453;
	wire [16-1:0] node7454;
	wire [16-1:0] node7455;
	wire [16-1:0] node7458;
	wire [16-1:0] node7461;
	wire [16-1:0] node7463;
	wire [16-1:0] node7466;
	wire [16-1:0] node7467;
	wire [16-1:0] node7468;
	wire [16-1:0] node7469;
	wire [16-1:0] node7470;
	wire [16-1:0] node7473;
	wire [16-1:0] node7476;
	wire [16-1:0] node7478;
	wire [16-1:0] node7480;
	wire [16-1:0] node7483;
	wire [16-1:0] node7484;
	wire [16-1:0] node7485;
	wire [16-1:0] node7486;
	wire [16-1:0] node7490;
	wire [16-1:0] node7493;
	wire [16-1:0] node7494;
	wire [16-1:0] node7498;
	wire [16-1:0] node7499;
	wire [16-1:0] node7500;
	wire [16-1:0] node7503;
	wire [16-1:0] node7504;
	wire [16-1:0] node7508;
	wire [16-1:0] node7509;
	wire [16-1:0] node7510;
	wire [16-1:0] node7514;
	wire [16-1:0] node7515;
	wire [16-1:0] node7517;
	wire [16-1:0] node7518;
	wire [16-1:0] node7523;
	wire [16-1:0] node7524;
	wire [16-1:0] node7525;
	wire [16-1:0] node7526;
	wire [16-1:0] node7527;
	wire [16-1:0] node7528;
	wire [16-1:0] node7530;
	wire [16-1:0] node7533;
	wire [16-1:0] node7534;
	wire [16-1:0] node7538;
	wire [16-1:0] node7539;
	wire [16-1:0] node7540;
	wire [16-1:0] node7541;
	wire [16-1:0] node7542;
	wire [16-1:0] node7547;
	wire [16-1:0] node7550;
	wire [16-1:0] node7551;
	wire [16-1:0] node7552;
	wire [16-1:0] node7554;
	wire [16-1:0] node7559;
	wire [16-1:0] node7560;
	wire [16-1:0] node7561;
	wire [16-1:0] node7562;
	wire [16-1:0] node7563;
	wire [16-1:0] node7567;
	wire [16-1:0] node7570;
	wire [16-1:0] node7571;
	wire [16-1:0] node7573;
	wire [16-1:0] node7574;
	wire [16-1:0] node7578;
	wire [16-1:0] node7579;
	wire [16-1:0] node7583;
	wire [16-1:0] node7585;
	wire [16-1:0] node7586;
	wire [16-1:0] node7588;
	wire [16-1:0] node7591;
	wire [16-1:0] node7594;
	wire [16-1:0] node7595;
	wire [16-1:0] node7596;
	wire [16-1:0] node7597;
	wire [16-1:0] node7598;
	wire [16-1:0] node7600;
	wire [16-1:0] node7601;
	wire [16-1:0] node7607;
	wire [16-1:0] node7608;
	wire [16-1:0] node7609;
	wire [16-1:0] node7611;
	wire [16-1:0] node7614;
	wire [16-1:0] node7617;
	wire [16-1:0] node7618;
	wire [16-1:0] node7621;
	wire [16-1:0] node7622;
	wire [16-1:0] node7626;
	wire [16-1:0] node7627;
	wire [16-1:0] node7628;
	wire [16-1:0] node7629;
	wire [16-1:0] node7632;
	wire [16-1:0] node7633;
	wire [16-1:0] node7635;
	wire [16-1:0] node7638;
	wire [16-1:0] node7640;
	wire [16-1:0] node7644;
	wire [16-1:0] node7645;
	wire [16-1:0] node7646;
	wire [16-1:0] node7649;
	wire [16-1:0] node7651;
	wire [16-1:0] node7654;
	wire [16-1:0] node7655;
	wire [16-1:0] node7659;
	wire [16-1:0] node7660;
	wire [16-1:0] node7661;
	wire [16-1:0] node7662;
	wire [16-1:0] node7663;
	wire [16-1:0] node7664;
	wire [16-1:0] node7666;
	wire [16-1:0] node7670;
	wire [16-1:0] node7671;
	wire [16-1:0] node7674;
	wire [16-1:0] node7676;
	wire [16-1:0] node7679;
	wire [16-1:0] node7680;
	wire [16-1:0] node7681;
	wire [16-1:0] node7684;
	wire [16-1:0] node7686;
	wire [16-1:0] node7689;
	wire [16-1:0] node7690;
	wire [16-1:0] node7692;
	wire [16-1:0] node7693;
	wire [16-1:0] node7697;
	wire [16-1:0] node7700;
	wire [16-1:0] node7701;
	wire [16-1:0] node7703;
	wire [16-1:0] node7704;
	wire [16-1:0] node7707;
	wire [16-1:0] node7710;
	wire [16-1:0] node7711;
	wire [16-1:0] node7713;
	wire [16-1:0] node7715;
	wire [16-1:0] node7718;
	wire [16-1:0] node7720;
	wire [16-1:0] node7723;
	wire [16-1:0] node7724;
	wire [16-1:0] node7725;
	wire [16-1:0] node7726;
	wire [16-1:0] node7727;
	wire [16-1:0] node7728;
	wire [16-1:0] node7732;
	wire [16-1:0] node7733;
	wire [16-1:0] node7735;
	wire [16-1:0] node7738;
	wire [16-1:0] node7740;
	wire [16-1:0] node7743;
	wire [16-1:0] node7745;
	wire [16-1:0] node7748;
	wire [16-1:0] node7749;
	wire [16-1:0] node7752;
	wire [16-1:0] node7755;
	wire [16-1:0] node7756;
	wire [16-1:0] node7757;
	wire [16-1:0] node7759;
	wire [16-1:0] node7761;
	wire [16-1:0] node7762;
	wire [16-1:0] node7766;
	wire [16-1:0] node7767;
	wire [16-1:0] node7770;
	wire [16-1:0] node7772;
	wire [16-1:0] node7775;
	wire [16-1:0] node7776;
	wire [16-1:0] node7777;
	wire [16-1:0] node7781;
	wire [16-1:0] node7782;
	wire [16-1:0] node7784;
	wire [16-1:0] node7787;
	wire [16-1:0] node7790;
	wire [16-1:0] node7791;
	wire [16-1:0] node7792;
	wire [16-1:0] node7793;
	wire [16-1:0] node7794;
	wire [16-1:0] node7795;
	wire [16-1:0] node7796;
	wire [16-1:0] node7797;
	wire [16-1:0] node7800;
	wire [16-1:0] node7801;
	wire [16-1:0] node7806;
	wire [16-1:0] node7807;
	wire [16-1:0] node7808;
	wire [16-1:0] node7809;
	wire [16-1:0] node7813;
	wire [16-1:0] node7815;
	wire [16-1:0] node7818;
	wire [16-1:0] node7819;
	wire [16-1:0] node7821;
	wire [16-1:0] node7822;
	wire [16-1:0] node7826;
	wire [16-1:0] node7827;
	wire [16-1:0] node7829;
	wire [16-1:0] node7833;
	wire [16-1:0] node7834;
	wire [16-1:0] node7835;
	wire [16-1:0] node7836;
	wire [16-1:0] node7839;
	wire [16-1:0] node7841;
	wire [16-1:0] node7844;
	wire [16-1:0] node7845;
	wire [16-1:0] node7846;
	wire [16-1:0] node7848;
	wire [16-1:0] node7853;
	wire [16-1:0] node7854;
	wire [16-1:0] node7855;
	wire [16-1:0] node7856;
	wire [16-1:0] node7858;
	wire [16-1:0] node7862;
	wire [16-1:0] node7865;
	wire [16-1:0] node7867;
	wire [16-1:0] node7870;
	wire [16-1:0] node7871;
	wire [16-1:0] node7872;
	wire [16-1:0] node7873;
	wire [16-1:0] node7874;
	wire [16-1:0] node7875;
	wire [16-1:0] node7876;
	wire [16-1:0] node7882;
	wire [16-1:0] node7883;
	wire [16-1:0] node7884;
	wire [16-1:0] node7888;
	wire [16-1:0] node7891;
	wire [16-1:0] node7892;
	wire [16-1:0] node7894;
	wire [16-1:0] node7896;
	wire [16-1:0] node7899;
	wire [16-1:0] node7900;
	wire [16-1:0] node7901;
	wire [16-1:0] node7906;
	wire [16-1:0] node7907;
	wire [16-1:0] node7908;
	wire [16-1:0] node7909;
	wire [16-1:0] node7912;
	wire [16-1:0] node7915;
	wire [16-1:0] node7916;
	wire [16-1:0] node7917;
	wire [16-1:0] node7919;
	wire [16-1:0] node7922;
	wire [16-1:0] node7923;
	wire [16-1:0] node7927;
	wire [16-1:0] node7930;
	wire [16-1:0] node7931;
	wire [16-1:0] node7932;
	wire [16-1:0] node7936;
	wire [16-1:0] node7937;
	wire [16-1:0] node7938;
	wire [16-1:0] node7939;
	wire [16-1:0] node7944;
	wire [16-1:0] node7946;
	wire [16-1:0] node7949;
	wire [16-1:0] node7950;
	wire [16-1:0] node7951;
	wire [16-1:0] node7952;
	wire [16-1:0] node7953;
	wire [16-1:0] node7955;
	wire [16-1:0] node7958;
	wire [16-1:0] node7959;
	wire [16-1:0] node7960;
	wire [16-1:0] node7962;
	wire [16-1:0] node7967;
	wire [16-1:0] node7969;
	wire [16-1:0] node7970;
	wire [16-1:0] node7971;
	wire [16-1:0] node7975;
	wire [16-1:0] node7978;
	wire [16-1:0] node7979;
	wire [16-1:0] node7980;
	wire [16-1:0] node7982;
	wire [16-1:0] node7983;
	wire [16-1:0] node7987;
	wire [16-1:0] node7988;
	wire [16-1:0] node7990;
	wire [16-1:0] node7991;
	wire [16-1:0] node7995;
	wire [16-1:0] node7998;
	wire [16-1:0] node7999;
	wire [16-1:0] node8000;
	wire [16-1:0] node8002;
	wire [16-1:0] node8005;
	wire [16-1:0] node8006;
	wire [16-1:0] node8010;
	wire [16-1:0] node8012;
	wire [16-1:0] node8013;
	wire [16-1:0] node8015;
	wire [16-1:0] node8019;
	wire [16-1:0] node8020;
	wire [16-1:0] node8021;
	wire [16-1:0] node8022;
	wire [16-1:0] node8023;
	wire [16-1:0] node8024;
	wire [16-1:0] node8028;
	wire [16-1:0] node8029;
	wire [16-1:0] node8033;
	wire [16-1:0] node8034;
	wire [16-1:0] node8037;
	wire [16-1:0] node8039;
	wire [16-1:0] node8040;
	wire [16-1:0] node8044;
	wire [16-1:0] node8045;
	wire [16-1:0] node8046;
	wire [16-1:0] node8049;
	wire [16-1:0] node8050;
	wire [16-1:0] node8052;
	wire [16-1:0] node8056;
	wire [16-1:0] node8057;
	wire [16-1:0] node8058;
	wire [16-1:0] node8062;
	wire [16-1:0] node8065;
	wire [16-1:0] node8066;
	wire [16-1:0] node8067;
	wire [16-1:0] node8068;
	wire [16-1:0] node8069;
	wire [16-1:0] node8074;
	wire [16-1:0] node8076;
	wire [16-1:0] node8078;
	wire [16-1:0] node8081;
	wire [16-1:0] node8082;
	wire [16-1:0] node8083;
	wire [16-1:0] node8086;
	wire [16-1:0] node8088;
	wire [16-1:0] node8091;
	wire [16-1:0] node8094;
	wire [16-1:0] node8095;
	wire [16-1:0] node8096;
	wire [16-1:0] node8097;
	wire [16-1:0] node8098;
	wire [16-1:0] node8099;
	wire [16-1:0] node8100;
	wire [16-1:0] node8101;
	wire [16-1:0] node8102;
	wire [16-1:0] node8107;
	wire [16-1:0] node8110;
	wire [16-1:0] node8113;
	wire [16-1:0] node8115;
	wire [16-1:0] node8116;
	wire [16-1:0] node8118;
	wire [16-1:0] node8122;
	wire [16-1:0] node8123;
	wire [16-1:0] node8124;
	wire [16-1:0] node8126;
	wire [16-1:0] node8127;
	wire [16-1:0] node8131;
	wire [16-1:0] node8132;
	wire [16-1:0] node8133;
	wire [16-1:0] node8135;
	wire [16-1:0] node8139;
	wire [16-1:0] node8142;
	wire [16-1:0] node8143;
	wire [16-1:0] node8144;
	wire [16-1:0] node8145;
	wire [16-1:0] node8147;
	wire [16-1:0] node8151;
	wire [16-1:0] node8154;
	wire [16-1:0] node8155;
	wire [16-1:0] node8158;
	wire [16-1:0] node8160;
	wire [16-1:0] node8163;
	wire [16-1:0] node8164;
	wire [16-1:0] node8165;
	wire [16-1:0] node8166;
	wire [16-1:0] node8167;
	wire [16-1:0] node8168;
	wire [16-1:0] node8170;
	wire [16-1:0] node8174;
	wire [16-1:0] node8176;
	wire [16-1:0] node8179;
	wire [16-1:0] node8180;
	wire [16-1:0] node8182;
	wire [16-1:0] node8183;
	wire [16-1:0] node8187;
	wire [16-1:0] node8188;
	wire [16-1:0] node8190;
	wire [16-1:0] node8193;
	wire [16-1:0] node8196;
	wire [16-1:0] node8197;
	wire [16-1:0] node8198;
	wire [16-1:0] node8201;
	wire [16-1:0] node8202;
	wire [16-1:0] node8206;
	wire [16-1:0] node8207;
	wire [16-1:0] node8211;
	wire [16-1:0] node8212;
	wire [16-1:0] node8213;
	wire [16-1:0] node8214;
	wire [16-1:0] node8218;
	wire [16-1:0] node8219;
	wire [16-1:0] node8220;
	wire [16-1:0] node8222;
	wire [16-1:0] node8225;
	wire [16-1:0] node8227;
	wire [16-1:0] node8230;
	wire [16-1:0] node8233;
	wire [16-1:0] node8234;
	wire [16-1:0] node8236;
	wire [16-1:0] node8239;
	wire [16-1:0] node8240;
	wire [16-1:0] node8244;
	wire [16-1:0] node8245;
	wire [16-1:0] node8246;
	wire [16-1:0] node8247;
	wire [16-1:0] node8248;
	wire [16-1:0] node8249;
	wire [16-1:0] node8251;
	wire [16-1:0] node8255;
	wire [16-1:0] node8256;
	wire [16-1:0] node8259;
	wire [16-1:0] node8262;
	wire [16-1:0] node8263;
	wire [16-1:0] node8265;
	wire [16-1:0] node8266;
	wire [16-1:0] node8268;
	wire [16-1:0] node8272;
	wire [16-1:0] node8275;
	wire [16-1:0] node8276;
	wire [16-1:0] node8277;
	wire [16-1:0] node8278;
	wire [16-1:0] node8282;
	wire [16-1:0] node8284;
	wire [16-1:0] node8285;
	wire [16-1:0] node8287;
	wire [16-1:0] node8291;
	wire [16-1:0] node8292;
	wire [16-1:0] node8294;
	wire [16-1:0] node8297;
	wire [16-1:0] node8298;
	wire [16-1:0] node8301;
	wire [16-1:0] node8303;
	wire [16-1:0] node8306;
	wire [16-1:0] node8307;
	wire [16-1:0] node8308;
	wire [16-1:0] node8309;
	wire [16-1:0] node8312;
	wire [16-1:0] node8313;
	wire [16-1:0] node8317;
	wire [16-1:0] node8318;
	wire [16-1:0] node8320;
	wire [16-1:0] node8321;
	wire [16-1:0] node8323;
	wire [16-1:0] node8327;
	wire [16-1:0] node8328;
	wire [16-1:0] node8329;
	wire [16-1:0] node8331;
	wire [16-1:0] node8335;
	wire [16-1:0] node8338;
	wire [16-1:0] node8339;
	wire [16-1:0] node8340;
	wire [16-1:0] node8341;
	wire [16-1:0] node8344;
	wire [16-1:0] node8345;
	wire [16-1:0] node8347;
	wire [16-1:0] node8351;
	wire [16-1:0] node8352;
	wire [16-1:0] node8354;
	wire [16-1:0] node8356;
	wire [16-1:0] node8360;
	wire [16-1:0] node8361;
	wire [16-1:0] node8363;
	wire [16-1:0] node8366;
	wire [16-1:0] node8368;
	wire [16-1:0] node8371;
	wire [16-1:0] node8372;
	wire [16-1:0] node8373;
	wire [16-1:0] node8374;
	wire [16-1:0] node8375;
	wire [16-1:0] node8376;
	wire [16-1:0] node8377;
	wire [16-1:0] node8378;
	wire [16-1:0] node8379;
	wire [16-1:0] node8380;
	wire [16-1:0] node8381;
	wire [16-1:0] node8382;
	wire [16-1:0] node8383;
	wire [16-1:0] node8384;
	wire [16-1:0] node8388;
	wire [16-1:0] node8391;
	wire [16-1:0] node8392;
	wire [16-1:0] node8393;
	wire [16-1:0] node8397;
	wire [16-1:0] node8400;
	wire [16-1:0] node8401;
	wire [16-1:0] node8402;
	wire [16-1:0] node8407;
	wire [16-1:0] node8408;
	wire [16-1:0] node8409;
	wire [16-1:0] node8411;
	wire [16-1:0] node8412;
	wire [16-1:0] node8416;
	wire [16-1:0] node8420;
	wire [16-1:0] node8421;
	wire [16-1:0] node8422;
	wire [16-1:0] node8423;
	wire [16-1:0] node8426;
	wire [16-1:0] node8428;
	wire [16-1:0] node8429;
	wire [16-1:0] node8433;
	wire [16-1:0] node8434;
	wire [16-1:0] node8438;
	wire [16-1:0] node8439;
	wire [16-1:0] node8440;
	wire [16-1:0] node8441;
	wire [16-1:0] node8443;
	wire [16-1:0] node8447;
	wire [16-1:0] node8449;
	wire [16-1:0] node8452;
	wire [16-1:0] node8453;
	wire [16-1:0] node8455;
	wire [16-1:0] node8458;
	wire [16-1:0] node8461;
	wire [16-1:0] node8462;
	wire [16-1:0] node8463;
	wire [16-1:0] node8464;
	wire [16-1:0] node8465;
	wire [16-1:0] node8467;
	wire [16-1:0] node8470;
	wire [16-1:0] node8473;
	wire [16-1:0] node8474;
	wire [16-1:0] node8478;
	wire [16-1:0] node8479;
	wire [16-1:0] node8480;
	wire [16-1:0] node8482;
	wire [16-1:0] node8485;
	wire [16-1:0] node8488;
	wire [16-1:0] node8489;
	wire [16-1:0] node8490;
	wire [16-1:0] node8495;
	wire [16-1:0] node8496;
	wire [16-1:0] node8497;
	wire [16-1:0] node8499;
	wire [16-1:0] node8502;
	wire [16-1:0] node8503;
	wire [16-1:0] node8507;
	wire [16-1:0] node8508;
	wire [16-1:0] node8509;
	wire [16-1:0] node8510;
	wire [16-1:0] node8512;
	wire [16-1:0] node8516;
	wire [16-1:0] node8517;
	wire [16-1:0] node8521;
	wire [16-1:0] node8523;
	wire [16-1:0] node8524;
	wire [16-1:0] node8525;
	wire [16-1:0] node8530;
	wire [16-1:0] node8531;
	wire [16-1:0] node8532;
	wire [16-1:0] node8533;
	wire [16-1:0] node8535;
	wire [16-1:0] node8536;
	wire [16-1:0] node8540;
	wire [16-1:0] node8541;
	wire [16-1:0] node8542;
	wire [16-1:0] node8545;
	wire [16-1:0] node8548;
	wire [16-1:0] node8551;
	wire [16-1:0] node8552;
	wire [16-1:0] node8553;
	wire [16-1:0] node8556;
	wire [16-1:0] node8557;
	wire [16-1:0] node8559;
	wire [16-1:0] node8560;
	wire [16-1:0] node8564;
	wire [16-1:0] node8566;
	wire [16-1:0] node8569;
	wire [16-1:0] node8571;
	wire [16-1:0] node8572;
	wire [16-1:0] node8574;
	wire [16-1:0] node8578;
	wire [16-1:0] node8579;
	wire [16-1:0] node8580;
	wire [16-1:0] node8581;
	wire [16-1:0] node8582;
	wire [16-1:0] node8583;
	wire [16-1:0] node8586;
	wire [16-1:0] node8587;
	wire [16-1:0] node8591;
	wire [16-1:0] node8593;
	wire [16-1:0] node8594;
	wire [16-1:0] node8597;
	wire [16-1:0] node8600;
	wire [16-1:0] node8601;
	wire [16-1:0] node8602;
	wire [16-1:0] node8607;
	wire [16-1:0] node8608;
	wire [16-1:0] node8610;
	wire [16-1:0] node8611;
	wire [16-1:0] node8613;
	wire [16-1:0] node8617;
	wire [16-1:0] node8620;
	wire [16-1:0] node8621;
	wire [16-1:0] node8622;
	wire [16-1:0] node8623;
	wire [16-1:0] node8626;
	wire [16-1:0] node8627;
	wire [16-1:0] node8632;
	wire [16-1:0] node8633;
	wire [16-1:0] node8635;
	wire [16-1:0] node8638;
	wire [16-1:0] node8639;
	wire [16-1:0] node8642;
	wire [16-1:0] node8643;
	wire [16-1:0] node8647;
	wire [16-1:0] node8648;
	wire [16-1:0] node8649;
	wire [16-1:0] node8650;
	wire [16-1:0] node8651;
	wire [16-1:0] node8652;
	wire [16-1:0] node8653;
	wire [16-1:0] node8657;
	wire [16-1:0] node8658;
	wire [16-1:0] node8661;
	wire [16-1:0] node8664;
	wire [16-1:0] node8665;
	wire [16-1:0] node8667;
	wire [16-1:0] node8670;
	wire [16-1:0] node8671;
	wire [16-1:0] node8673;
	wire [16-1:0] node8676;
	wire [16-1:0] node8679;
	wire [16-1:0] node8680;
	wire [16-1:0] node8681;
	wire [16-1:0] node8682;
	wire [16-1:0] node8683;
	wire [16-1:0] node8688;
	wire [16-1:0] node8689;
	wire [16-1:0] node8692;
	wire [16-1:0] node8695;
	wire [16-1:0] node8696;
	wire [16-1:0] node8697;
	wire [16-1:0] node8700;
	wire [16-1:0] node8702;
	wire [16-1:0] node8705;
	wire [16-1:0] node8706;
	wire [16-1:0] node8709;
	wire [16-1:0] node8712;
	wire [16-1:0] node8713;
	wire [16-1:0] node8714;
	wire [16-1:0] node8715;
	wire [16-1:0] node8716;
	wire [16-1:0] node8719;
	wire [16-1:0] node8721;
	wire [16-1:0] node8722;
	wire [16-1:0] node8726;
	wire [16-1:0] node8727;
	wire [16-1:0] node8728;
	wire [16-1:0] node8732;
	wire [16-1:0] node8735;
	wire [16-1:0] node8736;
	wire [16-1:0] node8738;
	wire [16-1:0] node8740;
	wire [16-1:0] node8743;
	wire [16-1:0] node8746;
	wire [16-1:0] node8747;
	wire [16-1:0] node8748;
	wire [16-1:0] node8750;
	wire [16-1:0] node8751;
	wire [16-1:0] node8755;
	wire [16-1:0] node8756;
	wire [16-1:0] node8759;
	wire [16-1:0] node8761;
	wire [16-1:0] node8764;
	wire [16-1:0] node8765;
	wire [16-1:0] node8766;
	wire [16-1:0] node8770;
	wire [16-1:0] node8773;
	wire [16-1:0] node8774;
	wire [16-1:0] node8775;
	wire [16-1:0] node8776;
	wire [16-1:0] node8777;
	wire [16-1:0] node8778;
	wire [16-1:0] node8779;
	wire [16-1:0] node8783;
	wire [16-1:0] node8785;
	wire [16-1:0] node8788;
	wire [16-1:0] node8789;
	wire [16-1:0] node8792;
	wire [16-1:0] node8795;
	wire [16-1:0] node8796;
	wire [16-1:0] node8798;
	wire [16-1:0] node8801;
	wire [16-1:0] node8802;
	wire [16-1:0] node8804;
	wire [16-1:0] node8808;
	wire [16-1:0] node8809;
	wire [16-1:0] node8810;
	wire [16-1:0] node8811;
	wire [16-1:0] node8812;
	wire [16-1:0] node8817;
	wire [16-1:0] node8820;
	wire [16-1:0] node8821;
	wire [16-1:0] node8822;
	wire [16-1:0] node8823;
	wire [16-1:0] node8827;
	wire [16-1:0] node8830;
	wire [16-1:0] node8831;
	wire [16-1:0] node8832;
	wire [16-1:0] node8837;
	wire [16-1:0] node8838;
	wire [16-1:0] node8839;
	wire [16-1:0] node8841;
	wire [16-1:0] node8842;
	wire [16-1:0] node8846;
	wire [16-1:0] node8847;
	wire [16-1:0] node8848;
	wire [16-1:0] node8852;
	wire [16-1:0] node8853;
	wire [16-1:0] node8855;
	wire [16-1:0] node8856;
	wire [16-1:0] node8861;
	wire [16-1:0] node8862;
	wire [16-1:0] node8863;
	wire [16-1:0] node8865;
	wire [16-1:0] node8868;
	wire [16-1:0] node8869;
	wire [16-1:0] node8873;
	wire [16-1:0] node8875;
	wire [16-1:0] node8876;
	wire [16-1:0] node8877;
	wire [16-1:0] node8879;
	wire [16-1:0] node8884;
	wire [16-1:0] node8885;
	wire [16-1:0] node8886;
	wire [16-1:0] node8887;
	wire [16-1:0] node8888;
	wire [16-1:0] node8889;
	wire [16-1:0] node8890;
	wire [16-1:0] node8891;
	wire [16-1:0] node8892;
	wire [16-1:0] node8897;
	wire [16-1:0] node8898;
	wire [16-1:0] node8901;
	wire [16-1:0] node8903;
	wire [16-1:0] node8906;
	wire [16-1:0] node8907;
	wire [16-1:0] node8908;
	wire [16-1:0] node8909;
	wire [16-1:0] node8913;
	wire [16-1:0] node8916;
	wire [16-1:0] node8919;
	wire [16-1:0] node8920;
	wire [16-1:0] node8921;
	wire [16-1:0] node8922;
	wire [16-1:0] node8923;
	wire [16-1:0] node8927;
	wire [16-1:0] node8929;
	wire [16-1:0] node8933;
	wire [16-1:0] node8934;
	wire [16-1:0] node8935;
	wire [16-1:0] node8936;
	wire [16-1:0] node8937;
	wire [16-1:0] node8942;
	wire [16-1:0] node8943;
	wire [16-1:0] node8944;
	wire [16-1:0] node8949;
	wire [16-1:0] node8950;
	wire [16-1:0] node8952;
	wire [16-1:0] node8953;
	wire [16-1:0] node8957;
	wire [16-1:0] node8960;
	wire [16-1:0] node8961;
	wire [16-1:0] node8962;
	wire [16-1:0] node8963;
	wire [16-1:0] node8964;
	wire [16-1:0] node8967;
	wire [16-1:0] node8969;
	wire [16-1:0] node8972;
	wire [16-1:0] node8975;
	wire [16-1:0] node8976;
	wire [16-1:0] node8977;
	wire [16-1:0] node8979;
	wire [16-1:0] node8980;
	wire [16-1:0] node8984;
	wire [16-1:0] node8987;
	wire [16-1:0] node8988;
	wire [16-1:0] node8989;
	wire [16-1:0] node8993;
	wire [16-1:0] node8995;
	wire [16-1:0] node8998;
	wire [16-1:0] node8999;
	wire [16-1:0] node9000;
	wire [16-1:0] node9002;
	wire [16-1:0] node9003;
	wire [16-1:0] node9005;
	wire [16-1:0] node9010;
	wire [16-1:0] node9011;
	wire [16-1:0] node9012;
	wire [16-1:0] node9015;
	wire [16-1:0] node9017;
	wire [16-1:0] node9021;
	wire [16-1:0] node9022;
	wire [16-1:0] node9023;
	wire [16-1:0] node9024;
	wire [16-1:0] node9025;
	wire [16-1:0] node9026;
	wire [16-1:0] node9030;
	wire [16-1:0] node9031;
	wire [16-1:0] node9035;
	wire [16-1:0] node9036;
	wire [16-1:0] node9038;
	wire [16-1:0] node9039;
	wire [16-1:0] node9041;
	wire [16-1:0] node9045;
	wire [16-1:0] node9046;
	wire [16-1:0] node9049;
	wire [16-1:0] node9050;
	wire [16-1:0] node9054;
	wire [16-1:0] node9055;
	wire [16-1:0] node9056;
	wire [16-1:0] node9057;
	wire [16-1:0] node9060;
	wire [16-1:0] node9063;
	wire [16-1:0] node9064;
	wire [16-1:0] node9066;
	wire [16-1:0] node9069;
	wire [16-1:0] node9070;
	wire [16-1:0] node9071;
	wire [16-1:0] node9076;
	wire [16-1:0] node9077;
	wire [16-1:0] node9078;
	wire [16-1:0] node9082;
	wire [16-1:0] node9084;
	wire [16-1:0] node9086;
	wire [16-1:0] node9089;
	wire [16-1:0] node9090;
	wire [16-1:0] node9091;
	wire [16-1:0] node9092;
	wire [16-1:0] node9093;
	wire [16-1:0] node9096;
	wire [16-1:0] node9097;
	wire [16-1:0] node9101;
	wire [16-1:0] node9102;
	wire [16-1:0] node9106;
	wire [16-1:0] node9107;
	wire [16-1:0] node9108;
	wire [16-1:0] node9109;
	wire [16-1:0] node9111;
	wire [16-1:0] node9115;
	wire [16-1:0] node9117;
	wire [16-1:0] node9118;
	wire [16-1:0] node9122;
	wire [16-1:0] node9123;
	wire [16-1:0] node9124;
	wire [16-1:0] node9128;
	wire [16-1:0] node9131;
	wire [16-1:0] node9132;
	wire [16-1:0] node9133;
	wire [16-1:0] node9135;
	wire [16-1:0] node9139;
	wire [16-1:0] node9140;
	wire [16-1:0] node9143;
	wire [16-1:0] node9145;
	wire [16-1:0] node9146;
	wire [16-1:0] node9150;
	wire [16-1:0] node9151;
	wire [16-1:0] node9152;
	wire [16-1:0] node9153;
	wire [16-1:0] node9154;
	wire [16-1:0] node9155;
	wire [16-1:0] node9156;
	wire [16-1:0] node9158;
	wire [16-1:0] node9159;
	wire [16-1:0] node9163;
	wire [16-1:0] node9166;
	wire [16-1:0] node9169;
	wire [16-1:0] node9170;
	wire [16-1:0] node9171;
	wire [16-1:0] node9174;
	wire [16-1:0] node9176;
	wire [16-1:0] node9179;
	wire [16-1:0] node9180;
	wire [16-1:0] node9181;
	wire [16-1:0] node9185;
	wire [16-1:0] node9186;
	wire [16-1:0] node9190;
	wire [16-1:0] node9191;
	wire [16-1:0] node9192;
	wire [16-1:0] node9195;
	wire [16-1:0] node9196;
	wire [16-1:0] node9199;
	wire [16-1:0] node9202;
	wire [16-1:0] node9204;
	wire [16-1:0] node9205;
	wire [16-1:0] node9206;
	wire [16-1:0] node9210;
	wire [16-1:0] node9213;
	wire [16-1:0] node9214;
	wire [16-1:0] node9215;
	wire [16-1:0] node9216;
	wire [16-1:0] node9217;
	wire [16-1:0] node9220;
	wire [16-1:0] node9221;
	wire [16-1:0] node9225;
	wire [16-1:0] node9227;
	wire [16-1:0] node9230;
	wire [16-1:0] node9231;
	wire [16-1:0] node9232;
	wire [16-1:0] node9233;
	wire [16-1:0] node9235;
	wire [16-1:0] node9239;
	wire [16-1:0] node9242;
	wire [16-1:0] node9243;
	wire [16-1:0] node9245;
	wire [16-1:0] node9246;
	wire [16-1:0] node9251;
	wire [16-1:0] node9252;
	wire [16-1:0] node9254;
	wire [16-1:0] node9255;
	wire [16-1:0] node9257;
	wire [16-1:0] node9259;
	wire [16-1:0] node9263;
	wire [16-1:0] node9264;
	wire [16-1:0] node9265;
	wire [16-1:0] node9267;
	wire [16-1:0] node9270;
	wire [16-1:0] node9274;
	wire [16-1:0] node9275;
	wire [16-1:0] node9276;
	wire [16-1:0] node9277;
	wire [16-1:0] node9278;
	wire [16-1:0] node9279;
	wire [16-1:0] node9281;
	wire [16-1:0] node9284;
	wire [16-1:0] node9287;
	wire [16-1:0] node9288;
	wire [16-1:0] node9292;
	wire [16-1:0] node9293;
	wire [16-1:0] node9294;
	wire [16-1:0] node9298;
	wire [16-1:0] node9300;
	wire [16-1:0] node9301;
	wire [16-1:0] node9302;
	wire [16-1:0] node9306;
	wire [16-1:0] node9309;
	wire [16-1:0] node9310;
	wire [16-1:0] node9311;
	wire [16-1:0] node9312;
	wire [16-1:0] node9313;
	wire [16-1:0] node9317;
	wire [16-1:0] node9318;
	wire [16-1:0] node9322;
	wire [16-1:0] node9325;
	wire [16-1:0] node9326;
	wire [16-1:0] node9328;
	wire [16-1:0] node9331;
	wire [16-1:0] node9334;
	wire [16-1:0] node9335;
	wire [16-1:0] node9336;
	wire [16-1:0] node9337;
	wire [16-1:0] node9338;
	wire [16-1:0] node9341;
	wire [16-1:0] node9343;
	wire [16-1:0] node9346;
	wire [16-1:0] node9348;
	wire [16-1:0] node9349;
	wire [16-1:0] node9351;
	wire [16-1:0] node9355;
	wire [16-1:0] node9356;
	wire [16-1:0] node9357;
	wire [16-1:0] node9360;
	wire [16-1:0] node9363;
	wire [16-1:0] node9364;
	wire [16-1:0] node9365;
	wire [16-1:0] node9370;
	wire [16-1:0] node9371;
	wire [16-1:0] node9372;
	wire [16-1:0] node9374;
	wire [16-1:0] node9376;
	wire [16-1:0] node9379;
	wire [16-1:0] node9381;
	wire [16-1:0] node9384;
	wire [16-1:0] node9385;
	wire [16-1:0] node9387;
	wire [16-1:0] node9389;
	wire [16-1:0] node9392;
	wire [16-1:0] node9393;
	wire [16-1:0] node9394;
	wire [16-1:0] node9398;
	wire [16-1:0] node9400;
	wire [16-1:0] node9402;
	wire [16-1:0] node9405;
	wire [16-1:0] node9406;
	wire [16-1:0] node9407;
	wire [16-1:0] node9408;
	wire [16-1:0] node9409;
	wire [16-1:0] node9410;
	wire [16-1:0] node9411;
	wire [16-1:0] node9412;
	wire [16-1:0] node9414;
	wire [16-1:0] node9416;
	wire [16-1:0] node9419;
	wire [16-1:0] node9420;
	wire [16-1:0] node9421;
	wire [16-1:0] node9426;
	wire [16-1:0] node9427;
	wire [16-1:0] node9429;
	wire [16-1:0] node9431;
	wire [16-1:0] node9432;
	wire [16-1:0] node9436;
	wire [16-1:0] node9437;
	wire [16-1:0] node9438;
	wire [16-1:0] node9440;
	wire [16-1:0] node9444;
	wire [16-1:0] node9447;
	wire [16-1:0] node9448;
	wire [16-1:0] node9449;
	wire [16-1:0] node9450;
	wire [16-1:0] node9451;
	wire [16-1:0] node9456;
	wire [16-1:0] node9457;
	wire [16-1:0] node9461;
	wire [16-1:0] node9462;
	wire [16-1:0] node9464;
	wire [16-1:0] node9465;
	wire [16-1:0] node9469;
	wire [16-1:0] node9470;
	wire [16-1:0] node9473;
	wire [16-1:0] node9475;
	wire [16-1:0] node9476;
	wire [16-1:0] node9480;
	wire [16-1:0] node9481;
	wire [16-1:0] node9482;
	wire [16-1:0] node9483;
	wire [16-1:0] node9484;
	wire [16-1:0] node9485;
	wire [16-1:0] node9490;
	wire [16-1:0] node9491;
	wire [16-1:0] node9492;
	wire [16-1:0] node9496;
	wire [16-1:0] node9499;
	wire [16-1:0] node9500;
	wire [16-1:0] node9502;
	wire [16-1:0] node9504;
	wire [16-1:0] node9505;
	wire [16-1:0] node9509;
	wire [16-1:0] node9510;
	wire [16-1:0] node9513;
	wire [16-1:0] node9514;
	wire [16-1:0] node9515;
	wire [16-1:0] node9520;
	wire [16-1:0] node9521;
	wire [16-1:0] node9522;
	wire [16-1:0] node9523;
	wire [16-1:0] node9527;
	wire [16-1:0] node9528;
	wire [16-1:0] node9529;
	wire [16-1:0] node9531;
	wire [16-1:0] node9535;
	wire [16-1:0] node9536;
	wire [16-1:0] node9540;
	wire [16-1:0] node9541;
	wire [16-1:0] node9543;
	wire [16-1:0] node9545;
	wire [16-1:0] node9546;
	wire [16-1:0] node9550;
	wire [16-1:0] node9551;
	wire [16-1:0] node9554;
	wire [16-1:0] node9557;
	wire [16-1:0] node9558;
	wire [16-1:0] node9559;
	wire [16-1:0] node9560;
	wire [16-1:0] node9561;
	wire [16-1:0] node9562;
	wire [16-1:0] node9565;
	wire [16-1:0] node9568;
	wire [16-1:0] node9569;
	wire [16-1:0] node9573;
	wire [16-1:0] node9574;
	wire [16-1:0] node9575;
	wire [16-1:0] node9578;
	wire [16-1:0] node9580;
	wire [16-1:0] node9583;
	wire [16-1:0] node9584;
	wire [16-1:0] node9586;
	wire [16-1:0] node9588;
	wire [16-1:0] node9591;
	wire [16-1:0] node9593;
	wire [16-1:0] node9596;
	wire [16-1:0] node9597;
	wire [16-1:0] node9598;
	wire [16-1:0] node9599;
	wire [16-1:0] node9602;
	wire [16-1:0] node9603;
	wire [16-1:0] node9605;
	wire [16-1:0] node9609;
	wire [16-1:0] node9610;
	wire [16-1:0] node9611;
	wire [16-1:0] node9615;
	wire [16-1:0] node9618;
	wire [16-1:0] node9619;
	wire [16-1:0] node9620;
	wire [16-1:0] node9623;
	wire [16-1:0] node9625;
	wire [16-1:0] node9628;
	wire [16-1:0] node9629;
	wire [16-1:0] node9633;
	wire [16-1:0] node9634;
	wire [16-1:0] node9635;
	wire [16-1:0] node9636;
	wire [16-1:0] node9638;
	wire [16-1:0] node9640;
	wire [16-1:0] node9641;
	wire [16-1:0] node9645;
	wire [16-1:0] node9646;
	wire [16-1:0] node9647;
	wire [16-1:0] node9651;
	wire [16-1:0] node9654;
	wire [16-1:0] node9655;
	wire [16-1:0] node9656;
	wire [16-1:0] node9659;
	wire [16-1:0] node9662;
	wire [16-1:0] node9663;
	wire [16-1:0] node9666;
	wire [16-1:0] node9669;
	wire [16-1:0] node9670;
	wire [16-1:0] node9671;
	wire [16-1:0] node9672;
	wire [16-1:0] node9675;
	wire [16-1:0] node9678;
	wire [16-1:0] node9679;
	wire [16-1:0] node9680;
	wire [16-1:0] node9682;
	wire [16-1:0] node9685;
	wire [16-1:0] node9688;
	wire [16-1:0] node9689;
	wire [16-1:0] node9691;
	wire [16-1:0] node9695;
	wire [16-1:0] node9696;
	wire [16-1:0] node9699;
	wire [16-1:0] node9702;
	wire [16-1:0] node9703;
	wire [16-1:0] node9704;
	wire [16-1:0] node9705;
	wire [16-1:0] node9706;
	wire [16-1:0] node9707;
	wire [16-1:0] node9708;
	wire [16-1:0] node9709;
	wire [16-1:0] node9710;
	wire [16-1:0] node9715;
	wire [16-1:0] node9717;
	wire [16-1:0] node9720;
	wire [16-1:0] node9721;
	wire [16-1:0] node9724;
	wire [16-1:0] node9726;
	wire [16-1:0] node9729;
	wire [16-1:0] node9730;
	wire [16-1:0] node9731;
	wire [16-1:0] node9734;
	wire [16-1:0] node9737;
	wire [16-1:0] node9739;
	wire [16-1:0] node9742;
	wire [16-1:0] node9743;
	wire [16-1:0] node9744;
	wire [16-1:0] node9745;
	wire [16-1:0] node9746;
	wire [16-1:0] node9748;
	wire [16-1:0] node9751;
	wire [16-1:0] node9753;
	wire [16-1:0] node9757;
	wire [16-1:0] node9758;
	wire [16-1:0] node9761;
	wire [16-1:0] node9763;
	wire [16-1:0] node9764;
	wire [16-1:0] node9768;
	wire [16-1:0] node9769;
	wire [16-1:0] node9770;
	wire [16-1:0] node9773;
	wire [16-1:0] node9776;
	wire [16-1:0] node9778;
	wire [16-1:0] node9781;
	wire [16-1:0] node9782;
	wire [16-1:0] node9783;
	wire [16-1:0] node9784;
	wire [16-1:0] node9787;
	wire [16-1:0] node9788;
	wire [16-1:0] node9792;
	wire [16-1:0] node9793;
	wire [16-1:0] node9794;
	wire [16-1:0] node9795;
	wire [16-1:0] node9799;
	wire [16-1:0] node9801;
	wire [16-1:0] node9802;
	wire [16-1:0] node9806;
	wire [16-1:0] node9809;
	wire [16-1:0] node9810;
	wire [16-1:0] node9811;
	wire [16-1:0] node9812;
	wire [16-1:0] node9815;
	wire [16-1:0] node9817;
	wire [16-1:0] node9820;
	wire [16-1:0] node9821;
	wire [16-1:0] node9822;
	wire [16-1:0] node9824;
	wire [16-1:0] node9829;
	wire [16-1:0] node9830;
	wire [16-1:0] node9832;
	wire [16-1:0] node9835;
	wire [16-1:0] node9836;
	wire [16-1:0] node9837;
	wire [16-1:0] node9841;
	wire [16-1:0] node9844;
	wire [16-1:0] node9845;
	wire [16-1:0] node9846;
	wire [16-1:0] node9847;
	wire [16-1:0] node9848;
	wire [16-1:0] node9849;
	wire [16-1:0] node9853;
	wire [16-1:0] node9854;
	wire [16-1:0] node9855;
	wire [16-1:0] node9857;
	wire [16-1:0] node9862;
	wire [16-1:0] node9863;
	wire [16-1:0] node9866;
	wire [16-1:0] node9867;
	wire [16-1:0] node9870;
	wire [16-1:0] node9873;
	wire [16-1:0] node9874;
	wire [16-1:0] node9875;
	wire [16-1:0] node9876;
	wire [16-1:0] node9878;
	wire [16-1:0] node9881;
	wire [16-1:0] node9884;
	wire [16-1:0] node9885;
	wire [16-1:0] node9887;
	wire [16-1:0] node9888;
	wire [16-1:0] node9893;
	wire [16-1:0] node9894;
	wire [16-1:0] node9895;
	wire [16-1:0] node9896;
	wire [16-1:0] node9900;
	wire [16-1:0] node9902;
	wire [16-1:0] node9905;
	wire [16-1:0] node9906;
	wire [16-1:0] node9907;
	wire [16-1:0] node9909;
	wire [16-1:0] node9913;
	wire [16-1:0] node9916;
	wire [16-1:0] node9917;
	wire [16-1:0] node9918;
	wire [16-1:0] node9919;
	wire [16-1:0] node9920;
	wire [16-1:0] node9922;
	wire [16-1:0] node9924;
	wire [16-1:0] node9929;
	wire [16-1:0] node9931;
	wire [16-1:0] node9932;
	wire [16-1:0] node9935;
	wire [16-1:0] node9938;
	wire [16-1:0] node9939;
	wire [16-1:0] node9940;
	wire [16-1:0] node9941;
	wire [16-1:0] node9944;
	wire [16-1:0] node9948;
	wire [16-1:0] node9949;
	wire [16-1:0] node9950;
	wire [16-1:0] node9953;
	wire [16-1:0] node9956;
	wire [16-1:0] node9958;
	wire [16-1:0] node9961;
	wire [16-1:0] node9962;
	wire [16-1:0] node9963;
	wire [16-1:0] node9964;
	wire [16-1:0] node9965;
	wire [16-1:0] node9966;
	wire [16-1:0] node9967;
	wire [16-1:0] node9968;
	wire [16-1:0] node9971;
	wire [16-1:0] node9974;
	wire [16-1:0] node9975;
	wire [16-1:0] node9978;
	wire [16-1:0] node9980;
	wire [16-1:0] node9983;
	wire [16-1:0] node9985;
	wire [16-1:0] node9986;
	wire [16-1:0] node9987;
	wire [16-1:0] node9988;
	wire [16-1:0] node9993;
	wire [16-1:0] node9994;
	wire [16-1:0] node9998;
	wire [16-1:0] node9999;
	wire [16-1:0] node10000;
	wire [16-1:0] node10001;
	wire [16-1:0] node10003;
	wire [16-1:0] node10006;
	wire [16-1:0] node10009;
	wire [16-1:0] node10010;
	wire [16-1:0] node10013;
	wire [16-1:0] node10016;
	wire [16-1:0] node10017;
	wire [16-1:0] node10019;
	wire [16-1:0] node10020;
	wire [16-1:0] node10024;
	wire [16-1:0] node10026;
	wire [16-1:0] node10029;
	wire [16-1:0] node10030;
	wire [16-1:0] node10031;
	wire [16-1:0] node10032;
	wire [16-1:0] node10033;
	wire [16-1:0] node10034;
	wire [16-1:0] node10038;
	wire [16-1:0] node10041;
	wire [16-1:0] node10044;
	wire [16-1:0] node10045;
	wire [16-1:0] node10046;
	wire [16-1:0] node10047;
	wire [16-1:0] node10049;
	wire [16-1:0] node10053;
	wire [16-1:0] node10056;
	wire [16-1:0] node10057;
	wire [16-1:0] node10060;
	wire [16-1:0] node10063;
	wire [16-1:0] node10064;
	wire [16-1:0] node10065;
	wire [16-1:0] node10067;
	wire [16-1:0] node10070;
	wire [16-1:0] node10071;
	wire [16-1:0] node10074;
	wire [16-1:0] node10077;
	wire [16-1:0] node10078;
	wire [16-1:0] node10079;
	wire [16-1:0] node10080;
	wire [16-1:0] node10084;
	wire [16-1:0] node10087;
	wire [16-1:0] node10090;
	wire [16-1:0] node10091;
	wire [16-1:0] node10092;
	wire [16-1:0] node10093;
	wire [16-1:0] node10094;
	wire [16-1:0] node10097;
	wire [16-1:0] node10098;
	wire [16-1:0] node10099;
	wire [16-1:0] node10101;
	wire [16-1:0] node10105;
	wire [16-1:0] node10108;
	wire [16-1:0] node10109;
	wire [16-1:0] node10110;
	wire [16-1:0] node10112;
	wire [16-1:0] node10115;
	wire [16-1:0] node10116;
	wire [16-1:0] node10120;
	wire [16-1:0] node10123;
	wire [16-1:0] node10124;
	wire [16-1:0] node10125;
	wire [16-1:0] node10127;
	wire [16-1:0] node10130;
	wire [16-1:0] node10131;
	wire [16-1:0] node10132;
	wire [16-1:0] node10136;
	wire [16-1:0] node10138;
	wire [16-1:0] node10141;
	wire [16-1:0] node10142;
	wire [16-1:0] node10144;
	wire [16-1:0] node10147;
	wire [16-1:0] node10150;
	wire [16-1:0] node10151;
	wire [16-1:0] node10152;
	wire [16-1:0] node10153;
	wire [16-1:0] node10155;
	wire [16-1:0] node10158;
	wire [16-1:0] node10161;
	wire [16-1:0] node10162;
	wire [16-1:0] node10163;
	wire [16-1:0] node10167;
	wire [16-1:0] node10168;
	wire [16-1:0] node10171;
	wire [16-1:0] node10173;
	wire [16-1:0] node10176;
	wire [16-1:0] node10177;
	wire [16-1:0] node10178;
	wire [16-1:0] node10181;
	wire [16-1:0] node10183;
	wire [16-1:0] node10184;
	wire [16-1:0] node10188;
	wire [16-1:0] node10189;
	wire [16-1:0] node10191;
	wire [16-1:0] node10193;
	wire [16-1:0] node10195;
	wire [16-1:0] node10198;
	wire [16-1:0] node10200;
	wire [16-1:0] node10201;
	wire [16-1:0] node10203;
	wire [16-1:0] node10206;
	wire [16-1:0] node10208;
	wire [16-1:0] node10211;
	wire [16-1:0] node10212;
	wire [16-1:0] node10213;
	wire [16-1:0] node10214;
	wire [16-1:0] node10215;
	wire [16-1:0] node10216;
	wire [16-1:0] node10219;
	wire [16-1:0] node10221;
	wire [16-1:0] node10222;
	wire [16-1:0] node10226;
	wire [16-1:0] node10227;
	wire [16-1:0] node10228;
	wire [16-1:0] node10229;
	wire [16-1:0] node10231;
	wire [16-1:0] node10235;
	wire [16-1:0] node10237;
	wire [16-1:0] node10240;
	wire [16-1:0] node10243;
	wire [16-1:0] node10244;
	wire [16-1:0] node10245;
	wire [16-1:0] node10247;
	wire [16-1:0] node10250;
	wire [16-1:0] node10251;
	wire [16-1:0] node10255;
	wire [16-1:0] node10256;
	wire [16-1:0] node10257;
	wire [16-1:0] node10261;
	wire [16-1:0] node10262;
	wire [16-1:0] node10265;
	wire [16-1:0] node10268;
	wire [16-1:0] node10269;
	wire [16-1:0] node10270;
	wire [16-1:0] node10271;
	wire [16-1:0] node10272;
	wire [16-1:0] node10275;
	wire [16-1:0] node10278;
	wire [16-1:0] node10279;
	wire [16-1:0] node10282;
	wire [16-1:0] node10284;
	wire [16-1:0] node10287;
	wire [16-1:0] node10288;
	wire [16-1:0] node10290;
	wire [16-1:0] node10291;
	wire [16-1:0] node10292;
	wire [16-1:0] node10295;
	wire [16-1:0] node10299;
	wire [16-1:0] node10301;
	wire [16-1:0] node10302;
	wire [16-1:0] node10306;
	wire [16-1:0] node10307;
	wire [16-1:0] node10308;
	wire [16-1:0] node10310;
	wire [16-1:0] node10313;
	wire [16-1:0] node10315;
	wire [16-1:0] node10316;
	wire [16-1:0] node10318;
	wire [16-1:0] node10322;
	wire [16-1:0] node10324;
	wire [16-1:0] node10325;
	wire [16-1:0] node10329;
	wire [16-1:0] node10330;
	wire [16-1:0] node10331;
	wire [16-1:0] node10332;
	wire [16-1:0] node10333;
	wire [16-1:0] node10334;
	wire [16-1:0] node10336;
	wire [16-1:0] node10339;
	wire [16-1:0] node10342;
	wire [16-1:0] node10343;
	wire [16-1:0] node10346;
	wire [16-1:0] node10349;
	wire [16-1:0] node10350;
	wire [16-1:0] node10353;
	wire [16-1:0] node10355;
	wire [16-1:0] node10358;
	wire [16-1:0] node10359;
	wire [16-1:0] node10360;
	wire [16-1:0] node10361;
	wire [16-1:0] node10363;
	wire [16-1:0] node10366;
	wire [16-1:0] node10369;
	wire [16-1:0] node10370;
	wire [16-1:0] node10371;
	wire [16-1:0] node10375;
	wire [16-1:0] node10378;
	wire [16-1:0] node10379;
	wire [16-1:0] node10380;
	wire [16-1:0] node10382;
	wire [16-1:0] node10385;
	wire [16-1:0] node10386;
	wire [16-1:0] node10388;
	wire [16-1:0] node10392;
	wire [16-1:0] node10393;
	wire [16-1:0] node10394;
	wire [16-1:0] node10398;
	wire [16-1:0] node10399;
	wire [16-1:0] node10401;
	wire [16-1:0] node10405;
	wire [16-1:0] node10406;
	wire [16-1:0] node10407;
	wire [16-1:0] node10409;
	wire [16-1:0] node10410;
	wire [16-1:0] node10412;
	wire [16-1:0] node10415;
	wire [16-1:0] node10416;
	wire [16-1:0] node10420;
	wire [16-1:0] node10421;
	wire [16-1:0] node10423;
	wire [16-1:0] node10426;
	wire [16-1:0] node10427;
	wire [16-1:0] node10428;
	wire [16-1:0] node10430;
	wire [16-1:0] node10434;
	wire [16-1:0] node10435;
	wire [16-1:0] node10437;
	wire [16-1:0] node10441;
	wire [16-1:0] node10442;
	wire [16-1:0] node10443;
	wire [16-1:0] node10445;
	wire [16-1:0] node10447;
	wire [16-1:0] node10448;
	wire [16-1:0] node10452;
	wire [16-1:0] node10453;
	wire [16-1:0] node10456;
	wire [16-1:0] node10457;
	wire [16-1:0] node10461;
	wire [16-1:0] node10462;
	wire [16-1:0] node10463;
	wire [16-1:0] node10464;
	wire [16-1:0] node10466;
	wire [16-1:0] node10469;
	wire [16-1:0] node10472;
	wire [16-1:0] node10473;
	wire [16-1:0] node10475;
	wire [16-1:0] node10479;
	wire [16-1:0] node10481;
	wire [16-1:0] node10482;
	wire [16-1:0] node10484;
	wire [16-1:0] node10488;
	wire [16-1:0] node10489;
	wire [16-1:0] node10490;
	wire [16-1:0] node10491;
	wire [16-1:0] node10492;
	wire [16-1:0] node10493;
	wire [16-1:0] node10494;
	wire [16-1:0] node10495;
	wire [16-1:0] node10496;
	wire [16-1:0] node10497;
	wire [16-1:0] node10501;
	wire [16-1:0] node10502;
	wire [16-1:0] node10506;
	wire [16-1:0] node10507;
	wire [16-1:0] node10510;
	wire [16-1:0] node10511;
	wire [16-1:0] node10515;
	wire [16-1:0] node10516;
	wire [16-1:0] node10517;
	wire [16-1:0] node10518;
	wire [16-1:0] node10521;
	wire [16-1:0] node10523;
	wire [16-1:0] node10524;
	wire [16-1:0] node10528;
	wire [16-1:0] node10529;
	wire [16-1:0] node10530;
	wire [16-1:0] node10535;
	wire [16-1:0] node10536;
	wire [16-1:0] node10537;
	wire [16-1:0] node10539;
	wire [16-1:0] node10540;
	wire [16-1:0] node10544;
	wire [16-1:0] node10547;
	wire [16-1:0] node10548;
	wire [16-1:0] node10549;
	wire [16-1:0] node10553;
	wire [16-1:0] node10555;
	wire [16-1:0] node10558;
	wire [16-1:0] node10559;
	wire [16-1:0] node10560;
	wire [16-1:0] node10561;
	wire [16-1:0] node10562;
	wire [16-1:0] node10566;
	wire [16-1:0] node10567;
	wire [16-1:0] node10570;
	wire [16-1:0] node10573;
	wire [16-1:0] node10574;
	wire [16-1:0] node10575;
	wire [16-1:0] node10576;
	wire [16-1:0] node10580;
	wire [16-1:0] node10581;
	wire [16-1:0] node10583;
	wire [16-1:0] node10587;
	wire [16-1:0] node10588;
	wire [16-1:0] node10589;
	wire [16-1:0] node10591;
	wire [16-1:0] node10595;
	wire [16-1:0] node10598;
	wire [16-1:0] node10599;
	wire [16-1:0] node10600;
	wire [16-1:0] node10601;
	wire [16-1:0] node10605;
	wire [16-1:0] node10606;
	wire [16-1:0] node10609;
	wire [16-1:0] node10612;
	wire [16-1:0] node10613;
	wire [16-1:0] node10615;
	wire [16-1:0] node10618;
	wire [16-1:0] node10619;
	wire [16-1:0] node10620;
	wire [16-1:0] node10622;
	wire [16-1:0] node10626;
	wire [16-1:0] node10628;
	wire [16-1:0] node10631;
	wire [16-1:0] node10632;
	wire [16-1:0] node10633;
	wire [16-1:0] node10634;
	wire [16-1:0] node10635;
	wire [16-1:0] node10636;
	wire [16-1:0] node10637;
	wire [16-1:0] node10638;
	wire [16-1:0] node10643;
	wire [16-1:0] node10646;
	wire [16-1:0] node10647;
	wire [16-1:0] node10650;
	wire [16-1:0] node10653;
	wire [16-1:0] node10654;
	wire [16-1:0] node10655;
	wire [16-1:0] node10658;
	wire [16-1:0] node10660;
	wire [16-1:0] node10663;
	wire [16-1:0] node10665;
	wire [16-1:0] node10668;
	wire [16-1:0] node10669;
	wire [16-1:0] node10670;
	wire [16-1:0] node10673;
	wire [16-1:0] node10675;
	wire [16-1:0] node10678;
	wire [16-1:0] node10679;
	wire [16-1:0] node10681;
	wire [16-1:0] node10684;
	wire [16-1:0] node10685;
	wire [16-1:0] node10688;
	wire [16-1:0] node10690;
	wire [16-1:0] node10693;
	wire [16-1:0] node10694;
	wire [16-1:0] node10695;
	wire [16-1:0] node10696;
	wire [16-1:0] node10698;
	wire [16-1:0] node10700;
	wire [16-1:0] node10703;
	wire [16-1:0] node10704;
	wire [16-1:0] node10706;
	wire [16-1:0] node10710;
	wire [16-1:0] node10711;
	wire [16-1:0] node10714;
	wire [16-1:0] node10715;
	wire [16-1:0] node10717;
	wire [16-1:0] node10720;
	wire [16-1:0] node10723;
	wire [16-1:0] node10724;
	wire [16-1:0] node10725;
	wire [16-1:0] node10726;
	wire [16-1:0] node10729;
	wire [16-1:0] node10730;
	wire [16-1:0] node10734;
	wire [16-1:0] node10736;
	wire [16-1:0] node10739;
	wire [16-1:0] node10740;
	wire [16-1:0] node10742;
	wire [16-1:0] node10744;
	wire [16-1:0] node10747;
	wire [16-1:0] node10748;
	wire [16-1:0] node10751;
	wire [16-1:0] node10754;
	wire [16-1:0] node10755;
	wire [16-1:0] node10756;
	wire [16-1:0] node10757;
	wire [16-1:0] node10758;
	wire [16-1:0] node10759;
	wire [16-1:0] node10760;
	wire [16-1:0] node10762;
	wire [16-1:0] node10763;
	wire [16-1:0] node10767;
	wire [16-1:0] node10770;
	wire [16-1:0] node10771;
	wire [16-1:0] node10772;
	wire [16-1:0] node10776;
	wire [16-1:0] node10779;
	wire [16-1:0] node10780;
	wire [16-1:0] node10781;
	wire [16-1:0] node10784;
	wire [16-1:0] node10786;
	wire [16-1:0] node10787;
	wire [16-1:0] node10791;
	wire [16-1:0] node10792;
	wire [16-1:0] node10794;
	wire [16-1:0] node10795;
	wire [16-1:0] node10799;
	wire [16-1:0] node10801;
	wire [16-1:0] node10804;
	wire [16-1:0] node10805;
	wire [16-1:0] node10806;
	wire [16-1:0] node10808;
	wire [16-1:0] node10811;
	wire [16-1:0] node10812;
	wire [16-1:0] node10815;
	wire [16-1:0] node10817;
	wire [16-1:0] node10820;
	wire [16-1:0] node10821;
	wire [16-1:0] node10822;
	wire [16-1:0] node10823;
	wire [16-1:0] node10825;
	wire [16-1:0] node10829;
	wire [16-1:0] node10832;
	wire [16-1:0] node10833;
	wire [16-1:0] node10837;
	wire [16-1:0] node10838;
	wire [16-1:0] node10839;
	wire [16-1:0] node10840;
	wire [16-1:0] node10842;
	wire [16-1:0] node10843;
	wire [16-1:0] node10847;
	wire [16-1:0] node10848;
	wire [16-1:0] node10851;
	wire [16-1:0] node10853;
	wire [16-1:0] node10856;
	wire [16-1:0] node10858;
	wire [16-1:0] node10859;
	wire [16-1:0] node10860;
	wire [16-1:0] node10865;
	wire [16-1:0] node10866;
	wire [16-1:0] node10867;
	wire [16-1:0] node10868;
	wire [16-1:0] node10871;
	wire [16-1:0] node10872;
	wire [16-1:0] node10874;
	wire [16-1:0] node10878;
	wire [16-1:0] node10879;
	wire [16-1:0] node10880;
	wire [16-1:0] node10885;
	wire [16-1:0] node10888;
	wire [16-1:0] node10889;
	wire [16-1:0] node10890;
	wire [16-1:0] node10891;
	wire [16-1:0] node10892;
	wire [16-1:0] node10893;
	wire [16-1:0] node10896;
	wire [16-1:0] node10897;
	wire [16-1:0] node10899;
	wire [16-1:0] node10903;
	wire [16-1:0] node10904;
	wire [16-1:0] node10907;
	wire [16-1:0] node10910;
	wire [16-1:0] node10911;
	wire [16-1:0] node10912;
	wire [16-1:0] node10915;
	wire [16-1:0] node10917;
	wire [16-1:0] node10920;
	wire [16-1:0] node10921;
	wire [16-1:0] node10925;
	wire [16-1:0] node10926;
	wire [16-1:0] node10927;
	wire [16-1:0] node10928;
	wire [16-1:0] node10930;
	wire [16-1:0] node10931;
	wire [16-1:0] node10935;
	wire [16-1:0] node10938;
	wire [16-1:0] node10939;
	wire [16-1:0] node10941;
	wire [16-1:0] node10942;
	wire [16-1:0] node10945;
	wire [16-1:0] node10948;
	wire [16-1:0] node10950;
	wire [16-1:0] node10953;
	wire [16-1:0] node10954;
	wire [16-1:0] node10955;
	wire [16-1:0] node10958;
	wire [16-1:0] node10960;
	wire [16-1:0] node10963;
	wire [16-1:0] node10964;
	wire [16-1:0] node10968;
	wire [16-1:0] node10969;
	wire [16-1:0] node10970;
	wire [16-1:0] node10971;
	wire [16-1:0] node10972;
	wire [16-1:0] node10974;
	wire [16-1:0] node10977;
	wire [16-1:0] node10980;
	wire [16-1:0] node10981;
	wire [16-1:0] node10984;
	wire [16-1:0] node10987;
	wire [16-1:0] node10988;
	wire [16-1:0] node10989;
	wire [16-1:0] node10992;
	wire [16-1:0] node10994;
	wire [16-1:0] node10997;
	wire [16-1:0] node10998;
	wire [16-1:0] node11002;
	wire [16-1:0] node11003;
	wire [16-1:0] node11004;
	wire [16-1:0] node11006;
	wire [16-1:0] node11008;
	wire [16-1:0] node11011;
	wire [16-1:0] node11012;
	wire [16-1:0] node11014;
	wire [16-1:0] node11017;
	wire [16-1:0] node11020;
	wire [16-1:0] node11021;
	wire [16-1:0] node11023;
	wire [16-1:0] node11026;
	wire [16-1:0] node11027;
	wire [16-1:0] node11028;
	wire [16-1:0] node11030;
	wire [16-1:0] node11034;
	wire [16-1:0] node11037;
	wire [16-1:0] node11038;
	wire [16-1:0] node11039;
	wire [16-1:0] node11040;
	wire [16-1:0] node11041;
	wire [16-1:0] node11042;
	wire [16-1:0] node11043;
	wire [16-1:0] node11044;
	wire [16-1:0] node11045;
	wire [16-1:0] node11046;
	wire [16-1:0] node11051;
	wire [16-1:0] node11054;
	wire [16-1:0] node11055;
	wire [16-1:0] node11059;
	wire [16-1:0] node11060;
	wire [16-1:0] node11061;
	wire [16-1:0] node11064;
	wire [16-1:0] node11066;
	wire [16-1:0] node11069;
	wire [16-1:0] node11070;
	wire [16-1:0] node11074;
	wire [16-1:0] node11075;
	wire [16-1:0] node11076;
	wire [16-1:0] node11077;
	wire [16-1:0] node11080;
	wire [16-1:0] node11083;
	wire [16-1:0] node11084;
	wire [16-1:0] node11088;
	wire [16-1:0] node11090;
	wire [16-1:0] node11091;
	wire [16-1:0] node11094;
	wire [16-1:0] node11096;
	wire [16-1:0] node11099;
	wire [16-1:0] node11100;
	wire [16-1:0] node11101;
	wire [16-1:0] node11104;
	wire [16-1:0] node11105;
	wire [16-1:0] node11106;
	wire [16-1:0] node11109;
	wire [16-1:0] node11110;
	wire [16-1:0] node11114;
	wire [16-1:0] node11115;
	wire [16-1:0] node11119;
	wire [16-1:0] node11120;
	wire [16-1:0] node11121;
	wire [16-1:0] node11122;
	wire [16-1:0] node11124;
	wire [16-1:0] node11125;
	wire [16-1:0] node11130;
	wire [16-1:0] node11131;
	wire [16-1:0] node11134;
	wire [16-1:0] node11135;
	wire [16-1:0] node11137;
	wire [16-1:0] node11141;
	wire [16-1:0] node11142;
	wire [16-1:0] node11144;
	wire [16-1:0] node11147;
	wire [16-1:0] node11149;
	wire [16-1:0] node11151;
	wire [16-1:0] node11154;
	wire [16-1:0] node11155;
	wire [16-1:0] node11156;
	wire [16-1:0] node11157;
	wire [16-1:0] node11158;
	wire [16-1:0] node11160;
	wire [16-1:0] node11161;
	wire [16-1:0] node11164;
	wire [16-1:0] node11167;
	wire [16-1:0] node11169;
	wire [16-1:0] node11171;
	wire [16-1:0] node11172;
	wire [16-1:0] node11176;
	wire [16-1:0] node11177;
	wire [16-1:0] node11179;
	wire [16-1:0] node11183;
	wire [16-1:0] node11184;
	wire [16-1:0] node11185;
	wire [16-1:0] node11186;
	wire [16-1:0] node11189;
	wire [16-1:0] node11192;
	wire [16-1:0] node11193;
	wire [16-1:0] node11194;
	wire [16-1:0] node11196;
	wire [16-1:0] node11200;
	wire [16-1:0] node11201;
	wire [16-1:0] node11203;
	wire [16-1:0] node11207;
	wire [16-1:0] node11208;
	wire [16-1:0] node11209;
	wire [16-1:0] node11212;
	wire [16-1:0] node11215;
	wire [16-1:0] node11216;
	wire [16-1:0] node11219;
	wire [16-1:0] node11222;
	wire [16-1:0] node11223;
	wire [16-1:0] node11224;
	wire [16-1:0] node11225;
	wire [16-1:0] node11227;
	wire [16-1:0] node11229;
	wire [16-1:0] node11230;
	wire [16-1:0] node11235;
	wire [16-1:0] node11236;
	wire [16-1:0] node11237;
	wire [16-1:0] node11240;
	wire [16-1:0] node11242;
	wire [16-1:0] node11245;
	wire [16-1:0] node11246;
	wire [16-1:0] node11249;
	wire [16-1:0] node11252;
	wire [16-1:0] node11253;
	wire [16-1:0] node11254;
	wire [16-1:0] node11256;
	wire [16-1:0] node11258;
	wire [16-1:0] node11259;
	wire [16-1:0] node11263;
	wire [16-1:0] node11264;
	wire [16-1:0] node11267;
	wire [16-1:0] node11270;
	wire [16-1:0] node11271;
	wire [16-1:0] node11272;
	wire [16-1:0] node11275;
	wire [16-1:0] node11277;
	wire [16-1:0] node11278;
	wire [16-1:0] node11283;
	wire [16-1:0] node11284;
	wire [16-1:0] node11285;
	wire [16-1:0] node11286;
	wire [16-1:0] node11287;
	wire [16-1:0] node11288;
	wire [16-1:0] node11290;
	wire [16-1:0] node11293;
	wire [16-1:0] node11295;
	wire [16-1:0] node11298;
	wire [16-1:0] node11299;
	wire [16-1:0] node11300;
	wire [16-1:0] node11304;
	wire [16-1:0] node11305;
	wire [16-1:0] node11308;
	wire [16-1:0] node11310;
	wire [16-1:0] node11313;
	wire [16-1:0] node11314;
	wire [16-1:0] node11315;
	wire [16-1:0] node11317;
	wire [16-1:0] node11320;
	wire [16-1:0] node11321;
	wire [16-1:0] node11324;
	wire [16-1:0] node11326;
	wire [16-1:0] node11329;
	wire [16-1:0] node11330;
	wire [16-1:0] node11331;
	wire [16-1:0] node11334;
	wire [16-1:0] node11337;
	wire [16-1:0] node11338;
	wire [16-1:0] node11340;
	wire [16-1:0] node11344;
	wire [16-1:0] node11345;
	wire [16-1:0] node11346;
	wire [16-1:0] node11347;
	wire [16-1:0] node11348;
	wire [16-1:0] node11349;
	wire [16-1:0] node11353;
	wire [16-1:0] node11356;
	wire [16-1:0] node11357;
	wire [16-1:0] node11360;
	wire [16-1:0] node11362;
	wire [16-1:0] node11365;
	wire [16-1:0] node11366;
	wire [16-1:0] node11367;
	wire [16-1:0] node11370;
	wire [16-1:0] node11371;
	wire [16-1:0] node11376;
	wire [16-1:0] node11377;
	wire [16-1:0] node11378;
	wire [16-1:0] node11380;
	wire [16-1:0] node11383;
	wire [16-1:0] node11384;
	wire [16-1:0] node11385;
	wire [16-1:0] node11389;
	wire [16-1:0] node11390;
	wire [16-1:0] node11392;
	wire [16-1:0] node11396;
	wire [16-1:0] node11397;
	wire [16-1:0] node11398;
	wire [16-1:0] node11401;
	wire [16-1:0] node11403;
	wire [16-1:0] node11406;
	wire [16-1:0] node11407;
	wire [16-1:0] node11410;
	wire [16-1:0] node11413;
	wire [16-1:0] node11414;
	wire [16-1:0] node11415;
	wire [16-1:0] node11416;
	wire [16-1:0] node11417;
	wire [16-1:0] node11419;
	wire [16-1:0] node11421;
	wire [16-1:0] node11422;
	wire [16-1:0] node11426;
	wire [16-1:0] node11429;
	wire [16-1:0] node11430;
	wire [16-1:0] node11431;
	wire [16-1:0] node11436;
	wire [16-1:0] node11437;
	wire [16-1:0] node11438;
	wire [16-1:0] node11440;
	wire [16-1:0] node11441;
	wire [16-1:0] node11444;
	wire [16-1:0] node11447;
	wire [16-1:0] node11448;
	wire [16-1:0] node11449;
	wire [16-1:0] node11453;
	wire [16-1:0] node11454;
	wire [16-1:0] node11456;
	wire [16-1:0] node11460;
	wire [16-1:0] node11461;
	wire [16-1:0] node11464;
	wire [16-1:0] node11466;
	wire [16-1:0] node11469;
	wire [16-1:0] node11470;
	wire [16-1:0] node11471;
	wire [16-1:0] node11472;
	wire [16-1:0] node11475;
	wire [16-1:0] node11476;
	wire [16-1:0] node11479;
	wire [16-1:0] node11481;
	wire [16-1:0] node11484;
	wire [16-1:0] node11485;
	wire [16-1:0] node11486;
	wire [16-1:0] node11489;
	wire [16-1:0] node11492;
	wire [16-1:0] node11493;
	wire [16-1:0] node11494;
	wire [16-1:0] node11499;
	wire [16-1:0] node11500;
	wire [16-1:0] node11501;
	wire [16-1:0] node11503;
	wire [16-1:0] node11506;
	wire [16-1:0] node11507;
	wire [16-1:0] node11510;
	wire [16-1:0] node11513;
	wire [16-1:0] node11514;
	wire [16-1:0] node11516;
	wire [16-1:0] node11519;
	wire [16-1:0] node11520;
	wire [16-1:0] node11523;
	wire [16-1:0] node11526;
	wire [16-1:0] node11527;
	wire [16-1:0] node11528;
	wire [16-1:0] node11529;
	wire [16-1:0] node11530;
	wire [16-1:0] node11531;
	wire [16-1:0] node11532;
	wire [16-1:0] node11533;
	wire [16-1:0] node11534;
	wire [16-1:0] node11538;
	wire [16-1:0] node11539;
	wire [16-1:0] node11543;
	wire [16-1:0] node11544;
	wire [16-1:0] node11547;
	wire [16-1:0] node11550;
	wire [16-1:0] node11551;
	wire [16-1:0] node11552;
	wire [16-1:0] node11555;
	wire [16-1:0] node11556;
	wire [16-1:0] node11560;
	wire [16-1:0] node11561;
	wire [16-1:0] node11562;
	wire [16-1:0] node11564;
	wire [16-1:0] node11567;
	wire [16-1:0] node11570;
	wire [16-1:0] node11571;
	wire [16-1:0] node11573;
	wire [16-1:0] node11577;
	wire [16-1:0] node11578;
	wire [16-1:0] node11579;
	wire [16-1:0] node11580;
	wire [16-1:0] node11582;
	wire [16-1:0] node11585;
	wire [16-1:0] node11586;
	wire [16-1:0] node11590;
	wire [16-1:0] node11591;
	wire [16-1:0] node11592;
	wire [16-1:0] node11593;
	wire [16-1:0] node11595;
	wire [16-1:0] node11598;
	wire [16-1:0] node11601;
	wire [16-1:0] node11603;
	wire [16-1:0] node11606;
	wire [16-1:0] node11607;
	wire [16-1:0] node11609;
	wire [16-1:0] node11610;
	wire [16-1:0] node11614;
	wire [16-1:0] node11617;
	wire [16-1:0] node11618;
	wire [16-1:0] node11620;
	wire [16-1:0] node11623;
	wire [16-1:0] node11624;
	wire [16-1:0] node11625;
	wire [16-1:0] node11628;
	wire [16-1:0] node11631;
	wire [16-1:0] node11633;
	wire [16-1:0] node11636;
	wire [16-1:0] node11637;
	wire [16-1:0] node11638;
	wire [16-1:0] node11639;
	wire [16-1:0] node11640;
	wire [16-1:0] node11641;
	wire [16-1:0] node11642;
	wire [16-1:0] node11643;
	wire [16-1:0] node11649;
	wire [16-1:0] node11651;
	wire [16-1:0] node11654;
	wire [16-1:0] node11655;
	wire [16-1:0] node11656;
	wire [16-1:0] node11657;
	wire [16-1:0] node11661;
	wire [16-1:0] node11663;
	wire [16-1:0] node11664;
	wire [16-1:0] node11668;
	wire [16-1:0] node11669;
	wire [16-1:0] node11670;
	wire [16-1:0] node11672;
	wire [16-1:0] node11676;
	wire [16-1:0] node11679;
	wire [16-1:0] node11680;
	wire [16-1:0] node11681;
	wire [16-1:0] node11682;
	wire [16-1:0] node11685;
	wire [16-1:0] node11687;
	wire [16-1:0] node11688;
	wire [16-1:0] node11692;
	wire [16-1:0] node11693;
	wire [16-1:0] node11694;
	wire [16-1:0] node11698;
	wire [16-1:0] node11700;
	wire [16-1:0] node11703;
	wire [16-1:0] node11704;
	wire [16-1:0] node11705;
	wire [16-1:0] node11706;
	wire [16-1:0] node11708;
	wire [16-1:0] node11713;
	wire [16-1:0] node11714;
	wire [16-1:0] node11715;
	wire [16-1:0] node11719;
	wire [16-1:0] node11722;
	wire [16-1:0] node11723;
	wire [16-1:0] node11724;
	wire [16-1:0] node11726;
	wire [16-1:0] node11727;
	wire [16-1:0] node11730;
	wire [16-1:0] node11733;
	wire [16-1:0] node11734;
	wire [16-1:0] node11735;
	wire [16-1:0] node11736;
	wire [16-1:0] node11740;
	wire [16-1:0] node11742;
	wire [16-1:0] node11745;
	wire [16-1:0] node11746;
	wire [16-1:0] node11748;
	wire [16-1:0] node11749;
	wire [16-1:0] node11753;
	wire [16-1:0] node11756;
	wire [16-1:0] node11757;
	wire [16-1:0] node11758;
	wire [16-1:0] node11759;
	wire [16-1:0] node11761;
	wire [16-1:0] node11764;
	wire [16-1:0] node11767;
	wire [16-1:0] node11770;
	wire [16-1:0] node11771;
	wire [16-1:0] node11773;
	wire [16-1:0] node11776;
	wire [16-1:0] node11778;
	wire [16-1:0] node11781;
	wire [16-1:0] node11782;
	wire [16-1:0] node11783;
	wire [16-1:0] node11784;
	wire [16-1:0] node11785;
	wire [16-1:0] node11788;
	wire [16-1:0] node11789;
	wire [16-1:0] node11791;
	wire [16-1:0] node11794;
	wire [16-1:0] node11795;
	wire [16-1:0] node11799;
	wire [16-1:0] node11800;
	wire [16-1:0] node11801;
	wire [16-1:0] node11802;
	wire [16-1:0] node11803;
	wire [16-1:0] node11806;
	wire [16-1:0] node11810;
	wire [16-1:0] node11811;
	wire [16-1:0] node11812;
	wire [16-1:0] node11816;
	wire [16-1:0] node11819;
	wire [16-1:0] node11820;
	wire [16-1:0] node11823;
	wire [16-1:0] node11825;
	wire [16-1:0] node11828;
	wire [16-1:0] node11829;
	wire [16-1:0] node11830;
	wire [16-1:0] node11831;
	wire [16-1:0] node11833;
	wire [16-1:0] node11836;
	wire [16-1:0] node11837;
	wire [16-1:0] node11838;
	wire [16-1:0] node11842;
	wire [16-1:0] node11845;
	wire [16-1:0] node11846;
	wire [16-1:0] node11847;
	wire [16-1:0] node11849;
	wire [16-1:0] node11851;
	wire [16-1:0] node11854;
	wire [16-1:0] node11856;
	wire [16-1:0] node11859;
	wire [16-1:0] node11860;
	wire [16-1:0] node11861;
	wire [16-1:0] node11863;
	wire [16-1:0] node11866;
	wire [16-1:0] node11867;
	wire [16-1:0] node11871;
	wire [16-1:0] node11874;
	wire [16-1:0] node11875;
	wire [16-1:0] node11877;
	wire [16-1:0] node11878;
	wire [16-1:0] node11881;
	wire [16-1:0] node11884;
	wire [16-1:0] node11885;
	wire [16-1:0] node11886;
	wire [16-1:0] node11890;
	wire [16-1:0] node11893;
	wire [16-1:0] node11894;
	wire [16-1:0] node11895;
	wire [16-1:0] node11896;
	wire [16-1:0] node11898;
	wire [16-1:0] node11899;
	wire [16-1:0] node11900;
	wire [16-1:0] node11905;
	wire [16-1:0] node11906;
	wire [16-1:0] node11907;
	wire [16-1:0] node11909;
	wire [16-1:0] node11912;
	wire [16-1:0] node11914;
	wire [16-1:0] node11917;
	wire [16-1:0] node11918;
	wire [16-1:0] node11922;
	wire [16-1:0] node11923;
	wire [16-1:0] node11924;
	wire [16-1:0] node11925;
	wire [16-1:0] node11929;
	wire [16-1:0] node11930;
	wire [16-1:0] node11932;
	wire [16-1:0] node11933;
	wire [16-1:0] node11937;
	wire [16-1:0] node11940;
	wire [16-1:0] node11941;
	wire [16-1:0] node11942;
	wire [16-1:0] node11945;
	wire [16-1:0] node11948;
	wire [16-1:0] node11949;
	wire [16-1:0] node11952;
	wire [16-1:0] node11955;
	wire [16-1:0] node11956;
	wire [16-1:0] node11957;
	wire [16-1:0] node11959;
	wire [16-1:0] node11962;
	wire [16-1:0] node11963;
	wire [16-1:0] node11965;
	wire [16-1:0] node11967;
	wire [16-1:0] node11970;
	wire [16-1:0] node11971;
	wire [16-1:0] node11974;
	wire [16-1:0] node11976;
	wire [16-1:0] node11979;
	wire [16-1:0] node11980;
	wire [16-1:0] node11982;
	wire [16-1:0] node11983;
	wire [16-1:0] node11985;
	wire [16-1:0] node11988;
	wire [16-1:0] node11989;
	wire [16-1:0] node11991;
	wire [16-1:0] node11995;
	wire [16-1:0] node11996;
	wire [16-1:0] node11998;
	wire [16-1:0] node12000;
	wire [16-1:0] node12001;
	wire [16-1:0] node12005;
	wire [16-1:0] node12006;
	wire [16-1:0] node12008;
	wire [16-1:0] node12009;
	wire [16-1:0] node12013;
	wire [16-1:0] node12016;
	wire [16-1:0] node12017;
	wire [16-1:0] node12018;
	wire [16-1:0] node12019;
	wire [16-1:0] node12020;
	wire [16-1:0] node12021;
	wire [16-1:0] node12022;
	wire [16-1:0] node12023;
	wire [16-1:0] node12024;
	wire [16-1:0] node12029;
	wire [16-1:0] node12030;
	wire [16-1:0] node12031;
	wire [16-1:0] node12035;
	wire [16-1:0] node12038;
	wire [16-1:0] node12039;
	wire [16-1:0] node12042;
	wire [16-1:0] node12044;
	wire [16-1:0] node12047;
	wire [16-1:0] node12048;
	wire [16-1:0] node12049;
	wire [16-1:0] node12051;
	wire [16-1:0] node12055;
	wire [16-1:0] node12056;
	wire [16-1:0] node12057;
	wire [16-1:0] node12061;
	wire [16-1:0] node12064;
	wire [16-1:0] node12065;
	wire [16-1:0] node12066;
	wire [16-1:0] node12068;
	wire [16-1:0] node12069;
	wire [16-1:0] node12071;
	wire [16-1:0] node12074;
	wire [16-1:0] node12077;
	wire [16-1:0] node12078;
	wire [16-1:0] node12080;
	wire [16-1:0] node12081;
	wire [16-1:0] node12085;
	wire [16-1:0] node12086;
	wire [16-1:0] node12089;
	wire [16-1:0] node12092;
	wire [16-1:0] node12093;
	wire [16-1:0] node12094;
	wire [16-1:0] node12095;
	wire [16-1:0] node12097;
	wire [16-1:0] node12100;
	wire [16-1:0] node12102;
	wire [16-1:0] node12103;
	wire [16-1:0] node12107;
	wire [16-1:0] node12108;
	wire [16-1:0] node12111;
	wire [16-1:0] node12112;
	wire [16-1:0] node12116;
	wire [16-1:0] node12117;
	wire [16-1:0] node12119;
	wire [16-1:0] node12120;
	wire [16-1:0] node12122;
	wire [16-1:0] node12126;
	wire [16-1:0] node12127;
	wire [16-1:0] node12131;
	wire [16-1:0] node12132;
	wire [16-1:0] node12133;
	wire [16-1:0] node12134;
	wire [16-1:0] node12136;
	wire [16-1:0] node12138;
	wire [16-1:0] node12141;
	wire [16-1:0] node12142;
	wire [16-1:0] node12144;
	wire [16-1:0] node12147;
	wire [16-1:0] node12149;
	wire [16-1:0] node12152;
	wire [16-1:0] node12153;
	wire [16-1:0] node12154;
	wire [16-1:0] node12155;
	wire [16-1:0] node12158;
	wire [16-1:0] node12161;
	wire [16-1:0] node12162;
	wire [16-1:0] node12165;
	wire [16-1:0] node12168;
	wire [16-1:0] node12169;
	wire [16-1:0] node12171;
	wire [16-1:0] node12172;
	wire [16-1:0] node12176;
	wire [16-1:0] node12178;
	wire [16-1:0] node12181;
	wire [16-1:0] node12182;
	wire [16-1:0] node12183;
	wire [16-1:0] node12184;
	wire [16-1:0] node12186;
	wire [16-1:0] node12189;
	wire [16-1:0] node12191;
	wire [16-1:0] node12193;
	wire [16-1:0] node12196;
	wire [16-1:0] node12197;
	wire [16-1:0] node12198;
	wire [16-1:0] node12200;
	wire [16-1:0] node12201;
	wire [16-1:0] node12205;
	wire [16-1:0] node12207;
	wire [16-1:0] node12208;
	wire [16-1:0] node12212;
	wire [16-1:0] node12213;
	wire [16-1:0] node12214;
	wire [16-1:0] node12216;
	wire [16-1:0] node12221;
	wire [16-1:0] node12222;
	wire [16-1:0] node12223;
	wire [16-1:0] node12225;
	wire [16-1:0] node12228;
	wire [16-1:0] node12230;
	wire [16-1:0] node12231;
	wire [16-1:0] node12235;
	wire [16-1:0] node12236;
	wire [16-1:0] node12239;
	wire [16-1:0] node12241;
	wire [16-1:0] node12243;
	wire [16-1:0] node12245;
	wire [16-1:0] node12248;
	wire [16-1:0] node12249;
	wire [16-1:0] node12250;
	wire [16-1:0] node12251;
	wire [16-1:0] node12252;
	wire [16-1:0] node12253;
	wire [16-1:0] node12254;
	wire [16-1:0] node12258;
	wire [16-1:0] node12259;
	wire [16-1:0] node12263;
	wire [16-1:0] node12265;
	wire [16-1:0] node12268;
	wire [16-1:0] node12269;
	wire [16-1:0] node12270;
	wire [16-1:0] node12271;
	wire [16-1:0] node12275;
	wire [16-1:0] node12276;
	wire [16-1:0] node12280;
	wire [16-1:0] node12281;
	wire [16-1:0] node12283;
	wire [16-1:0] node12286;
	wire [16-1:0] node12287;
	wire [16-1:0] node12291;
	wire [16-1:0] node12292;
	wire [16-1:0] node12293;
	wire [16-1:0] node12294;
	wire [16-1:0] node12295;
	wire [16-1:0] node12296;
	wire [16-1:0] node12297;
	wire [16-1:0] node12302;
	wire [16-1:0] node12305;
	wire [16-1:0] node12307;
	wire [16-1:0] node12309;
	wire [16-1:0] node12312;
	wire [16-1:0] node12313;
	wire [16-1:0] node12314;
	wire [16-1:0] node12317;
	wire [16-1:0] node12320;
	wire [16-1:0] node12322;
	wire [16-1:0] node12325;
	wire [16-1:0] node12326;
	wire [16-1:0] node12327;
	wire [16-1:0] node12328;
	wire [16-1:0] node12329;
	wire [16-1:0] node12332;
	wire [16-1:0] node12334;
	wire [16-1:0] node12338;
	wire [16-1:0] node12339;
	wire [16-1:0] node12342;
	wire [16-1:0] node12344;
	wire [16-1:0] node12347;
	wire [16-1:0] node12348;
	wire [16-1:0] node12349;
	wire [16-1:0] node12352;
	wire [16-1:0] node12354;
	wire [16-1:0] node12357;
	wire [16-1:0] node12358;
	wire [16-1:0] node12362;
	wire [16-1:0] node12363;
	wire [16-1:0] node12364;
	wire [16-1:0] node12365;
	wire [16-1:0] node12366;
	wire [16-1:0] node12367;
	wire [16-1:0] node12368;
	wire [16-1:0] node12372;
	wire [16-1:0] node12376;
	wire [16-1:0] node12377;
	wire [16-1:0] node12379;
	wire [16-1:0] node12382;
	wire [16-1:0] node12383;
	wire [16-1:0] node12386;
	wire [16-1:0] node12389;
	wire [16-1:0] node12390;
	wire [16-1:0] node12391;
	wire [16-1:0] node12394;
	wire [16-1:0] node12395;
	wire [16-1:0] node12399;
	wire [16-1:0] node12400;
	wire [16-1:0] node12401;
	wire [16-1:0] node12404;
	wire [16-1:0] node12407;
	wire [16-1:0] node12408;
	wire [16-1:0] node12411;
	wire [16-1:0] node12412;
	wire [16-1:0] node12414;
	wire [16-1:0] node12418;
	wire [16-1:0] node12419;
	wire [16-1:0] node12420;
	wire [16-1:0] node12422;
	wire [16-1:0] node12424;
	wire [16-1:0] node12425;
	wire [16-1:0] node12426;
	wire [16-1:0] node12431;
	wire [16-1:0] node12432;
	wire [16-1:0] node12433;
	wire [16-1:0] node12434;
	wire [16-1:0] node12436;
	wire [16-1:0] node12439;
	wire [16-1:0] node12441;
	wire [16-1:0] node12445;
	wire [16-1:0] node12446;
	wire [16-1:0] node12449;
	wire [16-1:0] node12452;
	wire [16-1:0] node12453;
	wire [16-1:0] node12454;
	wire [16-1:0] node12456;
	wire [16-1:0] node12459;
	wire [16-1:0] node12460;
	wire [16-1:0] node12463;
	wire [16-1:0] node12464;
	wire [16-1:0] node12466;
	wire [16-1:0] node12470;
	wire [16-1:0] node12471;
	wire [16-1:0] node12473;
	wire [16-1:0] node12475;
	wire [16-1:0] node12476;
	wire [16-1:0] node12480;
	wire [16-1:0] node12481;
	wire [16-1:0] node12484;
	wire [16-1:0] node12486;
	wire [16-1:0] node12489;
	wire [16-1:0] node12490;
	wire [16-1:0] node12491;
	wire [16-1:0] node12492;
	wire [16-1:0] node12493;
	wire [16-1:0] node12494;
	wire [16-1:0] node12495;
	wire [16-1:0] node12496;
	wire [16-1:0] node12497;
	wire [16-1:0] node12498;
	wire [16-1:0] node12499;
	wire [16-1:0] node12501;
	wire [16-1:0] node12502;
	wire [16-1:0] node12506;
	wire [16-1:0] node12508;
	wire [16-1:0] node12511;
	wire [16-1:0] node12512;
	wire [16-1:0] node12514;
	wire [16-1:0] node12518;
	wire [16-1:0] node12519;
	wire [16-1:0] node12520;
	wire [16-1:0] node12521;
	wire [16-1:0] node12522;
	wire [16-1:0] node12527;
	wire [16-1:0] node12529;
	wire [16-1:0] node12532;
	wire [16-1:0] node12533;
	wire [16-1:0] node12534;
	wire [16-1:0] node12539;
	wire [16-1:0] node12540;
	wire [16-1:0] node12541;
	wire [16-1:0] node12543;
	wire [16-1:0] node12544;
	wire [16-1:0] node12545;
	wire [16-1:0] node12550;
	wire [16-1:0] node12552;
	wire [16-1:0] node12555;
	wire [16-1:0] node12556;
	wire [16-1:0] node12557;
	wire [16-1:0] node12560;
	wire [16-1:0] node12563;
	wire [16-1:0] node12565;
	wire [16-1:0] node12568;
	wire [16-1:0] node12569;
	wire [16-1:0] node12570;
	wire [16-1:0] node12571;
	wire [16-1:0] node12573;
	wire [16-1:0] node12576;
	wire [16-1:0] node12579;
	wire [16-1:0] node12580;
	wire [16-1:0] node12581;
	wire [16-1:0] node12582;
	wire [16-1:0] node12587;
	wire [16-1:0] node12590;
	wire [16-1:0] node12591;
	wire [16-1:0] node12592;
	wire [16-1:0] node12595;
	wire [16-1:0] node12596;
	wire [16-1:0] node12598;
	wire [16-1:0] node12602;
	wire [16-1:0] node12603;
	wire [16-1:0] node12604;
	wire [16-1:0] node12605;
	wire [16-1:0] node12609;
	wire [16-1:0] node12612;
	wire [16-1:0] node12614;
	wire [16-1:0] node12617;
	wire [16-1:0] node12618;
	wire [16-1:0] node12619;
	wire [16-1:0] node12620;
	wire [16-1:0] node12621;
	wire [16-1:0] node12622;
	wire [16-1:0] node12625;
	wire [16-1:0] node12628;
	wire [16-1:0] node12629;
	wire [16-1:0] node12630;
	wire [16-1:0] node12632;
	wire [16-1:0] node12637;
	wire [16-1:0] node12638;
	wire [16-1:0] node12641;
	wire [16-1:0] node12642;
	wire [16-1:0] node12643;
	wire [16-1:0] node12648;
	wire [16-1:0] node12649;
	wire [16-1:0] node12650;
	wire [16-1:0] node12652;
	wire [16-1:0] node12655;
	wire [16-1:0] node12656;
	wire [16-1:0] node12660;
	wire [16-1:0] node12662;
	wire [16-1:0] node12663;
	wire [16-1:0] node12664;
	wire [16-1:0] node12665;
	wire [16-1:0] node12669;
	wire [16-1:0] node12670;
	wire [16-1:0] node12675;
	wire [16-1:0] node12676;
	wire [16-1:0] node12677;
	wire [16-1:0] node12678;
	wire [16-1:0] node12679;
	wire [16-1:0] node12683;
	wire [16-1:0] node12685;
	wire [16-1:0] node12688;
	wire [16-1:0] node12689;
	wire [16-1:0] node12690;
	wire [16-1:0] node12694;
	wire [16-1:0] node12696;
	wire [16-1:0] node12699;
	wire [16-1:0] node12700;
	wire [16-1:0] node12701;
	wire [16-1:0] node12702;
	wire [16-1:0] node12706;
	wire [16-1:0] node12707;
	wire [16-1:0] node12710;
	wire [16-1:0] node12711;
	wire [16-1:0] node12712;
	wire [16-1:0] node12716;
	wire [16-1:0] node12719;
	wire [16-1:0] node12720;
	wire [16-1:0] node12721;
	wire [16-1:0] node12723;
	wire [16-1:0] node12726;
	wire [16-1:0] node12728;
	wire [16-1:0] node12731;
	wire [16-1:0] node12732;
	wire [16-1:0] node12736;
	wire [16-1:0] node12737;
	wire [16-1:0] node12738;
	wire [16-1:0] node12739;
	wire [16-1:0] node12740;
	wire [16-1:0] node12741;
	wire [16-1:0] node12742;
	wire [16-1:0] node12746;
	wire [16-1:0] node12747;
	wire [16-1:0] node12748;
	wire [16-1:0] node12749;
	wire [16-1:0] node12755;
	wire [16-1:0] node12756;
	wire [16-1:0] node12757;
	wire [16-1:0] node12759;
	wire [16-1:0] node12761;
	wire [16-1:0] node12764;
	wire [16-1:0] node12767;
	wire [16-1:0] node12770;
	wire [16-1:0] node12771;
	wire [16-1:0] node12772;
	wire [16-1:0] node12774;
	wire [16-1:0] node12777;
	wire [16-1:0] node12778;
	wire [16-1:0] node12782;
	wire [16-1:0] node12783;
	wire [16-1:0] node12784;
	wire [16-1:0] node12787;
	wire [16-1:0] node12790;
	wire [16-1:0] node12791;
	wire [16-1:0] node12794;
	wire [16-1:0] node12795;
	wire [16-1:0] node12797;
	wire [16-1:0] node12801;
	wire [16-1:0] node12802;
	wire [16-1:0] node12803;
	wire [16-1:0] node12804;
	wire [16-1:0] node12805;
	wire [16-1:0] node12808;
	wire [16-1:0] node12812;
	wire [16-1:0] node12813;
	wire [16-1:0] node12814;
	wire [16-1:0] node12818;
	wire [16-1:0] node12819;
	wire [16-1:0] node12820;
	wire [16-1:0] node12824;
	wire [16-1:0] node12827;
	wire [16-1:0] node12828;
	wire [16-1:0] node12829;
	wire [16-1:0] node12831;
	wire [16-1:0] node12832;
	wire [16-1:0] node12836;
	wire [16-1:0] node12837;
	wire [16-1:0] node12840;
	wire [16-1:0] node12843;
	wire [16-1:0] node12844;
	wire [16-1:0] node12845;
	wire [16-1:0] node12847;
	wire [16-1:0] node12850;
	wire [16-1:0] node12853;
	wire [16-1:0] node12854;
	wire [16-1:0] node12855;
	wire [16-1:0] node12857;
	wire [16-1:0] node12861;
	wire [16-1:0] node12864;
	wire [16-1:0] node12865;
	wire [16-1:0] node12866;
	wire [16-1:0] node12867;
	wire [16-1:0] node12868;
	wire [16-1:0] node12870;
	wire [16-1:0] node12873;
	wire [16-1:0] node12874;
	wire [16-1:0] node12875;
	wire [16-1:0] node12877;
	wire [16-1:0] node12880;
	wire [16-1:0] node12883;
	wire [16-1:0] node12885;
	wire [16-1:0] node12888;
	wire [16-1:0] node12889;
	wire [16-1:0] node12891;
	wire [16-1:0] node12894;
	wire [16-1:0] node12895;
	wire [16-1:0] node12898;
	wire [16-1:0] node12899;
	wire [16-1:0] node12903;
	wire [16-1:0] node12904;
	wire [16-1:0] node12905;
	wire [16-1:0] node12906;
	wire [16-1:0] node12910;
	wire [16-1:0] node12911;
	wire [16-1:0] node12914;
	wire [16-1:0] node12915;
	wire [16-1:0] node12919;
	wire [16-1:0] node12921;
	wire [16-1:0] node12922;
	wire [16-1:0] node12925;
	wire [16-1:0] node12927;
	wire [16-1:0] node12928;
	wire [16-1:0] node12932;
	wire [16-1:0] node12933;
	wire [16-1:0] node12934;
	wire [16-1:0] node12936;
	wire [16-1:0] node12937;
	wire [16-1:0] node12938;
	wire [16-1:0] node12943;
	wire [16-1:0] node12944;
	wire [16-1:0] node12945;
	wire [16-1:0] node12948;
	wire [16-1:0] node12951;
	wire [16-1:0] node12952;
	wire [16-1:0] node12955;
	wire [16-1:0] node12958;
	wire [16-1:0] node12959;
	wire [16-1:0] node12960;
	wire [16-1:0] node12961;
	wire [16-1:0] node12965;
	wire [16-1:0] node12967;
	wire [16-1:0] node12970;
	wire [16-1:0] node12971;
	wire [16-1:0] node12972;
	wire [16-1:0] node12974;
	wire [16-1:0] node12978;
	wire [16-1:0] node12979;
	wire [16-1:0] node12983;
	wire [16-1:0] node12984;
	wire [16-1:0] node12985;
	wire [16-1:0] node12986;
	wire [16-1:0] node12987;
	wire [16-1:0] node12988;
	wire [16-1:0] node12989;
	wire [16-1:0] node12991;
	wire [16-1:0] node12992;
	wire [16-1:0] node12996;
	wire [16-1:0] node12998;
	wire [16-1:0] node12999;
	wire [16-1:0] node13003;
	wire [16-1:0] node13004;
	wire [16-1:0] node13005;
	wire [16-1:0] node13006;
	wire [16-1:0] node13010;
	wire [16-1:0] node13012;
	wire [16-1:0] node13016;
	wire [16-1:0] node13017;
	wire [16-1:0] node13018;
	wire [16-1:0] node13021;
	wire [16-1:0] node13023;
	wire [16-1:0] node13026;
	wire [16-1:0] node13027;
	wire [16-1:0] node13028;
	wire [16-1:0] node13031;
	wire [16-1:0] node13034;
	wire [16-1:0] node13035;
	wire [16-1:0] node13039;
	wire [16-1:0] node13040;
	wire [16-1:0] node13041;
	wire [16-1:0] node13042;
	wire [16-1:0] node13044;
	wire [16-1:0] node13047;
	wire [16-1:0] node13048;
	wire [16-1:0] node13050;
	wire [16-1:0] node13051;
	wire [16-1:0] node13055;
	wire [16-1:0] node13058;
	wire [16-1:0] node13059;
	wire [16-1:0] node13060;
	wire [16-1:0] node13061;
	wire [16-1:0] node13065;
	wire [16-1:0] node13066;
	wire [16-1:0] node13070;
	wire [16-1:0] node13073;
	wire [16-1:0] node13074;
	wire [16-1:0] node13076;
	wire [16-1:0] node13077;
	wire [16-1:0] node13078;
	wire [16-1:0] node13080;
	wire [16-1:0] node13085;
	wire [16-1:0] node13086;
	wire [16-1:0] node13088;
	wire [16-1:0] node13091;
	wire [16-1:0] node13092;
	wire [16-1:0] node13095;
	wire [16-1:0] node13096;
	wire [16-1:0] node13100;
	wire [16-1:0] node13101;
	wire [16-1:0] node13102;
	wire [16-1:0] node13103;
	wire [16-1:0] node13104;
	wire [16-1:0] node13106;
	wire [16-1:0] node13108;
	wire [16-1:0] node13111;
	wire [16-1:0] node13112;
	wire [16-1:0] node13113;
	wire [16-1:0] node13114;
	wire [16-1:0] node13120;
	wire [16-1:0] node13121;
	wire [16-1:0] node13124;
	wire [16-1:0] node13127;
	wire [16-1:0] node13128;
	wire [16-1:0] node13129;
	wire [16-1:0] node13132;
	wire [16-1:0] node13134;
	wire [16-1:0] node13136;
	wire [16-1:0] node13137;
	wire [16-1:0] node13141;
	wire [16-1:0] node13142;
	wire [16-1:0] node13143;
	wire [16-1:0] node13146;
	wire [16-1:0] node13147;
	wire [16-1:0] node13152;
	wire [16-1:0] node13153;
	wire [16-1:0] node13154;
	wire [16-1:0] node13155;
	wire [16-1:0] node13156;
	wire [16-1:0] node13159;
	wire [16-1:0] node13160;
	wire [16-1:0] node13162;
	wire [16-1:0] node13165;
	wire [16-1:0] node13169;
	wire [16-1:0] node13170;
	wire [16-1:0] node13173;
	wire [16-1:0] node13175;
	wire [16-1:0] node13178;
	wire [16-1:0] node13179;
	wire [16-1:0] node13180;
	wire [16-1:0] node13181;
	wire [16-1:0] node13183;
	wire [16-1:0] node13184;
	wire [16-1:0] node13189;
	wire [16-1:0] node13190;
	wire [16-1:0] node13191;
	wire [16-1:0] node13196;
	wire [16-1:0] node13197;
	wire [16-1:0] node13199;
	wire [16-1:0] node13200;
	wire [16-1:0] node13202;
	wire [16-1:0] node13206;
	wire [16-1:0] node13208;
	wire [16-1:0] node13211;
	wire [16-1:0] node13212;
	wire [16-1:0] node13213;
	wire [16-1:0] node13214;
	wire [16-1:0] node13215;
	wire [16-1:0] node13216;
	wire [16-1:0] node13217;
	wire [16-1:0] node13220;
	wire [16-1:0] node13221;
	wire [16-1:0] node13222;
	wire [16-1:0] node13227;
	wire [16-1:0] node13228;
	wire [16-1:0] node13231;
	wire [16-1:0] node13234;
	wire [16-1:0] node13235;
	wire [16-1:0] node13236;
	wire [16-1:0] node13239;
	wire [16-1:0] node13241;
	wire [16-1:0] node13244;
	wire [16-1:0] node13245;
	wire [16-1:0] node13249;
	wire [16-1:0] node13250;
	wire [16-1:0] node13251;
	wire [16-1:0] node13252;
	wire [16-1:0] node13256;
	wire [16-1:0] node13257;
	wire [16-1:0] node13260;
	wire [16-1:0] node13263;
	wire [16-1:0] node13265;
	wire [16-1:0] node13266;
	wire [16-1:0] node13269;
	wire [16-1:0] node13271;
	wire [16-1:0] node13272;
	wire [16-1:0] node13276;
	wire [16-1:0] node13277;
	wire [16-1:0] node13278;
	wire [16-1:0] node13279;
	wire [16-1:0] node13280;
	wire [16-1:0] node13284;
	wire [16-1:0] node13285;
	wire [16-1:0] node13288;
	wire [16-1:0] node13290;
	wire [16-1:0] node13293;
	wire [16-1:0] node13294;
	wire [16-1:0] node13295;
	wire [16-1:0] node13298;
	wire [16-1:0] node13301;
	wire [16-1:0] node13303;
	wire [16-1:0] node13306;
	wire [16-1:0] node13307;
	wire [16-1:0] node13308;
	wire [16-1:0] node13309;
	wire [16-1:0] node13310;
	wire [16-1:0] node13314;
	wire [16-1:0] node13315;
	wire [16-1:0] node13317;
	wire [16-1:0] node13320;
	wire [16-1:0] node13322;
	wire [16-1:0] node13325;
	wire [16-1:0] node13327;
	wire [16-1:0] node13330;
	wire [16-1:0] node13331;
	wire [16-1:0] node13332;
	wire [16-1:0] node13335;
	wire [16-1:0] node13338;
	wire [16-1:0] node13339;
	wire [16-1:0] node13342;
	wire [16-1:0] node13344;
	wire [16-1:0] node13347;
	wire [16-1:0] node13348;
	wire [16-1:0] node13349;
	wire [16-1:0] node13350;
	wire [16-1:0] node13351;
	wire [16-1:0] node13353;
	wire [16-1:0] node13356;
	wire [16-1:0] node13357;
	wire [16-1:0] node13358;
	wire [16-1:0] node13362;
	wire [16-1:0] node13364;
	wire [16-1:0] node13367;
	wire [16-1:0] node13368;
	wire [16-1:0] node13369;
	wire [16-1:0] node13372;
	wire [16-1:0] node13375;
	wire [16-1:0] node13377;
	wire [16-1:0] node13379;
	wire [16-1:0] node13381;
	wire [16-1:0] node13384;
	wire [16-1:0] node13385;
	wire [16-1:0] node13386;
	wire [16-1:0] node13388;
	wire [16-1:0] node13391;
	wire [16-1:0] node13392;
	wire [16-1:0] node13395;
	wire [16-1:0] node13397;
	wire [16-1:0] node13400;
	wire [16-1:0] node13401;
	wire [16-1:0] node13403;
	wire [16-1:0] node13406;
	wire [16-1:0] node13407;
	wire [16-1:0] node13409;
	wire [16-1:0] node13411;
	wire [16-1:0] node13415;
	wire [16-1:0] node13416;
	wire [16-1:0] node13417;
	wire [16-1:0] node13418;
	wire [16-1:0] node13419;
	wire [16-1:0] node13422;
	wire [16-1:0] node13425;
	wire [16-1:0] node13426;
	wire [16-1:0] node13429;
	wire [16-1:0] node13431;
	wire [16-1:0] node13432;
	wire [16-1:0] node13436;
	wire [16-1:0] node13437;
	wire [16-1:0] node13438;
	wire [16-1:0] node13439;
	wire [16-1:0] node13443;
	wire [16-1:0] node13445;
	wire [16-1:0] node13447;
	wire [16-1:0] node13450;
	wire [16-1:0] node13452;
	wire [16-1:0] node13454;
	wire [16-1:0] node13457;
	wire [16-1:0] node13458;
	wire [16-1:0] node13459;
	wire [16-1:0] node13462;
	wire [16-1:0] node13463;
	wire [16-1:0] node13464;
	wire [16-1:0] node13467;
	wire [16-1:0] node13469;
	wire [16-1:0] node13472;
	wire [16-1:0] node13473;
	wire [16-1:0] node13477;
	wire [16-1:0] node13478;
	wire [16-1:0] node13480;
	wire [16-1:0] node13481;
	wire [16-1:0] node13486;
	wire [16-1:0] node13487;
	wire [16-1:0] node13488;
	wire [16-1:0] node13489;
	wire [16-1:0] node13490;
	wire [16-1:0] node13491;
	wire [16-1:0] node13492;
	wire [16-1:0] node13493;
	wire [16-1:0] node13494;
	wire [16-1:0] node13498;
	wire [16-1:0] node13499;
	wire [16-1:0] node13501;
	wire [16-1:0] node13504;
	wire [16-1:0] node13507;
	wire [16-1:0] node13508;
	wire [16-1:0] node13509;
	wire [16-1:0] node13513;
	wire [16-1:0] node13514;
	wire [16-1:0] node13516;
	wire [16-1:0] node13517;
	wire [16-1:0] node13522;
	wire [16-1:0] node13523;
	wire [16-1:0] node13524;
	wire [16-1:0] node13525;
	wire [16-1:0] node13526;
	wire [16-1:0] node13528;
	wire [16-1:0] node13532;
	wire [16-1:0] node13535;
	wire [16-1:0] node13536;
	wire [16-1:0] node13539;
	wire [16-1:0] node13542;
	wire [16-1:0] node13543;
	wire [16-1:0] node13544;
	wire [16-1:0] node13547;
	wire [16-1:0] node13548;
	wire [16-1:0] node13550;
	wire [16-1:0] node13554;
	wire [16-1:0] node13555;
	wire [16-1:0] node13556;
	wire [16-1:0] node13558;
	wire [16-1:0] node13562;
	wire [16-1:0] node13565;
	wire [16-1:0] node13566;
	wire [16-1:0] node13567;
	wire [16-1:0] node13568;
	wire [16-1:0] node13570;
	wire [16-1:0] node13573;
	wire [16-1:0] node13574;
	wire [16-1:0] node13575;
	wire [16-1:0] node13579;
	wire [16-1:0] node13582;
	wire [16-1:0] node13583;
	wire [16-1:0] node13586;
	wire [16-1:0] node13588;
	wire [16-1:0] node13589;
	wire [16-1:0] node13590;
	wire [16-1:0] node13595;
	wire [16-1:0] node13596;
	wire [16-1:0] node13597;
	wire [16-1:0] node13598;
	wire [16-1:0] node13599;
	wire [16-1:0] node13603;
	wire [16-1:0] node13606;
	wire [16-1:0] node13607;
	wire [16-1:0] node13610;
	wire [16-1:0] node13613;
	wire [16-1:0] node13614;
	wire [16-1:0] node13618;
	wire [16-1:0] node13619;
	wire [16-1:0] node13620;
	wire [16-1:0] node13621;
	wire [16-1:0] node13622;
	wire [16-1:0] node13624;
	wire [16-1:0] node13627;
	wire [16-1:0] node13628;
	wire [16-1:0] node13632;
	wire [16-1:0] node13633;
	wire [16-1:0] node13634;
	wire [16-1:0] node13636;
	wire [16-1:0] node13640;
	wire [16-1:0] node13643;
	wire [16-1:0] node13644;
	wire [16-1:0] node13646;
	wire [16-1:0] node13648;
	wire [16-1:0] node13651;
	wire [16-1:0] node13652;
	wire [16-1:0] node13654;
	wire [16-1:0] node13657;
	wire [16-1:0] node13658;
	wire [16-1:0] node13660;
	wire [16-1:0] node13661;
	wire [16-1:0] node13665;
	wire [16-1:0] node13668;
	wire [16-1:0] node13669;
	wire [16-1:0] node13670;
	wire [16-1:0] node13671;
	wire [16-1:0] node13674;
	wire [16-1:0] node13675;
	wire [16-1:0] node13679;
	wire [16-1:0] node13680;
	wire [16-1:0] node13681;
	wire [16-1:0] node13684;
	wire [16-1:0] node13686;
	wire [16-1:0] node13689;
	wire [16-1:0] node13690;
	wire [16-1:0] node13694;
	wire [16-1:0] node13695;
	wire [16-1:0] node13696;
	wire [16-1:0] node13698;
	wire [16-1:0] node13701;
	wire [16-1:0] node13704;
	wire [16-1:0] node13705;
	wire [16-1:0] node13707;
	wire [16-1:0] node13709;
	wire [16-1:0] node13710;
	wire [16-1:0] node13714;
	wire [16-1:0] node13717;
	wire [16-1:0] node13718;
	wire [16-1:0] node13719;
	wire [16-1:0] node13720;
	wire [16-1:0] node13721;
	wire [16-1:0] node13722;
	wire [16-1:0] node13723;
	wire [16-1:0] node13725;
	wire [16-1:0] node13726;
	wire [16-1:0] node13730;
	wire [16-1:0] node13733;
	wire [16-1:0] node13734;
	wire [16-1:0] node13735;
	wire [16-1:0] node13737;
	wire [16-1:0] node13742;
	wire [16-1:0] node13743;
	wire [16-1:0] node13745;
	wire [16-1:0] node13747;
	wire [16-1:0] node13750;
	wire [16-1:0] node13753;
	wire [16-1:0] node13754;
	wire [16-1:0] node13755;
	wire [16-1:0] node13757;
	wire [16-1:0] node13758;
	wire [16-1:0] node13762;
	wire [16-1:0] node13763;
	wire [16-1:0] node13767;
	wire [16-1:0] node13768;
	wire [16-1:0] node13769;
	wire [16-1:0] node13772;
	wire [16-1:0] node13773;
	wire [16-1:0] node13774;
	wire [16-1:0] node13778;
	wire [16-1:0] node13781;
	wire [16-1:0] node13782;
	wire [16-1:0] node13785;
	wire [16-1:0] node13788;
	wire [16-1:0] node13789;
	wire [16-1:0] node13790;
	wire [16-1:0] node13791;
	wire [16-1:0] node13792;
	wire [16-1:0] node13795;
	wire [16-1:0] node13799;
	wire [16-1:0] node13800;
	wire [16-1:0] node13801;
	wire [16-1:0] node13804;
	wire [16-1:0] node13805;
	wire [16-1:0] node13809;
	wire [16-1:0] node13810;
	wire [16-1:0] node13813;
	wire [16-1:0] node13816;
	wire [16-1:0] node13817;
	wire [16-1:0] node13818;
	wire [16-1:0] node13820;
	wire [16-1:0] node13823;
	wire [16-1:0] node13824;
	wire [16-1:0] node13828;
	wire [16-1:0] node13829;
	wire [16-1:0] node13830;
	wire [16-1:0] node13834;
	wire [16-1:0] node13836;
	wire [16-1:0] node13839;
	wire [16-1:0] node13840;
	wire [16-1:0] node13841;
	wire [16-1:0] node13842;
	wire [16-1:0] node13843;
	wire [16-1:0] node13844;
	wire [16-1:0] node13845;
	wire [16-1:0] node13848;
	wire [16-1:0] node13852;
	wire [16-1:0] node13854;
	wire [16-1:0] node13855;
	wire [16-1:0] node13859;
	wire [16-1:0] node13860;
	wire [16-1:0] node13861;
	wire [16-1:0] node13863;
	wire [16-1:0] node13866;
	wire [16-1:0] node13868;
	wire [16-1:0] node13871;
	wire [16-1:0] node13872;
	wire [16-1:0] node13873;
	wire [16-1:0] node13875;
	wire [16-1:0] node13878;
	wire [16-1:0] node13879;
	wire [16-1:0] node13883;
	wire [16-1:0] node13886;
	wire [16-1:0] node13887;
	wire [16-1:0] node13888;
	wire [16-1:0] node13889;
	wire [16-1:0] node13891;
	wire [16-1:0] node13895;
	wire [16-1:0] node13897;
	wire [16-1:0] node13900;
	wire [16-1:0] node13901;
	wire [16-1:0] node13903;
	wire [16-1:0] node13904;
	wire [16-1:0] node13906;
	wire [16-1:0] node13910;
	wire [16-1:0] node13911;
	wire [16-1:0] node13914;
	wire [16-1:0] node13916;
	wire [16-1:0] node13919;
	wire [16-1:0] node13920;
	wire [16-1:0] node13921;
	wire [16-1:0] node13922;
	wire [16-1:0] node13923;
	wire [16-1:0] node13926;
	wire [16-1:0] node13927;
	wire [16-1:0] node13929;
	wire [16-1:0] node13933;
	wire [16-1:0] node13936;
	wire [16-1:0] node13937;
	wire [16-1:0] node13938;
	wire [16-1:0] node13942;
	wire [16-1:0] node13944;
	wire [16-1:0] node13947;
	wire [16-1:0] node13948;
	wire [16-1:0] node13950;
	wire [16-1:0] node13951;
	wire [16-1:0] node13954;
	wire [16-1:0] node13957;
	wire [16-1:0] node13958;
	wire [16-1:0] node13960;
	wire [16-1:0] node13963;
	wire [16-1:0] node13964;
	wire [16-1:0] node13965;
	wire [16-1:0] node13969;
	wire [16-1:0] node13971;
	wire [16-1:0] node13972;
	wire [16-1:0] node13976;
	wire [16-1:0] node13977;
	wire [16-1:0] node13978;
	wire [16-1:0] node13979;
	wire [16-1:0] node13980;
	wire [16-1:0] node13981;
	wire [16-1:0] node13982;
	wire [16-1:0] node13983;
	wire [16-1:0] node13984;
	wire [16-1:0] node13989;
	wire [16-1:0] node13992;
	wire [16-1:0] node13993;
	wire [16-1:0] node13994;
	wire [16-1:0] node13996;
	wire [16-1:0] node13999;
	wire [16-1:0] node14000;
	wire [16-1:0] node14001;
	wire [16-1:0] node14006;
	wire [16-1:0] node14007;
	wire [16-1:0] node14008;
	wire [16-1:0] node14010;
	wire [16-1:0] node14014;
	wire [16-1:0] node14017;
	wire [16-1:0] node14018;
	wire [16-1:0] node14019;
	wire [16-1:0] node14020;
	wire [16-1:0] node14022;
	wire [16-1:0] node14025;
	wire [16-1:0] node14028;
	wire [16-1:0] node14029;
	wire [16-1:0] node14030;
	wire [16-1:0] node14034;
	wire [16-1:0] node14036;
	wire [16-1:0] node14039;
	wire [16-1:0] node14040;
	wire [16-1:0] node14042;
	wire [16-1:0] node14044;
	wire [16-1:0] node14047;
	wire [16-1:0] node14048;
	wire [16-1:0] node14051;
	wire [16-1:0] node14054;
	wire [16-1:0] node14055;
	wire [16-1:0] node14056;
	wire [16-1:0] node14057;
	wire [16-1:0] node14058;
	wire [16-1:0] node14059;
	wire [16-1:0] node14063;
	wire [16-1:0] node14064;
	wire [16-1:0] node14069;
	wire [16-1:0] node14070;
	wire [16-1:0] node14071;
	wire [16-1:0] node14075;
	wire [16-1:0] node14077;
	wire [16-1:0] node14079;
	wire [16-1:0] node14081;
	wire [16-1:0] node14084;
	wire [16-1:0] node14085;
	wire [16-1:0] node14086;
	wire [16-1:0] node14087;
	wire [16-1:0] node14089;
	wire [16-1:0] node14092;
	wire [16-1:0] node14093;
	wire [16-1:0] node14097;
	wire [16-1:0] node14099;
	wire [16-1:0] node14100;
	wire [16-1:0] node14104;
	wire [16-1:0] node14105;
	wire [16-1:0] node14106;
	wire [16-1:0] node14109;
	wire [16-1:0] node14111;
	wire [16-1:0] node14114;
	wire [16-1:0] node14116;
	wire [16-1:0] node14119;
	wire [16-1:0] node14120;
	wire [16-1:0] node14121;
	wire [16-1:0] node14122;
	wire [16-1:0] node14123;
	wire [16-1:0] node14124;
	wire [16-1:0] node14125;
	wire [16-1:0] node14129;
	wire [16-1:0] node14132;
	wire [16-1:0] node14134;
	wire [16-1:0] node14137;
	wire [16-1:0] node14138;
	wire [16-1:0] node14139;
	wire [16-1:0] node14140;
	wire [16-1:0] node14142;
	wire [16-1:0] node14145;
	wire [16-1:0] node14147;
	wire [16-1:0] node14151;
	wire [16-1:0] node14153;
	wire [16-1:0] node14155;
	wire [16-1:0] node14156;
	wire [16-1:0] node14159;
	wire [16-1:0] node14162;
	wire [16-1:0] node14163;
	wire [16-1:0] node14164;
	wire [16-1:0] node14165;
	wire [16-1:0] node14167;
	wire [16-1:0] node14172;
	wire [16-1:0] node14173;
	wire [16-1:0] node14176;
	wire [16-1:0] node14178;
	wire [16-1:0] node14181;
	wire [16-1:0] node14182;
	wire [16-1:0] node14183;
	wire [16-1:0] node14184;
	wire [16-1:0] node14185;
	wire [16-1:0] node14189;
	wire [16-1:0] node14190;
	wire [16-1:0] node14191;
	wire [16-1:0] node14196;
	wire [16-1:0] node14197;
	wire [16-1:0] node14198;
	wire [16-1:0] node14199;
	wire [16-1:0] node14203;
	wire [16-1:0] node14206;
	wire [16-1:0] node14207;
	wire [16-1:0] node14208;
	wire [16-1:0] node14212;
	wire [16-1:0] node14213;
	wire [16-1:0] node14217;
	wire [16-1:0] node14218;
	wire [16-1:0] node14219;
	wire [16-1:0] node14220;
	wire [16-1:0] node14223;
	wire [16-1:0] node14224;
	wire [16-1:0] node14226;
	wire [16-1:0] node14230;
	wire [16-1:0] node14231;
	wire [16-1:0] node14234;
	wire [16-1:0] node14237;
	wire [16-1:0] node14238;
	wire [16-1:0] node14240;
	wire [16-1:0] node14242;
	wire [16-1:0] node14245;
	wire [16-1:0] node14247;
	wire [16-1:0] node14249;
	wire [16-1:0] node14252;
	wire [16-1:0] node14253;
	wire [16-1:0] node14254;
	wire [16-1:0] node14255;
	wire [16-1:0] node14256;
	wire [16-1:0] node14258;
	wire [16-1:0] node14259;
	wire [16-1:0] node14263;
	wire [16-1:0] node14264;
	wire [16-1:0] node14265;
	wire [16-1:0] node14266;
	wire [16-1:0] node14268;
	wire [16-1:0] node14272;
	wire [16-1:0] node14275;
	wire [16-1:0] node14276;
	wire [16-1:0] node14279;
	wire [16-1:0] node14282;
	wire [16-1:0] node14283;
	wire [16-1:0] node14285;
	wire [16-1:0] node14286;
	wire [16-1:0] node14288;
	wire [16-1:0] node14291;
	wire [16-1:0] node14294;
	wire [16-1:0] node14295;
	wire [16-1:0] node14298;
	wire [16-1:0] node14299;
	wire [16-1:0] node14303;
	wire [16-1:0] node14304;
	wire [16-1:0] node14305;
	wire [16-1:0] node14306;
	wire [16-1:0] node14307;
	wire [16-1:0] node14311;
	wire [16-1:0] node14312;
	wire [16-1:0] node14313;
	wire [16-1:0] node14317;
	wire [16-1:0] node14320;
	wire [16-1:0] node14321;
	wire [16-1:0] node14322;
	wire [16-1:0] node14324;
	wire [16-1:0] node14326;
	wire [16-1:0] node14329;
	wire [16-1:0] node14330;
	wire [16-1:0] node14334;
	wire [16-1:0] node14335;
	wire [16-1:0] node14337;
	wire [16-1:0] node14340;
	wire [16-1:0] node14341;
	wire [16-1:0] node14344;
	wire [16-1:0] node14346;
	wire [16-1:0] node14349;
	wire [16-1:0] node14350;
	wire [16-1:0] node14351;
	wire [16-1:0] node14352;
	wire [16-1:0] node14354;
	wire [16-1:0] node14356;
	wire [16-1:0] node14360;
	wire [16-1:0] node14361;
	wire [16-1:0] node14365;
	wire [16-1:0] node14366;
	wire [16-1:0] node14368;
	wire [16-1:0] node14369;
	wire [16-1:0] node14373;
	wire [16-1:0] node14376;
	wire [16-1:0] node14377;
	wire [16-1:0] node14378;
	wire [16-1:0] node14379;
	wire [16-1:0] node14380;
	wire [16-1:0] node14383;
	wire [16-1:0] node14386;
	wire [16-1:0] node14387;
	wire [16-1:0] node14388;
	wire [16-1:0] node14389;
	wire [16-1:0] node14394;
	wire [16-1:0] node14395;
	wire [16-1:0] node14396;
	wire [16-1:0] node14398;
	wire [16-1:0] node14402;
	wire [16-1:0] node14403;
	wire [16-1:0] node14407;
	wire [16-1:0] node14408;
	wire [16-1:0] node14409;
	wire [16-1:0] node14410;
	wire [16-1:0] node14412;
	wire [16-1:0] node14414;
	wire [16-1:0] node14417;
	wire [16-1:0] node14420;
	wire [16-1:0] node14422;
	wire [16-1:0] node14425;
	wire [16-1:0] node14426;
	wire [16-1:0] node14427;
	wire [16-1:0] node14430;
	wire [16-1:0] node14433;
	wire [16-1:0] node14434;
	wire [16-1:0] node14435;
	wire [16-1:0] node14439;
	wire [16-1:0] node14440;
	wire [16-1:0] node14444;
	wire [16-1:0] node14445;
	wire [16-1:0] node14446;
	wire [16-1:0] node14447;
	wire [16-1:0] node14449;
	wire [16-1:0] node14451;
	wire [16-1:0] node14454;
	wire [16-1:0] node14455;
	wire [16-1:0] node14458;
	wire [16-1:0] node14460;
	wire [16-1:0] node14463;
	wire [16-1:0] node14464;
	wire [16-1:0] node14466;
	wire [16-1:0] node14468;
	wire [16-1:0] node14471;
	wire [16-1:0] node14472;
	wire [16-1:0] node14473;
	wire [16-1:0] node14475;
	wire [16-1:0] node14479;
	wire [16-1:0] node14480;
	wire [16-1:0] node14484;
	wire [16-1:0] node14485;
	wire [16-1:0] node14486;
	wire [16-1:0] node14488;
	wire [16-1:0] node14491;
	wire [16-1:0] node14493;
	wire [16-1:0] node14494;
	wire [16-1:0] node14498;
	wire [16-1:0] node14499;
	wire [16-1:0] node14501;
	wire [16-1:0] node14502;
	wire [16-1:0] node14506;
	wire [16-1:0] node14508;
	wire [16-1:0] node14511;
	wire [16-1:0] node14512;
	wire [16-1:0] node14513;
	wire [16-1:0] node14514;
	wire [16-1:0] node14515;
	wire [16-1:0] node14516;
	wire [16-1:0] node14517;
	wire [16-1:0] node14518;
	wire [16-1:0] node14519;
	wire [16-1:0] node14520;
	wire [16-1:0] node14521;
	wire [16-1:0] node14525;
	wire [16-1:0] node14528;
	wire [16-1:0] node14529;
	wire [16-1:0] node14533;
	wire [16-1:0] node14535;
	wire [16-1:0] node14537;
	wire [16-1:0] node14539;
	wire [16-1:0] node14540;
	wire [16-1:0] node14544;
	wire [16-1:0] node14545;
	wire [16-1:0] node14546;
	wire [16-1:0] node14547;
	wire [16-1:0] node14548;
	wire [16-1:0] node14552;
	wire [16-1:0] node14555;
	wire [16-1:0] node14556;
	wire [16-1:0] node14557;
	wire [16-1:0] node14562;
	wire [16-1:0] node14563;
	wire [16-1:0] node14564;
	wire [16-1:0] node14565;
	wire [16-1:0] node14570;
	wire [16-1:0] node14571;
	wire [16-1:0] node14573;
	wire [16-1:0] node14574;
	wire [16-1:0] node14578;
	wire [16-1:0] node14581;
	wire [16-1:0] node14582;
	wire [16-1:0] node14583;
	wire [16-1:0] node14584;
	wire [16-1:0] node14586;
	wire [16-1:0] node14589;
	wire [16-1:0] node14591;
	wire [16-1:0] node14594;
	wire [16-1:0] node14596;
	wire [16-1:0] node14597;
	wire [16-1:0] node14598;
	wire [16-1:0] node14599;
	wire [16-1:0] node14604;
	wire [16-1:0] node14607;
	wire [16-1:0] node14608;
	wire [16-1:0] node14610;
	wire [16-1:0] node14611;
	wire [16-1:0] node14615;
	wire [16-1:0] node14616;
	wire [16-1:0] node14618;
	wire [16-1:0] node14619;
	wire [16-1:0] node14621;
	wire [16-1:0] node14625;
	wire [16-1:0] node14626;
	wire [16-1:0] node14629;
	wire [16-1:0] node14631;
	wire [16-1:0] node14634;
	wire [16-1:0] node14635;
	wire [16-1:0] node14636;
	wire [16-1:0] node14637;
	wire [16-1:0] node14638;
	wire [16-1:0] node14639;
	wire [16-1:0] node14642;
	wire [16-1:0] node14645;
	wire [16-1:0] node14647;
	wire [16-1:0] node14648;
	wire [16-1:0] node14650;
	wire [16-1:0] node14654;
	wire [16-1:0] node14656;
	wire [16-1:0] node14657;
	wire [16-1:0] node14659;
	wire [16-1:0] node14660;
	wire [16-1:0] node14665;
	wire [16-1:0] node14666;
	wire [16-1:0] node14667;
	wire [16-1:0] node14668;
	wire [16-1:0] node14671;
	wire [16-1:0] node14673;
	wire [16-1:0] node14676;
	wire [16-1:0] node14677;
	wire [16-1:0] node14680;
	wire [16-1:0] node14681;
	wire [16-1:0] node14685;
	wire [16-1:0] node14687;
	wire [16-1:0] node14688;
	wire [16-1:0] node14691;
	wire [16-1:0] node14692;
	wire [16-1:0] node14696;
	wire [16-1:0] node14697;
	wire [16-1:0] node14698;
	wire [16-1:0] node14699;
	wire [16-1:0] node14701;
	wire [16-1:0] node14702;
	wire [16-1:0] node14707;
	wire [16-1:0] node14708;
	wire [16-1:0] node14709;
	wire [16-1:0] node14712;
	wire [16-1:0] node14713;
	wire [16-1:0] node14718;
	wire [16-1:0] node14719;
	wire [16-1:0] node14720;
	wire [16-1:0] node14721;
	wire [16-1:0] node14722;
	wire [16-1:0] node14726;
	wire [16-1:0] node14729;
	wire [16-1:0] node14732;
	wire [16-1:0] node14733;
	wire [16-1:0] node14734;
	wire [16-1:0] node14736;
	wire [16-1:0] node14737;
	wire [16-1:0] node14741;
	wire [16-1:0] node14742;
	wire [16-1:0] node14746;
	wire [16-1:0] node14747;
	wire [16-1:0] node14750;
	wire [16-1:0] node14752;
	wire [16-1:0] node14755;
	wire [16-1:0] node14756;
	wire [16-1:0] node14757;
	wire [16-1:0] node14758;
	wire [16-1:0] node14759;
	wire [16-1:0] node14760;
	wire [16-1:0] node14761;
	wire [16-1:0] node14762;
	wire [16-1:0] node14764;
	wire [16-1:0] node14768;
	wire [16-1:0] node14769;
	wire [16-1:0] node14771;
	wire [16-1:0] node14775;
	wire [16-1:0] node14776;
	wire [16-1:0] node14780;
	wire [16-1:0] node14781;
	wire [16-1:0] node14782;
	wire [16-1:0] node14785;
	wire [16-1:0] node14787;
	wire [16-1:0] node14790;
	wire [16-1:0] node14791;
	wire [16-1:0] node14792;
	wire [16-1:0] node14794;
	wire [16-1:0] node14798;
	wire [16-1:0] node14799;
	wire [16-1:0] node14803;
	wire [16-1:0] node14804;
	wire [16-1:0] node14805;
	wire [16-1:0] node14806;
	wire [16-1:0] node14807;
	wire [16-1:0] node14809;
	wire [16-1:0] node14814;
	wire [16-1:0] node14815;
	wire [16-1:0] node14818;
	wire [16-1:0] node14820;
	wire [16-1:0] node14821;
	wire [16-1:0] node14825;
	wire [16-1:0] node14826;
	wire [16-1:0] node14827;
	wire [16-1:0] node14830;
	wire [16-1:0] node14833;
	wire [16-1:0] node14835;
	wire [16-1:0] node14838;
	wire [16-1:0] node14839;
	wire [16-1:0] node14840;
	wire [16-1:0] node14841;
	wire [16-1:0] node14842;
	wire [16-1:0] node14845;
	wire [16-1:0] node14847;
	wire [16-1:0] node14850;
	wire [16-1:0] node14851;
	wire [16-1:0] node14852;
	wire [16-1:0] node14856;
	wire [16-1:0] node14859;
	wire [16-1:0] node14860;
	wire [16-1:0] node14862;
	wire [16-1:0] node14865;
	wire [16-1:0] node14867;
	wire [16-1:0] node14868;
	wire [16-1:0] node14871;
	wire [16-1:0] node14874;
	wire [16-1:0] node14875;
	wire [16-1:0] node14876;
	wire [16-1:0] node14877;
	wire [16-1:0] node14880;
	wire [16-1:0] node14883;
	wire [16-1:0] node14884;
	wire [16-1:0] node14887;
	wire [16-1:0] node14889;
	wire [16-1:0] node14890;
	wire [16-1:0] node14894;
	wire [16-1:0] node14895;
	wire [16-1:0] node14897;
	wire [16-1:0] node14899;
	wire [16-1:0] node14902;
	wire [16-1:0] node14904;
	wire [16-1:0] node14907;
	wire [16-1:0] node14908;
	wire [16-1:0] node14909;
	wire [16-1:0] node14910;
	wire [16-1:0] node14911;
	wire [16-1:0] node14914;
	wire [16-1:0] node14915;
	wire [16-1:0] node14919;
	wire [16-1:0] node14920;
	wire [16-1:0] node14921;
	wire [16-1:0] node14925;
	wire [16-1:0] node14928;
	wire [16-1:0] node14929;
	wire [16-1:0] node14930;
	wire [16-1:0] node14933;
	wire [16-1:0] node14934;
	wire [16-1:0] node14938;
	wire [16-1:0] node14939;
	wire [16-1:0] node14941;
	wire [16-1:0] node14942;
	wire [16-1:0] node14946;
	wire [16-1:0] node14948;
	wire [16-1:0] node14950;
	wire [16-1:0] node14953;
	wire [16-1:0] node14954;
	wire [16-1:0] node14955;
	wire [16-1:0] node14956;
	wire [16-1:0] node14957;
	wire [16-1:0] node14958;
	wire [16-1:0] node14962;
	wire [16-1:0] node14965;
	wire [16-1:0] node14966;
	wire [16-1:0] node14969;
	wire [16-1:0] node14972;
	wire [16-1:0] node14973;
	wire [16-1:0] node14975;
	wire [16-1:0] node14978;
	wire [16-1:0] node14979;
	wire [16-1:0] node14980;
	wire [16-1:0] node14982;
	wire [16-1:0] node14986;
	wire [16-1:0] node14988;
	wire [16-1:0] node14991;
	wire [16-1:0] node14992;
	wire [16-1:0] node14993;
	wire [16-1:0] node14994;
	wire [16-1:0] node14995;
	wire [16-1:0] node14997;
	wire [16-1:0] node15001;
	wire [16-1:0] node15004;
	wire [16-1:0] node15006;
	wire [16-1:0] node15007;
	wire [16-1:0] node15011;
	wire [16-1:0] node15012;
	wire [16-1:0] node15013;
	wire [16-1:0] node15016;
	wire [16-1:0] node15017;
	wire [16-1:0] node15019;
	wire [16-1:0] node15023;
	wire [16-1:0] node15024;
	wire [16-1:0] node15025;
	wire [16-1:0] node15029;
	wire [16-1:0] node15032;
	wire [16-1:0] node15033;
	wire [16-1:0] node15034;
	wire [16-1:0] node15035;
	wire [16-1:0] node15036;
	wire [16-1:0] node15037;
	wire [16-1:0] node15038;
	wire [16-1:0] node15039;
	wire [16-1:0] node15040;
	wire [16-1:0] node15045;
	wire [16-1:0] node15046;
	wire [16-1:0] node15048;
	wire [16-1:0] node15052;
	wire [16-1:0] node15053;
	wire [16-1:0] node15054;
	wire [16-1:0] node15058;
	wire [16-1:0] node15061;
	wire [16-1:0] node15062;
	wire [16-1:0] node15064;
	wire [16-1:0] node15065;
	wire [16-1:0] node15067;
	wire [16-1:0] node15071;
	wire [16-1:0] node15072;
	wire [16-1:0] node15073;
	wire [16-1:0] node15077;
	wire [16-1:0] node15078;
	wire [16-1:0] node15081;
	wire [16-1:0] node15084;
	wire [16-1:0] node15085;
	wire [16-1:0] node15086;
	wire [16-1:0] node15087;
	wire [16-1:0] node15088;
	wire [16-1:0] node15089;
	wire [16-1:0] node15093;
	wire [16-1:0] node15096;
	wire [16-1:0] node15097;
	wire [16-1:0] node15098;
	wire [16-1:0] node15100;
	wire [16-1:0] node15104;
	wire [16-1:0] node15106;
	wire [16-1:0] node15109;
	wire [16-1:0] node15110;
	wire [16-1:0] node15112;
	wire [16-1:0] node15115;
	wire [16-1:0] node15116;
	wire [16-1:0] node15119;
	wire [16-1:0] node15122;
	wire [16-1:0] node15123;
	wire [16-1:0] node15124;
	wire [16-1:0] node15125;
	wire [16-1:0] node15127;
	wire [16-1:0] node15128;
	wire [16-1:0] node15132;
	wire [16-1:0] node15135;
	wire [16-1:0] node15136;
	wire [16-1:0] node15139;
	wire [16-1:0] node15140;
	wire [16-1:0] node15142;
	wire [16-1:0] node15146;
	wire [16-1:0] node15147;
	wire [16-1:0] node15149;
	wire [16-1:0] node15152;
	wire [16-1:0] node15153;
	wire [16-1:0] node15155;
	wire [16-1:0] node15156;
	wire [16-1:0] node15160;
	wire [16-1:0] node15163;
	wire [16-1:0] node15164;
	wire [16-1:0] node15165;
	wire [16-1:0] node15166;
	wire [16-1:0] node15167;
	wire [16-1:0] node15168;
	wire [16-1:0] node15171;
	wire [16-1:0] node15174;
	wire [16-1:0] node15175;
	wire [16-1:0] node15176;
	wire [16-1:0] node15181;
	wire [16-1:0] node15182;
	wire [16-1:0] node15183;
	wire [16-1:0] node15184;
	wire [16-1:0] node15186;
	wire [16-1:0] node15191;
	wire [16-1:0] node15193;
	wire [16-1:0] node15194;
	wire [16-1:0] node15196;
	wire [16-1:0] node15199;
	wire [16-1:0] node15202;
	wire [16-1:0] node15203;
	wire [16-1:0] node15204;
	wire [16-1:0] node15205;
	wire [16-1:0] node15209;
	wire [16-1:0] node15210;
	wire [16-1:0] node15212;
	wire [16-1:0] node15213;
	wire [16-1:0] node15217;
	wire [16-1:0] node15218;
	wire [16-1:0] node15222;
	wire [16-1:0] node15223;
	wire [16-1:0] node15224;
	wire [16-1:0] node15225;
	wire [16-1:0] node15230;
	wire [16-1:0] node15231;
	wire [16-1:0] node15233;
	wire [16-1:0] node15236;
	wire [16-1:0] node15237;
	wire [16-1:0] node15238;
	wire [16-1:0] node15243;
	wire [16-1:0] node15244;
	wire [16-1:0] node15245;
	wire [16-1:0] node15246;
	wire [16-1:0] node15247;
	wire [16-1:0] node15251;
	wire [16-1:0] node15252;
	wire [16-1:0] node15254;
	wire [16-1:0] node15255;
	wire [16-1:0] node15259;
	wire [16-1:0] node15262;
	wire [16-1:0] node15264;
	wire [16-1:0] node15265;
	wire [16-1:0] node15266;
	wire [16-1:0] node15270;
	wire [16-1:0] node15272;
	wire [16-1:0] node15273;
	wire [16-1:0] node15277;
	wire [16-1:0] node15278;
	wire [16-1:0] node15280;
	wire [16-1:0] node15281;
	wire [16-1:0] node15283;
	wire [16-1:0] node15287;
	wire [16-1:0] node15288;
	wire [16-1:0] node15289;
	wire [16-1:0] node15293;
	wire [16-1:0] node15294;
	wire [16-1:0] node15295;
	wire [16-1:0] node15296;
	wire [16-1:0] node15302;
	wire [16-1:0] node15303;
	wire [16-1:0] node15304;
	wire [16-1:0] node15305;
	wire [16-1:0] node15306;
	wire [16-1:0] node15308;
	wire [16-1:0] node15309;
	wire [16-1:0] node15311;
	wire [16-1:0] node15315;
	wire [16-1:0] node15316;
	wire [16-1:0] node15317;
	wire [16-1:0] node15320;
	wire [16-1:0] node15323;
	wire [16-1:0] node15324;
	wire [16-1:0] node15328;
	wire [16-1:0] node15329;
	wire [16-1:0] node15330;
	wire [16-1:0] node15332;
	wire [16-1:0] node15334;
	wire [16-1:0] node15337;
	wire [16-1:0] node15338;
	wire [16-1:0] node15341;
	wire [16-1:0] node15343;
	wire [16-1:0] node15346;
	wire [16-1:0] node15347;
	wire [16-1:0] node15348;
	wire [16-1:0] node15352;
	wire [16-1:0] node15353;
	wire [16-1:0] node15355;
	wire [16-1:0] node15359;
	wire [16-1:0] node15360;
	wire [16-1:0] node15361;
	wire [16-1:0] node15362;
	wire [16-1:0] node15363;
	wire [16-1:0] node15365;
	wire [16-1:0] node15366;
	wire [16-1:0] node15371;
	wire [16-1:0] node15372;
	wire [16-1:0] node15374;
	wire [16-1:0] node15377;
	wire [16-1:0] node15380;
	wire [16-1:0] node15381;
	wire [16-1:0] node15383;
	wire [16-1:0] node15384;
	wire [16-1:0] node15386;
	wire [16-1:0] node15389;
	wire [16-1:0] node15390;
	wire [16-1:0] node15394;
	wire [16-1:0] node15395;
	wire [16-1:0] node15399;
	wire [16-1:0] node15400;
	wire [16-1:0] node15401;
	wire [16-1:0] node15403;
	wire [16-1:0] node15406;
	wire [16-1:0] node15407;
	wire [16-1:0] node15408;
	wire [16-1:0] node15410;
	wire [16-1:0] node15415;
	wire [16-1:0] node15416;
	wire [16-1:0] node15418;
	wire [16-1:0] node15421;
	wire [16-1:0] node15423;
	wire [16-1:0] node15424;
	wire [16-1:0] node15425;
	wire [16-1:0] node15430;
	wire [16-1:0] node15431;
	wire [16-1:0] node15432;
	wire [16-1:0] node15433;
	wire [16-1:0] node15434;
	wire [16-1:0] node15435;
	wire [16-1:0] node15436;
	wire [16-1:0] node15440;
	wire [16-1:0] node15443;
	wire [16-1:0] node15444;
	wire [16-1:0] node15448;
	wire [16-1:0] node15449;
	wire [16-1:0] node15450;
	wire [16-1:0] node15453;
	wire [16-1:0] node15454;
	wire [16-1:0] node15456;
	wire [16-1:0] node15460;
	wire [16-1:0] node15461;
	wire [16-1:0] node15465;
	wire [16-1:0] node15466;
	wire [16-1:0] node15467;
	wire [16-1:0] node15468;
	wire [16-1:0] node15471;
	wire [16-1:0] node15473;
	wire [16-1:0] node15474;
	wire [16-1:0] node15478;
	wire [16-1:0] node15479;
	wire [16-1:0] node15480;
	wire [16-1:0] node15483;
	wire [16-1:0] node15484;
	wire [16-1:0] node15488;
	wire [16-1:0] node15489;
	wire [16-1:0] node15490;
	wire [16-1:0] node15493;
	wire [16-1:0] node15496;
	wire [16-1:0] node15497;
	wire [16-1:0] node15501;
	wire [16-1:0] node15502;
	wire [16-1:0] node15503;
	wire [16-1:0] node15506;
	wire [16-1:0] node15507;
	wire [16-1:0] node15509;
	wire [16-1:0] node15512;
	wire [16-1:0] node15513;
	wire [16-1:0] node15517;
	wire [16-1:0] node15518;
	wire [16-1:0] node15520;
	wire [16-1:0] node15522;
	wire [16-1:0] node15526;
	wire [16-1:0] node15527;
	wire [16-1:0] node15528;
	wire [16-1:0] node15529;
	wire [16-1:0] node15530;
	wire [16-1:0] node15533;
	wire [16-1:0] node15536;
	wire [16-1:0] node15537;
	wire [16-1:0] node15540;
	wire [16-1:0] node15541;
	wire [16-1:0] node15543;
	wire [16-1:0] node15547;
	wire [16-1:0] node15548;
	wire [16-1:0] node15550;
	wire [16-1:0] node15551;
	wire [16-1:0] node15553;
	wire [16-1:0] node15557;
	wire [16-1:0] node15558;
	wire [16-1:0] node15560;
	wire [16-1:0] node15561;
	wire [16-1:0] node15565;
	wire [16-1:0] node15568;
	wire [16-1:0] node15569;
	wire [16-1:0] node15570;
	wire [16-1:0] node15571;
	wire [16-1:0] node15573;
	wire [16-1:0] node15576;
	wire [16-1:0] node15577;
	wire [16-1:0] node15581;
	wire [16-1:0] node15583;
	wire [16-1:0] node15586;
	wire [16-1:0] node15587;
	wire [16-1:0] node15589;
	wire [16-1:0] node15590;
	wire [16-1:0] node15594;
	wire [16-1:0] node15596;
	wire [16-1:0] node15597;
	wire [16-1:0] node15601;
	wire [16-1:0] node15602;
	wire [16-1:0] node15603;
	wire [16-1:0] node15604;
	wire [16-1:0] node15605;
	wire [16-1:0] node15606;
	wire [16-1:0] node15607;
	wire [16-1:0] node15608;
	wire [16-1:0] node15609;
	wire [16-1:0] node15612;
	wire [16-1:0] node15614;
	wire [16-1:0] node15615;
	wire [16-1:0] node15619;
	wire [16-1:0] node15620;
	wire [16-1:0] node15622;
	wire [16-1:0] node15625;
	wire [16-1:0] node15627;
	wire [16-1:0] node15630;
	wire [16-1:0] node15631;
	wire [16-1:0] node15632;
	wire [16-1:0] node15634;
	wire [16-1:0] node15637;
	wire [16-1:0] node15640;
	wire [16-1:0] node15641;
	wire [16-1:0] node15644;
	wire [16-1:0] node15647;
	wire [16-1:0] node15648;
	wire [16-1:0] node15649;
	wire [16-1:0] node15651;
	wire [16-1:0] node15652;
	wire [16-1:0] node15655;
	wire [16-1:0] node15658;
	wire [16-1:0] node15659;
	wire [16-1:0] node15661;
	wire [16-1:0] node15662;
	wire [16-1:0] node15667;
	wire [16-1:0] node15668;
	wire [16-1:0] node15669;
	wire [16-1:0] node15672;
	wire [16-1:0] node15673;
	wire [16-1:0] node15675;
	wire [16-1:0] node15679;
	wire [16-1:0] node15681;
	wire [16-1:0] node15683;
	wire [16-1:0] node15686;
	wire [16-1:0] node15687;
	wire [16-1:0] node15688;
	wire [16-1:0] node15689;
	wire [16-1:0] node15690;
	wire [16-1:0] node15694;
	wire [16-1:0] node15695;
	wire [16-1:0] node15696;
	wire [16-1:0] node15698;
	wire [16-1:0] node15703;
	wire [16-1:0] node15704;
	wire [16-1:0] node15706;
	wire [16-1:0] node15709;
	wire [16-1:0] node15710;
	wire [16-1:0] node15711;
	wire [16-1:0] node15715;
	wire [16-1:0] node15717;
	wire [16-1:0] node15720;
	wire [16-1:0] node15722;
	wire [16-1:0] node15723;
	wire [16-1:0] node15724;
	wire [16-1:0] node15725;
	wire [16-1:0] node15727;
	wire [16-1:0] node15730;
	wire [16-1:0] node15732;
	wire [16-1:0] node15736;
	wire [16-1:0] node15737;
	wire [16-1:0] node15740;
	wire [16-1:0] node15741;
	wire [16-1:0] node15743;
	wire [16-1:0] node15747;
	wire [16-1:0] node15748;
	wire [16-1:0] node15749;
	wire [16-1:0] node15750;
	wire [16-1:0] node15751;
	wire [16-1:0] node15753;
	wire [16-1:0] node15755;
	wire [16-1:0] node15758;
	wire [16-1:0] node15759;
	wire [16-1:0] node15761;
	wire [16-1:0] node15765;
	wire [16-1:0] node15766;
	wire [16-1:0] node15768;
	wire [16-1:0] node15771;
	wire [16-1:0] node15772;
	wire [16-1:0] node15773;
	wire [16-1:0] node15775;
	wire [16-1:0] node15779;
	wire [16-1:0] node15781;
	wire [16-1:0] node15784;
	wire [16-1:0] node15785;
	wire [16-1:0] node15786;
	wire [16-1:0] node15788;
	wire [16-1:0] node15790;
	wire [16-1:0] node15793;
	wire [16-1:0] node15794;
	wire [16-1:0] node15797;
	wire [16-1:0] node15800;
	wire [16-1:0] node15801;
	wire [16-1:0] node15802;
	wire [16-1:0] node15805;
	wire [16-1:0] node15807;
	wire [16-1:0] node15808;
	wire [16-1:0] node15812;
	wire [16-1:0] node15814;
	wire [16-1:0] node15817;
	wire [16-1:0] node15818;
	wire [16-1:0] node15819;
	wire [16-1:0] node15820;
	wire [16-1:0] node15822;
	wire [16-1:0] node15825;
	wire [16-1:0] node15827;
	wire [16-1:0] node15829;
	wire [16-1:0] node15832;
	wire [16-1:0] node15833;
	wire [16-1:0] node15834;
	wire [16-1:0] node15838;
	wire [16-1:0] node15839;
	wire [16-1:0] node15841;
	wire [16-1:0] node15842;
	wire [16-1:0] node15847;
	wire [16-1:0] node15848;
	wire [16-1:0] node15849;
	wire [16-1:0] node15851;
	wire [16-1:0] node15854;
	wire [16-1:0] node15856;
	wire [16-1:0] node15859;
	wire [16-1:0] node15861;
	wire [16-1:0] node15863;
	wire [16-1:0] node15865;
	wire [16-1:0] node15867;
	wire [16-1:0] node15870;
	wire [16-1:0] node15871;
	wire [16-1:0] node15872;
	wire [16-1:0] node15873;
	wire [16-1:0] node15874;
	wire [16-1:0] node15875;
	wire [16-1:0] node15876;
	wire [16-1:0] node15880;
	wire [16-1:0] node15881;
	wire [16-1:0] node15885;
	wire [16-1:0] node15886;
	wire [16-1:0] node15890;
	wire [16-1:0] node15891;
	wire [16-1:0] node15893;
	wire [16-1:0] node15894;
	wire [16-1:0] node15896;
	wire [16-1:0] node15899;
	wire [16-1:0] node15902;
	wire [16-1:0] node15903;
	wire [16-1:0] node15906;
	wire [16-1:0] node15907;
	wire [16-1:0] node15909;
	wire [16-1:0] node15913;
	wire [16-1:0] node15914;
	wire [16-1:0] node15915;
	wire [16-1:0] node15916;
	wire [16-1:0] node15917;
	wire [16-1:0] node15919;
	wire [16-1:0] node15923;
	wire [16-1:0] node15925;
	wire [16-1:0] node15928;
	wire [16-1:0] node15929;
	wire [16-1:0] node15930;
	wire [16-1:0] node15932;
	wire [16-1:0] node15935;
	wire [16-1:0] node15937;
	wire [16-1:0] node15940;
	wire [16-1:0] node15941;
	wire [16-1:0] node15944;
	wire [16-1:0] node15947;
	wire [16-1:0] node15948;
	wire [16-1:0] node15949;
	wire [16-1:0] node15951;
	wire [16-1:0] node15952;
	wire [16-1:0] node15953;
	wire [16-1:0] node15959;
	wire [16-1:0] node15960;
	wire [16-1:0] node15961;
	wire [16-1:0] node15962;
	wire [16-1:0] node15966;
	wire [16-1:0] node15969;
	wire [16-1:0] node15970;
	wire [16-1:0] node15973;
	wire [16-1:0] node15975;
	wire [16-1:0] node15978;
	wire [16-1:0] node15979;
	wire [16-1:0] node15980;
	wire [16-1:0] node15981;
	wire [16-1:0] node15982;
	wire [16-1:0] node15984;
	wire [16-1:0] node15987;
	wire [16-1:0] node15989;
	wire [16-1:0] node15992;
	wire [16-1:0] node15993;
	wire [16-1:0] node15994;
	wire [16-1:0] node15997;
	wire [16-1:0] node16000;
	wire [16-1:0] node16001;
	wire [16-1:0] node16005;
	wire [16-1:0] node16006;
	wire [16-1:0] node16007;
	wire [16-1:0] node16008;
	wire [16-1:0] node16011;
	wire [16-1:0] node16013;
	wire [16-1:0] node16016;
	wire [16-1:0] node16018;
	wire [16-1:0] node16020;
	wire [16-1:0] node16021;
	wire [16-1:0] node16025;
	wire [16-1:0] node16026;
	wire [16-1:0] node16027;
	wire [16-1:0] node16030;
	wire [16-1:0] node16033;
	wire [16-1:0] node16034;
	wire [16-1:0] node16036;
	wire [16-1:0] node16037;
	wire [16-1:0] node16041;
	wire [16-1:0] node16043;
	wire [16-1:0] node16046;
	wire [16-1:0] node16047;
	wire [16-1:0] node16048;
	wire [16-1:0] node16049;
	wire [16-1:0] node16050;
	wire [16-1:0] node16051;
	wire [16-1:0] node16053;
	wire [16-1:0] node16057;
	wire [16-1:0] node16060;
	wire [16-1:0] node16061;
	wire [16-1:0] node16064;
	wire [16-1:0] node16066;
	wire [16-1:0] node16069;
	wire [16-1:0] node16070;
	wire [16-1:0] node16071;
	wire [16-1:0] node16074;
	wire [16-1:0] node16075;
	wire [16-1:0] node16079;
	wire [16-1:0] node16080;
	wire [16-1:0] node16082;
	wire [16-1:0] node16085;
	wire [16-1:0] node16087;
	wire [16-1:0] node16089;
	wire [16-1:0] node16092;
	wire [16-1:0] node16093;
	wire [16-1:0] node16095;
	wire [16-1:0] node16096;
	wire [16-1:0] node16099;
	wire [16-1:0] node16101;
	wire [16-1:0] node16103;
	wire [16-1:0] node16106;
	wire [16-1:0] node16107;
	wire [16-1:0] node16109;
	wire [16-1:0] node16110;
	wire [16-1:0] node16112;
	wire [16-1:0] node16115;
	wire [16-1:0] node16118;
	wire [16-1:0] node16119;
	wire [16-1:0] node16120;
	wire [16-1:0] node16124;
	wire [16-1:0] node16125;
	wire [16-1:0] node16127;
	wire [16-1:0] node16131;
	wire [16-1:0] node16132;
	wire [16-1:0] node16133;
	wire [16-1:0] node16134;
	wire [16-1:0] node16135;
	wire [16-1:0] node16136;
	wire [16-1:0] node16137;
	wire [16-1:0] node16138;
	wire [16-1:0] node16139;
	wire [16-1:0] node16143;
	wire [16-1:0] node16146;
	wire [16-1:0] node16147;
	wire [16-1:0] node16151;
	wire [16-1:0] node16154;
	wire [16-1:0] node16155;
	wire [16-1:0] node16156;
	wire [16-1:0] node16158;
	wire [16-1:0] node16161;
	wire [16-1:0] node16164;
	wire [16-1:0] node16165;
	wire [16-1:0] node16166;
	wire [16-1:0] node16168;
	wire [16-1:0] node16171;
	wire [16-1:0] node16174;
	wire [16-1:0] node16175;
	wire [16-1:0] node16179;
	wire [16-1:0] node16180;
	wire [16-1:0] node16181;
	wire [16-1:0] node16182;
	wire [16-1:0] node16183;
	wire [16-1:0] node16186;
	wire [16-1:0] node16189;
	wire [16-1:0] node16191;
	wire [16-1:0] node16192;
	wire [16-1:0] node16196;
	wire [16-1:0] node16198;
	wire [16-1:0] node16201;
	wire [16-1:0] node16202;
	wire [16-1:0] node16203;
	wire [16-1:0] node16204;
	wire [16-1:0] node16206;
	wire [16-1:0] node16207;
	wire [16-1:0] node16211;
	wire [16-1:0] node16214;
	wire [16-1:0] node16215;
	wire [16-1:0] node16216;
	wire [16-1:0] node16219;
	wire [16-1:0] node16222;
	wire [16-1:0] node16225;
	wire [16-1:0] node16226;
	wire [16-1:0] node16227;
	wire [16-1:0] node16228;
	wire [16-1:0] node16232;
	wire [16-1:0] node16233;
	wire [16-1:0] node16237;
	wire [16-1:0] node16238;
	wire [16-1:0] node16239;
	wire [16-1:0] node16241;
	wire [16-1:0] node16245;
	wire [16-1:0] node16246;
	wire [16-1:0] node16250;
	wire [16-1:0] node16251;
	wire [16-1:0] node16252;
	wire [16-1:0] node16253;
	wire [16-1:0] node16254;
	wire [16-1:0] node16256;
	wire [16-1:0] node16259;
	wire [16-1:0] node16260;
	wire [16-1:0] node16263;
	wire [16-1:0] node16265;
	wire [16-1:0] node16266;
	wire [16-1:0] node16270;
	wire [16-1:0] node16272;
	wire [16-1:0] node16274;
	wire [16-1:0] node16277;
	wire [16-1:0] node16278;
	wire [16-1:0] node16279;
	wire [16-1:0] node16280;
	wire [16-1:0] node16281;
	wire [16-1:0] node16285;
	wire [16-1:0] node16287;
	wire [16-1:0] node16290;
	wire [16-1:0] node16291;
	wire [16-1:0] node16292;
	wire [16-1:0] node16296;
	wire [16-1:0] node16299;
	wire [16-1:0] node16300;
	wire [16-1:0] node16303;
	wire [16-1:0] node16305;
	wire [16-1:0] node16308;
	wire [16-1:0] node16309;
	wire [16-1:0] node16310;
	wire [16-1:0] node16311;
	wire [16-1:0] node16314;
	wire [16-1:0] node16315;
	wire [16-1:0] node16317;
	wire [16-1:0] node16318;
	wire [16-1:0] node16322;
	wire [16-1:0] node16323;
	wire [16-1:0] node16327;
	wire [16-1:0] node16328;
	wire [16-1:0] node16329;
	wire [16-1:0] node16332;
	wire [16-1:0] node16334;
	wire [16-1:0] node16337;
	wire [16-1:0] node16338;
	wire [16-1:0] node16341;
	wire [16-1:0] node16342;
	wire [16-1:0] node16344;
	wire [16-1:0] node16348;
	wire [16-1:0] node16349;
	wire [16-1:0] node16350;
	wire [16-1:0] node16352;
	wire [16-1:0] node16353;
	wire [16-1:0] node16354;
	wire [16-1:0] node16358;
	wire [16-1:0] node16359;
	wire [16-1:0] node16362;
	wire [16-1:0] node16366;
	wire [16-1:0] node16367;
	wire [16-1:0] node16368;
	wire [16-1:0] node16369;
	wire [16-1:0] node16371;
	wire [16-1:0] node16374;
	wire [16-1:0] node16375;
	wire [16-1:0] node16378;
	wire [16-1:0] node16381;
	wire [16-1:0] node16383;
	wire [16-1:0] node16384;
	wire [16-1:0] node16388;
	wire [16-1:0] node16389;
	wire [16-1:0] node16390;
	wire [16-1:0] node16392;
	wire [16-1:0] node16396;
	wire [16-1:0] node16399;
	wire [16-1:0] node16400;
	wire [16-1:0] node16401;
	wire [16-1:0] node16402;
	wire [16-1:0] node16403;
	wire [16-1:0] node16404;
	wire [16-1:0] node16405;
	wire [16-1:0] node16408;
	wire [16-1:0] node16411;
	wire [16-1:0] node16412;
	wire [16-1:0] node16416;
	wire [16-1:0] node16417;
	wire [16-1:0] node16419;
	wire [16-1:0] node16420;
	wire [16-1:0] node16422;
	wire [16-1:0] node16425;
	wire [16-1:0] node16428;
	wire [16-1:0] node16430;
	wire [16-1:0] node16433;
	wire [16-1:0] node16434;
	wire [16-1:0] node16435;
	wire [16-1:0] node16437;
	wire [16-1:0] node16440;
	wire [16-1:0] node16441;
	wire [16-1:0] node16444;
	wire [16-1:0] node16446;
	wire [16-1:0] node16447;
	wire [16-1:0] node16451;
	wire [16-1:0] node16452;
	wire [16-1:0] node16453;
	wire [16-1:0] node16456;
	wire [16-1:0] node16457;
	wire [16-1:0] node16461;
	wire [16-1:0] node16463;
	wire [16-1:0] node16464;
	wire [16-1:0] node16468;
	wire [16-1:0] node16469;
	wire [16-1:0] node16470;
	wire [16-1:0] node16471;
	wire [16-1:0] node16473;
	wire [16-1:0] node16477;
	wire [16-1:0] node16478;
	wire [16-1:0] node16480;
	wire [16-1:0] node16483;
	wire [16-1:0] node16485;
	wire [16-1:0] node16488;
	wire [16-1:0] node16489;
	wire [16-1:0] node16490;
	wire [16-1:0] node16492;
	wire [16-1:0] node16495;
	wire [16-1:0] node16496;
	wire [16-1:0] node16498;
	wire [16-1:0] node16501;
	wire [16-1:0] node16503;
	wire [16-1:0] node16506;
	wire [16-1:0] node16507;
	wire [16-1:0] node16508;
	wire [16-1:0] node16509;
	wire [16-1:0] node16513;
	wire [16-1:0] node16515;
	wire [16-1:0] node16518;
	wire [16-1:0] node16519;
	wire [16-1:0] node16522;
	wire [16-1:0] node16524;
	wire [16-1:0] node16527;
	wire [16-1:0] node16528;
	wire [16-1:0] node16529;
	wire [16-1:0] node16530;
	wire [16-1:0] node16532;
	wire [16-1:0] node16533;
	wire [16-1:0] node16534;
	wire [16-1:0] node16538;
	wire [16-1:0] node16541;
	wire [16-1:0] node16542;
	wire [16-1:0] node16543;
	wire [16-1:0] node16546;
	wire [16-1:0] node16547;
	wire [16-1:0] node16549;
	wire [16-1:0] node16553;
	wire [16-1:0] node16555;
	wire [16-1:0] node16558;
	wire [16-1:0] node16559;
	wire [16-1:0] node16560;
	wire [16-1:0] node16562;
	wire [16-1:0] node16563;
	wire [16-1:0] node16567;
	wire [16-1:0] node16568;
	wire [16-1:0] node16571;
	wire [16-1:0] node16574;
	wire [16-1:0] node16575;
	wire [16-1:0] node16577;
	wire [16-1:0] node16580;
	wire [16-1:0] node16581;
	wire [16-1:0] node16584;
	wire [16-1:0] node16585;
	wire [16-1:0] node16589;
	wire [16-1:0] node16590;
	wire [16-1:0] node16591;
	wire [16-1:0] node16592;
	wire [16-1:0] node16594;
	wire [16-1:0] node16597;
	wire [16-1:0] node16598;
	wire [16-1:0] node16601;
	wire [16-1:0] node16603;
	wire [16-1:0] node16606;
	wire [16-1:0] node16607;
	wire [16-1:0] node16609;
	wire [16-1:0] node16611;
	wire [16-1:0] node16614;
	wire [16-1:0] node16615;
	wire [16-1:0] node16618;
	wire [16-1:0] node16621;
	wire [16-1:0] node16622;
	wire [16-1:0] node16623;
	wire [16-1:0] node16625;
	wire [16-1:0] node16628;
	wire [16-1:0] node16631;
	wire [16-1:0] node16632;
	wire [16-1:0] node16633;
	wire [16-1:0] node16635;
	wire [16-1:0] node16639;
	wire [16-1:0] node16642;
	wire [16-1:0] node16643;
	wire [16-1:0] node16644;
	wire [16-1:0] node16645;
	wire [16-1:0] node16646;
	wire [16-1:0] node16647;
	wire [16-1:0] node16648;
	wire [16-1:0] node16649;
	wire [16-1:0] node16650;
	wire [16-1:0] node16651;
	wire [16-1:0] node16652;
	wire [16-1:0] node16653;
	wire [16-1:0] node16654;
	wire [16-1:0] node16658;
	wire [16-1:0] node16659;
	wire [16-1:0] node16660;
	wire [16-1:0] node16661;
	wire [16-1:0] node16665;
	wire [16-1:0] node16666;
	wire [16-1:0] node16671;
	wire [16-1:0] node16672;
	wire [16-1:0] node16673;
	wire [16-1:0] node16675;
	wire [16-1:0] node16676;
	wire [16-1:0] node16681;
	wire [16-1:0] node16682;
	wire [16-1:0] node16686;
	wire [16-1:0] node16687;
	wire [16-1:0] node16688;
	wire [16-1:0] node16689;
	wire [16-1:0] node16690;
	wire [16-1:0] node16694;
	wire [16-1:0] node16697;
	wire [16-1:0] node16698;
	wire [16-1:0] node16699;
	wire [16-1:0] node16702;
	wire [16-1:0] node16705;
	wire [16-1:0] node16708;
	wire [16-1:0] node16709;
	wire [16-1:0] node16710;
	wire [16-1:0] node16712;
	wire [16-1:0] node16715;
	wire [16-1:0] node16717;
	wire [16-1:0] node16720;
	wire [16-1:0] node16721;
	wire [16-1:0] node16722;
	wire [16-1:0] node16727;
	wire [16-1:0] node16728;
	wire [16-1:0] node16729;
	wire [16-1:0] node16730;
	wire [16-1:0] node16731;
	wire [16-1:0] node16732;
	wire [16-1:0] node16733;
	wire [16-1:0] node16738;
	wire [16-1:0] node16741;
	wire [16-1:0] node16742;
	wire [16-1:0] node16746;
	wire [16-1:0] node16747;
	wire [16-1:0] node16748;
	wire [16-1:0] node16750;
	wire [16-1:0] node16751;
	wire [16-1:0] node16755;
	wire [16-1:0] node16758;
	wire [16-1:0] node16759;
	wire [16-1:0] node16762;
	wire [16-1:0] node16765;
	wire [16-1:0] node16766;
	wire [16-1:0] node16767;
	wire [16-1:0] node16768;
	wire [16-1:0] node16770;
	wire [16-1:0] node16771;
	wire [16-1:0] node16775;
	wire [16-1:0] node16777;
	wire [16-1:0] node16780;
	wire [16-1:0] node16781;
	wire [16-1:0] node16784;
	wire [16-1:0] node16787;
	wire [16-1:0] node16788;
	wire [16-1:0] node16790;
	wire [16-1:0] node16793;
	wire [16-1:0] node16794;
	wire [16-1:0] node16797;
	wire [16-1:0] node16799;
	wire [16-1:0] node16802;
	wire [16-1:0] node16803;
	wire [16-1:0] node16804;
	wire [16-1:0] node16805;
	wire [16-1:0] node16806;
	wire [16-1:0] node16807;
	wire [16-1:0] node16810;
	wire [16-1:0] node16813;
	wire [16-1:0] node16814;
	wire [16-1:0] node16815;
	wire [16-1:0] node16817;
	wire [16-1:0] node16821;
	wire [16-1:0] node16824;
	wire [16-1:0] node16825;
	wire [16-1:0] node16828;
	wire [16-1:0] node16830;
	wire [16-1:0] node16833;
	wire [16-1:0] node16834;
	wire [16-1:0] node16835;
	wire [16-1:0] node16836;
	wire [16-1:0] node16837;
	wire [16-1:0] node16840;
	wire [16-1:0] node16843;
	wire [16-1:0] node16845;
	wire [16-1:0] node16848;
	wire [16-1:0] node16849;
	wire [16-1:0] node16850;
	wire [16-1:0] node16854;
	wire [16-1:0] node16857;
	wire [16-1:0] node16858;
	wire [16-1:0] node16860;
	wire [16-1:0] node16863;
	wire [16-1:0] node16864;
	wire [16-1:0] node16865;
	wire [16-1:0] node16869;
	wire [16-1:0] node16872;
	wire [16-1:0] node16873;
	wire [16-1:0] node16874;
	wire [16-1:0] node16875;
	wire [16-1:0] node16876;
	wire [16-1:0] node16878;
	wire [16-1:0] node16881;
	wire [16-1:0] node16882;
	wire [16-1:0] node16883;
	wire [16-1:0] node16889;
	wire [16-1:0] node16890;
	wire [16-1:0] node16891;
	wire [16-1:0] node16895;
	wire [16-1:0] node16896;
	wire [16-1:0] node16897;
	wire [16-1:0] node16898;
	wire [16-1:0] node16903;
	wire [16-1:0] node16904;
	wire [16-1:0] node16906;
	wire [16-1:0] node16910;
	wire [16-1:0] node16911;
	wire [16-1:0] node16912;
	wire [16-1:0] node16914;
	wire [16-1:0] node16916;
	wire [16-1:0] node16919;
	wire [16-1:0] node16922;
	wire [16-1:0] node16923;
	wire [16-1:0] node16926;
	wire [16-1:0] node16928;
	wire [16-1:0] node16930;
	wire [16-1:0] node16933;
	wire [16-1:0] node16934;
	wire [16-1:0] node16935;
	wire [16-1:0] node16936;
	wire [16-1:0] node16937;
	wire [16-1:0] node16938;
	wire [16-1:0] node16940;
	wire [16-1:0] node16941;
	wire [16-1:0] node16945;
	wire [16-1:0] node16946;
	wire [16-1:0] node16947;
	wire [16-1:0] node16948;
	wire [16-1:0] node16952;
	wire [16-1:0] node16955;
	wire [16-1:0] node16957;
	wire [16-1:0] node16960;
	wire [16-1:0] node16961;
	wire [16-1:0] node16962;
	wire [16-1:0] node16964;
	wire [16-1:0] node16965;
	wire [16-1:0] node16969;
	wire [16-1:0] node16972;
	wire [16-1:0] node16974;
	wire [16-1:0] node16977;
	wire [16-1:0] node16978;
	wire [16-1:0] node16979;
	wire [16-1:0] node16980;
	wire [16-1:0] node16983;
	wire [16-1:0] node16986;
	wire [16-1:0] node16987;
	wire [16-1:0] node16990;
	wire [16-1:0] node16991;
	wire [16-1:0] node16995;
	wire [16-1:0] node16996;
	wire [16-1:0] node16997;
	wire [16-1:0] node16999;
	wire [16-1:0] node17003;
	wire [16-1:0] node17005;
	wire [16-1:0] node17008;
	wire [16-1:0] node17009;
	wire [16-1:0] node17010;
	wire [16-1:0] node17011;
	wire [16-1:0] node17012;
	wire [16-1:0] node17014;
	wire [16-1:0] node17015;
	wire [16-1:0] node17020;
	wire [16-1:0] node17021;
	wire [16-1:0] node17023;
	wire [16-1:0] node17024;
	wire [16-1:0] node17028;
	wire [16-1:0] node17030;
	wire [16-1:0] node17033;
	wire [16-1:0] node17034;
	wire [16-1:0] node17035;
	wire [16-1:0] node17038;
	wire [16-1:0] node17040;
	wire [16-1:0] node17043;
	wire [16-1:0] node17044;
	wire [16-1:0] node17048;
	wire [16-1:0] node17049;
	wire [16-1:0] node17050;
	wire [16-1:0] node17051;
	wire [16-1:0] node17054;
	wire [16-1:0] node17057;
	wire [16-1:0] node17058;
	wire [16-1:0] node17059;
	wire [16-1:0] node17062;
	wire [16-1:0] node17065;
	wire [16-1:0] node17067;
	wire [16-1:0] node17068;
	wire [16-1:0] node17072;
	wire [16-1:0] node17073;
	wire [16-1:0] node17075;
	wire [16-1:0] node17076;
	wire [16-1:0] node17080;
	wire [16-1:0] node17081;
	wire [16-1:0] node17083;
	wire [16-1:0] node17087;
	wire [16-1:0] node17088;
	wire [16-1:0] node17089;
	wire [16-1:0] node17090;
	wire [16-1:0] node17091;
	wire [16-1:0] node17092;
	wire [16-1:0] node17094;
	wire [16-1:0] node17097;
	wire [16-1:0] node17100;
	wire [16-1:0] node17103;
	wire [16-1:0] node17104;
	wire [16-1:0] node17105;
	wire [16-1:0] node17106;
	wire [16-1:0] node17111;
	wire [16-1:0] node17112;
	wire [16-1:0] node17114;
	wire [16-1:0] node17118;
	wire [16-1:0] node17119;
	wire [16-1:0] node17120;
	wire [16-1:0] node17122;
	wire [16-1:0] node17124;
	wire [16-1:0] node17127;
	wire [16-1:0] node17128;
	wire [16-1:0] node17131;
	wire [16-1:0] node17134;
	wire [16-1:0] node17135;
	wire [16-1:0] node17136;
	wire [16-1:0] node17138;
	wire [16-1:0] node17141;
	wire [16-1:0] node17143;
	wire [16-1:0] node17146;
	wire [16-1:0] node17147;
	wire [16-1:0] node17149;
	wire [16-1:0] node17150;
	wire [16-1:0] node17154;
	wire [16-1:0] node17157;
	wire [16-1:0] node17158;
	wire [16-1:0] node17159;
	wire [16-1:0] node17160;
	wire [16-1:0] node17161;
	wire [16-1:0] node17163;
	wire [16-1:0] node17166;
	wire [16-1:0] node17168;
	wire [16-1:0] node17169;
	wire [16-1:0] node17173;
	wire [16-1:0] node17174;
	wire [16-1:0] node17178;
	wire [16-1:0] node17180;
	wire [16-1:0] node17181;
	wire [16-1:0] node17184;
	wire [16-1:0] node17187;
	wire [16-1:0] node17188;
	wire [16-1:0] node17189;
	wire [16-1:0] node17190;
	wire [16-1:0] node17192;
	wire [16-1:0] node17195;
	wire [16-1:0] node17198;
	wire [16-1:0] node17200;
	wire [16-1:0] node17203;
	wire [16-1:0] node17204;
	wire [16-1:0] node17205;
	wire [16-1:0] node17208;
	wire [16-1:0] node17211;
	wire [16-1:0] node17212;
	wire [16-1:0] node17215;
	wire [16-1:0] node17216;
	wire [16-1:0] node17220;
	wire [16-1:0] node17221;
	wire [16-1:0] node17222;
	wire [16-1:0] node17223;
	wire [16-1:0] node17224;
	wire [16-1:0] node17225;
	wire [16-1:0] node17226;
	wire [16-1:0] node17228;
	wire [16-1:0] node17230;
	wire [16-1:0] node17233;
	wire [16-1:0] node17234;
	wire [16-1:0] node17237;
	wire [16-1:0] node17240;
	wire [16-1:0] node17241;
	wire [16-1:0] node17242;
	wire [16-1:0] node17244;
	wire [16-1:0] node17245;
	wire [16-1:0] node17249;
	wire [16-1:0] node17251;
	wire [16-1:0] node17252;
	wire [16-1:0] node17256;
	wire [16-1:0] node17257;
	wire [16-1:0] node17260;
	wire [16-1:0] node17263;
	wire [16-1:0] node17264;
	wire [16-1:0] node17265;
	wire [16-1:0] node17266;
	wire [16-1:0] node17267;
	wire [16-1:0] node17271;
	wire [16-1:0] node17274;
	wire [16-1:0] node17275;
	wire [16-1:0] node17276;
	wire [16-1:0] node17278;
	wire [16-1:0] node17282;
	wire [16-1:0] node17284;
	wire [16-1:0] node17286;
	wire [16-1:0] node17289;
	wire [16-1:0] node17290;
	wire [16-1:0] node17291;
	wire [16-1:0] node17294;
	wire [16-1:0] node17295;
	wire [16-1:0] node17299;
	wire [16-1:0] node17300;
	wire [16-1:0] node17303;
	wire [16-1:0] node17304;
	wire [16-1:0] node17308;
	wire [16-1:0] node17309;
	wire [16-1:0] node17310;
	wire [16-1:0] node17311;
	wire [16-1:0] node17312;
	wire [16-1:0] node17315;
	wire [16-1:0] node17318;
	wire [16-1:0] node17319;
	wire [16-1:0] node17320;
	wire [16-1:0] node17324;
	wire [16-1:0] node17325;
	wire [16-1:0] node17327;
	wire [16-1:0] node17331;
	wire [16-1:0] node17332;
	wire [16-1:0] node17334;
	wire [16-1:0] node17336;
	wire [16-1:0] node17339;
	wire [16-1:0] node17340;
	wire [16-1:0] node17341;
	wire [16-1:0] node17346;
	wire [16-1:0] node17347;
	wire [16-1:0] node17348;
	wire [16-1:0] node17349;
	wire [16-1:0] node17350;
	wire [16-1:0] node17354;
	wire [16-1:0] node17357;
	wire [16-1:0] node17358;
	wire [16-1:0] node17360;
	wire [16-1:0] node17361;
	wire [16-1:0] node17366;
	wire [16-1:0] node17367;
	wire [16-1:0] node17368;
	wire [16-1:0] node17369;
	wire [16-1:0] node17373;
	wire [16-1:0] node17376;
	wire [16-1:0] node17377;
	wire [16-1:0] node17381;
	wire [16-1:0] node17382;
	wire [16-1:0] node17383;
	wire [16-1:0] node17384;
	wire [16-1:0] node17385;
	wire [16-1:0] node17386;
	wire [16-1:0] node17387;
	wire [16-1:0] node17388;
	wire [16-1:0] node17392;
	wire [16-1:0] node17395;
	wire [16-1:0] node17397;
	wire [16-1:0] node17400;
	wire [16-1:0] node17401;
	wire [16-1:0] node17405;
	wire [16-1:0] node17406;
	wire [16-1:0] node17407;
	wire [16-1:0] node17408;
	wire [16-1:0] node17411;
	wire [16-1:0] node17415;
	wire [16-1:0] node17416;
	wire [16-1:0] node17417;
	wire [16-1:0] node17419;
	wire [16-1:0] node17423;
	wire [16-1:0] node17424;
	wire [16-1:0] node17426;
	wire [16-1:0] node17430;
	wire [16-1:0] node17431;
	wire [16-1:0] node17432;
	wire [16-1:0] node17433;
	wire [16-1:0] node17437;
	wire [16-1:0] node17438;
	wire [16-1:0] node17441;
	wire [16-1:0] node17443;
	wire [16-1:0] node17446;
	wire [16-1:0] node17447;
	wire [16-1:0] node17448;
	wire [16-1:0] node17451;
	wire [16-1:0] node17452;
	wire [16-1:0] node17453;
	wire [16-1:0] node17458;
	wire [16-1:0] node17459;
	wire [16-1:0] node17463;
	wire [16-1:0] node17464;
	wire [16-1:0] node17465;
	wire [16-1:0] node17466;
	wire [16-1:0] node17468;
	wire [16-1:0] node17470;
	wire [16-1:0] node17473;
	wire [16-1:0] node17474;
	wire [16-1:0] node17478;
	wire [16-1:0] node17479;
	wire [16-1:0] node17481;
	wire [16-1:0] node17483;
	wire [16-1:0] node17486;
	wire [16-1:0] node17487;
	wire [16-1:0] node17489;
	wire [16-1:0] node17492;
	wire [16-1:0] node17493;
	wire [16-1:0] node17497;
	wire [16-1:0] node17498;
	wire [16-1:0] node17499;
	wire [16-1:0] node17500;
	wire [16-1:0] node17502;
	wire [16-1:0] node17505;
	wire [16-1:0] node17508;
	wire [16-1:0] node17509;
	wire [16-1:0] node17511;
	wire [16-1:0] node17512;
	wire [16-1:0] node17516;
	wire [16-1:0] node17519;
	wire [16-1:0] node17520;
	wire [16-1:0] node17521;
	wire [16-1:0] node17522;
	wire [16-1:0] node17526;
	wire [16-1:0] node17529;
	wire [16-1:0] node17530;
	wire [16-1:0] node17533;
	wire [16-1:0] node17536;
	wire [16-1:0] node17537;
	wire [16-1:0] node17538;
	wire [16-1:0] node17539;
	wire [16-1:0] node17540;
	wire [16-1:0] node17541;
	wire [16-1:0] node17542;
	wire [16-1:0] node17545;
	wire [16-1:0] node17548;
	wire [16-1:0] node17549;
	wire [16-1:0] node17551;
	wire [16-1:0] node17555;
	wire [16-1:0] node17556;
	wire [16-1:0] node17557;
	wire [16-1:0] node17560;
	wire [16-1:0] node17563;
	wire [16-1:0] node17564;
	wire [16-1:0] node17568;
	wire [16-1:0] node17569;
	wire [16-1:0] node17570;
	wire [16-1:0] node17571;
	wire [16-1:0] node17575;
	wire [16-1:0] node17578;
	wire [16-1:0] node17579;
	wire [16-1:0] node17581;
	wire [16-1:0] node17584;
	wire [16-1:0] node17585;
	wire [16-1:0] node17586;
	wire [16-1:0] node17591;
	wire [16-1:0] node17592;
	wire [16-1:0] node17593;
	wire [16-1:0] node17594;
	wire [16-1:0] node17595;
	wire [16-1:0] node17598;
	wire [16-1:0] node17600;
	wire [16-1:0] node17601;
	wire [16-1:0] node17605;
	wire [16-1:0] node17606;
	wire [16-1:0] node17610;
	wire [16-1:0] node17612;
	wire [16-1:0] node17613;
	wire [16-1:0] node17616;
	wire [16-1:0] node17619;
	wire [16-1:0] node17620;
	wire [16-1:0] node17621;
	wire [16-1:0] node17622;
	wire [16-1:0] node17623;
	wire [16-1:0] node17627;
	wire [16-1:0] node17628;
	wire [16-1:0] node17630;
	wire [16-1:0] node17634;
	wire [16-1:0] node17635;
	wire [16-1:0] node17638;
	wire [16-1:0] node17641;
	wire [16-1:0] node17642;
	wire [16-1:0] node17644;
	wire [16-1:0] node17645;
	wire [16-1:0] node17650;
	wire [16-1:0] node17651;
	wire [16-1:0] node17652;
	wire [16-1:0] node17653;
	wire [16-1:0] node17654;
	wire [16-1:0] node17655;
	wire [16-1:0] node17659;
	wire [16-1:0] node17660;
	wire [16-1:0] node17662;
	wire [16-1:0] node17666;
	wire [16-1:0] node17667;
	wire [16-1:0] node17668;
	wire [16-1:0] node17670;
	wire [16-1:0] node17671;
	wire [16-1:0] node17676;
	wire [16-1:0] node17677;
	wire [16-1:0] node17681;
	wire [16-1:0] node17682;
	wire [16-1:0] node17683;
	wire [16-1:0] node17684;
	wire [16-1:0] node17687;
	wire [16-1:0] node17690;
	wire [16-1:0] node17691;
	wire [16-1:0] node17693;
	wire [16-1:0] node17697;
	wire [16-1:0] node17698;
	wire [16-1:0] node17700;
	wire [16-1:0] node17701;
	wire [16-1:0] node17703;
	wire [16-1:0] node17708;
	wire [16-1:0] node17709;
	wire [16-1:0] node17710;
	wire [16-1:0] node17711;
	wire [16-1:0] node17712;
	wire [16-1:0] node17715;
	wire [16-1:0] node17717;
	wire [16-1:0] node17720;
	wire [16-1:0] node17721;
	wire [16-1:0] node17725;
	wire [16-1:0] node17726;
	wire [16-1:0] node17727;
	wire [16-1:0] node17731;
	wire [16-1:0] node17732;
	wire [16-1:0] node17733;
	wire [16-1:0] node17737;
	wire [16-1:0] node17740;
	wire [16-1:0] node17741;
	wire [16-1:0] node17742;
	wire [16-1:0] node17743;
	wire [16-1:0] node17746;
	wire [16-1:0] node17747;
	wire [16-1:0] node17751;
	wire [16-1:0] node17752;
	wire [16-1:0] node17753;
	wire [16-1:0] node17758;
	wire [16-1:0] node17759;
	wire [16-1:0] node17761;
	wire [16-1:0] node17764;
	wire [16-1:0] node17766;
	wire [16-1:0] node17767;
	wire [16-1:0] node17769;
	wire [16-1:0] node17773;
	wire [16-1:0] node17774;
	wire [16-1:0] node17775;
	wire [16-1:0] node17776;
	wire [16-1:0] node17777;
	wire [16-1:0] node17778;
	wire [16-1:0] node17779;
	wire [16-1:0] node17780;
	wire [16-1:0] node17781;
	wire [16-1:0] node17782;
	wire [16-1:0] node17785;
	wire [16-1:0] node17786;
	wire [16-1:0] node17790;
	wire [16-1:0] node17791;
	wire [16-1:0] node17792;
	wire [16-1:0] node17797;
	wire [16-1:0] node17798;
	wire [16-1:0] node17802;
	wire [16-1:0] node17803;
	wire [16-1:0] node17805;
	wire [16-1:0] node17807;
	wire [16-1:0] node17810;
	wire [16-1:0] node17812;
	wire [16-1:0] node17814;
	wire [16-1:0] node17817;
	wire [16-1:0] node17818;
	wire [16-1:0] node17820;
	wire [16-1:0] node17821;
	wire [16-1:0] node17825;
	wire [16-1:0] node17826;
	wire [16-1:0] node17828;
	wire [16-1:0] node17831;
	wire [16-1:0] node17834;
	wire [16-1:0] node17835;
	wire [16-1:0] node17836;
	wire [16-1:0] node17837;
	wire [16-1:0] node17838;
	wire [16-1:0] node17840;
	wire [16-1:0] node17843;
	wire [16-1:0] node17846;
	wire [16-1:0] node17848;
	wire [16-1:0] node17849;
	wire [16-1:0] node17853;
	wire [16-1:0] node17854;
	wire [16-1:0] node17855;
	wire [16-1:0] node17858;
	wire [16-1:0] node17859;
	wire [16-1:0] node17863;
	wire [16-1:0] node17865;
	wire [16-1:0] node17868;
	wire [16-1:0] node17869;
	wire [16-1:0] node17870;
	wire [16-1:0] node17872;
	wire [16-1:0] node17875;
	wire [16-1:0] node17876;
	wire [16-1:0] node17879;
	wire [16-1:0] node17880;
	wire [16-1:0] node17881;
	wire [16-1:0] node17886;
	wire [16-1:0] node17887;
	wire [16-1:0] node17888;
	wire [16-1:0] node17890;
	wire [16-1:0] node17892;
	wire [16-1:0] node17895;
	wire [16-1:0] node17898;
	wire [16-1:0] node17899;
	wire [16-1:0] node17902;
	wire [16-1:0] node17904;
	wire [16-1:0] node17907;
	wire [16-1:0] node17908;
	wire [16-1:0] node17909;
	wire [16-1:0] node17910;
	wire [16-1:0] node17911;
	wire [16-1:0] node17913;
	wire [16-1:0] node17915;
	wire [16-1:0] node17916;
	wire [16-1:0] node17920;
	wire [16-1:0] node17921;
	wire [16-1:0] node17925;
	wire [16-1:0] node17927;
	wire [16-1:0] node17928;
	wire [16-1:0] node17931;
	wire [16-1:0] node17934;
	wire [16-1:0] node17935;
	wire [16-1:0] node17936;
	wire [16-1:0] node17937;
	wire [16-1:0] node17939;
	wire [16-1:0] node17942;
	wire [16-1:0] node17943;
	wire [16-1:0] node17945;
	wire [16-1:0] node17949;
	wire [16-1:0] node17950;
	wire [16-1:0] node17953;
	wire [16-1:0] node17956;
	wire [16-1:0] node17958;
	wire [16-1:0] node17960;
	wire [16-1:0] node17963;
	wire [16-1:0] node17964;
	wire [16-1:0] node17965;
	wire [16-1:0] node17966;
	wire [16-1:0] node17967;
	wire [16-1:0] node17968;
	wire [16-1:0] node17972;
	wire [16-1:0] node17975;
	wire [16-1:0] node17976;
	wire [16-1:0] node17980;
	wire [16-1:0] node17981;
	wire [16-1:0] node17982;
	wire [16-1:0] node17983;
	wire [16-1:0] node17985;
	wire [16-1:0] node17989;
	wire [16-1:0] node17991;
	wire [16-1:0] node17994;
	wire [16-1:0] node17997;
	wire [16-1:0] node17998;
	wire [16-1:0] node17999;
	wire [16-1:0] node18000;
	wire [16-1:0] node18001;
	wire [16-1:0] node18003;
	wire [16-1:0] node18006;
	wire [16-1:0] node18009;
	wire [16-1:0] node18011;
	wire [16-1:0] node18014;
	wire [16-1:0] node18015;
	wire [16-1:0] node18018;
	wire [16-1:0] node18021;
	wire [16-1:0] node18022;
	wire [16-1:0] node18023;
	wire [16-1:0] node18026;
	wire [16-1:0] node18029;
	wire [16-1:0] node18030;
	wire [16-1:0] node18033;
	wire [16-1:0] node18036;
	wire [16-1:0] node18037;
	wire [16-1:0] node18038;
	wire [16-1:0] node18039;
	wire [16-1:0] node18040;
	wire [16-1:0] node18041;
	wire [16-1:0] node18042;
	wire [16-1:0] node18045;
	wire [16-1:0] node18047;
	wire [16-1:0] node18050;
	wire [16-1:0] node18051;
	wire [16-1:0] node18055;
	wire [16-1:0] node18057;
	wire [16-1:0] node18058;
	wire [16-1:0] node18062;
	wire [16-1:0] node18063;
	wire [16-1:0] node18064;
	wire [16-1:0] node18065;
	wire [16-1:0] node18066;
	wire [16-1:0] node18070;
	wire [16-1:0] node18073;
	wire [16-1:0] node18074;
	wire [16-1:0] node18078;
	wire [16-1:0] node18079;
	wire [16-1:0] node18081;
	wire [16-1:0] node18083;
	wire [16-1:0] node18087;
	wire [16-1:0] node18088;
	wire [16-1:0] node18089;
	wire [16-1:0] node18090;
	wire [16-1:0] node18091;
	wire [16-1:0] node18094;
	wire [16-1:0] node18096;
	wire [16-1:0] node18099;
	wire [16-1:0] node18101;
	wire [16-1:0] node18104;
	wire [16-1:0] node18106;
	wire [16-1:0] node18107;
	wire [16-1:0] node18108;
	wire [16-1:0] node18109;
	wire [16-1:0] node18114;
	wire [16-1:0] node18117;
	wire [16-1:0] node18118;
	wire [16-1:0] node18120;
	wire [16-1:0] node18121;
	wire [16-1:0] node18122;
	wire [16-1:0] node18124;
	wire [16-1:0] node18129;
	wire [16-1:0] node18130;
	wire [16-1:0] node18131;
	wire [16-1:0] node18134;
	wire [16-1:0] node18137;
	wire [16-1:0] node18138;
	wire [16-1:0] node18141;
	wire [16-1:0] node18143;
	wire [16-1:0] node18145;
	wire [16-1:0] node18148;
	wire [16-1:0] node18149;
	wire [16-1:0] node18150;
	wire [16-1:0] node18151;
	wire [16-1:0] node18152;
	wire [16-1:0] node18153;
	wire [16-1:0] node18155;
	wire [16-1:0] node18159;
	wire [16-1:0] node18160;
	wire [16-1:0] node18162;
	wire [16-1:0] node18163;
	wire [16-1:0] node18167;
	wire [16-1:0] node18170;
	wire [16-1:0] node18171;
	wire [16-1:0] node18172;
	wire [16-1:0] node18175;
	wire [16-1:0] node18178;
	wire [16-1:0] node18179;
	wire [16-1:0] node18181;
	wire [16-1:0] node18182;
	wire [16-1:0] node18186;
	wire [16-1:0] node18188;
	wire [16-1:0] node18191;
	wire [16-1:0] node18192;
	wire [16-1:0] node18193;
	wire [16-1:0] node18194;
	wire [16-1:0] node18196;
	wire [16-1:0] node18201;
	wire [16-1:0] node18202;
	wire [16-1:0] node18203;
	wire [16-1:0] node18205;
	wire [16-1:0] node18208;
	wire [16-1:0] node18209;
	wire [16-1:0] node18211;
	wire [16-1:0] node18215;
	wire [16-1:0] node18217;
	wire [16-1:0] node18220;
	wire [16-1:0] node18221;
	wire [16-1:0] node18222;
	wire [16-1:0] node18223;
	wire [16-1:0] node18224;
	wire [16-1:0] node18227;
	wire [16-1:0] node18231;
	wire [16-1:0] node18232;
	wire [16-1:0] node18233;
	wire [16-1:0] node18236;
	wire [16-1:0] node18238;
	wire [16-1:0] node18239;
	wire [16-1:0] node18243;
	wire [16-1:0] node18246;
	wire [16-1:0] node18247;
	wire [16-1:0] node18248;
	wire [16-1:0] node18249;
	wire [16-1:0] node18252;
	wire [16-1:0] node18255;
	wire [16-1:0] node18256;
	wire [16-1:0] node18260;
	wire [16-1:0] node18261;
	wire [16-1:0] node18262;
	wire [16-1:0] node18263;
	wire [16-1:0] node18267;
	wire [16-1:0] node18269;
	wire [16-1:0] node18273;
	wire [16-1:0] node18274;
	wire [16-1:0] node18275;
	wire [16-1:0] node18276;
	wire [16-1:0] node18277;
	wire [16-1:0] node18278;
	wire [16-1:0] node18279;
	wire [16-1:0] node18280;
	wire [16-1:0] node18283;
	wire [16-1:0] node18286;
	wire [16-1:0] node18287;
	wire [16-1:0] node18290;
	wire [16-1:0] node18293;
	wire [16-1:0] node18294;
	wire [16-1:0] node18295;
	wire [16-1:0] node18298;
	wire [16-1:0] node18301;
	wire [16-1:0] node18302;
	wire [16-1:0] node18303;
	wire [16-1:0] node18307;
	wire [16-1:0] node18310;
	wire [16-1:0] node18311;
	wire [16-1:0] node18312;
	wire [16-1:0] node18313;
	wire [16-1:0] node18316;
	wire [16-1:0] node18318;
	wire [16-1:0] node18321;
	wire [16-1:0] node18322;
	wire [16-1:0] node18323;
	wire [16-1:0] node18327;
	wire [16-1:0] node18328;
	wire [16-1:0] node18332;
	wire [16-1:0] node18333;
	wire [16-1:0] node18335;
	wire [16-1:0] node18338;
	wire [16-1:0] node18339;
	wire [16-1:0] node18343;
	wire [16-1:0] node18344;
	wire [16-1:0] node18345;
	wire [16-1:0] node18347;
	wire [16-1:0] node18348;
	wire [16-1:0] node18352;
	wire [16-1:0] node18353;
	wire [16-1:0] node18354;
	wire [16-1:0] node18355;
	wire [16-1:0] node18360;
	wire [16-1:0] node18362;
	wire [16-1:0] node18365;
	wire [16-1:0] node18366;
	wire [16-1:0] node18367;
	wire [16-1:0] node18368;
	wire [16-1:0] node18372;
	wire [16-1:0] node18373;
	wire [16-1:0] node18376;
	wire [16-1:0] node18379;
	wire [16-1:0] node18380;
	wire [16-1:0] node18381;
	wire [16-1:0] node18385;
	wire [16-1:0] node18386;
	wire [16-1:0] node18387;
	wire [16-1:0] node18392;
	wire [16-1:0] node18393;
	wire [16-1:0] node18394;
	wire [16-1:0] node18395;
	wire [16-1:0] node18396;
	wire [16-1:0] node18398;
	wire [16-1:0] node18402;
	wire [16-1:0] node18403;
	wire [16-1:0] node18405;
	wire [16-1:0] node18406;
	wire [16-1:0] node18411;
	wire [16-1:0] node18412;
	wire [16-1:0] node18413;
	wire [16-1:0] node18414;
	wire [16-1:0] node18417;
	wire [16-1:0] node18419;
	wire [16-1:0] node18422;
	wire [16-1:0] node18423;
	wire [16-1:0] node18426;
	wire [16-1:0] node18429;
	wire [16-1:0] node18430;
	wire [16-1:0] node18431;
	wire [16-1:0] node18433;
	wire [16-1:0] node18434;
	wire [16-1:0] node18438;
	wire [16-1:0] node18441;
	wire [16-1:0] node18442;
	wire [16-1:0] node18445;
	wire [16-1:0] node18446;
	wire [16-1:0] node18450;
	wire [16-1:0] node18451;
	wire [16-1:0] node18452;
	wire [16-1:0] node18453;
	wire [16-1:0] node18456;
	wire [16-1:0] node18457;
	wire [16-1:0] node18460;
	wire [16-1:0] node18463;
	wire [16-1:0] node18464;
	wire [16-1:0] node18465;
	wire [16-1:0] node18468;
	wire [16-1:0] node18471;
	wire [16-1:0] node18472;
	wire [16-1:0] node18475;
	wire [16-1:0] node18477;
	wire [16-1:0] node18480;
	wire [16-1:0] node18481;
	wire [16-1:0] node18482;
	wire [16-1:0] node18483;
	wire [16-1:0] node18486;
	wire [16-1:0] node18490;
	wire [16-1:0] node18491;
	wire [16-1:0] node18494;
	wire [16-1:0] node18495;
	wire [16-1:0] node18496;
	wire [16-1:0] node18500;
	wire [16-1:0] node18503;
	wire [16-1:0] node18504;
	wire [16-1:0] node18505;
	wire [16-1:0] node18506;
	wire [16-1:0] node18507;
	wire [16-1:0] node18508;
	wire [16-1:0] node18510;
	wire [16-1:0] node18514;
	wire [16-1:0] node18515;
	wire [16-1:0] node18516;
	wire [16-1:0] node18518;
	wire [16-1:0] node18520;
	wire [16-1:0] node18523;
	wire [16-1:0] node18527;
	wire [16-1:0] node18528;
	wire [16-1:0] node18529;
	wire [16-1:0] node18532;
	wire [16-1:0] node18533;
	wire [16-1:0] node18536;
	wire [16-1:0] node18539;
	wire [16-1:0] node18540;
	wire [16-1:0] node18541;
	wire [16-1:0] node18542;
	wire [16-1:0] node18546;
	wire [16-1:0] node18547;
	wire [16-1:0] node18548;
	wire [16-1:0] node18553;
	wire [16-1:0] node18554;
	wire [16-1:0] node18557;
	wire [16-1:0] node18560;
	wire [16-1:0] node18561;
	wire [16-1:0] node18562;
	wire [16-1:0] node18565;
	wire [16-1:0] node18567;
	wire [16-1:0] node18568;
	wire [16-1:0] node18572;
	wire [16-1:0] node18573;
	wire [16-1:0] node18576;
	wire [16-1:0] node18577;
	wire [16-1:0] node18578;
	wire [16-1:0] node18583;
	wire [16-1:0] node18584;
	wire [16-1:0] node18585;
	wire [16-1:0] node18586;
	wire [16-1:0] node18587;
	wire [16-1:0] node18588;
	wire [16-1:0] node18589;
	wire [16-1:0] node18593;
	wire [16-1:0] node18597;
	wire [16-1:0] node18598;
	wire [16-1:0] node18599;
	wire [16-1:0] node18602;
	wire [16-1:0] node18605;
	wire [16-1:0] node18606;
	wire [16-1:0] node18607;
	wire [16-1:0] node18612;
	wire [16-1:0] node18613;
	wire [16-1:0] node18615;
	wire [16-1:0] node18617;
	wire [16-1:0] node18618;
	wire [16-1:0] node18619;
	wire [16-1:0] node18624;
	wire [16-1:0] node18625;
	wire [16-1:0] node18628;
	wire [16-1:0] node18629;
	wire [16-1:0] node18632;
	wire [16-1:0] node18635;
	wire [16-1:0] node18636;
	wire [16-1:0] node18637;
	wire [16-1:0] node18638;
	wire [16-1:0] node18639;
	wire [16-1:0] node18643;
	wire [16-1:0] node18644;
	wire [16-1:0] node18646;
	wire [16-1:0] node18647;
	wire [16-1:0] node18651;
	wire [16-1:0] node18652;
	wire [16-1:0] node18655;
	wire [16-1:0] node18658;
	wire [16-1:0] node18659;
	wire [16-1:0] node18661;
	wire [16-1:0] node18664;
	wire [16-1:0] node18665;
	wire [16-1:0] node18666;
	wire [16-1:0] node18670;
	wire [16-1:0] node18673;
	wire [16-1:0] node18674;
	wire [16-1:0] node18675;
	wire [16-1:0] node18677;
	wire [16-1:0] node18680;
	wire [16-1:0] node18682;
	wire [16-1:0] node18685;
	wire [16-1:0] node18686;
	wire [16-1:0] node18688;
	wire [16-1:0] node18689;
	wire [16-1:0] node18693;
	wire [16-1:0] node18694;
	wire [16-1:0] node18696;
	wire [16-1:0] node18698;
	wire [16-1:0] node18701;
	wire [16-1:0] node18703;
	wire [16-1:0] node18706;
	wire [16-1:0] node18707;
	wire [16-1:0] node18708;
	wire [16-1:0] node18709;
	wire [16-1:0] node18710;
	wire [16-1:0] node18711;
	wire [16-1:0] node18712;
	wire [16-1:0] node18713;
	wire [16-1:0] node18714;
	wire [16-1:0] node18715;
	wire [16-1:0] node18717;
	wire [16-1:0] node18718;
	wire [16-1:0] node18722;
	wire [16-1:0] node18723;
	wire [16-1:0] node18727;
	wire [16-1:0] node18728;
	wire [16-1:0] node18729;
	wire [16-1:0] node18734;
	wire [16-1:0] node18735;
	wire [16-1:0] node18737;
	wire [16-1:0] node18740;
	wire [16-1:0] node18741;
	wire [16-1:0] node18745;
	wire [16-1:0] node18746;
	wire [16-1:0] node18747;
	wire [16-1:0] node18749;
	wire [16-1:0] node18752;
	wire [16-1:0] node18753;
	wire [16-1:0] node18755;
	wire [16-1:0] node18759;
	wire [16-1:0] node18760;
	wire [16-1:0] node18761;
	wire [16-1:0] node18763;
	wire [16-1:0] node18766;
	wire [16-1:0] node18769;
	wire [16-1:0] node18770;
	wire [16-1:0] node18773;
	wire [16-1:0] node18775;
	wire [16-1:0] node18778;
	wire [16-1:0] node18779;
	wire [16-1:0] node18780;
	wire [16-1:0] node18781;
	wire [16-1:0] node18782;
	wire [16-1:0] node18783;
	wire [16-1:0] node18788;
	wire [16-1:0] node18790;
	wire [16-1:0] node18793;
	wire [16-1:0] node18794;
	wire [16-1:0] node18795;
	wire [16-1:0] node18798;
	wire [16-1:0] node18801;
	wire [16-1:0] node18802;
	wire [16-1:0] node18805;
	wire [16-1:0] node18807;
	wire [16-1:0] node18810;
	wire [16-1:0] node18811;
	wire [16-1:0] node18812;
	wire [16-1:0] node18813;
	wire [16-1:0] node18816;
	wire [16-1:0] node18817;
	wire [16-1:0] node18818;
	wire [16-1:0] node18823;
	wire [16-1:0] node18824;
	wire [16-1:0] node18826;
	wire [16-1:0] node18829;
	wire [16-1:0] node18831;
	wire [16-1:0] node18832;
	wire [16-1:0] node18836;
	wire [16-1:0] node18837;
	wire [16-1:0] node18838;
	wire [16-1:0] node18839;
	wire [16-1:0] node18841;
	wire [16-1:0] node18844;
	wire [16-1:0] node18846;
	wire [16-1:0] node18849;
	wire [16-1:0] node18853;
	wire [16-1:0] node18854;
	wire [16-1:0] node18855;
	wire [16-1:0] node18856;
	wire [16-1:0] node18857;
	wire [16-1:0] node18859;
	wire [16-1:0] node18861;
	wire [16-1:0] node18864;
	wire [16-1:0] node18865;
	wire [16-1:0] node18867;
	wire [16-1:0] node18871;
	wire [16-1:0] node18872;
	wire [16-1:0] node18873;
	wire [16-1:0] node18875;
	wire [16-1:0] node18879;
	wire [16-1:0] node18880;
	wire [16-1:0] node18881;
	wire [16-1:0] node18885;
	wire [16-1:0] node18888;
	wire [16-1:0] node18889;
	wire [16-1:0] node18890;
	wire [16-1:0] node18893;
	wire [16-1:0] node18894;
	wire [16-1:0] node18897;
	wire [16-1:0] node18899;
	wire [16-1:0] node18902;
	wire [16-1:0] node18903;
	wire [16-1:0] node18904;
	wire [16-1:0] node18906;
	wire [16-1:0] node18909;
	wire [16-1:0] node18912;
	wire [16-1:0] node18913;
	wire [16-1:0] node18914;
	wire [16-1:0] node18916;
	wire [16-1:0] node18920;
	wire [16-1:0] node18923;
	wire [16-1:0] node18924;
	wire [16-1:0] node18925;
	wire [16-1:0] node18926;
	wire [16-1:0] node18928;
	wire [16-1:0] node18929;
	wire [16-1:0] node18933;
	wire [16-1:0] node18934;
	wire [16-1:0] node18937;
	wire [16-1:0] node18939;
	wire [16-1:0] node18942;
	wire [16-1:0] node18944;
	wire [16-1:0] node18945;
	wire [16-1:0] node18947;
	wire [16-1:0] node18948;
	wire [16-1:0] node18952;
	wire [16-1:0] node18954;
	wire [16-1:0] node18957;
	wire [16-1:0] node18958;
	wire [16-1:0] node18959;
	wire [16-1:0] node18960;
	wire [16-1:0] node18964;
	wire [16-1:0] node18965;
	wire [16-1:0] node18968;
	wire [16-1:0] node18970;
	wire [16-1:0] node18973;
	wire [16-1:0] node18974;
	wire [16-1:0] node18975;
	wire [16-1:0] node18978;
	wire [16-1:0] node18981;
	wire [16-1:0] node18982;
	wire [16-1:0] node18984;
	wire [16-1:0] node18987;
	wire [16-1:0] node18989;
	wire [16-1:0] node18992;
	wire [16-1:0] node18993;
	wire [16-1:0] node18994;
	wire [16-1:0] node18995;
	wire [16-1:0] node18996;
	wire [16-1:0] node18997;
	wire [16-1:0] node18998;
	wire [16-1:0] node18999;
	wire [16-1:0] node19003;
	wire [16-1:0] node19004;
	wire [16-1:0] node19006;
	wire [16-1:0] node19011;
	wire [16-1:0] node19012;
	wire [16-1:0] node19013;
	wire [16-1:0] node19014;
	wire [16-1:0] node19018;
	wire [16-1:0] node19021;
	wire [16-1:0] node19022;
	wire [16-1:0] node19026;
	wire [16-1:0] node19027;
	wire [16-1:0] node19028;
	wire [16-1:0] node19029;
	wire [16-1:0] node19031;
	wire [16-1:0] node19035;
	wire [16-1:0] node19036;
	wire [16-1:0] node19040;
	wire [16-1:0] node19041;
	wire [16-1:0] node19042;
	wire [16-1:0] node19045;
	wire [16-1:0] node19048;
	wire [16-1:0] node19049;
	wire [16-1:0] node19052;
	wire [16-1:0] node19054;
	wire [16-1:0] node19055;
	wire [16-1:0] node19059;
	wire [16-1:0] node19060;
	wire [16-1:0] node19061;
	wire [16-1:0] node19062;
	wire [16-1:0] node19064;
	wire [16-1:0] node19066;
	wire [16-1:0] node19069;
	wire [16-1:0] node19070;
	wire [16-1:0] node19071;
	wire [16-1:0] node19076;
	wire [16-1:0] node19078;
	wire [16-1:0] node19081;
	wire [16-1:0] node19082;
	wire [16-1:0] node19083;
	wire [16-1:0] node19084;
	wire [16-1:0] node19087;
	wire [16-1:0] node19088;
	wire [16-1:0] node19092;
	wire [16-1:0] node19093;
	wire [16-1:0] node19094;
	wire [16-1:0] node19098;
	wire [16-1:0] node19099;
	wire [16-1:0] node19100;
	wire [16-1:0] node19105;
	wire [16-1:0] node19106;
	wire [16-1:0] node19107;
	wire [16-1:0] node19110;
	wire [16-1:0] node19112;
	wire [16-1:0] node19113;
	wire [16-1:0] node19117;
	wire [16-1:0] node19118;
	wire [16-1:0] node19119;
	wire [16-1:0] node19124;
	wire [16-1:0] node19125;
	wire [16-1:0] node19126;
	wire [16-1:0] node19127;
	wire [16-1:0] node19128;
	wire [16-1:0] node19131;
	wire [16-1:0] node19133;
	wire [16-1:0] node19136;
	wire [16-1:0] node19137;
	wire [16-1:0] node19139;
	wire [16-1:0] node19140;
	wire [16-1:0] node19144;
	wire [16-1:0] node19146;
	wire [16-1:0] node19149;
	wire [16-1:0] node19150;
	wire [16-1:0] node19151;
	wire [16-1:0] node19153;
	wire [16-1:0] node19156;
	wire [16-1:0] node19158;
	wire [16-1:0] node19159;
	wire [16-1:0] node19163;
	wire [16-1:0] node19164;
	wire [16-1:0] node19165;
	wire [16-1:0] node19168;
	wire [16-1:0] node19172;
	wire [16-1:0] node19173;
	wire [16-1:0] node19174;
	wire [16-1:0] node19175;
	wire [16-1:0] node19177;
	wire [16-1:0] node19181;
	wire [16-1:0] node19182;
	wire [16-1:0] node19183;
	wire [16-1:0] node19186;
	wire [16-1:0] node19187;
	wire [16-1:0] node19191;
	wire [16-1:0] node19192;
	wire [16-1:0] node19195;
	wire [16-1:0] node19198;
	wire [16-1:0] node19199;
	wire [16-1:0] node19200;
	wire [16-1:0] node19202;
	wire [16-1:0] node19205;
	wire [16-1:0] node19206;
	wire [16-1:0] node19207;
	wire [16-1:0] node19212;
	wire [16-1:0] node19213;
	wire [16-1:0] node19215;
	wire [16-1:0] node19218;
	wire [16-1:0] node19219;
	wire [16-1:0] node19220;
	wire [16-1:0] node19225;
	wire [16-1:0] node19226;
	wire [16-1:0] node19227;
	wire [16-1:0] node19228;
	wire [16-1:0] node19229;
	wire [16-1:0] node19230;
	wire [16-1:0] node19231;
	wire [16-1:0] node19232;
	wire [16-1:0] node19236;
	wire [16-1:0] node19237;
	wire [16-1:0] node19240;
	wire [16-1:0] node19243;
	wire [16-1:0] node19244;
	wire [16-1:0] node19245;
	wire [16-1:0] node19248;
	wire [16-1:0] node19250;
	wire [16-1:0] node19251;
	wire [16-1:0] node19255;
	wire [16-1:0] node19256;
	wire [16-1:0] node19258;
	wire [16-1:0] node19259;
	wire [16-1:0] node19263;
	wire [16-1:0] node19266;
	wire [16-1:0] node19267;
	wire [16-1:0] node19269;
	wire [16-1:0] node19270;
	wire [16-1:0] node19273;
	wire [16-1:0] node19276;
	wire [16-1:0] node19278;
	wire [16-1:0] node19279;
	wire [16-1:0] node19280;
	wire [16-1:0] node19281;
	wire [16-1:0] node19285;
	wire [16-1:0] node19286;
	wire [16-1:0] node19290;
	wire [16-1:0] node19293;
	wire [16-1:0] node19294;
	wire [16-1:0] node19295;
	wire [16-1:0] node19296;
	wire [16-1:0] node19297;
	wire [16-1:0] node19300;
	wire [16-1:0] node19303;
	wire [16-1:0] node19304;
	wire [16-1:0] node19305;
	wire [16-1:0] node19307;
	wire [16-1:0] node19310;
	wire [16-1:0] node19314;
	wire [16-1:0] node19315;
	wire [16-1:0] node19316;
	wire [16-1:0] node19319;
	wire [16-1:0] node19321;
	wire [16-1:0] node19324;
	wire [16-1:0] node19325;
	wire [16-1:0] node19327;
	wire [16-1:0] node19331;
	wire [16-1:0] node19332;
	wire [16-1:0] node19333;
	wire [16-1:0] node19334;
	wire [16-1:0] node19337;
	wire [16-1:0] node19341;
	wire [16-1:0] node19342;
	wire [16-1:0] node19343;
	wire [16-1:0] node19345;
	wire [16-1:0] node19346;
	wire [16-1:0] node19350;
	wire [16-1:0] node19353;
	wire [16-1:0] node19355;
	wire [16-1:0] node19358;
	wire [16-1:0] node19359;
	wire [16-1:0] node19360;
	wire [16-1:0] node19361;
	wire [16-1:0] node19362;
	wire [16-1:0] node19363;
	wire [16-1:0] node19365;
	wire [16-1:0] node19366;
	wire [16-1:0] node19370;
	wire [16-1:0] node19373;
	wire [16-1:0] node19374;
	wire [16-1:0] node19375;
	wire [16-1:0] node19378;
	wire [16-1:0] node19381;
	wire [16-1:0] node19383;
	wire [16-1:0] node19384;
	wire [16-1:0] node19388;
	wire [16-1:0] node19389;
	wire [16-1:0] node19390;
	wire [16-1:0] node19393;
	wire [16-1:0] node19394;
	wire [16-1:0] node19396;
	wire [16-1:0] node19399;
	wire [16-1:0] node19400;
	wire [16-1:0] node19404;
	wire [16-1:0] node19407;
	wire [16-1:0] node19408;
	wire [16-1:0] node19409;
	wire [16-1:0] node19410;
	wire [16-1:0] node19413;
	wire [16-1:0] node19416;
	wire [16-1:0] node19417;
	wire [16-1:0] node19420;
	wire [16-1:0] node19422;
	wire [16-1:0] node19425;
	wire [16-1:0] node19426;
	wire [16-1:0] node19428;
	wire [16-1:0] node19430;
	wire [16-1:0] node19433;
	wire [16-1:0] node19434;
	wire [16-1:0] node19436;
	wire [16-1:0] node19439;
	wire [16-1:0] node19441;
	wire [16-1:0] node19444;
	wire [16-1:0] node19445;
	wire [16-1:0] node19446;
	wire [16-1:0] node19447;
	wire [16-1:0] node19449;
	wire [16-1:0] node19451;
	wire [16-1:0] node19455;
	wire [16-1:0] node19456;
	wire [16-1:0] node19459;
	wire [16-1:0] node19460;
	wire [16-1:0] node19464;
	wire [16-1:0] node19465;
	wire [16-1:0] node19466;
	wire [16-1:0] node19467;
	wire [16-1:0] node19471;
	wire [16-1:0] node19472;
	wire [16-1:0] node19475;
	wire [16-1:0] node19477;
	wire [16-1:0] node19478;
	wire [16-1:0] node19482;
	wire [16-1:0] node19483;
	wire [16-1:0] node19485;
	wire [16-1:0] node19487;
	wire [16-1:0] node19489;
	wire [16-1:0] node19492;
	wire [16-1:0] node19495;
	wire [16-1:0] node19496;
	wire [16-1:0] node19497;
	wire [16-1:0] node19498;
	wire [16-1:0] node19499;
	wire [16-1:0] node19500;
	wire [16-1:0] node19503;
	wire [16-1:0] node19505;
	wire [16-1:0] node19506;
	wire [16-1:0] node19510;
	wire [16-1:0] node19511;
	wire [16-1:0] node19512;
	wire [16-1:0] node19516;
	wire [16-1:0] node19518;
	wire [16-1:0] node19521;
	wire [16-1:0] node19522;
	wire [16-1:0] node19524;
	wire [16-1:0] node19525;
	wire [16-1:0] node19526;
	wire [16-1:0] node19528;
	wire [16-1:0] node19533;
	wire [16-1:0] node19534;
	wire [16-1:0] node19535;
	wire [16-1:0] node19538;
	wire [16-1:0] node19541;
	wire [16-1:0] node19542;
	wire [16-1:0] node19544;
	wire [16-1:0] node19545;
	wire [16-1:0] node19550;
	wire [16-1:0] node19551;
	wire [16-1:0] node19552;
	wire [16-1:0] node19553;
	wire [16-1:0] node19554;
	wire [16-1:0] node19558;
	wire [16-1:0] node19560;
	wire [16-1:0] node19562;
	wire [16-1:0] node19565;
	wire [16-1:0] node19566;
	wire [16-1:0] node19568;
	wire [16-1:0] node19569;
	wire [16-1:0] node19571;
	wire [16-1:0] node19575;
	wire [16-1:0] node19577;
	wire [16-1:0] node19580;
	wire [16-1:0] node19581;
	wire [16-1:0] node19583;
	wire [16-1:0] node19584;
	wire [16-1:0] node19585;
	wire [16-1:0] node19587;
	wire [16-1:0] node19591;
	wire [16-1:0] node19594;
	wire [16-1:0] node19595;
	wire [16-1:0] node19597;
	wire [16-1:0] node19598;
	wire [16-1:0] node19603;
	wire [16-1:0] node19604;
	wire [16-1:0] node19605;
	wire [16-1:0] node19606;
	wire [16-1:0] node19607;
	wire [16-1:0] node19608;
	wire [16-1:0] node19612;
	wire [16-1:0] node19613;
	wire [16-1:0] node19617;
	wire [16-1:0] node19619;
	wire [16-1:0] node19620;
	wire [16-1:0] node19623;
	wire [16-1:0] node19626;
	wire [16-1:0] node19627;
	wire [16-1:0] node19628;
	wire [16-1:0] node19629;
	wire [16-1:0] node19631;
	wire [16-1:0] node19633;
	wire [16-1:0] node19636;
	wire [16-1:0] node19637;
	wire [16-1:0] node19641;
	wire [16-1:0] node19642;
	wire [16-1:0] node19644;
	wire [16-1:0] node19646;
	wire [16-1:0] node19650;
	wire [16-1:0] node19651;
	wire [16-1:0] node19652;
	wire [16-1:0] node19655;
	wire [16-1:0] node19658;
	wire [16-1:0] node19659;
	wire [16-1:0] node19661;
	wire [16-1:0] node19663;
	wire [16-1:0] node19667;
	wire [16-1:0] node19668;
	wire [16-1:0] node19669;
	wire [16-1:0] node19670;
	wire [16-1:0] node19672;
	wire [16-1:0] node19674;
	wire [16-1:0] node19675;
	wire [16-1:0] node19679;
	wire [16-1:0] node19680;
	wire [16-1:0] node19684;
	wire [16-1:0] node19686;
	wire [16-1:0] node19687;
	wire [16-1:0] node19688;
	wire [16-1:0] node19690;
	wire [16-1:0] node19694;
	wire [16-1:0] node19696;
	wire [16-1:0] node19699;
	wire [16-1:0] node19700;
	wire [16-1:0] node19701;
	wire [16-1:0] node19704;
	wire [16-1:0] node19707;
	wire [16-1:0] node19708;
	wire [16-1:0] node19710;
	wire [16-1:0] node19713;
	wire [16-1:0] node19716;
	wire [16-1:0] node19717;
	wire [16-1:0] node19718;
	wire [16-1:0] node19719;
	wire [16-1:0] node19720;
	wire [16-1:0] node19721;
	wire [16-1:0] node19722;
	wire [16-1:0] node19723;
	wire [16-1:0] node19724;
	wire [16-1:0] node19726;
	wire [16-1:0] node19727;
	wire [16-1:0] node19732;
	wire [16-1:0] node19733;
	wire [16-1:0] node19737;
	wire [16-1:0] node19738;
	wire [16-1:0] node19739;
	wire [16-1:0] node19740;
	wire [16-1:0] node19742;
	wire [16-1:0] node19746;
	wire [16-1:0] node19749;
	wire [16-1:0] node19752;
	wire [16-1:0] node19753;
	wire [16-1:0] node19754;
	wire [16-1:0] node19757;
	wire [16-1:0] node19758;
	wire [16-1:0] node19759;
	wire [16-1:0] node19763;
	wire [16-1:0] node19766;
	wire [16-1:0] node19767;
	wire [16-1:0] node19768;
	wire [16-1:0] node19769;
	wire [16-1:0] node19773;
	wire [16-1:0] node19775;
	wire [16-1:0] node19778;
	wire [16-1:0] node19779;
	wire [16-1:0] node19780;
	wire [16-1:0] node19784;
	wire [16-1:0] node19787;
	wire [16-1:0] node19788;
	wire [16-1:0] node19789;
	wire [16-1:0] node19790;
	wire [16-1:0] node19791;
	wire [16-1:0] node19794;
	wire [16-1:0] node19795;
	wire [16-1:0] node19799;
	wire [16-1:0] node19800;
	wire [16-1:0] node19801;
	wire [16-1:0] node19806;
	wire [16-1:0] node19807;
	wire [16-1:0] node19808;
	wire [16-1:0] node19809;
	wire [16-1:0] node19813;
	wire [16-1:0] node19814;
	wire [16-1:0] node19816;
	wire [16-1:0] node19820;
	wire [16-1:0] node19821;
	wire [16-1:0] node19822;
	wire [16-1:0] node19826;
	wire [16-1:0] node19829;
	wire [16-1:0] node19830;
	wire [16-1:0] node19831;
	wire [16-1:0] node19832;
	wire [16-1:0] node19834;
	wire [16-1:0] node19838;
	wire [16-1:0] node19839;
	wire [16-1:0] node19842;
	wire [16-1:0] node19845;
	wire [16-1:0] node19846;
	wire [16-1:0] node19848;
	wire [16-1:0] node19849;
	wire [16-1:0] node19853;
	wire [16-1:0] node19855;
	wire [16-1:0] node19856;
	wire [16-1:0] node19860;
	wire [16-1:0] node19861;
	wire [16-1:0] node19862;
	wire [16-1:0] node19863;
	wire [16-1:0] node19864;
	wire [16-1:0] node19865;
	wire [16-1:0] node19868;
	wire [16-1:0] node19871;
	wire [16-1:0] node19872;
	wire [16-1:0] node19873;
	wire [16-1:0] node19877;
	wire [16-1:0] node19880;
	wire [16-1:0] node19881;
	wire [16-1:0] node19882;
	wire [16-1:0] node19883;
	wire [16-1:0] node19887;
	wire [16-1:0] node19888;
	wire [16-1:0] node19890;
	wire [16-1:0] node19894;
	wire [16-1:0] node19897;
	wire [16-1:0] node19898;
	wire [16-1:0] node19900;
	wire [16-1:0] node19901;
	wire [16-1:0] node19904;
	wire [16-1:0] node19906;
	wire [16-1:0] node19909;
	wire [16-1:0] node19911;
	wire [16-1:0] node19912;
	wire [16-1:0] node19914;
	wire [16-1:0] node19915;
	wire [16-1:0] node19920;
	wire [16-1:0] node19921;
	wire [16-1:0] node19922;
	wire [16-1:0] node19923;
	wire [16-1:0] node19925;
	wire [16-1:0] node19928;
	wire [16-1:0] node19929;
	wire [16-1:0] node19930;
	wire [16-1:0] node19934;
	wire [16-1:0] node19937;
	wire [16-1:0] node19938;
	wire [16-1:0] node19939;
	wire [16-1:0] node19940;
	wire [16-1:0] node19944;
	wire [16-1:0] node19946;
	wire [16-1:0] node19947;
	wire [16-1:0] node19951;
	wire [16-1:0] node19953;
	wire [16-1:0] node19956;
	wire [16-1:0] node19957;
	wire [16-1:0] node19958;
	wire [16-1:0] node19961;
	wire [16-1:0] node19962;
	wire [16-1:0] node19964;
	wire [16-1:0] node19967;
	wire [16-1:0] node19970;
	wire [16-1:0] node19971;
	wire [16-1:0] node19974;
	wire [16-1:0] node19976;
	wire [16-1:0] node19978;
	wire [16-1:0] node19980;
	wire [16-1:0] node19983;
	wire [16-1:0] node19984;
	wire [16-1:0] node19985;
	wire [16-1:0] node19986;
	wire [16-1:0] node19987;
	wire [16-1:0] node19988;
	wire [16-1:0] node19990;
	wire [16-1:0] node19993;
	wire [16-1:0] node19994;
	wire [16-1:0] node19995;
	wire [16-1:0] node19999;
	wire [16-1:0] node20002;
	wire [16-1:0] node20003;
	wire [16-1:0] node20005;
	wire [16-1:0] node20008;
	wire [16-1:0] node20009;
	wire [16-1:0] node20011;
	wire [16-1:0] node20012;
	wire [16-1:0] node20017;
	wire [16-1:0] node20018;
	wire [16-1:0] node20019;
	wire [16-1:0] node20021;
	wire [16-1:0] node20024;
	wire [16-1:0] node20025;
	wire [16-1:0] node20029;
	wire [16-1:0] node20030;
	wire [16-1:0] node20031;
	wire [16-1:0] node20032;
	wire [16-1:0] node20036;
	wire [16-1:0] node20039;
	wire [16-1:0] node20042;
	wire [16-1:0] node20043;
	wire [16-1:0] node20044;
	wire [16-1:0] node20045;
	wire [16-1:0] node20047;
	wire [16-1:0] node20048;
	wire [16-1:0] node20052;
	wire [16-1:0] node20053;
	wire [16-1:0] node20057;
	wire [16-1:0] node20058;
	wire [16-1:0] node20059;
	wire [16-1:0] node20062;
	wire [16-1:0] node20063;
	wire [16-1:0] node20068;
	wire [16-1:0] node20069;
	wire [16-1:0] node20070;
	wire [16-1:0] node20072;
	wire [16-1:0] node20075;
	wire [16-1:0] node20076;
	wire [16-1:0] node20077;
	wire [16-1:0] node20079;
	wire [16-1:0] node20083;
	wire [16-1:0] node20086;
	wire [16-1:0] node20088;
	wire [16-1:0] node20089;
	wire [16-1:0] node20093;
	wire [16-1:0] node20094;
	wire [16-1:0] node20095;
	wire [16-1:0] node20096;
	wire [16-1:0] node20097;
	wire [16-1:0] node20098;
	wire [16-1:0] node20099;
	wire [16-1:0] node20104;
	wire [16-1:0] node20105;
	wire [16-1:0] node20106;
	wire [16-1:0] node20110;
	wire [16-1:0] node20112;
	wire [16-1:0] node20115;
	wire [16-1:0] node20116;
	wire [16-1:0] node20117;
	wire [16-1:0] node20121;
	wire [16-1:0] node20122;
	wire [16-1:0] node20126;
	wire [16-1:0] node20127;
	wire [16-1:0] node20128;
	wire [16-1:0] node20129;
	wire [16-1:0] node20132;
	wire [16-1:0] node20135;
	wire [16-1:0] node20137;
	wire [16-1:0] node20140;
	wire [16-1:0] node20141;
	wire [16-1:0] node20143;
	wire [16-1:0] node20146;
	wire [16-1:0] node20147;
	wire [16-1:0] node20151;
	wire [16-1:0] node20152;
	wire [16-1:0] node20153;
	wire [16-1:0] node20154;
	wire [16-1:0] node20155;
	wire [16-1:0] node20159;
	wire [16-1:0] node20160;
	wire [16-1:0] node20161;
	wire [16-1:0] node20164;
	wire [16-1:0] node20165;
	wire [16-1:0] node20169;
	wire [16-1:0] node20172;
	wire [16-1:0] node20173;
	wire [16-1:0] node20174;
	wire [16-1:0] node20177;
	wire [16-1:0] node20178;
	wire [16-1:0] node20180;
	wire [16-1:0] node20184;
	wire [16-1:0] node20185;
	wire [16-1:0] node20186;
	wire [16-1:0] node20190;
	wire [16-1:0] node20192;
	wire [16-1:0] node20195;
	wire [16-1:0] node20196;
	wire [16-1:0] node20197;
	wire [16-1:0] node20199;
	wire [16-1:0] node20200;
	wire [16-1:0] node20202;
	wire [16-1:0] node20206;
	wire [16-1:0] node20207;
	wire [16-1:0] node20208;
	wire [16-1:0] node20212;
	wire [16-1:0] node20215;
	wire [16-1:0] node20216;
	wire [16-1:0] node20217;
	wire [16-1:0] node20220;
	wire [16-1:0] node20222;
	wire [16-1:0] node20223;
	wire [16-1:0] node20227;
	wire [16-1:0] node20228;
	wire [16-1:0] node20232;
	wire [16-1:0] node20233;
	wire [16-1:0] node20234;
	wire [16-1:0] node20235;
	wire [16-1:0] node20236;
	wire [16-1:0] node20237;
	wire [16-1:0] node20238;
	wire [16-1:0] node20239;
	wire [16-1:0] node20243;
	wire [16-1:0] node20244;
	wire [16-1:0] node20246;
	wire [16-1:0] node20247;
	wire [16-1:0] node20251;
	wire [16-1:0] node20254;
	wire [16-1:0] node20255;
	wire [16-1:0] node20256;
	wire [16-1:0] node20257;
	wire [16-1:0] node20261;
	wire [16-1:0] node20263;
	wire [16-1:0] node20266;
	wire [16-1:0] node20267;
	wire [16-1:0] node20270;
	wire [16-1:0] node20273;
	wire [16-1:0] node20274;
	wire [16-1:0] node20275;
	wire [16-1:0] node20278;
	wire [16-1:0] node20279;
	wire [16-1:0] node20281;
	wire [16-1:0] node20284;
	wire [16-1:0] node20286;
	wire [16-1:0] node20289;
	wire [16-1:0] node20290;
	wire [16-1:0] node20291;
	wire [16-1:0] node20294;
	wire [16-1:0] node20297;
	wire [16-1:0] node20298;
	wire [16-1:0] node20301;
	wire [16-1:0] node20304;
	wire [16-1:0] node20305;
	wire [16-1:0] node20306;
	wire [16-1:0] node20308;
	wire [16-1:0] node20309;
	wire [16-1:0] node20311;
	wire [16-1:0] node20315;
	wire [16-1:0] node20316;
	wire [16-1:0] node20317;
	wire [16-1:0] node20320;
	wire [16-1:0] node20323;
	wire [16-1:0] node20324;
	wire [16-1:0] node20325;
	wire [16-1:0] node20329;
	wire [16-1:0] node20332;
	wire [16-1:0] node20333;
	wire [16-1:0] node20334;
	wire [16-1:0] node20336;
	wire [16-1:0] node20339;
	wire [16-1:0] node20340;
	wire [16-1:0] node20343;
	wire [16-1:0] node20346;
	wire [16-1:0] node20347;
	wire [16-1:0] node20348;
	wire [16-1:0] node20349;
	wire [16-1:0] node20353;
	wire [16-1:0] node20356;
	wire [16-1:0] node20358;
	wire [16-1:0] node20361;
	wire [16-1:0] node20362;
	wire [16-1:0] node20363;
	wire [16-1:0] node20364;
	wire [16-1:0] node20365;
	wire [16-1:0] node20366;
	wire [16-1:0] node20367;
	wire [16-1:0] node20370;
	wire [16-1:0] node20371;
	wire [16-1:0] node20375;
	wire [16-1:0] node20377;
	wire [16-1:0] node20380;
	wire [16-1:0] node20381;
	wire [16-1:0] node20382;
	wire [16-1:0] node20384;
	wire [16-1:0] node20388;
	wire [16-1:0] node20389;
	wire [16-1:0] node20393;
	wire [16-1:0] node20394;
	wire [16-1:0] node20395;
	wire [16-1:0] node20399;
	wire [16-1:0] node20400;
	wire [16-1:0] node20403;
	wire [16-1:0] node20404;
	wire [16-1:0] node20408;
	wire [16-1:0] node20409;
	wire [16-1:0] node20410;
	wire [16-1:0] node20412;
	wire [16-1:0] node20415;
	wire [16-1:0] node20416;
	wire [16-1:0] node20419;
	wire [16-1:0] node20422;
	wire [16-1:0] node20423;
	wire [16-1:0] node20425;
	wire [16-1:0] node20428;
	wire [16-1:0] node20429;
	wire [16-1:0] node20432;
	wire [16-1:0] node20434;
	wire [16-1:0] node20436;
	wire [16-1:0] node20439;
	wire [16-1:0] node20440;
	wire [16-1:0] node20441;
	wire [16-1:0] node20442;
	wire [16-1:0] node20443;
	wire [16-1:0] node20447;
	wire [16-1:0] node20448;
	wire [16-1:0] node20451;
	wire [16-1:0] node20454;
	wire [16-1:0] node20455;
	wire [16-1:0] node20456;
	wire [16-1:0] node20460;
	wire [16-1:0] node20462;
	wire [16-1:0] node20463;
	wire [16-1:0] node20464;
	wire [16-1:0] node20468;
	wire [16-1:0] node20471;
	wire [16-1:0] node20472;
	wire [16-1:0] node20473;
	wire [16-1:0] node20474;
	wire [16-1:0] node20477;
	wire [16-1:0] node20478;
	wire [16-1:0] node20480;
	wire [16-1:0] node20483;
	wire [16-1:0] node20486;
	wire [16-1:0] node20487;
	wire [16-1:0] node20491;
	wire [16-1:0] node20492;
	wire [16-1:0] node20493;
	wire [16-1:0] node20494;
	wire [16-1:0] node20498;
	wire [16-1:0] node20501;
	wire [16-1:0] node20502;
	wire [16-1:0] node20505;
	wire [16-1:0] node20507;
	wire [16-1:0] node20510;
	wire [16-1:0] node20511;
	wire [16-1:0] node20512;
	wire [16-1:0] node20513;
	wire [16-1:0] node20514;
	wire [16-1:0] node20516;
	wire [16-1:0] node20517;
	wire [16-1:0] node20521;
	wire [16-1:0] node20522;
	wire [16-1:0] node20523;
	wire [16-1:0] node20526;
	wire [16-1:0] node20528;
	wire [16-1:0] node20531;
	wire [16-1:0] node20532;
	wire [16-1:0] node20536;
	wire [16-1:0] node20537;
	wire [16-1:0] node20538;
	wire [16-1:0] node20539;
	wire [16-1:0] node20542;
	wire [16-1:0] node20544;
	wire [16-1:0] node20545;
	wire [16-1:0] node20549;
	wire [16-1:0] node20551;
	wire [16-1:0] node20554;
	wire [16-1:0] node20555;
	wire [16-1:0] node20557;
	wire [16-1:0] node20558;
	wire [16-1:0] node20560;
	wire [16-1:0] node20564;
	wire [16-1:0] node20565;
	wire [16-1:0] node20568;
	wire [16-1:0] node20569;
	wire [16-1:0] node20571;
	wire [16-1:0] node20575;
	wire [16-1:0] node20576;
	wire [16-1:0] node20577;
	wire [16-1:0] node20578;
	wire [16-1:0] node20581;
	wire [16-1:0] node20582;
	wire [16-1:0] node20586;
	wire [16-1:0] node20587;
	wire [16-1:0] node20589;
	wire [16-1:0] node20591;
	wire [16-1:0] node20594;
	wire [16-1:0] node20595;
	wire [16-1:0] node20597;
	wire [16-1:0] node20600;
	wire [16-1:0] node20603;
	wire [16-1:0] node20604;
	wire [16-1:0] node20606;
	wire [16-1:0] node20607;
	wire [16-1:0] node20609;
	wire [16-1:0] node20612;
	wire [16-1:0] node20615;
	wire [16-1:0] node20616;
	wire [16-1:0] node20618;
	wire [16-1:0] node20620;
	wire [16-1:0] node20623;
	wire [16-1:0] node20624;
	wire [16-1:0] node20625;
	wire [16-1:0] node20630;
	wire [16-1:0] node20631;
	wire [16-1:0] node20632;
	wire [16-1:0] node20633;
	wire [16-1:0] node20634;
	wire [16-1:0] node20635;
	wire [16-1:0] node20638;
	wire [16-1:0] node20639;
	wire [16-1:0] node20643;
	wire [16-1:0] node20644;
	wire [16-1:0] node20647;
	wire [16-1:0] node20650;
	wire [16-1:0] node20651;
	wire [16-1:0] node20652;
	wire [16-1:0] node20655;
	wire [16-1:0] node20658;
	wire [16-1:0] node20660;
	wire [16-1:0] node20663;
	wire [16-1:0] node20664;
	wire [16-1:0] node20665;
	wire [16-1:0] node20667;
	wire [16-1:0] node20669;
	wire [16-1:0] node20670;
	wire [16-1:0] node20674;
	wire [16-1:0] node20676;
	wire [16-1:0] node20677;
	wire [16-1:0] node20679;
	wire [16-1:0] node20683;
	wire [16-1:0] node20684;
	wire [16-1:0] node20686;
	wire [16-1:0] node20687;
	wire [16-1:0] node20691;
	wire [16-1:0] node20694;
	wire [16-1:0] node20695;
	wire [16-1:0] node20696;
	wire [16-1:0] node20697;
	wire [16-1:0] node20699;
	wire [16-1:0] node20702;
	wire [16-1:0] node20704;
	wire [16-1:0] node20706;
	wire [16-1:0] node20707;
	wire [16-1:0] node20711;
	wire [16-1:0] node20712;
	wire [16-1:0] node20713;
	wire [16-1:0] node20716;
	wire [16-1:0] node20717;
	wire [16-1:0] node20719;
	wire [16-1:0] node20723;
	wire [16-1:0] node20724;
	wire [16-1:0] node20725;
	wire [16-1:0] node20729;
	wire [16-1:0] node20732;
	wire [16-1:0] node20733;
	wire [16-1:0] node20734;
	wire [16-1:0] node20735;
	wire [16-1:0] node20738;
	wire [16-1:0] node20740;
	wire [16-1:0] node20742;
	wire [16-1:0] node20745;
	wire [16-1:0] node20747;
	wire [16-1:0] node20750;
	wire [16-1:0] node20751;
	wire [16-1:0] node20753;
	wire [16-1:0] node20755;
	wire [16-1:0] node20758;
	wire [16-1:0] node20759;
	wire [16-1:0] node20761;
	wire [16-1:0] node20764;
	wire [16-1:0] node20766;
	wire [16-1:0] node20768;
	wire [16-1:0] node20771;
	wire [16-1:0] node20772;
	wire [16-1:0] node20773;
	wire [16-1:0] node20774;
	wire [16-1:0] node20775;
	wire [16-1:0] node20776;
	wire [16-1:0] node20777;
	wire [16-1:0] node20778;
	wire [16-1:0] node20779;
	wire [16-1:0] node20780;
	wire [16-1:0] node20781;
	wire [16-1:0] node20782;
	wire [16-1:0] node20786;
	wire [16-1:0] node20788;
	wire [16-1:0] node20790;
	wire [16-1:0] node20793;
	wire [16-1:0] node20794;
	wire [16-1:0] node20795;
	wire [16-1:0] node20799;
	wire [16-1:0] node20802;
	wire [16-1:0] node20803;
	wire [16-1:0] node20805;
	wire [16-1:0] node20808;
	wire [16-1:0] node20809;
	wire [16-1:0] node20811;
	wire [16-1:0] node20814;
	wire [16-1:0] node20817;
	wire [16-1:0] node20818;
	wire [16-1:0] node20819;
	wire [16-1:0] node20821;
	wire [16-1:0] node20823;
	wire [16-1:0] node20826;
	wire [16-1:0] node20827;
	wire [16-1:0] node20828;
	wire [16-1:0] node20833;
	wire [16-1:0] node20835;
	wire [16-1:0] node20836;
	wire [16-1:0] node20838;
	wire [16-1:0] node20842;
	wire [16-1:0] node20843;
	wire [16-1:0] node20844;
	wire [16-1:0] node20845;
	wire [16-1:0] node20846;
	wire [16-1:0] node20848;
	wire [16-1:0] node20851;
	wire [16-1:0] node20852;
	wire [16-1:0] node20856;
	wire [16-1:0] node20857;
	wire [16-1:0] node20858;
	wire [16-1:0] node20862;
	wire [16-1:0] node20864;
	wire [16-1:0] node20865;
	wire [16-1:0] node20869;
	wire [16-1:0] node20870;
	wire [16-1:0] node20871;
	wire [16-1:0] node20874;
	wire [16-1:0] node20876;
	wire [16-1:0] node20879;
	wire [16-1:0] node20880;
	wire [16-1:0] node20882;
	wire [16-1:0] node20885;
	wire [16-1:0] node20887;
	wire [16-1:0] node20889;
	wire [16-1:0] node20892;
	wire [16-1:0] node20893;
	wire [16-1:0] node20894;
	wire [16-1:0] node20895;
	wire [16-1:0] node20899;
	wire [16-1:0] node20900;
	wire [16-1:0] node20904;
	wire [16-1:0] node20905;
	wire [16-1:0] node20906;
	wire [16-1:0] node20909;
	wire [16-1:0] node20912;
	wire [16-1:0] node20914;
	wire [16-1:0] node20917;
	wire [16-1:0] node20918;
	wire [16-1:0] node20919;
	wire [16-1:0] node20920;
	wire [16-1:0] node20921;
	wire [16-1:0] node20923;
	wire [16-1:0] node20924;
	wire [16-1:0] node20925;
	wire [16-1:0] node20930;
	wire [16-1:0] node20933;
	wire [16-1:0] node20934;
	wire [16-1:0] node20935;
	wire [16-1:0] node20937;
	wire [16-1:0] node20940;
	wire [16-1:0] node20943;
	wire [16-1:0] node20944;
	wire [16-1:0] node20946;
	wire [16-1:0] node20950;
	wire [16-1:0] node20951;
	wire [16-1:0] node20952;
	wire [16-1:0] node20953;
	wire [16-1:0] node20954;
	wire [16-1:0] node20958;
	wire [16-1:0] node20959;
	wire [16-1:0] node20961;
	wire [16-1:0] node20965;
	wire [16-1:0] node20966;
	wire [16-1:0] node20969;
	wire [16-1:0] node20970;
	wire [16-1:0] node20971;
	wire [16-1:0] node20976;
	wire [16-1:0] node20977;
	wire [16-1:0] node20978;
	wire [16-1:0] node20979;
	wire [16-1:0] node20983;
	wire [16-1:0] node20986;
	wire [16-1:0] node20988;
	wire [16-1:0] node20990;
	wire [16-1:0] node20992;
	wire [16-1:0] node20995;
	wire [16-1:0] node20996;
	wire [16-1:0] node20997;
	wire [16-1:0] node20998;
	wire [16-1:0] node20999;
	wire [16-1:0] node21000;
	wire [16-1:0] node21004;
	wire [16-1:0] node21008;
	wire [16-1:0] node21010;
	wire [16-1:0] node21012;
	wire [16-1:0] node21013;
	wire [16-1:0] node21014;
	wire [16-1:0] node21019;
	wire [16-1:0] node21020;
	wire [16-1:0] node21021;
	wire [16-1:0] node21022;
	wire [16-1:0] node21025;
	wire [16-1:0] node21028;
	wire [16-1:0] node21029;
	wire [16-1:0] node21032;
	wire [16-1:0] node21033;
	wire [16-1:0] node21037;
	wire [16-1:0] node21038;
	wire [16-1:0] node21039;
	wire [16-1:0] node21040;
	wire [16-1:0] node21045;
	wire [16-1:0] node21046;
	wire [16-1:0] node21047;
	wire [16-1:0] node21049;
	wire [16-1:0] node21053;
	wire [16-1:0] node21055;
	wire [16-1:0] node21056;
	wire [16-1:0] node21060;
	wire [16-1:0] node21061;
	wire [16-1:0] node21062;
	wire [16-1:0] node21063;
	wire [16-1:0] node21064;
	wire [16-1:0] node21065;
	wire [16-1:0] node21066;
	wire [16-1:0] node21068;
	wire [16-1:0] node21072;
	wire [16-1:0] node21074;
	wire [16-1:0] node21077;
	wire [16-1:0] node21078;
	wire [16-1:0] node21079;
	wire [16-1:0] node21082;
	wire [16-1:0] node21085;
	wire [16-1:0] node21087;
	wire [16-1:0] node21090;
	wire [16-1:0] node21091;
	wire [16-1:0] node21092;
	wire [16-1:0] node21094;
	wire [16-1:0] node21096;
	wire [16-1:0] node21100;
	wire [16-1:0] node21101;
	wire [16-1:0] node21102;
	wire [16-1:0] node21106;
	wire [16-1:0] node21107;
	wire [16-1:0] node21111;
	wire [16-1:0] node21112;
	wire [16-1:0] node21113;
	wire [16-1:0] node21114;
	wire [16-1:0] node21115;
	wire [16-1:0] node21116;
	wire [16-1:0] node21118;
	wire [16-1:0] node21122;
	wire [16-1:0] node21125;
	wire [16-1:0] node21126;
	wire [16-1:0] node21127;
	wire [16-1:0] node21131;
	wire [16-1:0] node21134;
	wire [16-1:0] node21136;
	wire [16-1:0] node21138;
	wire [16-1:0] node21141;
	wire [16-1:0] node21142;
	wire [16-1:0] node21144;
	wire [16-1:0] node21145;
	wire [16-1:0] node21147;
	wire [16-1:0] node21148;
	wire [16-1:0] node21152;
	wire [16-1:0] node21155;
	wire [16-1:0] node21156;
	wire [16-1:0] node21157;
	wire [16-1:0] node21160;
	wire [16-1:0] node21161;
	wire [16-1:0] node21165;
	wire [16-1:0] node21166;
	wire [16-1:0] node21170;
	wire [16-1:0] node21171;
	wire [16-1:0] node21172;
	wire [16-1:0] node21173;
	wire [16-1:0] node21174;
	wire [16-1:0] node21175;
	wire [16-1:0] node21178;
	wire [16-1:0] node21181;
	wire [16-1:0] node21182;
	wire [16-1:0] node21183;
	wire [16-1:0] node21188;
	wire [16-1:0] node21189;
	wire [16-1:0] node21191;
	wire [16-1:0] node21192;
	wire [16-1:0] node21196;
	wire [16-1:0] node21198;
	wire [16-1:0] node21200;
	wire [16-1:0] node21202;
	wire [16-1:0] node21205;
	wire [16-1:0] node21206;
	wire [16-1:0] node21207;
	wire [16-1:0] node21208;
	wire [16-1:0] node21211;
	wire [16-1:0] node21214;
	wire [16-1:0] node21215;
	wire [16-1:0] node21219;
	wire [16-1:0] node21220;
	wire [16-1:0] node21221;
	wire [16-1:0] node21222;
	wire [16-1:0] node21226;
	wire [16-1:0] node21227;
	wire [16-1:0] node21228;
	wire [16-1:0] node21231;
	wire [16-1:0] node21235;
	wire [16-1:0] node21236;
	wire [16-1:0] node21238;
	wire [16-1:0] node21241;
	wire [16-1:0] node21242;
	wire [16-1:0] node21246;
	wire [16-1:0] node21247;
	wire [16-1:0] node21248;
	wire [16-1:0] node21249;
	wire [16-1:0] node21250;
	wire [16-1:0] node21253;
	wire [16-1:0] node21256;
	wire [16-1:0] node21257;
	wire [16-1:0] node21260;
	wire [16-1:0] node21263;
	wire [16-1:0] node21264;
	wire [16-1:0] node21265;
	wire [16-1:0] node21266;
	wire [16-1:0] node21270;
	wire [16-1:0] node21271;
	wire [16-1:0] node21275;
	wire [16-1:0] node21277;
	wire [16-1:0] node21280;
	wire [16-1:0] node21281;
	wire [16-1:0] node21282;
	wire [16-1:0] node21283;
	wire [16-1:0] node21285;
	wire [16-1:0] node21288;
	wire [16-1:0] node21289;
	wire [16-1:0] node21294;
	wire [16-1:0] node21295;
	wire [16-1:0] node21298;
	wire [16-1:0] node21300;
	wire [16-1:0] node21302;
	wire [16-1:0] node21304;
	wire [16-1:0] node21307;
	wire [16-1:0] node21308;
	wire [16-1:0] node21309;
	wire [16-1:0] node21310;
	wire [16-1:0] node21311;
	wire [16-1:0] node21312;
	wire [16-1:0] node21314;
	wire [16-1:0] node21315;
	wire [16-1:0] node21319;
	wire [16-1:0] node21320;
	wire [16-1:0] node21321;
	wire [16-1:0] node21323;
	wire [16-1:0] node21324;
	wire [16-1:0] node21328;
	wire [16-1:0] node21329;
	wire [16-1:0] node21331;
	wire [16-1:0] node21336;
	wire [16-1:0] node21337;
	wire [16-1:0] node21339;
	wire [16-1:0] node21340;
	wire [16-1:0] node21344;
	wire [16-1:0] node21345;
	wire [16-1:0] node21346;
	wire [16-1:0] node21348;
	wire [16-1:0] node21351;
	wire [16-1:0] node21354;
	wire [16-1:0] node21357;
	wire [16-1:0] node21358;
	wire [16-1:0] node21359;
	wire [16-1:0] node21360;
	wire [16-1:0] node21361;
	wire [16-1:0] node21364;
	wire [16-1:0] node21367;
	wire [16-1:0] node21369;
	wire [16-1:0] node21370;
	wire [16-1:0] node21372;
	wire [16-1:0] node21376;
	wire [16-1:0] node21378;
	wire [16-1:0] node21379;
	wire [16-1:0] node21381;
	wire [16-1:0] node21385;
	wire [16-1:0] node21386;
	wire [16-1:0] node21387;
	wire [16-1:0] node21389;
	wire [16-1:0] node21391;
	wire [16-1:0] node21394;
	wire [16-1:0] node21396;
	wire [16-1:0] node21397;
	wire [16-1:0] node21398;
	wire [16-1:0] node21403;
	wire [16-1:0] node21404;
	wire [16-1:0] node21405;
	wire [16-1:0] node21409;
	wire [16-1:0] node21411;
	wire [16-1:0] node21414;
	wire [16-1:0] node21415;
	wire [16-1:0] node21416;
	wire [16-1:0] node21417;
	wire [16-1:0] node21418;
	wire [16-1:0] node21421;
	wire [16-1:0] node21422;
	wire [16-1:0] node21424;
	wire [16-1:0] node21428;
	wire [16-1:0] node21429;
	wire [16-1:0] node21432;
	wire [16-1:0] node21433;
	wire [16-1:0] node21434;
	wire [16-1:0] node21438;
	wire [16-1:0] node21441;
	wire [16-1:0] node21442;
	wire [16-1:0] node21443;
	wire [16-1:0] node21445;
	wire [16-1:0] node21448;
	wire [16-1:0] node21449;
	wire [16-1:0] node21452;
	wire [16-1:0] node21454;
	wire [16-1:0] node21457;
	wire [16-1:0] node21458;
	wire [16-1:0] node21459;
	wire [16-1:0] node21462;
	wire [16-1:0] node21465;
	wire [16-1:0] node21467;
	wire [16-1:0] node21470;
	wire [16-1:0] node21471;
	wire [16-1:0] node21472;
	wire [16-1:0] node21473;
	wire [16-1:0] node21474;
	wire [16-1:0] node21475;
	wire [16-1:0] node21479;
	wire [16-1:0] node21481;
	wire [16-1:0] node21482;
	wire [16-1:0] node21487;
	wire [16-1:0] node21488;
	wire [16-1:0] node21490;
	wire [16-1:0] node21492;
	wire [16-1:0] node21495;
	wire [16-1:0] node21496;
	wire [16-1:0] node21497;
	wire [16-1:0] node21502;
	wire [16-1:0] node21503;
	wire [16-1:0] node21504;
	wire [16-1:0] node21505;
	wire [16-1:0] node21508;
	wire [16-1:0] node21511;
	wire [16-1:0] node21512;
	wire [16-1:0] node21515;
	wire [16-1:0] node21518;
	wire [16-1:0] node21519;
	wire [16-1:0] node21520;
	wire [16-1:0] node21521;
	wire [16-1:0] node21525;
	wire [16-1:0] node21528;
	wire [16-1:0] node21529;
	wire [16-1:0] node21531;
	wire [16-1:0] node21532;
	wire [16-1:0] node21536;
	wire [16-1:0] node21539;
	wire [16-1:0] node21540;
	wire [16-1:0] node21541;
	wire [16-1:0] node21542;
	wire [16-1:0] node21543;
	wire [16-1:0] node21544;
	wire [16-1:0] node21546;
	wire [16-1:0] node21548;
	wire [16-1:0] node21551;
	wire [16-1:0] node21552;
	wire [16-1:0] node21556;
	wire [16-1:0] node21557;
	wire [16-1:0] node21558;
	wire [16-1:0] node21562;
	wire [16-1:0] node21563;
	wire [16-1:0] node21565;
	wire [16-1:0] node21566;
	wire [16-1:0] node21570;
	wire [16-1:0] node21573;
	wire [16-1:0] node21574;
	wire [16-1:0] node21575;
	wire [16-1:0] node21577;
	wire [16-1:0] node21578;
	wire [16-1:0] node21580;
	wire [16-1:0] node21585;
	wire [16-1:0] node21586;
	wire [16-1:0] node21589;
	wire [16-1:0] node21592;
	wire [16-1:0] node21593;
	wire [16-1:0] node21594;
	wire [16-1:0] node21595;
	wire [16-1:0] node21596;
	wire [16-1:0] node21598;
	wire [16-1:0] node21602;
	wire [16-1:0] node21603;
	wire [16-1:0] node21605;
	wire [16-1:0] node21606;
	wire [16-1:0] node21610;
	wire [16-1:0] node21612;
	wire [16-1:0] node21615;
	wire [16-1:0] node21616;
	wire [16-1:0] node21617;
	wire [16-1:0] node21618;
	wire [16-1:0] node21620;
	wire [16-1:0] node21624;
	wire [16-1:0] node21626;
	wire [16-1:0] node21629;
	wire [16-1:0] node21631;
	wire [16-1:0] node21634;
	wire [16-1:0] node21635;
	wire [16-1:0] node21636;
	wire [16-1:0] node21637;
	wire [16-1:0] node21642;
	wire [16-1:0] node21643;
	wire [16-1:0] node21645;
	wire [16-1:0] node21646;
	wire [16-1:0] node21648;
	wire [16-1:0] node21652;
	wire [16-1:0] node21654;
	wire [16-1:0] node21657;
	wire [16-1:0] node21658;
	wire [16-1:0] node21659;
	wire [16-1:0] node21660;
	wire [16-1:0] node21661;
	wire [16-1:0] node21662;
	wire [16-1:0] node21665;
	wire [16-1:0] node21667;
	wire [16-1:0] node21668;
	wire [16-1:0] node21672;
	wire [16-1:0] node21673;
	wire [16-1:0] node21674;
	wire [16-1:0] node21679;
	wire [16-1:0] node21680;
	wire [16-1:0] node21681;
	wire [16-1:0] node21685;
	wire [16-1:0] node21686;
	wire [16-1:0] node21687;
	wire [16-1:0] node21691;
	wire [16-1:0] node21694;
	wire [16-1:0] node21695;
	wire [16-1:0] node21696;
	wire [16-1:0] node21697;
	wire [16-1:0] node21700;
	wire [16-1:0] node21702;
	wire [16-1:0] node21703;
	wire [16-1:0] node21707;
	wire [16-1:0] node21708;
	wire [16-1:0] node21711;
	wire [16-1:0] node21712;
	wire [16-1:0] node21714;
	wire [16-1:0] node21717;
	wire [16-1:0] node21720;
	wire [16-1:0] node21721;
	wire [16-1:0] node21722;
	wire [16-1:0] node21726;
	wire [16-1:0] node21727;
	wire [16-1:0] node21728;
	wire [16-1:0] node21732;
	wire [16-1:0] node21735;
	wire [16-1:0] node21736;
	wire [16-1:0] node21737;
	wire [16-1:0] node21738;
	wire [16-1:0] node21740;
	wire [16-1:0] node21743;
	wire [16-1:0] node21745;
	wire [16-1:0] node21748;
	wire [16-1:0] node21749;
	wire [16-1:0] node21750;
	wire [16-1:0] node21753;
	wire [16-1:0] node21754;
	wire [16-1:0] node21758;
	wire [16-1:0] node21759;
	wire [16-1:0] node21762;
	wire [16-1:0] node21765;
	wire [16-1:0] node21766;
	wire [16-1:0] node21767;
	wire [16-1:0] node21769;
	wire [16-1:0] node21772;
	wire [16-1:0] node21775;
	wire [16-1:0] node21776;
	wire [16-1:0] node21778;
	wire [16-1:0] node21781;
	wire [16-1:0] node21783;
	wire [16-1:0] node21786;
	wire [16-1:0] node21787;
	wire [16-1:0] node21788;
	wire [16-1:0] node21789;
	wire [16-1:0] node21790;
	wire [16-1:0] node21791;
	wire [16-1:0] node21792;
	wire [16-1:0] node21793;
	wire [16-1:0] node21795;
	wire [16-1:0] node21796;
	wire [16-1:0] node21800;
	wire [16-1:0] node21801;
	wire [16-1:0] node21802;
	wire [16-1:0] node21803;
	wire [16-1:0] node21808;
	wire [16-1:0] node21809;
	wire [16-1:0] node21810;
	wire [16-1:0] node21815;
	wire [16-1:0] node21816;
	wire [16-1:0] node21817;
	wire [16-1:0] node21819;
	wire [16-1:0] node21820;
	wire [16-1:0] node21824;
	wire [16-1:0] node21827;
	wire [16-1:0] node21828;
	wire [16-1:0] node21830;
	wire [16-1:0] node21831;
	wire [16-1:0] node21836;
	wire [16-1:0] node21837;
	wire [16-1:0] node21838;
	wire [16-1:0] node21841;
	wire [16-1:0] node21842;
	wire [16-1:0] node21843;
	wire [16-1:0] node21846;
	wire [16-1:0] node21850;
	wire [16-1:0] node21851;
	wire [16-1:0] node21852;
	wire [16-1:0] node21854;
	wire [16-1:0] node21855;
	wire [16-1:0] node21860;
	wire [16-1:0] node21863;
	wire [16-1:0] node21864;
	wire [16-1:0] node21865;
	wire [16-1:0] node21867;
	wire [16-1:0] node21868;
	wire [16-1:0] node21869;
	wire [16-1:0] node21872;
	wire [16-1:0] node21876;
	wire [16-1:0] node21877;
	wire [16-1:0] node21878;
	wire [16-1:0] node21881;
	wire [16-1:0] node21884;
	wire [16-1:0] node21885;
	wire [16-1:0] node21887;
	wire [16-1:0] node21888;
	wire [16-1:0] node21892;
	wire [16-1:0] node21895;
	wire [16-1:0] node21896;
	wire [16-1:0] node21897;
	wire [16-1:0] node21899;
	wire [16-1:0] node21900;
	wire [16-1:0] node21904;
	wire [16-1:0] node21905;
	wire [16-1:0] node21908;
	wire [16-1:0] node21911;
	wire [16-1:0] node21912;
	wire [16-1:0] node21914;
	wire [16-1:0] node21917;
	wire [16-1:0] node21918;
	wire [16-1:0] node21922;
	wire [16-1:0] node21923;
	wire [16-1:0] node21924;
	wire [16-1:0] node21925;
	wire [16-1:0] node21926;
	wire [16-1:0] node21927;
	wire [16-1:0] node21930;
	wire [16-1:0] node21931;
	wire [16-1:0] node21932;
	wire [16-1:0] node21936;
	wire [16-1:0] node21939;
	wire [16-1:0] node21941;
	wire [16-1:0] node21944;
	wire [16-1:0] node21945;
	wire [16-1:0] node21946;
	wire [16-1:0] node21949;
	wire [16-1:0] node21952;
	wire [16-1:0] node21953;
	wire [16-1:0] node21955;
	wire [16-1:0] node21959;
	wire [16-1:0] node21960;
	wire [16-1:0] node21961;
	wire [16-1:0] node21963;
	wire [16-1:0] node21966;
	wire [16-1:0] node21967;
	wire [16-1:0] node21971;
	wire [16-1:0] node21972;
	wire [16-1:0] node21973;
	wire [16-1:0] node21974;
	wire [16-1:0] node21979;
	wire [16-1:0] node21980;
	wire [16-1:0] node21981;
	wire [16-1:0] node21986;
	wire [16-1:0] node21987;
	wire [16-1:0] node21988;
	wire [16-1:0] node21989;
	wire [16-1:0] node21990;
	wire [16-1:0] node21993;
	wire [16-1:0] node21995;
	wire [16-1:0] node21998;
	wire [16-1:0] node21999;
	wire [16-1:0] node22000;
	wire [16-1:0] node22005;
	wire [16-1:0] node22006;
	wire [16-1:0] node22007;
	wire [16-1:0] node22008;
	wire [16-1:0] node22012;
	wire [16-1:0] node22015;
	wire [16-1:0] node22017;
	wire [16-1:0] node22020;
	wire [16-1:0] node22021;
	wire [16-1:0] node22022;
	wire [16-1:0] node22023;
	wire [16-1:0] node22025;
	wire [16-1:0] node22029;
	wire [16-1:0] node22031;
	wire [16-1:0] node22034;
	wire [16-1:0] node22035;
	wire [16-1:0] node22036;
	wire [16-1:0] node22037;
	wire [16-1:0] node22041;
	wire [16-1:0] node22042;
	wire [16-1:0] node22043;
	wire [16-1:0] node22046;
	wire [16-1:0] node22050;
	wire [16-1:0] node22051;
	wire [16-1:0] node22054;
	wire [16-1:0] node22055;
	wire [16-1:0] node22057;
	wire [16-1:0] node22061;
	wire [16-1:0] node22062;
	wire [16-1:0] node22063;
	wire [16-1:0] node22064;
	wire [16-1:0] node22065;
	wire [16-1:0] node22066;
	wire [16-1:0] node22067;
	wire [16-1:0] node22068;
	wire [16-1:0] node22072;
	wire [16-1:0] node22076;
	wire [16-1:0] node22077;
	wire [16-1:0] node22078;
	wire [16-1:0] node22080;
	wire [16-1:0] node22083;
	wire [16-1:0] node22086;
	wire [16-1:0] node22087;
	wire [16-1:0] node22090;
	wire [16-1:0] node22092;
	wire [16-1:0] node22095;
	wire [16-1:0] node22096;
	wire [16-1:0] node22097;
	wire [16-1:0] node22098;
	wire [16-1:0] node22101;
	wire [16-1:0] node22102;
	wire [16-1:0] node22107;
	wire [16-1:0] node22108;
	wire [16-1:0] node22109;
	wire [16-1:0] node22111;
	wire [16-1:0] node22114;
	wire [16-1:0] node22115;
	wire [16-1:0] node22119;
	wire [16-1:0] node22120;
	wire [16-1:0] node22123;
	wire [16-1:0] node22126;
	wire [16-1:0] node22127;
	wire [16-1:0] node22128;
	wire [16-1:0] node22129;
	wire [16-1:0] node22130;
	wire [16-1:0] node22134;
	wire [16-1:0] node22135;
	wire [16-1:0] node22139;
	wire [16-1:0] node22140;
	wire [16-1:0] node22142;
	wire [16-1:0] node22143;
	wire [16-1:0] node22144;
	wire [16-1:0] node22149;
	wire [16-1:0] node22151;
	wire [16-1:0] node22154;
	wire [16-1:0] node22155;
	wire [16-1:0] node22157;
	wire [16-1:0] node22158;
	wire [16-1:0] node22161;
	wire [16-1:0] node22164;
	wire [16-1:0] node22165;
	wire [16-1:0] node22166;
	wire [16-1:0] node22169;
	wire [16-1:0] node22170;
	wire [16-1:0] node22174;
	wire [16-1:0] node22175;
	wire [16-1:0] node22178;
	wire [16-1:0] node22179;
	wire [16-1:0] node22183;
	wire [16-1:0] node22184;
	wire [16-1:0] node22185;
	wire [16-1:0] node22186;
	wire [16-1:0] node22187;
	wire [16-1:0] node22189;
	wire [16-1:0] node22190;
	wire [16-1:0] node22194;
	wire [16-1:0] node22195;
	wire [16-1:0] node22197;
	wire [16-1:0] node22201;
	wire [16-1:0] node22202;
	wire [16-1:0] node22203;
	wire [16-1:0] node22206;
	wire [16-1:0] node22207;
	wire [16-1:0] node22212;
	wire [16-1:0] node22213;
	wire [16-1:0] node22214;
	wire [16-1:0] node22215;
	wire [16-1:0] node22217;
	wire [16-1:0] node22220;
	wire [16-1:0] node22221;
	wire [16-1:0] node22223;
	wire [16-1:0] node22227;
	wire [16-1:0] node22230;
	wire [16-1:0] node22231;
	wire [16-1:0] node22232;
	wire [16-1:0] node22235;
	wire [16-1:0] node22238;
	wire [16-1:0] node22241;
	wire [16-1:0] node22242;
	wire [16-1:0] node22243;
	wire [16-1:0] node22244;
	wire [16-1:0] node22245;
	wire [16-1:0] node22247;
	wire [16-1:0] node22250;
	wire [16-1:0] node22251;
	wire [16-1:0] node22253;
	wire [16-1:0] node22257;
	wire [16-1:0] node22258;
	wire [16-1:0] node22261;
	wire [16-1:0] node22262;
	wire [16-1:0] node22266;
	wire [16-1:0] node22268;
	wire [16-1:0] node22269;
	wire [16-1:0] node22270;
	wire [16-1:0] node22273;
	wire [16-1:0] node22274;
	wire [16-1:0] node22278;
	wire [16-1:0] node22281;
	wire [16-1:0] node22282;
	wire [16-1:0] node22283;
	wire [16-1:0] node22284;
	wire [16-1:0] node22287;
	wire [16-1:0] node22288;
	wire [16-1:0] node22290;
	wire [16-1:0] node22293;
	wire [16-1:0] node22294;
	wire [16-1:0] node22299;
	wire [16-1:0] node22300;
	wire [16-1:0] node22301;
	wire [16-1:0] node22302;
	wire [16-1:0] node22305;
	wire [16-1:0] node22306;
	wire [16-1:0] node22310;
	wire [16-1:0] node22311;
	wire [16-1:0] node22315;
	wire [16-1:0] node22316;
	wire [16-1:0] node22319;
	wire [16-1:0] node22321;
	wire [16-1:0] node22322;
	wire [16-1:0] node22326;
	wire [16-1:0] node22327;
	wire [16-1:0] node22328;
	wire [16-1:0] node22329;
	wire [16-1:0] node22330;
	wire [16-1:0] node22331;
	wire [16-1:0] node22332;
	wire [16-1:0] node22333;
	wire [16-1:0] node22336;
	wire [16-1:0] node22338;
	wire [16-1:0] node22341;
	wire [16-1:0] node22342;
	wire [16-1:0] node22345;
	wire [16-1:0] node22348;
	wire [16-1:0] node22349;
	wire [16-1:0] node22350;
	wire [16-1:0] node22351;
	wire [16-1:0] node22353;
	wire [16-1:0] node22357;
	wire [16-1:0] node22360;
	wire [16-1:0] node22361;
	wire [16-1:0] node22365;
	wire [16-1:0] node22366;
	wire [16-1:0] node22368;
	wire [16-1:0] node22369;
	wire [16-1:0] node22372;
	wire [16-1:0] node22374;
	wire [16-1:0] node22377;
	wire [16-1:0] node22378;
	wire [16-1:0] node22379;
	wire [16-1:0] node22382;
	wire [16-1:0] node22384;
	wire [16-1:0] node22388;
	wire [16-1:0] node22389;
	wire [16-1:0] node22390;
	wire [16-1:0] node22391;
	wire [16-1:0] node22392;
	wire [16-1:0] node22393;
	wire [16-1:0] node22397;
	wire [16-1:0] node22400;
	wire [16-1:0] node22401;
	wire [16-1:0] node22402;
	wire [16-1:0] node22404;
	wire [16-1:0] node22408;
	wire [16-1:0] node22410;
	wire [16-1:0] node22413;
	wire [16-1:0] node22414;
	wire [16-1:0] node22415;
	wire [16-1:0] node22418;
	wire [16-1:0] node22421;
	wire [16-1:0] node22422;
	wire [16-1:0] node22424;
	wire [16-1:0] node22425;
	wire [16-1:0] node22430;
	wire [16-1:0] node22431;
	wire [16-1:0] node22432;
	wire [16-1:0] node22433;
	wire [16-1:0] node22436;
	wire [16-1:0] node22440;
	wire [16-1:0] node22441;
	wire [16-1:0] node22443;
	wire [16-1:0] node22446;
	wire [16-1:0] node22447;
	wire [16-1:0] node22450;
	wire [16-1:0] node22453;
	wire [16-1:0] node22454;
	wire [16-1:0] node22455;
	wire [16-1:0] node22456;
	wire [16-1:0] node22457;
	wire [16-1:0] node22460;
	wire [16-1:0] node22461;
	wire [16-1:0] node22463;
	wire [16-1:0] node22466;
	wire [16-1:0] node22469;
	wire [16-1:0] node22470;
	wire [16-1:0] node22471;
	wire [16-1:0] node22472;
	wire [16-1:0] node22474;
	wire [16-1:0] node22479;
	wire [16-1:0] node22480;
	wire [16-1:0] node22482;
	wire [16-1:0] node22483;
	wire [16-1:0] node22487;
	wire [16-1:0] node22490;
	wire [16-1:0] node22491;
	wire [16-1:0] node22492;
	wire [16-1:0] node22493;
	wire [16-1:0] node22494;
	wire [16-1:0] node22498;
	wire [16-1:0] node22500;
	wire [16-1:0] node22503;
	wire [16-1:0] node22504;
	wire [16-1:0] node22507;
	wire [16-1:0] node22509;
	wire [16-1:0] node22512;
	wire [16-1:0] node22513;
	wire [16-1:0] node22515;
	wire [16-1:0] node22517;
	wire [16-1:0] node22520;
	wire [16-1:0] node22521;
	wire [16-1:0] node22522;
	wire [16-1:0] node22524;
	wire [16-1:0] node22528;
	wire [16-1:0] node22530;
	wire [16-1:0] node22531;
	wire [16-1:0] node22535;
	wire [16-1:0] node22536;
	wire [16-1:0] node22537;
	wire [16-1:0] node22539;
	wire [16-1:0] node22541;
	wire [16-1:0] node22542;
	wire [16-1:0] node22546;
	wire [16-1:0] node22547;
	wire [16-1:0] node22549;
	wire [16-1:0] node22550;
	wire [16-1:0] node22552;
	wire [16-1:0] node22556;
	wire [16-1:0] node22558;
	wire [16-1:0] node22560;
	wire [16-1:0] node22563;
	wire [16-1:0] node22564;
	wire [16-1:0] node22565;
	wire [16-1:0] node22568;
	wire [16-1:0] node22569;
	wire [16-1:0] node22571;
	wire [16-1:0] node22575;
	wire [16-1:0] node22576;
	wire [16-1:0] node22577;
	wire [16-1:0] node22579;
	wire [16-1:0] node22583;
	wire [16-1:0] node22585;
	wire [16-1:0] node22587;
	wire [16-1:0] node22590;
	wire [16-1:0] node22591;
	wire [16-1:0] node22592;
	wire [16-1:0] node22593;
	wire [16-1:0] node22594;
	wire [16-1:0] node22595;
	wire [16-1:0] node22596;
	wire [16-1:0] node22597;
	wire [16-1:0] node22598;
	wire [16-1:0] node22603;
	wire [16-1:0] node22606;
	wire [16-1:0] node22607;
	wire [16-1:0] node22611;
	wire [16-1:0] node22612;
	wire [16-1:0] node22613;
	wire [16-1:0] node22617;
	wire [16-1:0] node22618;
	wire [16-1:0] node22620;
	wire [16-1:0] node22623;
	wire [16-1:0] node22626;
	wire [16-1:0] node22627;
	wire [16-1:0] node22628;
	wire [16-1:0] node22629;
	wire [16-1:0] node22633;
	wire [16-1:0] node22634;
	wire [16-1:0] node22635;
	wire [16-1:0] node22637;
	wire [16-1:0] node22641;
	wire [16-1:0] node22644;
	wire [16-1:0] node22645;
	wire [16-1:0] node22647;
	wire [16-1:0] node22650;
	wire [16-1:0] node22652;
	wire [16-1:0] node22654;
	wire [16-1:0] node22657;
	wire [16-1:0] node22658;
	wire [16-1:0] node22659;
	wire [16-1:0] node22660;
	wire [16-1:0] node22661;
	wire [16-1:0] node22664;
	wire [16-1:0] node22667;
	wire [16-1:0] node22668;
	wire [16-1:0] node22670;
	wire [16-1:0] node22672;
	wire [16-1:0] node22675;
	wire [16-1:0] node22676;
	wire [16-1:0] node22680;
	wire [16-1:0] node22681;
	wire [16-1:0] node22683;
	wire [16-1:0] node22686;
	wire [16-1:0] node22687;
	wire [16-1:0] node22688;
	wire [16-1:0] node22690;
	wire [16-1:0] node22693;
	wire [16-1:0] node22694;
	wire [16-1:0] node22699;
	wire [16-1:0] node22700;
	wire [16-1:0] node22701;
	wire [16-1:0] node22703;
	wire [16-1:0] node22705;
	wire [16-1:0] node22708;
	wire [16-1:0] node22709;
	wire [16-1:0] node22711;
	wire [16-1:0] node22714;
	wire [16-1:0] node22716;
	wire [16-1:0] node22717;
	wire [16-1:0] node22721;
	wire [16-1:0] node22722;
	wire [16-1:0] node22723;
	wire [16-1:0] node22727;
	wire [16-1:0] node22728;
	wire [16-1:0] node22730;
	wire [16-1:0] node22734;
	wire [16-1:0] node22735;
	wire [16-1:0] node22736;
	wire [16-1:0] node22737;
	wire [16-1:0] node22738;
	wire [16-1:0] node22739;
	wire [16-1:0] node22742;
	wire [16-1:0] node22744;
	wire [16-1:0] node22747;
	wire [16-1:0] node22748;
	wire [16-1:0] node22749;
	wire [16-1:0] node22753;
	wire [16-1:0] node22754;
	wire [16-1:0] node22758;
	wire [16-1:0] node22759;
	wire [16-1:0] node22760;
	wire [16-1:0] node22763;
	wire [16-1:0] node22764;
	wire [16-1:0] node22766;
	wire [16-1:0] node22769;
	wire [16-1:0] node22772;
	wire [16-1:0] node22774;
	wire [16-1:0] node22777;
	wire [16-1:0] node22778;
	wire [16-1:0] node22779;
	wire [16-1:0] node22781;
	wire [16-1:0] node22782;
	wire [16-1:0] node22786;
	wire [16-1:0] node22788;
	wire [16-1:0] node22791;
	wire [16-1:0] node22792;
	wire [16-1:0] node22793;
	wire [16-1:0] node22794;
	wire [16-1:0] node22798;
	wire [16-1:0] node22801;
	wire [16-1:0] node22802;
	wire [16-1:0] node22805;
	wire [16-1:0] node22808;
	wire [16-1:0] node22809;
	wire [16-1:0] node22810;
	wire [16-1:0] node22811;
	wire [16-1:0] node22812;
	wire [16-1:0] node22813;
	wire [16-1:0] node22817;
	wire [16-1:0] node22819;
	wire [16-1:0] node22822;
	wire [16-1:0] node22823;
	wire [16-1:0] node22824;
	wire [16-1:0] node22826;
	wire [16-1:0] node22830;
	wire [16-1:0] node22831;
	wire [16-1:0] node22833;
	wire [16-1:0] node22837;
	wire [16-1:0] node22838;
	wire [16-1:0] node22839;
	wire [16-1:0] node22841;
	wire [16-1:0] node22843;
	wire [16-1:0] node22846;
	wire [16-1:0] node22847;
	wire [16-1:0] node22851;
	wire [16-1:0] node22852;
	wire [16-1:0] node22854;
	wire [16-1:0] node22856;
	wire [16-1:0] node22860;
	wire [16-1:0] node22861;
	wire [16-1:0] node22862;
	wire [16-1:0] node22864;
	wire [16-1:0] node22865;
	wire [16-1:0] node22870;
	wire [16-1:0] node22871;
	wire [16-1:0] node22873;
	wire [16-1:0] node22876;
	wire [16-1:0] node22877;
	wire [16-1:0] node22878;
	wire [16-1:0] node22880;
	wire [16-1:0] node22884;
	wire [16-1:0] node22885;
	wire [16-1:0] node22889;
	wire [16-1:0] node22890;
	wire [16-1:0] node22891;
	wire [16-1:0] node22892;
	wire [16-1:0] node22893;
	wire [16-1:0] node22894;
	wire [16-1:0] node22895;
	wire [16-1:0] node22896;
	wire [16-1:0] node22897;
	wire [16-1:0] node22898;
	wire [16-1:0] node22901;
	wire [16-1:0] node22903;
	wire [16-1:0] node22904;
	wire [16-1:0] node22908;
	wire [16-1:0] node22909;
	wire [16-1:0] node22911;
	wire [16-1:0] node22914;
	wire [16-1:0] node22917;
	wire [16-1:0] node22918;
	wire [16-1:0] node22920;
	wire [16-1:0] node22923;
	wire [16-1:0] node22924;
	wire [16-1:0] node22925;
	wire [16-1:0] node22927;
	wire [16-1:0] node22932;
	wire [16-1:0] node22933;
	wire [16-1:0] node22934;
	wire [16-1:0] node22935;
	wire [16-1:0] node22937;
	wire [16-1:0] node22940;
	wire [16-1:0] node22941;
	wire [16-1:0] node22946;
	wire [16-1:0] node22947;
	wire [16-1:0] node22948;
	wire [16-1:0] node22950;
	wire [16-1:0] node22953;
	wire [16-1:0] node22956;
	wire [16-1:0] node22957;
	wire [16-1:0] node22960;
	wire [16-1:0] node22963;
	wire [16-1:0] node22964;
	wire [16-1:0] node22965;
	wire [16-1:0] node22966;
	wire [16-1:0] node22967;
	wire [16-1:0] node22971;
	wire [16-1:0] node22972;
	wire [16-1:0] node22974;
	wire [16-1:0] node22975;
	wire [16-1:0] node22979;
	wire [16-1:0] node22981;
	wire [16-1:0] node22984;
	wire [16-1:0] node22985;
	wire [16-1:0] node22986;
	wire [16-1:0] node22990;
	wire [16-1:0] node22992;
	wire [16-1:0] node22993;
	wire [16-1:0] node22997;
	wire [16-1:0] node22998;
	wire [16-1:0] node22999;
	wire [16-1:0] node23001;
	wire [16-1:0] node23004;
	wire [16-1:0] node23007;
	wire [16-1:0] node23008;
	wire [16-1:0] node23009;
	wire [16-1:0] node23012;
	wire [16-1:0] node23015;
	wire [16-1:0] node23017;
	wire [16-1:0] node23020;
	wire [16-1:0] node23021;
	wire [16-1:0] node23022;
	wire [16-1:0] node23023;
	wire [16-1:0] node23024;
	wire [16-1:0] node23025;
	wire [16-1:0] node23026;
	wire [16-1:0] node23029;
	wire [16-1:0] node23032;
	wire [16-1:0] node23033;
	wire [16-1:0] node23037;
	wire [16-1:0] node23038;
	wire [16-1:0] node23039;
	wire [16-1:0] node23044;
	wire [16-1:0] node23045;
	wire [16-1:0] node23046;
	wire [16-1:0] node23048;
	wire [16-1:0] node23050;
	wire [16-1:0] node23054;
	wire [16-1:0] node23056;
	wire [16-1:0] node23057;
	wire [16-1:0] node23061;
	wire [16-1:0] node23062;
	wire [16-1:0] node23063;
	wire [16-1:0] node23064;
	wire [16-1:0] node23065;
	wire [16-1:0] node23069;
	wire [16-1:0] node23072;
	wire [16-1:0] node23075;
	wire [16-1:0] node23076;
	wire [16-1:0] node23077;
	wire [16-1:0] node23081;
	wire [16-1:0] node23082;
	wire [16-1:0] node23085;
	wire [16-1:0] node23088;
	wire [16-1:0] node23089;
	wire [16-1:0] node23090;
	wire [16-1:0] node23091;
	wire [16-1:0] node23093;
	wire [16-1:0] node23096;
	wire [16-1:0] node23097;
	wire [16-1:0] node23099;
	wire [16-1:0] node23103;
	wire [16-1:0] node23104;
	wire [16-1:0] node23106;
	wire [16-1:0] node23108;
	wire [16-1:0] node23111;
	wire [16-1:0] node23112;
	wire [16-1:0] node23113;
	wire [16-1:0] node23117;
	wire [16-1:0] node23119;
	wire [16-1:0] node23122;
	wire [16-1:0] node23123;
	wire [16-1:0] node23124;
	wire [16-1:0] node23125;
	wire [16-1:0] node23128;
	wire [16-1:0] node23131;
	wire [16-1:0] node23132;
	wire [16-1:0] node23134;
	wire [16-1:0] node23135;
	wire [16-1:0] node23140;
	wire [16-1:0] node23141;
	wire [16-1:0] node23142;
	wire [16-1:0] node23146;
	wire [16-1:0] node23147;
	wire [16-1:0] node23148;
	wire [16-1:0] node23153;
	wire [16-1:0] node23154;
	wire [16-1:0] node23155;
	wire [16-1:0] node23156;
	wire [16-1:0] node23157;
	wire [16-1:0] node23158;
	wire [16-1:0] node23159;
	wire [16-1:0] node23160;
	wire [16-1:0] node23162;
	wire [16-1:0] node23167;
	wire [16-1:0] node23168;
	wire [16-1:0] node23170;
	wire [16-1:0] node23173;
	wire [16-1:0] node23175;
	wire [16-1:0] node23178;
	wire [16-1:0] node23179;
	wire [16-1:0] node23182;
	wire [16-1:0] node23183;
	wire [16-1:0] node23185;
	wire [16-1:0] node23189;
	wire [16-1:0] node23190;
	wire [16-1:0] node23191;
	wire [16-1:0] node23192;
	wire [16-1:0] node23193;
	wire [16-1:0] node23197;
	wire [16-1:0] node23199;
	wire [16-1:0] node23202;
	wire [16-1:0] node23203;
	wire [16-1:0] node23204;
	wire [16-1:0] node23208;
	wire [16-1:0] node23209;
	wire [16-1:0] node23211;
	wire [16-1:0] node23215;
	wire [16-1:0] node23216;
	wire [16-1:0] node23217;
	wire [16-1:0] node23220;
	wire [16-1:0] node23223;
	wire [16-1:0] node23224;
	wire [16-1:0] node23227;
	wire [16-1:0] node23229;
	wire [16-1:0] node23232;
	wire [16-1:0] node23233;
	wire [16-1:0] node23234;
	wire [16-1:0] node23235;
	wire [16-1:0] node23238;
	wire [16-1:0] node23241;
	wire [16-1:0] node23242;
	wire [16-1:0] node23244;
	wire [16-1:0] node23247;
	wire [16-1:0] node23249;
	wire [16-1:0] node23252;
	wire [16-1:0] node23253;
	wire [16-1:0] node23254;
	wire [16-1:0] node23255;
	wire [16-1:0] node23258;
	wire [16-1:0] node23261;
	wire [16-1:0] node23262;
	wire [16-1:0] node23265;
	wire [16-1:0] node23268;
	wire [16-1:0] node23269;
	wire [16-1:0] node23271;
	wire [16-1:0] node23272;
	wire [16-1:0] node23274;
	wire [16-1:0] node23278;
	wire [16-1:0] node23280;
	wire [16-1:0] node23281;
	wire [16-1:0] node23285;
	wire [16-1:0] node23286;
	wire [16-1:0] node23287;
	wire [16-1:0] node23288;
	wire [16-1:0] node23289;
	wire [16-1:0] node23291;
	wire [16-1:0] node23292;
	wire [16-1:0] node23297;
	wire [16-1:0] node23298;
	wire [16-1:0] node23300;
	wire [16-1:0] node23302;
	wire [16-1:0] node23305;
	wire [16-1:0] node23306;
	wire [16-1:0] node23308;
	wire [16-1:0] node23311;
	wire [16-1:0] node23314;
	wire [16-1:0] node23315;
	wire [16-1:0] node23316;
	wire [16-1:0] node23317;
	wire [16-1:0] node23319;
	wire [16-1:0] node23323;
	wire [16-1:0] node23324;
	wire [16-1:0] node23326;
	wire [16-1:0] node23327;
	wire [16-1:0] node23331;
	wire [16-1:0] node23332;
	wire [16-1:0] node23336;
	wire [16-1:0] node23337;
	wire [16-1:0] node23338;
	wire [16-1:0] node23341;
	wire [16-1:0] node23343;
	wire [16-1:0] node23344;
	wire [16-1:0] node23348;
	wire [16-1:0] node23349;
	wire [16-1:0] node23353;
	wire [16-1:0] node23354;
	wire [16-1:0] node23355;
	wire [16-1:0] node23356;
	wire [16-1:0] node23357;
	wire [16-1:0] node23358;
	wire [16-1:0] node23362;
	wire [16-1:0] node23363;
	wire [16-1:0] node23365;
	wire [16-1:0] node23369;
	wire [16-1:0] node23371;
	wire [16-1:0] node23372;
	wire [16-1:0] node23376;
	wire [16-1:0] node23377;
	wire [16-1:0] node23378;
	wire [16-1:0] node23379;
	wire [16-1:0] node23383;
	wire [16-1:0] node23384;
	wire [16-1:0] node23386;
	wire [16-1:0] node23390;
	wire [16-1:0] node23391;
	wire [16-1:0] node23394;
	wire [16-1:0] node23397;
	wire [16-1:0] node23398;
	wire [16-1:0] node23399;
	wire [16-1:0] node23400;
	wire [16-1:0] node23403;
	wire [16-1:0] node23404;
	wire [16-1:0] node23406;
	wire [16-1:0] node23410;
	wire [16-1:0] node23411;
	wire [16-1:0] node23414;
	wire [16-1:0] node23417;
	wire [16-1:0] node23418;
	wire [16-1:0] node23419;
	wire [16-1:0] node23422;
	wire [16-1:0] node23423;
	wire [16-1:0] node23425;
	wire [16-1:0] node23428;
	wire [16-1:0] node23430;
	wire [16-1:0] node23434;
	wire [16-1:0] node23435;
	wire [16-1:0] node23436;
	wire [16-1:0] node23437;
	wire [16-1:0] node23438;
	wire [16-1:0] node23439;
	wire [16-1:0] node23440;
	wire [16-1:0] node23441;
	wire [16-1:0] node23443;
	wire [16-1:0] node23447;
	wire [16-1:0] node23448;
	wire [16-1:0] node23449;
	wire [16-1:0] node23453;
	wire [16-1:0] node23454;
	wire [16-1:0] node23458;
	wire [16-1:0] node23459;
	wire [16-1:0] node23462;
	wire [16-1:0] node23463;
	wire [16-1:0] node23466;
	wire [16-1:0] node23468;
	wire [16-1:0] node23471;
	wire [16-1:0] node23472;
	wire [16-1:0] node23473;
	wire [16-1:0] node23475;
	wire [16-1:0] node23476;
	wire [16-1:0] node23480;
	wire [16-1:0] node23481;
	wire [16-1:0] node23485;
	wire [16-1:0] node23486;
	wire [16-1:0] node23488;
	wire [16-1:0] node23491;
	wire [16-1:0] node23492;
	wire [16-1:0] node23496;
	wire [16-1:0] node23497;
	wire [16-1:0] node23498;
	wire [16-1:0] node23499;
	wire [16-1:0] node23502;
	wire [16-1:0] node23503;
	wire [16-1:0] node23506;
	wire [16-1:0] node23508;
	wire [16-1:0] node23511;
	wire [16-1:0] node23513;
	wire [16-1:0] node23514;
	wire [16-1:0] node23516;
	wire [16-1:0] node23520;
	wire [16-1:0] node23521;
	wire [16-1:0] node23522;
	wire [16-1:0] node23524;
	wire [16-1:0] node23525;
	wire [16-1:0] node23529;
	wire [16-1:0] node23530;
	wire [16-1:0] node23531;
	wire [16-1:0] node23533;
	wire [16-1:0] node23538;
	wire [16-1:0] node23539;
	wire [16-1:0] node23540;
	wire [16-1:0] node23543;
	wire [16-1:0] node23546;
	wire [16-1:0] node23547;
	wire [16-1:0] node23550;
	wire [16-1:0] node23553;
	wire [16-1:0] node23554;
	wire [16-1:0] node23555;
	wire [16-1:0] node23556;
	wire [16-1:0] node23557;
	wire [16-1:0] node23558;
	wire [16-1:0] node23559;
	wire [16-1:0] node23564;
	wire [16-1:0] node23565;
	wire [16-1:0] node23566;
	wire [16-1:0] node23568;
	wire [16-1:0] node23573;
	wire [16-1:0] node23574;
	wire [16-1:0] node23576;
	wire [16-1:0] node23578;
	wire [16-1:0] node23581;
	wire [16-1:0] node23582;
	wire [16-1:0] node23584;
	wire [16-1:0] node23585;
	wire [16-1:0] node23589;
	wire [16-1:0] node23592;
	wire [16-1:0] node23593;
	wire [16-1:0] node23594;
	wire [16-1:0] node23595;
	wire [16-1:0] node23598;
	wire [16-1:0] node23599;
	wire [16-1:0] node23601;
	wire [16-1:0] node23604;
	wire [16-1:0] node23605;
	wire [16-1:0] node23609;
	wire [16-1:0] node23610;
	wire [16-1:0] node23613;
	wire [16-1:0] node23615;
	wire [16-1:0] node23618;
	wire [16-1:0] node23619;
	wire [16-1:0] node23620;
	wire [16-1:0] node23623;
	wire [16-1:0] node23625;
	wire [16-1:0] node23628;
	wire [16-1:0] node23629;
	wire [16-1:0] node23630;
	wire [16-1:0] node23634;
	wire [16-1:0] node23637;
	wire [16-1:0] node23638;
	wire [16-1:0] node23639;
	wire [16-1:0] node23640;
	wire [16-1:0] node23642;
	wire [16-1:0] node23645;
	wire [16-1:0] node23646;
	wire [16-1:0] node23647;
	wire [16-1:0] node23649;
	wire [16-1:0] node23652;
	wire [16-1:0] node23654;
	wire [16-1:0] node23657;
	wire [16-1:0] node23660;
	wire [16-1:0] node23661;
	wire [16-1:0] node23662;
	wire [16-1:0] node23663;
	wire [16-1:0] node23666;
	wire [16-1:0] node23670;
	wire [16-1:0] node23672;
	wire [16-1:0] node23675;
	wire [16-1:0] node23676;
	wire [16-1:0] node23677;
	wire [16-1:0] node23680;
	wire [16-1:0] node23681;
	wire [16-1:0] node23684;
	wire [16-1:0] node23687;
	wire [16-1:0] node23688;
	wire [16-1:0] node23690;
	wire [16-1:0] node23693;
	wire [16-1:0] node23694;
	wire [16-1:0] node23696;
	wire [16-1:0] node23697;
	wire [16-1:0] node23701;
	wire [16-1:0] node23703;
	wire [16-1:0] node23706;
	wire [16-1:0] node23707;
	wire [16-1:0] node23708;
	wire [16-1:0] node23709;
	wire [16-1:0] node23710;
	wire [16-1:0] node23711;
	wire [16-1:0] node23712;
	wire [16-1:0] node23714;
	wire [16-1:0] node23718;
	wire [16-1:0] node23719;
	wire [16-1:0] node23720;
	wire [16-1:0] node23725;
	wire [16-1:0] node23726;
	wire [16-1:0] node23727;
	wire [16-1:0] node23731;
	wire [16-1:0] node23733;
	wire [16-1:0] node23735;
	wire [16-1:0] node23738;
	wire [16-1:0] node23739;
	wire [16-1:0] node23740;
	wire [16-1:0] node23742;
	wire [16-1:0] node23743;
	wire [16-1:0] node23747;
	wire [16-1:0] node23748;
	wire [16-1:0] node23749;
	wire [16-1:0] node23753;
	wire [16-1:0] node23756;
	wire [16-1:0] node23757;
	wire [16-1:0] node23759;
	wire [16-1:0] node23762;
	wire [16-1:0] node23764;
	wire [16-1:0] node23767;
	wire [16-1:0] node23768;
	wire [16-1:0] node23769;
	wire [16-1:0] node23770;
	wire [16-1:0] node23772;
	wire [16-1:0] node23773;
	wire [16-1:0] node23777;
	wire [16-1:0] node23778;
	wire [16-1:0] node23779;
	wire [16-1:0] node23783;
	wire [16-1:0] node23784;
	wire [16-1:0] node23788;
	wire [16-1:0] node23789;
	wire [16-1:0] node23790;
	wire [16-1:0] node23794;
	wire [16-1:0] node23795;
	wire [16-1:0] node23797;
	wire [16-1:0] node23799;
	wire [16-1:0] node23803;
	wire [16-1:0] node23804;
	wire [16-1:0] node23805;
	wire [16-1:0] node23806;
	wire [16-1:0] node23809;
	wire [16-1:0] node23812;
	wire [16-1:0] node23813;
	wire [16-1:0] node23814;
	wire [16-1:0] node23816;
	wire [16-1:0] node23820;
	wire [16-1:0] node23821;
	wire [16-1:0] node23823;
	wire [16-1:0] node23827;
	wire [16-1:0] node23828;
	wire [16-1:0] node23829;
	wire [16-1:0] node23831;
	wire [16-1:0] node23833;
	wire [16-1:0] node23837;
	wire [16-1:0] node23838;
	wire [16-1:0] node23841;
	wire [16-1:0] node23843;
	wire [16-1:0] node23844;
	wire [16-1:0] node23848;
	wire [16-1:0] node23849;
	wire [16-1:0] node23850;
	wire [16-1:0] node23851;
	wire [16-1:0] node23852;
	wire [16-1:0] node23853;
	wire [16-1:0] node23857;
	wire [16-1:0] node23858;
	wire [16-1:0] node23862;
	wire [16-1:0] node23863;
	wire [16-1:0] node23864;
	wire [16-1:0] node23865;
	wire [16-1:0] node23869;
	wire [16-1:0] node23870;
	wire [16-1:0] node23874;
	wire [16-1:0] node23876;
	wire [16-1:0] node23879;
	wire [16-1:0] node23880;
	wire [16-1:0] node23881;
	wire [16-1:0] node23883;
	wire [16-1:0] node23885;
	wire [16-1:0] node23886;
	wire [16-1:0] node23890;
	wire [16-1:0] node23892;
	wire [16-1:0] node23895;
	wire [16-1:0] node23896;
	wire [16-1:0] node23899;
	wire [16-1:0] node23901;
	wire [16-1:0] node23903;
	wire [16-1:0] node23904;
	wire [16-1:0] node23908;
	wire [16-1:0] node23909;
	wire [16-1:0] node23910;
	wire [16-1:0] node23911;
	wire [16-1:0] node23913;
	wire [16-1:0] node23916;
	wire [16-1:0] node23917;
	wire [16-1:0] node23920;
	wire [16-1:0] node23923;
	wire [16-1:0] node23924;
	wire [16-1:0] node23926;
	wire [16-1:0] node23927;
	wire [16-1:0] node23931;
	wire [16-1:0] node23932;
	wire [16-1:0] node23933;
	wire [16-1:0] node23938;
	wire [16-1:0] node23939;
	wire [16-1:0] node23940;
	wire [16-1:0] node23941;
	wire [16-1:0] node23942;
	wire [16-1:0] node23945;
	wire [16-1:0] node23946;
	wire [16-1:0] node23950;
	wire [16-1:0] node23953;
	wire [16-1:0] node23955;
	wire [16-1:0] node23956;
	wire [16-1:0] node23960;
	wire [16-1:0] node23961;
	wire [16-1:0] node23963;
	wire [16-1:0] node23964;
	wire [16-1:0] node23968;
	wire [16-1:0] node23970;
	wire [16-1:0] node23971;
	wire [16-1:0] node23973;
	wire [16-1:0] node23976;
	wire [16-1:0] node23977;
	wire [16-1:0] node23981;
	wire [16-1:0] node23982;
	wire [16-1:0] node23983;
	wire [16-1:0] node23984;
	wire [16-1:0] node23985;
	wire [16-1:0] node23986;
	wire [16-1:0] node23987;
	wire [16-1:0] node23988;
	wire [16-1:0] node23989;
	wire [16-1:0] node23993;
	wire [16-1:0] node23996;
	wire [16-1:0] node23998;
	wire [16-1:0] node24001;
	wire [16-1:0] node24002;
	wire [16-1:0] node24003;
	wire [16-1:0] node24004;
	wire [16-1:0] node24006;
	wire [16-1:0] node24010;
	wire [16-1:0] node24011;
	wire [16-1:0] node24015;
	wire [16-1:0] node24017;
	wire [16-1:0] node24018;
	wire [16-1:0] node24021;
	wire [16-1:0] node24023;
	wire [16-1:0] node24026;
	wire [16-1:0] node24027;
	wire [16-1:0] node24028;
	wire [16-1:0] node24029;
	wire [16-1:0] node24030;
	wire [16-1:0] node24033;
	wire [16-1:0] node24035;
	wire [16-1:0] node24038;
	wire [16-1:0] node24041;
	wire [16-1:0] node24042;
	wire [16-1:0] node24043;
	wire [16-1:0] node24044;
	wire [16-1:0] node24048;
	wire [16-1:0] node24051;
	wire [16-1:0] node24052;
	wire [16-1:0] node24055;
	wire [16-1:0] node24057;
	wire [16-1:0] node24060;
	wire [16-1:0] node24061;
	wire [16-1:0] node24063;
	wire [16-1:0] node24066;
	wire [16-1:0] node24067;
	wire [16-1:0] node24068;
	wire [16-1:0] node24071;
	wire [16-1:0] node24074;
	wire [16-1:0] node24075;
	wire [16-1:0] node24076;
	wire [16-1:0] node24080;
	wire [16-1:0] node24083;
	wire [16-1:0] node24084;
	wire [16-1:0] node24085;
	wire [16-1:0] node24086;
	wire [16-1:0] node24087;
	wire [16-1:0] node24090;
	wire [16-1:0] node24091;
	wire [16-1:0] node24093;
	wire [16-1:0] node24094;
	wire [16-1:0] node24099;
	wire [16-1:0] node24100;
	wire [16-1:0] node24102;
	wire [16-1:0] node24103;
	wire [16-1:0] node24104;
	wire [16-1:0] node24109;
	wire [16-1:0] node24110;
	wire [16-1:0] node24111;
	wire [16-1:0] node24116;
	wire [16-1:0] node24117;
	wire [16-1:0] node24118;
	wire [16-1:0] node24119;
	wire [16-1:0] node24120;
	wire [16-1:0] node24122;
	wire [16-1:0] node24125;
	wire [16-1:0] node24128;
	wire [16-1:0] node24130;
	wire [16-1:0] node24133;
	wire [16-1:0] node24134;
	wire [16-1:0] node24136;
	wire [16-1:0] node24139;
	wire [16-1:0] node24140;
	wire [16-1:0] node24144;
	wire [16-1:0] node24145;
	wire [16-1:0] node24147;
	wire [16-1:0] node24149;
	wire [16-1:0] node24152;
	wire [16-1:0] node24153;
	wire [16-1:0] node24155;
	wire [16-1:0] node24158;
	wire [16-1:0] node24161;
	wire [16-1:0] node24162;
	wire [16-1:0] node24163;
	wire [16-1:0] node24164;
	wire [16-1:0] node24165;
	wire [16-1:0] node24167;
	wire [16-1:0] node24170;
	wire [16-1:0] node24172;
	wire [16-1:0] node24175;
	wire [16-1:0] node24176;
	wire [16-1:0] node24179;
	wire [16-1:0] node24180;
	wire [16-1:0] node24182;
	wire [16-1:0] node24186;
	wire [16-1:0] node24187;
	wire [16-1:0] node24189;
	wire [16-1:0] node24192;
	wire [16-1:0] node24193;
	wire [16-1:0] node24194;
	wire [16-1:0] node24198;
	wire [16-1:0] node24201;
	wire [16-1:0] node24202;
	wire [16-1:0] node24203;
	wire [16-1:0] node24204;
	wire [16-1:0] node24207;
	wire [16-1:0] node24210;
	wire [16-1:0] node24211;
	wire [16-1:0] node24214;
	wire [16-1:0] node24217;
	wire [16-1:0] node24218;
	wire [16-1:0] node24219;
	wire [16-1:0] node24220;
	wire [16-1:0] node24223;
	wire [16-1:0] node24227;
	wire [16-1:0] node24230;
	wire [16-1:0] node24231;
	wire [16-1:0] node24232;
	wire [16-1:0] node24233;
	wire [16-1:0] node24234;
	wire [16-1:0] node24235;
	wire [16-1:0] node24236;
	wire [16-1:0] node24237;
	wire [16-1:0] node24242;
	wire [16-1:0] node24244;
	wire [16-1:0] node24247;
	wire [16-1:0] node24249;
	wire [16-1:0] node24250;
	wire [16-1:0] node24252;
	wire [16-1:0] node24256;
	wire [16-1:0] node24257;
	wire [16-1:0] node24258;
	wire [16-1:0] node24259;
	wire [16-1:0] node24262;
	wire [16-1:0] node24264;
	wire [16-1:0] node24267;
	wire [16-1:0] node24268;
	wire [16-1:0] node24269;
	wire [16-1:0] node24271;
	wire [16-1:0] node24275;
	wire [16-1:0] node24278;
	wire [16-1:0] node24279;
	wire [16-1:0] node24280;
	wire [16-1:0] node24283;
	wire [16-1:0] node24285;
	wire [16-1:0] node24286;
	wire [16-1:0] node24290;
	wire [16-1:0] node24292;
	wire [16-1:0] node24295;
	wire [16-1:0] node24296;
	wire [16-1:0] node24297;
	wire [16-1:0] node24298;
	wire [16-1:0] node24299;
	wire [16-1:0] node24301;
	wire [16-1:0] node24302;
	wire [16-1:0] node24306;
	wire [16-1:0] node24309;
	wire [16-1:0] node24310;
	wire [16-1:0] node24313;
	wire [16-1:0] node24315;
	wire [16-1:0] node24318;
	wire [16-1:0] node24319;
	wire [16-1:0] node24321;
	wire [16-1:0] node24322;
	wire [16-1:0] node24326;
	wire [16-1:0] node24327;
	wire [16-1:0] node24330;
	wire [16-1:0] node24332;
	wire [16-1:0] node24335;
	wire [16-1:0] node24336;
	wire [16-1:0] node24337;
	wire [16-1:0] node24338;
	wire [16-1:0] node24341;
	wire [16-1:0] node24344;
	wire [16-1:0] node24346;
	wire [16-1:0] node24347;
	wire [16-1:0] node24349;
	wire [16-1:0] node24353;
	wire [16-1:0] node24354;
	wire [16-1:0] node24356;
	wire [16-1:0] node24359;
	wire [16-1:0] node24360;
	wire [16-1:0] node24363;
	wire [16-1:0] node24365;
	wire [16-1:0] node24368;
	wire [16-1:0] node24369;
	wire [16-1:0] node24370;
	wire [16-1:0] node24371;
	wire [16-1:0] node24372;
	wire [16-1:0] node24375;
	wire [16-1:0] node24376;
	wire [16-1:0] node24380;
	wire [16-1:0] node24382;
	wire [16-1:0] node24385;
	wire [16-1:0] node24386;
	wire [16-1:0] node24387;
	wire [16-1:0] node24389;
	wire [16-1:0] node24393;
	wire [16-1:0] node24394;
	wire [16-1:0] node24395;
	wire [16-1:0] node24399;
	wire [16-1:0] node24401;
	wire [16-1:0] node24402;
	wire [16-1:0] node24406;
	wire [16-1:0] node24407;
	wire [16-1:0] node24408;
	wire [16-1:0] node24409;
	wire [16-1:0] node24410;
	wire [16-1:0] node24411;
	wire [16-1:0] node24416;
	wire [16-1:0] node24417;
	wire [16-1:0] node24420;
	wire [16-1:0] node24422;
	wire [16-1:0] node24425;
	wire [16-1:0] node24426;
	wire [16-1:0] node24427;
	wire [16-1:0] node24428;
	wire [16-1:0] node24433;
	wire [16-1:0] node24434;
	wire [16-1:0] node24437;
	wire [16-1:0] node24439;
	wire [16-1:0] node24442;
	wire [16-1:0] node24443;
	wire [16-1:0] node24444;
	wire [16-1:0] node24447;
	wire [16-1:0] node24449;
	wire [16-1:0] node24452;
	wire [16-1:0] node24453;
	wire [16-1:0] node24454;
	wire [16-1:0] node24457;
	wire [16-1:0] node24459;
	wire [16-1:0] node24462;
	wire [16-1:0] node24463;
	wire [16-1:0] node24465;
	wire [16-1:0] node24467;
	wire [16-1:0] node24470;
	wire [16-1:0] node24471;
	wire [16-1:0] node24475;
	wire [16-1:0] node24476;
	wire [16-1:0] node24477;
	wire [16-1:0] node24478;
	wire [16-1:0] node24479;
	wire [16-1:0] node24480;
	wire [16-1:0] node24481;
	wire [16-1:0] node24482;
	wire [16-1:0] node24486;
	wire [16-1:0] node24487;
	wire [16-1:0] node24491;
	wire [16-1:0] node24492;
	wire [16-1:0] node24493;
	wire [16-1:0] node24496;
	wire [16-1:0] node24497;
	wire [16-1:0] node24501;
	wire [16-1:0] node24502;
	wire [16-1:0] node24503;
	wire [16-1:0] node24508;
	wire [16-1:0] node24509;
	wire [16-1:0] node24510;
	wire [16-1:0] node24511;
	wire [16-1:0] node24513;
	wire [16-1:0] node24515;
	wire [16-1:0] node24518;
	wire [16-1:0] node24519;
	wire [16-1:0] node24523;
	wire [16-1:0] node24524;
	wire [16-1:0] node24527;
	wire [16-1:0] node24529;
	wire [16-1:0] node24532;
	wire [16-1:0] node24533;
	wire [16-1:0] node24534;
	wire [16-1:0] node24535;
	wire [16-1:0] node24540;
	wire [16-1:0] node24543;
	wire [16-1:0] node24544;
	wire [16-1:0] node24545;
	wire [16-1:0] node24546;
	wire [16-1:0] node24547;
	wire [16-1:0] node24551;
	wire [16-1:0] node24552;
	wire [16-1:0] node24553;
	wire [16-1:0] node24556;
	wire [16-1:0] node24557;
	wire [16-1:0] node24561;
	wire [16-1:0] node24563;
	wire [16-1:0] node24564;
	wire [16-1:0] node24568;
	wire [16-1:0] node24569;
	wire [16-1:0] node24570;
	wire [16-1:0] node24571;
	wire [16-1:0] node24575;
	wire [16-1:0] node24577;
	wire [16-1:0] node24579;
	wire [16-1:0] node24582;
	wire [16-1:0] node24583;
	wire [16-1:0] node24585;
	wire [16-1:0] node24589;
	wire [16-1:0] node24590;
	wire [16-1:0] node24591;
	wire [16-1:0] node24593;
	wire [16-1:0] node24595;
	wire [16-1:0] node24596;
	wire [16-1:0] node24600;
	wire [16-1:0] node24601;
	wire [16-1:0] node24604;
	wire [16-1:0] node24606;
	wire [16-1:0] node24607;
	wire [16-1:0] node24611;
	wire [16-1:0] node24613;
	wire [16-1:0] node24615;
	wire [16-1:0] node24616;
	wire [16-1:0] node24618;
	wire [16-1:0] node24622;
	wire [16-1:0] node24623;
	wire [16-1:0] node24624;
	wire [16-1:0] node24625;
	wire [16-1:0] node24626;
	wire [16-1:0] node24627;
	wire [16-1:0] node24630;
	wire [16-1:0] node24633;
	wire [16-1:0] node24634;
	wire [16-1:0] node24638;
	wire [16-1:0] node24639;
	wire [16-1:0] node24640;
	wire [16-1:0] node24642;
	wire [16-1:0] node24644;
	wire [16-1:0] node24647;
	wire [16-1:0] node24648;
	wire [16-1:0] node24653;
	wire [16-1:0] node24654;
	wire [16-1:0] node24655;
	wire [16-1:0] node24656;
	wire [16-1:0] node24658;
	wire [16-1:0] node24660;
	wire [16-1:0] node24664;
	wire [16-1:0] node24665;
	wire [16-1:0] node24669;
	wire [16-1:0] node24670;
	wire [16-1:0] node24671;
	wire [16-1:0] node24673;
	wire [16-1:0] node24675;
	wire [16-1:0] node24678;
	wire [16-1:0] node24681;
	wire [16-1:0] node24682;
	wire [16-1:0] node24683;
	wire [16-1:0] node24687;
	wire [16-1:0] node24688;
	wire [16-1:0] node24692;
	wire [16-1:0] node24693;
	wire [16-1:0] node24694;
	wire [16-1:0] node24695;
	wire [16-1:0] node24697;
	wire [16-1:0] node24698;
	wire [16-1:0] node24703;
	wire [16-1:0] node24704;
	wire [16-1:0] node24705;
	wire [16-1:0] node24708;
	wire [16-1:0] node24711;
	wire [16-1:0] node24713;
	wire [16-1:0] node24716;
	wire [16-1:0] node24717;
	wire [16-1:0] node24718;
	wire [16-1:0] node24719;
	wire [16-1:0] node24722;
	wire [16-1:0] node24725;
	wire [16-1:0] node24726;
	wire [16-1:0] node24730;
	wire [16-1:0] node24731;
	wire [16-1:0] node24733;
	wire [16-1:0] node24734;
	wire [16-1:0] node24736;
	wire [16-1:0] node24740;
	wire [16-1:0] node24741;
	wire [16-1:0] node24744;
	wire [16-1:0] node24745;
	wire [16-1:0] node24747;
	wire [16-1:0] node24750;
	wire [16-1:0] node24753;
	wire [16-1:0] node24754;
	wire [16-1:0] node24755;
	wire [16-1:0] node24756;
	wire [16-1:0] node24757;
	wire [16-1:0] node24758;
	wire [16-1:0] node24759;
	wire [16-1:0] node24763;
	wire [16-1:0] node24764;
	wire [16-1:0] node24765;
	wire [16-1:0] node24769;
	wire [16-1:0] node24772;
	wire [16-1:0] node24773;
	wire [16-1:0] node24774;
	wire [16-1:0] node24779;
	wire [16-1:0] node24780;
	wire [16-1:0] node24781;
	wire [16-1:0] node24783;
	wire [16-1:0] node24785;
	wire [16-1:0] node24789;
	wire [16-1:0] node24790;
	wire [16-1:0] node24791;
	wire [16-1:0] node24795;
	wire [16-1:0] node24796;
	wire [16-1:0] node24799;
	wire [16-1:0] node24802;
	wire [16-1:0] node24803;
	wire [16-1:0] node24804;
	wire [16-1:0] node24805;
	wire [16-1:0] node24806;
	wire [16-1:0] node24807;
	wire [16-1:0] node24809;
	wire [16-1:0] node24814;
	wire [16-1:0] node24815;
	wire [16-1:0] node24816;
	wire [16-1:0] node24820;
	wire [16-1:0] node24822;
	wire [16-1:0] node24825;
	wire [16-1:0] node24826;
	wire [16-1:0] node24828;
	wire [16-1:0] node24829;
	wire [16-1:0] node24834;
	wire [16-1:0] node24836;
	wire [16-1:0] node24837;
	wire [16-1:0] node24838;
	wire [16-1:0] node24841;
	wire [16-1:0] node24844;
	wire [16-1:0] node24845;
	wire [16-1:0] node24848;
	wire [16-1:0] node24849;
	wire [16-1:0] node24853;
	wire [16-1:0] node24854;
	wire [16-1:0] node24855;
	wire [16-1:0] node24856;
	wire [16-1:0] node24857;
	wire [16-1:0] node24858;
	wire [16-1:0] node24861;
	wire [16-1:0] node24864;
	wire [16-1:0] node24865;
	wire [16-1:0] node24868;
	wire [16-1:0] node24869;
	wire [16-1:0] node24871;
	wire [16-1:0] node24875;
	wire [16-1:0] node24876;
	wire [16-1:0] node24877;
	wire [16-1:0] node24879;
	wire [16-1:0] node24882;
	wire [16-1:0] node24883;
	wire [16-1:0] node24887;
	wire [16-1:0] node24888;
	wire [16-1:0] node24891;
	wire [16-1:0] node24893;
	wire [16-1:0] node24894;
	wire [16-1:0] node24898;
	wire [16-1:0] node24899;
	wire [16-1:0] node24900;
	wire [16-1:0] node24901;
	wire [16-1:0] node24905;
	wire [16-1:0] node24906;
	wire [16-1:0] node24909;
	wire [16-1:0] node24911;
	wire [16-1:0] node24914;
	wire [16-1:0] node24915;
	wire [16-1:0] node24916;
	wire [16-1:0] node24919;
	wire [16-1:0] node24922;
	wire [16-1:0] node24923;
	wire [16-1:0] node24924;
	wire [16-1:0] node24929;
	wire [16-1:0] node24930;
	wire [16-1:0] node24931;
	wire [16-1:0] node24933;
	wire [16-1:0] node24936;
	wire [16-1:0] node24937;
	wire [16-1:0] node24938;
	wire [16-1:0] node24940;
	wire [16-1:0] node24942;
	wire [16-1:0] node24946;
	wire [16-1:0] node24949;
	wire [16-1:0] node24950;
	wire [16-1:0] node24951;
	wire [16-1:0] node24954;
	wire [16-1:0] node24956;
	wire [16-1:0] node24959;
	wire [16-1:0] node24960;
	wire [16-1:0] node24961;
	wire [16-1:0] node24963;
	wire [16-1:0] node24966;
	wire [16-1:0] node24969;
	wire [16-1:0] node24971;
	wire [16-1:0] node24972;
	wire [16-1:0] node24973;
	wire [16-1:0] node24976;
	wire [16-1:0] node24980;
	wire [16-1:0] node24981;
	wire [16-1:0] node24982;
	wire [16-1:0] node24983;
	wire [16-1:0] node24984;
	wire [16-1:0] node24985;
	wire [16-1:0] node24986;
	wire [16-1:0] node24987;
	wire [16-1:0] node24988;
	wire [16-1:0] node24989;
	wire [16-1:0] node24990;
	wire [16-1:0] node24991;
	wire [16-1:0] node24995;
	wire [16-1:0] node24998;
	wire [16-1:0] node24999;
	wire [16-1:0] node25000;
	wire [16-1:0] node25002;
	wire [16-1:0] node25006;
	wire [16-1:0] node25007;
	wire [16-1:0] node25008;
	wire [16-1:0] node25012;
	wire [16-1:0] node25013;
	wire [16-1:0] node25017;
	wire [16-1:0] node25018;
	wire [16-1:0] node25019;
	wire [16-1:0] node25020;
	wire [16-1:0] node25024;
	wire [16-1:0] node25025;
	wire [16-1:0] node25028;
	wire [16-1:0] node25030;
	wire [16-1:0] node25033;
	wire [16-1:0] node25034;
	wire [16-1:0] node25035;
	wire [16-1:0] node25037;
	wire [16-1:0] node25038;
	wire [16-1:0] node25043;
	wire [16-1:0] node25044;
	wire [16-1:0] node25048;
	wire [16-1:0] node25049;
	wire [16-1:0] node25050;
	wire [16-1:0] node25051;
	wire [16-1:0] node25053;
	wire [16-1:0] node25054;
	wire [16-1:0] node25058;
	wire [16-1:0] node25059;
	wire [16-1:0] node25060;
	wire [16-1:0] node25064;
	wire [16-1:0] node25066;
	wire [16-1:0] node25067;
	wire [16-1:0] node25071;
	wire [16-1:0] node25072;
	wire [16-1:0] node25073;
	wire [16-1:0] node25076;
	wire [16-1:0] node25079;
	wire [16-1:0] node25080;
	wire [16-1:0] node25081;
	wire [16-1:0] node25083;
	wire [16-1:0] node25086;
	wire [16-1:0] node25088;
	wire [16-1:0] node25092;
	wire [16-1:0] node25093;
	wire [16-1:0] node25094;
	wire [16-1:0] node25096;
	wire [16-1:0] node25099;
	wire [16-1:0] node25100;
	wire [16-1:0] node25101;
	wire [16-1:0] node25105;
	wire [16-1:0] node25108;
	wire [16-1:0] node25109;
	wire [16-1:0] node25111;
	wire [16-1:0] node25112;
	wire [16-1:0] node25114;
	wire [16-1:0] node25119;
	wire [16-1:0] node25120;
	wire [16-1:0] node25121;
	wire [16-1:0] node25122;
	wire [16-1:0] node25123;
	wire [16-1:0] node25124;
	wire [16-1:0] node25125;
	wire [16-1:0] node25129;
	wire [16-1:0] node25132;
	wire [16-1:0] node25133;
	wire [16-1:0] node25137;
	wire [16-1:0] node25139;
	wire [16-1:0] node25140;
	wire [16-1:0] node25144;
	wire [16-1:0] node25145;
	wire [16-1:0] node25146;
	wire [16-1:0] node25147;
	wire [16-1:0] node25149;
	wire [16-1:0] node25152;
	wire [16-1:0] node25153;
	wire [16-1:0] node25157;
	wire [16-1:0] node25158;
	wire [16-1:0] node25161;
	wire [16-1:0] node25163;
	wire [16-1:0] node25166;
	wire [16-1:0] node25167;
	wire [16-1:0] node25170;
	wire [16-1:0] node25172;
	wire [16-1:0] node25175;
	wire [16-1:0] node25176;
	wire [16-1:0] node25177;
	wire [16-1:0] node25180;
	wire [16-1:0] node25181;
	wire [16-1:0] node25182;
	wire [16-1:0] node25185;
	wire [16-1:0] node25187;
	wire [16-1:0] node25190;
	wire [16-1:0] node25191;
	wire [16-1:0] node25193;
	wire [16-1:0] node25194;
	wire [16-1:0] node25199;
	wire [16-1:0] node25200;
	wire [16-1:0] node25201;
	wire [16-1:0] node25202;
	wire [16-1:0] node25206;
	wire [16-1:0] node25207;
	wire [16-1:0] node25208;
	wire [16-1:0] node25210;
	wire [16-1:0] node25214;
	wire [16-1:0] node25217;
	wire [16-1:0] node25218;
	wire [16-1:0] node25219;
	wire [16-1:0] node25220;
	wire [16-1:0] node25224;
	wire [16-1:0] node25226;
	wire [16-1:0] node25229;
	wire [16-1:0] node25231;
	wire [16-1:0] node25232;
	wire [16-1:0] node25236;
	wire [16-1:0] node25237;
	wire [16-1:0] node25238;
	wire [16-1:0] node25239;
	wire [16-1:0] node25240;
	wire [16-1:0] node25241;
	wire [16-1:0] node25242;
	wire [16-1:0] node25245;
	wire [16-1:0] node25248;
	wire [16-1:0] node25249;
	wire [16-1:0] node25250;
	wire [16-1:0] node25254;
	wire [16-1:0] node25257;
	wire [16-1:0] node25258;
	wire [16-1:0] node25259;
	wire [16-1:0] node25260;
	wire [16-1:0] node25262;
	wire [16-1:0] node25265;
	wire [16-1:0] node25267;
	wire [16-1:0] node25270;
	wire [16-1:0] node25271;
	wire [16-1:0] node25275;
	wire [16-1:0] node25276;
	wire [16-1:0] node25280;
	wire [16-1:0] node25281;
	wire [16-1:0] node25282;
	wire [16-1:0] node25283;
	wire [16-1:0] node25285;
	wire [16-1:0] node25286;
	wire [16-1:0] node25290;
	wire [16-1:0] node25293;
	wire [16-1:0] node25294;
	wire [16-1:0] node25295;
	wire [16-1:0] node25297;
	wire [16-1:0] node25301;
	wire [16-1:0] node25304;
	wire [16-1:0] node25305;
	wire [16-1:0] node25306;
	wire [16-1:0] node25309;
	wire [16-1:0] node25311;
	wire [16-1:0] node25314;
	wire [16-1:0] node25315;
	wire [16-1:0] node25316;
	wire [16-1:0] node25318;
	wire [16-1:0] node25322;
	wire [16-1:0] node25325;
	wire [16-1:0] node25326;
	wire [16-1:0] node25327;
	wire [16-1:0] node25328;
	wire [16-1:0] node25329;
	wire [16-1:0] node25330;
	wire [16-1:0] node25334;
	wire [16-1:0] node25337;
	wire [16-1:0] node25338;
	wire [16-1:0] node25339;
	wire [16-1:0] node25343;
	wire [16-1:0] node25346;
	wire [16-1:0] node25348;
	wire [16-1:0] node25349;
	wire [16-1:0] node25352;
	wire [16-1:0] node25355;
	wire [16-1:0] node25356;
	wire [16-1:0] node25358;
	wire [16-1:0] node25359;
	wire [16-1:0] node25360;
	wire [16-1:0] node25362;
	wire [16-1:0] node25367;
	wire [16-1:0] node25368;
	wire [16-1:0] node25370;
	wire [16-1:0] node25372;
	wire [16-1:0] node25375;
	wire [16-1:0] node25376;
	wire [16-1:0] node25378;
	wire [16-1:0] node25379;
	wire [16-1:0] node25384;
	wire [16-1:0] node25385;
	wire [16-1:0] node25386;
	wire [16-1:0] node25387;
	wire [16-1:0] node25388;
	wire [16-1:0] node25389;
	wire [16-1:0] node25391;
	wire [16-1:0] node25392;
	wire [16-1:0] node25396;
	wire [16-1:0] node25399;
	wire [16-1:0] node25400;
	wire [16-1:0] node25401;
	wire [16-1:0] node25405;
	wire [16-1:0] node25408;
	wire [16-1:0] node25409;
	wire [16-1:0] node25410;
	wire [16-1:0] node25414;
	wire [16-1:0] node25416;
	wire [16-1:0] node25417;
	wire [16-1:0] node25421;
	wire [16-1:0] node25422;
	wire [16-1:0] node25423;
	wire [16-1:0] node25425;
	wire [16-1:0] node25426;
	wire [16-1:0] node25430;
	wire [16-1:0] node25431;
	wire [16-1:0] node25432;
	wire [16-1:0] node25437;
	wire [16-1:0] node25438;
	wire [16-1:0] node25439;
	wire [16-1:0] node25443;
	wire [16-1:0] node25444;
	wire [16-1:0] node25447;
	wire [16-1:0] node25450;
	wire [16-1:0] node25451;
	wire [16-1:0] node25452;
	wire [16-1:0] node25453;
	wire [16-1:0] node25454;
	wire [16-1:0] node25459;
	wire [16-1:0] node25460;
	wire [16-1:0] node25461;
	wire [16-1:0] node25464;
	wire [16-1:0] node25467;
	wire [16-1:0] node25468;
	wire [16-1:0] node25471;
	wire [16-1:0] node25473;
	wire [16-1:0] node25476;
	wire [16-1:0] node25477;
	wire [16-1:0] node25479;
	wire [16-1:0] node25480;
	wire [16-1:0] node25484;
	wire [16-1:0] node25485;
	wire [16-1:0] node25486;
	wire [16-1:0] node25487;
	wire [16-1:0] node25491;
	wire [16-1:0] node25493;
	wire [16-1:0] node25495;
	wire [16-1:0] node25498;
	wire [16-1:0] node25500;
	wire [16-1:0] node25502;
	wire [16-1:0] node25505;
	wire [16-1:0] node25506;
	wire [16-1:0] node25507;
	wire [16-1:0] node25508;
	wire [16-1:0] node25509;
	wire [16-1:0] node25510;
	wire [16-1:0] node25511;
	wire [16-1:0] node25513;
	wire [16-1:0] node25514;
	wire [16-1:0] node25517;
	wire [16-1:0] node25518;
	wire [16-1:0] node25522;
	wire [16-1:0] node25525;
	wire [16-1:0] node25526;
	wire [16-1:0] node25528;
	wire [16-1:0] node25531;
	wire [16-1:0] node25534;
	wire [16-1:0] node25535;
	wire [16-1:0] node25536;
	wire [16-1:0] node25538;
	wire [16-1:0] node25541;
	wire [16-1:0] node25542;
	wire [16-1:0] node25546;
	wire [16-1:0] node25547;
	wire [16-1:0] node25548;
	wire [16-1:0] node25552;
	wire [16-1:0] node25553;
	wire [16-1:0] node25556;
	wire [16-1:0] node25559;
	wire [16-1:0] node25560;
	wire [16-1:0] node25561;
	wire [16-1:0] node25563;
	wire [16-1:0] node25564;
	wire [16-1:0] node25567;
	wire [16-1:0] node25570;
	wire [16-1:0] node25571;
	wire [16-1:0] node25572;
	wire [16-1:0] node25576;
	wire [16-1:0] node25577;
	wire [16-1:0] node25580;
	wire [16-1:0] node25583;
	wire [16-1:0] node25584;
	wire [16-1:0] node25585;
	wire [16-1:0] node25586;
	wire [16-1:0] node25588;
	wire [16-1:0] node25589;
	wire [16-1:0] node25593;
	wire [16-1:0] node25594;
	wire [16-1:0] node25598;
	wire [16-1:0] node25600;
	wire [16-1:0] node25603;
	wire [16-1:0] node25605;
	wire [16-1:0] node25606;
	wire [16-1:0] node25610;
	wire [16-1:0] node25611;
	wire [16-1:0] node25612;
	wire [16-1:0] node25613;
	wire [16-1:0] node25614;
	wire [16-1:0] node25615;
	wire [16-1:0] node25619;
	wire [16-1:0] node25620;
	wire [16-1:0] node25622;
	wire [16-1:0] node25623;
	wire [16-1:0] node25628;
	wire [16-1:0] node25629;
	wire [16-1:0] node25631;
	wire [16-1:0] node25634;
	wire [16-1:0] node25637;
	wire [16-1:0] node25638;
	wire [16-1:0] node25639;
	wire [16-1:0] node25640;
	wire [16-1:0] node25641;
	wire [16-1:0] node25642;
	wire [16-1:0] node25646;
	wire [16-1:0] node25649;
	wire [16-1:0] node25652;
	wire [16-1:0] node25654;
	wire [16-1:0] node25657;
	wire [16-1:0] node25658;
	wire [16-1:0] node25659;
	wire [16-1:0] node25660;
	wire [16-1:0] node25665;
	wire [16-1:0] node25666;
	wire [16-1:0] node25669;
	wire [16-1:0] node25672;
	wire [16-1:0] node25673;
	wire [16-1:0] node25674;
	wire [16-1:0] node25676;
	wire [16-1:0] node25677;
	wire [16-1:0] node25681;
	wire [16-1:0] node25682;
	wire [16-1:0] node25683;
	wire [16-1:0] node25684;
	wire [16-1:0] node25686;
	wire [16-1:0] node25690;
	wire [16-1:0] node25692;
	wire [16-1:0] node25693;
	wire [16-1:0] node25698;
	wire [16-1:0] node25699;
	wire [16-1:0] node25700;
	wire [16-1:0] node25701;
	wire [16-1:0] node25704;
	wire [16-1:0] node25706;
	wire [16-1:0] node25707;
	wire [16-1:0] node25711;
	wire [16-1:0] node25712;
	wire [16-1:0] node25714;
	wire [16-1:0] node25718;
	wire [16-1:0] node25719;
	wire [16-1:0] node25722;
	wire [16-1:0] node25723;
	wire [16-1:0] node25726;
	wire [16-1:0] node25728;
	wire [16-1:0] node25730;
	wire [16-1:0] node25733;
	wire [16-1:0] node25734;
	wire [16-1:0] node25735;
	wire [16-1:0] node25736;
	wire [16-1:0] node25737;
	wire [16-1:0] node25738;
	wire [16-1:0] node25739;
	wire [16-1:0] node25740;
	wire [16-1:0] node25745;
	wire [16-1:0] node25747;
	wire [16-1:0] node25749;
	wire [16-1:0] node25752;
	wire [16-1:0] node25753;
	wire [16-1:0] node25754;
	wire [16-1:0] node25757;
	wire [16-1:0] node25759;
	wire [16-1:0] node25760;
	wire [16-1:0] node25764;
	wire [16-1:0] node25765;
	wire [16-1:0] node25768;
	wire [16-1:0] node25769;
	wire [16-1:0] node25772;
	wire [16-1:0] node25775;
	wire [16-1:0] node25776;
	wire [16-1:0] node25777;
	wire [16-1:0] node25779;
	wire [16-1:0] node25781;
	wire [16-1:0] node25784;
	wire [16-1:0] node25785;
	wire [16-1:0] node25788;
	wire [16-1:0] node25791;
	wire [16-1:0] node25792;
	wire [16-1:0] node25795;
	wire [16-1:0] node25796;
	wire [16-1:0] node25798;
	wire [16-1:0] node25800;
	wire [16-1:0] node25803;
	wire [16-1:0] node25806;
	wire [16-1:0] node25807;
	wire [16-1:0] node25808;
	wire [16-1:0] node25809;
	wire [16-1:0] node25810;
	wire [16-1:0] node25812;
	wire [16-1:0] node25816;
	wire [16-1:0] node25817;
	wire [16-1:0] node25818;
	wire [16-1:0] node25823;
	wire [16-1:0] node25824;
	wire [16-1:0] node25825;
	wire [16-1:0] node25827;
	wire [16-1:0] node25830;
	wire [16-1:0] node25833;
	wire [16-1:0] node25834;
	wire [16-1:0] node25835;
	wire [16-1:0] node25837;
	wire [16-1:0] node25841;
	wire [16-1:0] node25843;
	wire [16-1:0] node25846;
	wire [16-1:0] node25847;
	wire [16-1:0] node25849;
	wire [16-1:0] node25850;
	wire [16-1:0] node25854;
	wire [16-1:0] node25855;
	wire [16-1:0] node25859;
	wire [16-1:0] node25860;
	wire [16-1:0] node25861;
	wire [16-1:0] node25862;
	wire [16-1:0] node25863;
	wire [16-1:0] node25865;
	wire [16-1:0] node25868;
	wire [16-1:0] node25869;
	wire [16-1:0] node25872;
	wire [16-1:0] node25875;
	wire [16-1:0] node25876;
	wire [16-1:0] node25877;
	wire [16-1:0] node25878;
	wire [16-1:0] node25881;
	wire [16-1:0] node25882;
	wire [16-1:0] node25886;
	wire [16-1:0] node25889;
	wire [16-1:0] node25890;
	wire [16-1:0] node25894;
	wire [16-1:0] node25895;
	wire [16-1:0] node25896;
	wire [16-1:0] node25897;
	wire [16-1:0] node25901;
	wire [16-1:0] node25903;
	wire [16-1:0] node25905;
	wire [16-1:0] node25908;
	wire [16-1:0] node25909;
	wire [16-1:0] node25911;
	wire [16-1:0] node25914;
	wire [16-1:0] node25915;
	wire [16-1:0] node25916;
	wire [16-1:0] node25921;
	wire [16-1:0] node25922;
	wire [16-1:0] node25923;
	wire [16-1:0] node25925;
	wire [16-1:0] node25926;
	wire [16-1:0] node25929;
	wire [16-1:0] node25932;
	wire [16-1:0] node25934;
	wire [16-1:0] node25936;
	wire [16-1:0] node25939;
	wire [16-1:0] node25940;
	wire [16-1:0] node25941;
	wire [16-1:0] node25942;
	wire [16-1:0] node25943;
	wire [16-1:0] node25948;
	wire [16-1:0] node25950;
	wire [16-1:0] node25951;
	wire [16-1:0] node25953;
	wire [16-1:0] node25957;
	wire [16-1:0] node25958;
	wire [16-1:0] node25960;
	wire [16-1:0] node25963;
	wire [16-1:0] node25964;
	wire [16-1:0] node25967;
	wire [16-1:0] node25969;
	wire [16-1:0] node25972;
	wire [16-1:0] node25973;
	wire [16-1:0] node25974;
	wire [16-1:0] node25975;
	wire [16-1:0] node25976;
	wire [16-1:0] node25977;
	wire [16-1:0] node25978;
	wire [16-1:0] node25979;
	wire [16-1:0] node25980;
	wire [16-1:0] node25982;
	wire [16-1:0] node25983;
	wire [16-1:0] node25987;
	wire [16-1:0] node25988;
	wire [16-1:0] node25990;
	wire [16-1:0] node25994;
	wire [16-1:0] node25995;
	wire [16-1:0] node25998;
	wire [16-1:0] node25999;
	wire [16-1:0] node26001;
	wire [16-1:0] node26005;
	wire [16-1:0] node26006;
	wire [16-1:0] node26008;
	wire [16-1:0] node26012;
	wire [16-1:0] node26013;
	wire [16-1:0] node26014;
	wire [16-1:0] node26015;
	wire [16-1:0] node26018;
	wire [16-1:0] node26021;
	wire [16-1:0] node26022;
	wire [16-1:0] node26025;
	wire [16-1:0] node26028;
	wire [16-1:0] node26029;
	wire [16-1:0] node26031;
	wire [16-1:0] node26032;
	wire [16-1:0] node26034;
	wire [16-1:0] node26038;
	wire [16-1:0] node26039;
	wire [16-1:0] node26042;
	wire [16-1:0] node26045;
	wire [16-1:0] node26046;
	wire [16-1:0] node26047;
	wire [16-1:0] node26048;
	wire [16-1:0] node26050;
	wire [16-1:0] node26051;
	wire [16-1:0] node26055;
	wire [16-1:0] node26057;
	wire [16-1:0] node26060;
	wire [16-1:0] node26061;
	wire [16-1:0] node26062;
	wire [16-1:0] node26064;
	wire [16-1:0] node26066;
	wire [16-1:0] node26069;
	wire [16-1:0] node26070;
	wire [16-1:0] node26074;
	wire [16-1:0] node26075;
	wire [16-1:0] node26079;
	wire [16-1:0] node26080;
	wire [16-1:0] node26081;
	wire [16-1:0] node26083;
	wire [16-1:0] node26084;
	wire [16-1:0] node26088;
	wire [16-1:0] node26089;
	wire [16-1:0] node26093;
	wire [16-1:0] node26095;
	wire [16-1:0] node26096;
	wire [16-1:0] node26098;
	wire [16-1:0] node26101;
	wire [16-1:0] node26102;
	wire [16-1:0] node26103;
	wire [16-1:0] node26108;
	wire [16-1:0] node26109;
	wire [16-1:0] node26110;
	wire [16-1:0] node26111;
	wire [16-1:0] node26112;
	wire [16-1:0] node26113;
	wire [16-1:0] node26117;
	wire [16-1:0] node26119;
	wire [16-1:0] node26122;
	wire [16-1:0] node26123;
	wire [16-1:0] node26124;
	wire [16-1:0] node26127;
	wire [16-1:0] node26129;
	wire [16-1:0] node26132;
	wire [16-1:0] node26133;
	wire [16-1:0] node26137;
	wire [16-1:0] node26138;
	wire [16-1:0] node26139;
	wire [16-1:0] node26140;
	wire [16-1:0] node26141;
	wire [16-1:0] node26145;
	wire [16-1:0] node26148;
	wire [16-1:0] node26149;
	wire [16-1:0] node26150;
	wire [16-1:0] node26154;
	wire [16-1:0] node26157;
	wire [16-1:0] node26158;
	wire [16-1:0] node26159;
	wire [16-1:0] node26162;
	wire [16-1:0] node26164;
	wire [16-1:0] node26168;
	wire [16-1:0] node26169;
	wire [16-1:0] node26170;
	wire [16-1:0] node26171;
	wire [16-1:0] node26173;
	wire [16-1:0] node26175;
	wire [16-1:0] node26178;
	wire [16-1:0] node26179;
	wire [16-1:0] node26183;
	wire [16-1:0] node26184;
	wire [16-1:0] node26185;
	wire [16-1:0] node26187;
	wire [16-1:0] node26190;
	wire [16-1:0] node26191;
	wire [16-1:0] node26195;
	wire [16-1:0] node26196;
	wire [16-1:0] node26199;
	wire [16-1:0] node26202;
	wire [16-1:0] node26203;
	wire [16-1:0] node26204;
	wire [16-1:0] node26206;
	wire [16-1:0] node26209;
	wire [16-1:0] node26210;
	wire [16-1:0] node26213;
	wire [16-1:0] node26215;
	wire [16-1:0] node26218;
	wire [16-1:0] node26219;
	wire [16-1:0] node26221;
	wire [16-1:0] node26224;
	wire [16-1:0] node26227;
	wire [16-1:0] node26228;
	wire [16-1:0] node26229;
	wire [16-1:0] node26230;
	wire [16-1:0] node26231;
	wire [16-1:0] node26232;
	wire [16-1:0] node26233;
	wire [16-1:0] node26236;
	wire [16-1:0] node26237;
	wire [16-1:0] node26241;
	wire [16-1:0] node26242;
	wire [16-1:0] node26245;
	wire [16-1:0] node26248;
	wire [16-1:0] node26249;
	wire [16-1:0] node26250;
	wire [16-1:0] node26251;
	wire [16-1:0] node26255;
	wire [16-1:0] node26258;
	wire [16-1:0] node26259;
	wire [16-1:0] node26260;
	wire [16-1:0] node26265;
	wire [16-1:0] node26266;
	wire [16-1:0] node26267;
	wire [16-1:0] node26268;
	wire [16-1:0] node26271;
	wire [16-1:0] node26274;
	wire [16-1:0] node26275;
	wire [16-1:0] node26278;
	wire [16-1:0] node26281;
	wire [16-1:0] node26282;
	wire [16-1:0] node26284;
	wire [16-1:0] node26287;
	wire [16-1:0] node26290;
	wire [16-1:0] node26291;
	wire [16-1:0] node26292;
	wire [16-1:0] node26293;
	wire [16-1:0] node26295;
	wire [16-1:0] node26296;
	wire [16-1:0] node26300;
	wire [16-1:0] node26301;
	wire [16-1:0] node26304;
	wire [16-1:0] node26307;
	wire [16-1:0] node26308;
	wire [16-1:0] node26309;
	wire [16-1:0] node26313;
	wire [16-1:0] node26314;
	wire [16-1:0] node26318;
	wire [16-1:0] node26319;
	wire [16-1:0] node26320;
	wire [16-1:0] node26321;
	wire [16-1:0] node26324;
	wire [16-1:0] node26327;
	wire [16-1:0] node26328;
	wire [16-1:0] node26330;
	wire [16-1:0] node26331;
	wire [16-1:0] node26335;
	wire [16-1:0] node26337;
	wire [16-1:0] node26340;
	wire [16-1:0] node26341;
	wire [16-1:0] node26343;
	wire [16-1:0] node26344;
	wire [16-1:0] node26345;
	wire [16-1:0] node26350;
	wire [16-1:0] node26351;
	wire [16-1:0] node26353;
	wire [16-1:0] node26354;
	wire [16-1:0] node26358;
	wire [16-1:0] node26361;
	wire [16-1:0] node26362;
	wire [16-1:0] node26363;
	wire [16-1:0] node26364;
	wire [16-1:0] node26365;
	wire [16-1:0] node26366;
	wire [16-1:0] node26370;
	wire [16-1:0] node26371;
	wire [16-1:0] node26375;
	wire [16-1:0] node26376;
	wire [16-1:0] node26377;
	wire [16-1:0] node26379;
	wire [16-1:0] node26382;
	wire [16-1:0] node26383;
	wire [16-1:0] node26387;
	wire [16-1:0] node26389;
	wire [16-1:0] node26390;
	wire [16-1:0] node26394;
	wire [16-1:0] node26395;
	wire [16-1:0] node26396;
	wire [16-1:0] node26398;
	wire [16-1:0] node26399;
	wire [16-1:0] node26401;
	wire [16-1:0] node26405;
	wire [16-1:0] node26406;
	wire [16-1:0] node26410;
	wire [16-1:0] node26411;
	wire [16-1:0] node26414;
	wire [16-1:0] node26416;
	wire [16-1:0] node26417;
	wire [16-1:0] node26419;
	wire [16-1:0] node26423;
	wire [16-1:0] node26424;
	wire [16-1:0] node26425;
	wire [16-1:0] node26426;
	wire [16-1:0] node26427;
	wire [16-1:0] node26428;
	wire [16-1:0] node26433;
	wire [16-1:0] node26436;
	wire [16-1:0] node26437;
	wire [16-1:0] node26439;
	wire [16-1:0] node26440;
	wire [16-1:0] node26444;
	wire [16-1:0] node26446;
	wire [16-1:0] node26447;
	wire [16-1:0] node26451;
	wire [16-1:0] node26452;
	wire [16-1:0] node26453;
	wire [16-1:0] node26455;
	wire [16-1:0] node26456;
	wire [16-1:0] node26458;
	wire [16-1:0] node26462;
	wire [16-1:0] node26464;
	wire [16-1:0] node26466;
	wire [16-1:0] node26469;
	wire [16-1:0] node26470;
	wire [16-1:0] node26471;
	wire [16-1:0] node26472;
	wire [16-1:0] node26476;
	wire [16-1:0] node26479;
	wire [16-1:0] node26480;
	wire [16-1:0] node26483;
	wire [16-1:0] node26486;
	wire [16-1:0] node26487;
	wire [16-1:0] node26488;
	wire [16-1:0] node26489;
	wire [16-1:0] node26490;
	wire [16-1:0] node26491;
	wire [16-1:0] node26492;
	wire [16-1:0] node26493;
	wire [16-1:0] node26494;
	wire [16-1:0] node26498;
	wire [16-1:0] node26501;
	wire [16-1:0] node26502;
	wire [16-1:0] node26505;
	wire [16-1:0] node26507;
	wire [16-1:0] node26510;
	wire [16-1:0] node26511;
	wire [16-1:0] node26512;
	wire [16-1:0] node26513;
	wire [16-1:0] node26515;
	wire [16-1:0] node26519;
	wire [16-1:0] node26521;
	wire [16-1:0] node26524;
	wire [16-1:0] node26525;
	wire [16-1:0] node26529;
	wire [16-1:0] node26530;
	wire [16-1:0] node26531;
	wire [16-1:0] node26532;
	wire [16-1:0] node26536;
	wire [16-1:0] node26537;
	wire [16-1:0] node26539;
	wire [16-1:0] node26542;
	wire [16-1:0] node26545;
	wire [16-1:0] node26546;
	wire [16-1:0] node26548;
	wire [16-1:0] node26550;
	wire [16-1:0] node26553;
	wire [16-1:0] node26554;
	wire [16-1:0] node26558;
	wire [16-1:0] node26559;
	wire [16-1:0] node26560;
	wire [16-1:0] node26562;
	wire [16-1:0] node26563;
	wire [16-1:0] node26564;
	wire [16-1:0] node26565;
	wire [16-1:0] node26570;
	wire [16-1:0] node26573;
	wire [16-1:0] node26574;
	wire [16-1:0] node26575;
	wire [16-1:0] node26576;
	wire [16-1:0] node26581;
	wire [16-1:0] node26583;
	wire [16-1:0] node26586;
	wire [16-1:0] node26587;
	wire [16-1:0] node26588;
	wire [16-1:0] node26590;
	wire [16-1:0] node26593;
	wire [16-1:0] node26594;
	wire [16-1:0] node26597;
	wire [16-1:0] node26600;
	wire [16-1:0] node26601;
	wire [16-1:0] node26602;
	wire [16-1:0] node26605;
	wire [16-1:0] node26608;
	wire [16-1:0] node26611;
	wire [16-1:0] node26612;
	wire [16-1:0] node26613;
	wire [16-1:0] node26614;
	wire [16-1:0] node26615;
	wire [16-1:0] node26616;
	wire [16-1:0] node26621;
	wire [16-1:0] node26622;
	wire [16-1:0] node26623;
	wire [16-1:0] node26626;
	wire [16-1:0] node26628;
	wire [16-1:0] node26631;
	wire [16-1:0] node26632;
	wire [16-1:0] node26635;
	wire [16-1:0] node26638;
	wire [16-1:0] node26639;
	wire [16-1:0] node26640;
	wire [16-1:0] node26641;
	wire [16-1:0] node26643;
	wire [16-1:0] node26647;
	wire [16-1:0] node26648;
	wire [16-1:0] node26649;
	wire [16-1:0] node26653;
	wire [16-1:0] node26654;
	wire [16-1:0] node26658;
	wire [16-1:0] node26659;
	wire [16-1:0] node26660;
	wire [16-1:0] node26661;
	wire [16-1:0] node26665;
	wire [16-1:0] node26667;
	wire [16-1:0] node26668;
	wire [16-1:0] node26671;
	wire [16-1:0] node26675;
	wire [16-1:0] node26676;
	wire [16-1:0] node26677;
	wire [16-1:0] node26680;
	wire [16-1:0] node26681;
	wire [16-1:0] node26682;
	wire [16-1:0] node26686;
	wire [16-1:0] node26687;
	wire [16-1:0] node26689;
	wire [16-1:0] node26692;
	wire [16-1:0] node26695;
	wire [16-1:0] node26696;
	wire [16-1:0] node26697;
	wire [16-1:0] node26698;
	wire [16-1:0] node26699;
	wire [16-1:0] node26704;
	wire [16-1:0] node26705;
	wire [16-1:0] node26706;
	wire [16-1:0] node26710;
	wire [16-1:0] node26713;
	wire [16-1:0] node26714;
	wire [16-1:0] node26715;
	wire [16-1:0] node26719;
	wire [16-1:0] node26720;
	wire [16-1:0] node26721;
	wire [16-1:0] node26724;
	wire [16-1:0] node26728;
	wire [16-1:0] node26729;
	wire [16-1:0] node26730;
	wire [16-1:0] node26731;
	wire [16-1:0] node26732;
	wire [16-1:0] node26733;
	wire [16-1:0] node26734;
	wire [16-1:0] node26738;
	wire [16-1:0] node26739;
	wire [16-1:0] node26742;
	wire [16-1:0] node26743;
	wire [16-1:0] node26745;
	wire [16-1:0] node26749;
	wire [16-1:0] node26750;
	wire [16-1:0] node26752;
	wire [16-1:0] node26754;
	wire [16-1:0] node26755;
	wire [16-1:0] node26760;
	wire [16-1:0] node26761;
	wire [16-1:0] node26762;
	wire [16-1:0] node26763;
	wire [16-1:0] node26766;
	wire [16-1:0] node26769;
	wire [16-1:0] node26770;
	wire [16-1:0] node26771;
	wire [16-1:0] node26773;
	wire [16-1:0] node26776;
	wire [16-1:0] node26778;
	wire [16-1:0] node26782;
	wire [16-1:0] node26783;
	wire [16-1:0] node26784;
	wire [16-1:0] node26787;
	wire [16-1:0] node26790;
	wire [16-1:0] node26791;
	wire [16-1:0] node26792;
	wire [16-1:0] node26796;
	wire [16-1:0] node26799;
	wire [16-1:0] node26800;
	wire [16-1:0] node26801;
	wire [16-1:0] node26802;
	wire [16-1:0] node26803;
	wire [16-1:0] node26806;
	wire [16-1:0] node26809;
	wire [16-1:0] node26811;
	wire [16-1:0] node26814;
	wire [16-1:0] node26816;
	wire [16-1:0] node26817;
	wire [16-1:0] node26818;
	wire [16-1:0] node26820;
	wire [16-1:0] node26825;
	wire [16-1:0] node26826;
	wire [16-1:0] node26828;
	wire [16-1:0] node26831;
	wire [16-1:0] node26832;
	wire [16-1:0] node26833;
	wire [16-1:0] node26835;
	wire [16-1:0] node26836;
	wire [16-1:0] node26840;
	wire [16-1:0] node26843;
	wire [16-1:0] node26845;
	wire [16-1:0] node26847;
	wire [16-1:0] node26850;
	wire [16-1:0] node26851;
	wire [16-1:0] node26852;
	wire [16-1:0] node26853;
	wire [16-1:0] node26854;
	wire [16-1:0] node26855;
	wire [16-1:0] node26857;
	wire [16-1:0] node26861;
	wire [16-1:0] node26862;
	wire [16-1:0] node26866;
	wire [16-1:0] node26867;
	wire [16-1:0] node26869;
	wire [16-1:0] node26870;
	wire [16-1:0] node26872;
	wire [16-1:0] node26877;
	wire [16-1:0] node26878;
	wire [16-1:0] node26879;
	wire [16-1:0] node26881;
	wire [16-1:0] node26884;
	wire [16-1:0] node26885;
	wire [16-1:0] node26886;
	wire [16-1:0] node26889;
	wire [16-1:0] node26890;
	wire [16-1:0] node26894;
	wire [16-1:0] node26897;
	wire [16-1:0] node26898;
	wire [16-1:0] node26899;
	wire [16-1:0] node26902;
	wire [16-1:0] node26905;
	wire [16-1:0] node26906;
	wire [16-1:0] node26907;
	wire [16-1:0] node26909;
	wire [16-1:0] node26912;
	wire [16-1:0] node26913;
	wire [16-1:0] node26917;
	wire [16-1:0] node26919;
	wire [16-1:0] node26922;
	wire [16-1:0] node26923;
	wire [16-1:0] node26924;
	wire [16-1:0] node26925;
	wire [16-1:0] node26927;
	wire [16-1:0] node26930;
	wire [16-1:0] node26931;
	wire [16-1:0] node26933;
	wire [16-1:0] node26936;
	wire [16-1:0] node26939;
	wire [16-1:0] node26940;
	wire [16-1:0] node26941;
	wire [16-1:0] node26944;
	wire [16-1:0] node26946;
	wire [16-1:0] node26948;
	wire [16-1:0] node26951;
	wire [16-1:0] node26953;
	wire [16-1:0] node26955;
	wire [16-1:0] node26958;
	wire [16-1:0] node26959;
	wire [16-1:0] node26960;
	wire [16-1:0] node26961;
	wire [16-1:0] node26964;
	wire [16-1:0] node26965;
	wire [16-1:0] node26969;
	wire [16-1:0] node26970;
	wire [16-1:0] node26974;
	wire [16-1:0] node26975;
	wire [16-1:0] node26977;
	wire [16-1:0] node26979;
	wire [16-1:0] node26982;
	wire [16-1:0] node26984;
	wire [16-1:0] node26985;
	wire [16-1:0] node26989;
	wire [16-1:0] node26990;
	wire [16-1:0] node26991;
	wire [16-1:0] node26992;
	wire [16-1:0] node26993;
	wire [16-1:0] node26994;
	wire [16-1:0] node26995;
	wire [16-1:0] node26996;
	wire [16-1:0] node26997;
	wire [16-1:0] node26998;
	wire [16-1:0] node27001;
	wire [16-1:0] node27002;
	wire [16-1:0] node27004;
	wire [16-1:0] node27008;
	wire [16-1:0] node27009;
	wire [16-1:0] node27012;
	wire [16-1:0] node27015;
	wire [16-1:0] node27016;
	wire [16-1:0] node27017;
	wire [16-1:0] node27020;
	wire [16-1:0] node27023;
	wire [16-1:0] node27024;
	wire [16-1:0] node27027;
	wire [16-1:0] node27029;
	wire [16-1:0] node27032;
	wire [16-1:0] node27033;
	wire [16-1:0] node27034;
	wire [16-1:0] node27035;
	wire [16-1:0] node27039;
	wire [16-1:0] node27040;
	wire [16-1:0] node27043;
	wire [16-1:0] node27046;
	wire [16-1:0] node27047;
	wire [16-1:0] node27048;
	wire [16-1:0] node27051;
	wire [16-1:0] node27054;
	wire [16-1:0] node27055;
	wire [16-1:0] node27056;
	wire [16-1:0] node27060;
	wire [16-1:0] node27063;
	wire [16-1:0] node27064;
	wire [16-1:0] node27065;
	wire [16-1:0] node27066;
	wire [16-1:0] node27067;
	wire [16-1:0] node27071;
	wire [16-1:0] node27073;
	wire [16-1:0] node27076;
	wire [16-1:0] node27078;
	wire [16-1:0] node27079;
	wire [16-1:0] node27082;
	wire [16-1:0] node27083;
	wire [16-1:0] node27084;
	wire [16-1:0] node27089;
	wire [16-1:0] node27090;
	wire [16-1:0] node27091;
	wire [16-1:0] node27093;
	wire [16-1:0] node27096;
	wire [16-1:0] node27097;
	wire [16-1:0] node27101;
	wire [16-1:0] node27102;
	wire [16-1:0] node27103;
	wire [16-1:0] node27106;
	wire [16-1:0] node27109;
	wire [16-1:0] node27110;
	wire [16-1:0] node27113;
	wire [16-1:0] node27116;
	wire [16-1:0] node27117;
	wire [16-1:0] node27118;
	wire [16-1:0] node27119;
	wire [16-1:0] node27121;
	wire [16-1:0] node27122;
	wire [16-1:0] node27125;
	wire [16-1:0] node27127;
	wire [16-1:0] node27130;
	wire [16-1:0] node27131;
	wire [16-1:0] node27132;
	wire [16-1:0] node27133;
	wire [16-1:0] node27137;
	wire [16-1:0] node27139;
	wire [16-1:0] node27142;
	wire [16-1:0] node27143;
	wire [16-1:0] node27145;
	wire [16-1:0] node27149;
	wire [16-1:0] node27150;
	wire [16-1:0] node27151;
	wire [16-1:0] node27154;
	wire [16-1:0] node27155;
	wire [16-1:0] node27156;
	wire [16-1:0] node27158;
	wire [16-1:0] node27163;
	wire [16-1:0] node27164;
	wire [16-1:0] node27166;
	wire [16-1:0] node27167;
	wire [16-1:0] node27171;
	wire [16-1:0] node27172;
	wire [16-1:0] node27174;
	wire [16-1:0] node27178;
	wire [16-1:0] node27179;
	wire [16-1:0] node27180;
	wire [16-1:0] node27181;
	wire [16-1:0] node27182;
	wire [16-1:0] node27184;
	wire [16-1:0] node27188;
	wire [16-1:0] node27189;
	wire [16-1:0] node27191;
	wire [16-1:0] node27194;
	wire [16-1:0] node27196;
	wire [16-1:0] node27199;
	wire [16-1:0] node27201;
	wire [16-1:0] node27202;
	wire [16-1:0] node27203;
	wire [16-1:0] node27207;
	wire [16-1:0] node27208;
	wire [16-1:0] node27212;
	wire [16-1:0] node27213;
	wire [16-1:0] node27214;
	wire [16-1:0] node27215;
	wire [16-1:0] node27218;
	wire [16-1:0] node27221;
	wire [16-1:0] node27222;
	wire [16-1:0] node27224;
	wire [16-1:0] node27225;
	wire [16-1:0] node27229;
	wire [16-1:0] node27232;
	wire [16-1:0] node27233;
	wire [16-1:0] node27235;
	wire [16-1:0] node27237;
	wire [16-1:0] node27240;
	wire [16-1:0] node27242;
	wire [16-1:0] node27245;
	wire [16-1:0] node27246;
	wire [16-1:0] node27247;
	wire [16-1:0] node27248;
	wire [16-1:0] node27249;
	wire [16-1:0] node27250;
	wire [16-1:0] node27251;
	wire [16-1:0] node27254;
	wire [16-1:0] node27257;
	wire [16-1:0] node27258;
	wire [16-1:0] node27261;
	wire [16-1:0] node27264;
	wire [16-1:0] node27266;
	wire [16-1:0] node27268;
	wire [16-1:0] node27269;
	wire [16-1:0] node27273;
	wire [16-1:0] node27274;
	wire [16-1:0] node27275;
	wire [16-1:0] node27277;
	wire [16-1:0] node27280;
	wire [16-1:0] node27283;
	wire [16-1:0] node27284;
	wire [16-1:0] node27285;
	wire [16-1:0] node27288;
	wire [16-1:0] node27291;
	wire [16-1:0] node27292;
	wire [16-1:0] node27295;
	wire [16-1:0] node27296;
	wire [16-1:0] node27298;
	wire [16-1:0] node27302;
	wire [16-1:0] node27303;
	wire [16-1:0] node27304;
	wire [16-1:0] node27305;
	wire [16-1:0] node27306;
	wire [16-1:0] node27307;
	wire [16-1:0] node27312;
	wire [16-1:0] node27313;
	wire [16-1:0] node27314;
	wire [16-1:0] node27318;
	wire [16-1:0] node27321;
	wire [16-1:0] node27323;
	wire [16-1:0] node27324;
	wire [16-1:0] node27327;
	wire [16-1:0] node27329;
	wire [16-1:0] node27332;
	wire [16-1:0] node27333;
	wire [16-1:0] node27334;
	wire [16-1:0] node27335;
	wire [16-1:0] node27336;
	wire [16-1:0] node27340;
	wire [16-1:0] node27341;
	wire [16-1:0] node27345;
	wire [16-1:0] node27348;
	wire [16-1:0] node27350;
	wire [16-1:0] node27351;
	wire [16-1:0] node27352;
	wire [16-1:0] node27354;
	wire [16-1:0] node27357;
	wire [16-1:0] node27358;
	wire [16-1:0] node27362;
	wire [16-1:0] node27365;
	wire [16-1:0] node27366;
	wire [16-1:0] node27367;
	wire [16-1:0] node27368;
	wire [16-1:0] node27369;
	wire [16-1:0] node27371;
	wire [16-1:0] node27374;
	wire [16-1:0] node27376;
	wire [16-1:0] node27379;
	wire [16-1:0] node27380;
	wire [16-1:0] node27381;
	wire [16-1:0] node27382;
	wire [16-1:0] node27386;
	wire [16-1:0] node27388;
	wire [16-1:0] node27389;
	wire [16-1:0] node27394;
	wire [16-1:0] node27395;
	wire [16-1:0] node27396;
	wire [16-1:0] node27397;
	wire [16-1:0] node27400;
	wire [16-1:0] node27401;
	wire [16-1:0] node27403;
	wire [16-1:0] node27406;
	wire [16-1:0] node27407;
	wire [16-1:0] node27411;
	wire [16-1:0] node27412;
	wire [16-1:0] node27413;
	wire [16-1:0] node27418;
	wire [16-1:0] node27419;
	wire [16-1:0] node27420;
	wire [16-1:0] node27422;
	wire [16-1:0] node27425;
	wire [16-1:0] node27426;
	wire [16-1:0] node27430;
	wire [16-1:0] node27432;
	wire [16-1:0] node27434;
	wire [16-1:0] node27437;
	wire [16-1:0] node27438;
	wire [16-1:0] node27439;
	wire [16-1:0] node27440;
	wire [16-1:0] node27443;
	wire [16-1:0] node27445;
	wire [16-1:0] node27447;
	wire [16-1:0] node27450;
	wire [16-1:0] node27451;
	wire [16-1:0] node27452;
	wire [16-1:0] node27455;
	wire [16-1:0] node27459;
	wire [16-1:0] node27460;
	wire [16-1:0] node27461;
	wire [16-1:0] node27463;
	wire [16-1:0] node27466;
	wire [16-1:0] node27467;
	wire [16-1:0] node27470;
	wire [16-1:0] node27472;
	wire [16-1:0] node27475;
	wire [16-1:0] node27476;
	wire [16-1:0] node27479;
	wire [16-1:0] node27481;
	wire [16-1:0] node27482;
	wire [16-1:0] node27486;
	wire [16-1:0] node27487;
	wire [16-1:0] node27488;
	wire [16-1:0] node27489;
	wire [16-1:0] node27490;
	wire [16-1:0] node27491;
	wire [16-1:0] node27492;
	wire [16-1:0] node27493;
	wire [16-1:0] node27495;
	wire [16-1:0] node27498;
	wire [16-1:0] node27499;
	wire [16-1:0] node27500;
	wire [16-1:0] node27505;
	wire [16-1:0] node27507;
	wire [16-1:0] node27510;
	wire [16-1:0] node27511;
	wire [16-1:0] node27513;
	wire [16-1:0] node27514;
	wire [16-1:0] node27515;
	wire [16-1:0] node27520;
	wire [16-1:0] node27521;
	wire [16-1:0] node27522;
	wire [16-1:0] node27527;
	wire [16-1:0] node27528;
	wire [16-1:0] node27529;
	wire [16-1:0] node27530;
	wire [16-1:0] node27532;
	wire [16-1:0] node27534;
	wire [16-1:0] node27537;
	wire [16-1:0] node27538;
	wire [16-1:0] node27542;
	wire [16-1:0] node27543;
	wire [16-1:0] node27544;
	wire [16-1:0] node27549;
	wire [16-1:0] node27550;
	wire [16-1:0] node27552;
	wire [16-1:0] node27555;
	wire [16-1:0] node27556;
	wire [16-1:0] node27557;
	wire [16-1:0] node27562;
	wire [16-1:0] node27563;
	wire [16-1:0] node27564;
	wire [16-1:0] node27565;
	wire [16-1:0] node27567;
	wire [16-1:0] node27569;
	wire [16-1:0] node27570;
	wire [16-1:0] node27574;
	wire [16-1:0] node27575;
	wire [16-1:0] node27579;
	wire [16-1:0] node27580;
	wire [16-1:0] node27582;
	wire [16-1:0] node27584;
	wire [16-1:0] node27585;
	wire [16-1:0] node27589;
	wire [16-1:0] node27590;
	wire [16-1:0] node27593;
	wire [16-1:0] node27595;
	wire [16-1:0] node27598;
	wire [16-1:0] node27599;
	wire [16-1:0] node27600;
	wire [16-1:0] node27601;
	wire [16-1:0] node27604;
	wire [16-1:0] node27607;
	wire [16-1:0] node27608;
	wire [16-1:0] node27611;
	wire [16-1:0] node27614;
	wire [16-1:0] node27615;
	wire [16-1:0] node27616;
	wire [16-1:0] node27619;
	wire [16-1:0] node27621;
	wire [16-1:0] node27624;
	wire [16-1:0] node27626;
	wire [16-1:0] node27629;
	wire [16-1:0] node27630;
	wire [16-1:0] node27631;
	wire [16-1:0] node27632;
	wire [16-1:0] node27633;
	wire [16-1:0] node27634;
	wire [16-1:0] node27638;
	wire [16-1:0] node27639;
	wire [16-1:0] node27642;
	wire [16-1:0] node27645;
	wire [16-1:0] node27646;
	wire [16-1:0] node27647;
	wire [16-1:0] node27648;
	wire [16-1:0] node27652;
	wire [16-1:0] node27655;
	wire [16-1:0] node27656;
	wire [16-1:0] node27660;
	wire [16-1:0] node27661;
	wire [16-1:0] node27663;
	wire [16-1:0] node27666;
	wire [16-1:0] node27667;
	wire [16-1:0] node27668;
	wire [16-1:0] node27670;
	wire [16-1:0] node27672;
	wire [16-1:0] node27675;
	wire [16-1:0] node27678;
	wire [16-1:0] node27679;
	wire [16-1:0] node27682;
	wire [16-1:0] node27685;
	wire [16-1:0] node27686;
	wire [16-1:0] node27687;
	wire [16-1:0] node27688;
	wire [16-1:0] node27689;
	wire [16-1:0] node27691;
	wire [16-1:0] node27693;
	wire [16-1:0] node27697;
	wire [16-1:0] node27698;
	wire [16-1:0] node27701;
	wire [16-1:0] node27704;
	wire [16-1:0] node27705;
	wire [16-1:0] node27706;
	wire [16-1:0] node27709;
	wire [16-1:0] node27710;
	wire [16-1:0] node27715;
	wire [16-1:0] node27716;
	wire [16-1:0] node27717;
	wire [16-1:0] node27718;
	wire [16-1:0] node27719;
	wire [16-1:0] node27723;
	wire [16-1:0] node27726;
	wire [16-1:0] node27727;
	wire [16-1:0] node27728;
	wire [16-1:0] node27732;
	wire [16-1:0] node27735;
	wire [16-1:0] node27736;
	wire [16-1:0] node27738;
	wire [16-1:0] node27739;
	wire [16-1:0] node27743;
	wire [16-1:0] node27745;
	wire [16-1:0] node27747;
	wire [16-1:0] node27750;
	wire [16-1:0] node27751;
	wire [16-1:0] node27752;
	wire [16-1:0] node27753;
	wire [16-1:0] node27754;
	wire [16-1:0] node27755;
	wire [16-1:0] node27757;
	wire [16-1:0] node27760;
	wire [16-1:0] node27761;
	wire [16-1:0] node27763;
	wire [16-1:0] node27766;
	wire [16-1:0] node27769;
	wire [16-1:0] node27770;
	wire [16-1:0] node27772;
	wire [16-1:0] node27774;
	wire [16-1:0] node27777;
	wire [16-1:0] node27778;
	wire [16-1:0] node27780;
	wire [16-1:0] node27781;
	wire [16-1:0] node27785;
	wire [16-1:0] node27788;
	wire [16-1:0] node27789;
	wire [16-1:0] node27790;
	wire [16-1:0] node27792;
	wire [16-1:0] node27794;
	wire [16-1:0] node27797;
	wire [16-1:0] node27798;
	wire [16-1:0] node27801;
	wire [16-1:0] node27804;
	wire [16-1:0] node27805;
	wire [16-1:0] node27807;
	wire [16-1:0] node27808;
	wire [16-1:0] node27812;
	wire [16-1:0] node27815;
	wire [16-1:0] node27816;
	wire [16-1:0] node27817;
	wire [16-1:0] node27818;
	wire [16-1:0] node27819;
	wire [16-1:0] node27820;
	wire [16-1:0] node27824;
	wire [16-1:0] node27827;
	wire [16-1:0] node27828;
	wire [16-1:0] node27829;
	wire [16-1:0] node27831;
	wire [16-1:0] node27835;
	wire [16-1:0] node27838;
	wire [16-1:0] node27839;
	wire [16-1:0] node27840;
	wire [16-1:0] node27841;
	wire [16-1:0] node27843;
	wire [16-1:0] node27847;
	wire [16-1:0] node27850;
	wire [16-1:0] node27851;
	wire [16-1:0] node27852;
	wire [16-1:0] node27857;
	wire [16-1:0] node27858;
	wire [16-1:0] node27859;
	wire [16-1:0] node27860;
	wire [16-1:0] node27861;
	wire [16-1:0] node27865;
	wire [16-1:0] node27868;
	wire [16-1:0] node27869;
	wire [16-1:0] node27871;
	wire [16-1:0] node27872;
	wire [16-1:0] node27876;
	wire [16-1:0] node27877;
	wire [16-1:0] node27880;
	wire [16-1:0] node27881;
	wire [16-1:0] node27885;
	wire [16-1:0] node27886;
	wire [16-1:0] node27887;
	wire [16-1:0] node27891;
	wire [16-1:0] node27892;
	wire [16-1:0] node27895;
	wire [16-1:0] node27897;
	wire [16-1:0] node27900;
	wire [16-1:0] node27901;
	wire [16-1:0] node27902;
	wire [16-1:0] node27903;
	wire [16-1:0] node27905;
	wire [16-1:0] node27906;
	wire [16-1:0] node27909;
	wire [16-1:0] node27912;
	wire [16-1:0] node27913;
	wire [16-1:0] node27915;
	wire [16-1:0] node27918;
	wire [16-1:0] node27919;
	wire [16-1:0] node27922;
	wire [16-1:0] node27925;
	wire [16-1:0] node27926;
	wire [16-1:0] node27927;
	wire [16-1:0] node27929;
	wire [16-1:0] node27931;
	wire [16-1:0] node27934;
	wire [16-1:0] node27936;
	wire [16-1:0] node27939;
	wire [16-1:0] node27940;
	wire [16-1:0] node27942;
	wire [16-1:0] node27943;
	wire [16-1:0] node27947;
	wire [16-1:0] node27949;
	wire [16-1:0] node27950;
	wire [16-1:0] node27952;
	wire [16-1:0] node27956;
	wire [16-1:0] node27957;
	wire [16-1:0] node27958;
	wire [16-1:0] node27960;
	wire [16-1:0] node27961;
	wire [16-1:0] node27962;
	wire [16-1:0] node27964;
	wire [16-1:0] node27968;
	wire [16-1:0] node27970;
	wire [16-1:0] node27972;
	wire [16-1:0] node27975;
	wire [16-1:0] node27976;
	wire [16-1:0] node27977;
	wire [16-1:0] node27979;
	wire [16-1:0] node27983;
	wire [16-1:0] node27985;
	wire [16-1:0] node27986;
	wire [16-1:0] node27990;
	wire [16-1:0] node27991;
	wire [16-1:0] node27992;
	wire [16-1:0] node27993;
	wire [16-1:0] node27995;
	wire [16-1:0] node27999;
	wire [16-1:0] node28002;
	wire [16-1:0] node28003;
	wire [16-1:0] node28004;
	wire [16-1:0] node28008;
	wire [16-1:0] node28010;
	wire [16-1:0] node28011;
	wire [16-1:0] node28014;
	wire [16-1:0] node28017;
	wire [16-1:0] node28018;
	wire [16-1:0] node28019;
	wire [16-1:0] node28020;
	wire [16-1:0] node28021;
	wire [16-1:0] node28022;
	wire [16-1:0] node28023;
	wire [16-1:0] node28024;
	wire [16-1:0] node28025;
	wire [16-1:0] node28029;
	wire [16-1:0] node28030;
	wire [16-1:0] node28033;
	wire [16-1:0] node28036;
	wire [16-1:0] node28037;
	wire [16-1:0] node28039;
	wire [16-1:0] node28041;
	wire [16-1:0] node28044;
	wire [16-1:0] node28045;
	wire [16-1:0] node28047;
	wire [16-1:0] node28048;
	wire [16-1:0] node28052;
	wire [16-1:0] node28054;
	wire [16-1:0] node28057;
	wire [16-1:0] node28058;
	wire [16-1:0] node28059;
	wire [16-1:0] node28060;
	wire [16-1:0] node28062;
	wire [16-1:0] node28065;
	wire [16-1:0] node28067;
	wire [16-1:0] node28070;
	wire [16-1:0] node28071;
	wire [16-1:0] node28075;
	wire [16-1:0] node28076;
	wire [16-1:0] node28077;
	wire [16-1:0] node28078;
	wire [16-1:0] node28082;
	wire [16-1:0] node28085;
	wire [16-1:0] node28086;
	wire [16-1:0] node28090;
	wire [16-1:0] node28091;
	wire [16-1:0] node28092;
	wire [16-1:0] node28093;
	wire [16-1:0] node28094;
	wire [16-1:0] node28097;
	wire [16-1:0] node28100;
	wire [16-1:0] node28101;
	wire [16-1:0] node28104;
	wire [16-1:0] node28107;
	wire [16-1:0] node28109;
	wire [16-1:0] node28110;
	wire [16-1:0] node28111;
	wire [16-1:0] node28116;
	wire [16-1:0] node28117;
	wire [16-1:0] node28118;
	wire [16-1:0] node28119;
	wire [16-1:0] node28120;
	wire [16-1:0] node28124;
	wire [16-1:0] node28126;
	wire [16-1:0] node28127;
	wire [16-1:0] node28131;
	wire [16-1:0] node28132;
	wire [16-1:0] node28135;
	wire [16-1:0] node28138;
	wire [16-1:0] node28139;
	wire [16-1:0] node28140;
	wire [16-1:0] node28144;
	wire [16-1:0] node28145;
	wire [16-1:0] node28148;
	wire [16-1:0] node28150;
	wire [16-1:0] node28151;
	wire [16-1:0] node28155;
	wire [16-1:0] node28156;
	wire [16-1:0] node28157;
	wire [16-1:0] node28158;
	wire [16-1:0] node28159;
	wire [16-1:0] node28160;
	wire [16-1:0] node28164;
	wire [16-1:0] node28165;
	wire [16-1:0] node28168;
	wire [16-1:0] node28171;
	wire [16-1:0] node28172;
	wire [16-1:0] node28173;
	wire [16-1:0] node28177;
	wire [16-1:0] node28178;
	wire [16-1:0] node28182;
	wire [16-1:0] node28183;
	wire [16-1:0] node28184;
	wire [16-1:0] node28185;
	wire [16-1:0] node28186;
	wire [16-1:0] node28191;
	wire [16-1:0] node28192;
	wire [16-1:0] node28195;
	wire [16-1:0] node28198;
	wire [16-1:0] node28199;
	wire [16-1:0] node28201;
	wire [16-1:0] node28204;
	wire [16-1:0] node28205;
	wire [16-1:0] node28209;
	wire [16-1:0] node28210;
	wire [16-1:0] node28211;
	wire [16-1:0] node28212;
	wire [16-1:0] node28213;
	wire [16-1:0] node28216;
	wire [16-1:0] node28219;
	wire [16-1:0] node28220;
	wire [16-1:0] node28221;
	wire [16-1:0] node28226;
	wire [16-1:0] node28227;
	wire [16-1:0] node28228;
	wire [16-1:0] node28231;
	wire [16-1:0] node28234;
	wire [16-1:0] node28235;
	wire [16-1:0] node28237;
	wire [16-1:0] node28241;
	wire [16-1:0] node28242;
	wire [16-1:0] node28243;
	wire [16-1:0] node28244;
	wire [16-1:0] node28247;
	wire [16-1:0] node28248;
	wire [16-1:0] node28250;
	wire [16-1:0] node28254;
	wire [16-1:0] node28255;
	wire [16-1:0] node28257;
	wire [16-1:0] node28261;
	wire [16-1:0] node28262;
	wire [16-1:0] node28264;
	wire [16-1:0] node28267;
	wire [16-1:0] node28268;
	wire [16-1:0] node28269;
	wire [16-1:0] node28272;
	wire [16-1:0] node28274;
	wire [16-1:0] node28278;
	wire [16-1:0] node28279;
	wire [16-1:0] node28280;
	wire [16-1:0] node28281;
	wire [16-1:0] node28282;
	wire [16-1:0] node28283;
	wire [16-1:0] node28285;
	wire [16-1:0] node28287;
	wire [16-1:0] node28290;
	wire [16-1:0] node28291;
	wire [16-1:0] node28292;
	wire [16-1:0] node28297;
	wire [16-1:0] node28298;
	wire [16-1:0] node28299;
	wire [16-1:0] node28302;
	wire [16-1:0] node28303;
	wire [16-1:0] node28304;
	wire [16-1:0] node28308;
	wire [16-1:0] node28309;
	wire [16-1:0] node28313;
	wire [16-1:0] node28314;
	wire [16-1:0] node28317;
	wire [16-1:0] node28320;
	wire [16-1:0] node28321;
	wire [16-1:0] node28322;
	wire [16-1:0] node28323;
	wire [16-1:0] node28327;
	wire [16-1:0] node28328;
	wire [16-1:0] node28329;
	wire [16-1:0] node28331;
	wire [16-1:0] node28336;
	wire [16-1:0] node28337;
	wire [16-1:0] node28338;
	wire [16-1:0] node28341;
	wire [16-1:0] node28344;
	wire [16-1:0] node28346;
	wire [16-1:0] node28347;
	wire [16-1:0] node28351;
	wire [16-1:0] node28352;
	wire [16-1:0] node28353;
	wire [16-1:0] node28354;
	wire [16-1:0] node28355;
	wire [16-1:0] node28359;
	wire [16-1:0] node28360;
	wire [16-1:0] node28363;
	wire [16-1:0] node28364;
	wire [16-1:0] node28367;
	wire [16-1:0] node28368;
	wire [16-1:0] node28372;
	wire [16-1:0] node28373;
	wire [16-1:0] node28375;
	wire [16-1:0] node28378;
	wire [16-1:0] node28379;
	wire [16-1:0] node28382;
	wire [16-1:0] node28385;
	wire [16-1:0] node28386;
	wire [16-1:0] node28387;
	wire [16-1:0] node28388;
	wire [16-1:0] node28390;
	wire [16-1:0] node28393;
	wire [16-1:0] node28395;
	wire [16-1:0] node28398;
	wire [16-1:0] node28399;
	wire [16-1:0] node28400;
	wire [16-1:0] node28404;
	wire [16-1:0] node28407;
	wire [16-1:0] node28408;
	wire [16-1:0] node28411;
	wire [16-1:0] node28412;
	wire [16-1:0] node28415;
	wire [16-1:0] node28418;
	wire [16-1:0] node28419;
	wire [16-1:0] node28420;
	wire [16-1:0] node28421;
	wire [16-1:0] node28422;
	wire [16-1:0] node28423;
	wire [16-1:0] node28425;
	wire [16-1:0] node28428;
	wire [16-1:0] node28429;
	wire [16-1:0] node28433;
	wire [16-1:0] node28434;
	wire [16-1:0] node28437;
	wire [16-1:0] node28438;
	wire [16-1:0] node28442;
	wire [16-1:0] node28443;
	wire [16-1:0] node28444;
	wire [16-1:0] node28445;
	wire [16-1:0] node28447;
	wire [16-1:0] node28451;
	wire [16-1:0] node28452;
	wire [16-1:0] node28454;
	wire [16-1:0] node28458;
	wire [16-1:0] node28459;
	wire [16-1:0] node28461;
	wire [16-1:0] node28465;
	wire [16-1:0] node28466;
	wire [16-1:0] node28468;
	wire [16-1:0] node28469;
	wire [16-1:0] node28471;
	wire [16-1:0] node28475;
	wire [16-1:0] node28476;
	wire [16-1:0] node28477;
	wire [16-1:0] node28478;
	wire [16-1:0] node28482;
	wire [16-1:0] node28485;
	wire [16-1:0] node28486;
	wire [16-1:0] node28489;
	wire [16-1:0] node28491;
	wire [16-1:0] node28492;
	wire [16-1:0] node28496;
	wire [16-1:0] node28497;
	wire [16-1:0] node28498;
	wire [16-1:0] node28499;
	wire [16-1:0] node28500;
	wire [16-1:0] node28501;
	wire [16-1:0] node28505;
	wire [16-1:0] node28506;
	wire [16-1:0] node28510;
	wire [16-1:0] node28511;
	wire [16-1:0] node28515;
	wire [16-1:0] node28516;
	wire [16-1:0] node28517;
	wire [16-1:0] node28520;
	wire [16-1:0] node28522;
	wire [16-1:0] node28525;
	wire [16-1:0] node28527;
	wire [16-1:0] node28529;
	wire [16-1:0] node28530;
	wire [16-1:0] node28534;
	wire [16-1:0] node28535;
	wire [16-1:0] node28536;
	wire [16-1:0] node28537;
	wire [16-1:0] node28540;
	wire [16-1:0] node28543;
	wire [16-1:0] node28545;
	wire [16-1:0] node28548;
	wire [16-1:0] node28549;
	wire [16-1:0] node28550;
	wire [16-1:0] node28553;
	wire [16-1:0] node28556;
	wire [16-1:0] node28557;
	wire [16-1:0] node28559;
	wire [16-1:0] node28561;
	wire [16-1:0] node28565;
	wire [16-1:0] node28566;
	wire [16-1:0] node28567;
	wire [16-1:0] node28568;
	wire [16-1:0] node28569;
	wire [16-1:0] node28570;
	wire [16-1:0] node28571;
	wire [16-1:0] node28572;
	wire [16-1:0] node28576;
	wire [16-1:0] node28578;
	wire [16-1:0] node28580;
	wire [16-1:0] node28583;
	wire [16-1:0] node28584;
	wire [16-1:0] node28586;
	wire [16-1:0] node28587;
	wire [16-1:0] node28588;
	wire [16-1:0] node28591;
	wire [16-1:0] node28594;
	wire [16-1:0] node28595;
	wire [16-1:0] node28599;
	wire [16-1:0] node28600;
	wire [16-1:0] node28604;
	wire [16-1:0] node28605;
	wire [16-1:0] node28608;
	wire [16-1:0] node28609;
	wire [16-1:0] node28610;
	wire [16-1:0] node28613;
	wire [16-1:0] node28615;
	wire [16-1:0] node28618;
	wire [16-1:0] node28619;
	wire [16-1:0] node28622;
	wire [16-1:0] node28624;
	wire [16-1:0] node28627;
	wire [16-1:0] node28628;
	wire [16-1:0] node28629;
	wire [16-1:0] node28630;
	wire [16-1:0] node28632;
	wire [16-1:0] node28635;
	wire [16-1:0] node28636;
	wire [16-1:0] node28639;
	wire [16-1:0] node28642;
	wire [16-1:0] node28643;
	wire [16-1:0] node28644;
	wire [16-1:0] node28645;
	wire [16-1:0] node28647;
	wire [16-1:0] node28651;
	wire [16-1:0] node28654;
	wire [16-1:0] node28656;
	wire [16-1:0] node28659;
	wire [16-1:0] node28660;
	wire [16-1:0] node28661;
	wire [16-1:0] node28662;
	wire [16-1:0] node28665;
	wire [16-1:0] node28669;
	wire [16-1:0] node28670;
	wire [16-1:0] node28671;
	wire [16-1:0] node28673;
	wire [16-1:0] node28677;
	wire [16-1:0] node28678;
	wire [16-1:0] node28682;
	wire [16-1:0] node28683;
	wire [16-1:0] node28684;
	wire [16-1:0] node28685;
	wire [16-1:0] node28686;
	wire [16-1:0] node28688;
	wire [16-1:0] node28691;
	wire [16-1:0] node28692;
	wire [16-1:0] node28695;
	wire [16-1:0] node28697;
	wire [16-1:0] node28698;
	wire [16-1:0] node28702;
	wire [16-1:0] node28703;
	wire [16-1:0] node28704;
	wire [16-1:0] node28707;
	wire [16-1:0] node28710;
	wire [16-1:0] node28712;
	wire [16-1:0] node28714;
	wire [16-1:0] node28717;
	wire [16-1:0] node28718;
	wire [16-1:0] node28720;
	wire [16-1:0] node28721;
	wire [16-1:0] node28723;
	wire [16-1:0] node28727;
	wire [16-1:0] node28728;
	wire [16-1:0] node28729;
	wire [16-1:0] node28730;
	wire [16-1:0] node28734;
	wire [16-1:0] node28735;
	wire [16-1:0] node28738;
	wire [16-1:0] node28739;
	wire [16-1:0] node28743;
	wire [16-1:0] node28744;
	wire [16-1:0] node28745;
	wire [16-1:0] node28747;
	wire [16-1:0] node28752;
	wire [16-1:0] node28753;
	wire [16-1:0] node28754;
	wire [16-1:0] node28755;
	wire [16-1:0] node28756;
	wire [16-1:0] node28757;
	wire [16-1:0] node28761;
	wire [16-1:0] node28764;
	wire [16-1:0] node28765;
	wire [16-1:0] node28768;
	wire [16-1:0] node28770;
	wire [16-1:0] node28773;
	wire [16-1:0] node28775;
	wire [16-1:0] node28776;
	wire [16-1:0] node28779;
	wire [16-1:0] node28782;
	wire [16-1:0] node28783;
	wire [16-1:0] node28784;
	wire [16-1:0] node28785;
	wire [16-1:0] node28789;
	wire [16-1:0] node28791;
	wire [16-1:0] node28793;
	wire [16-1:0] node28795;
	wire [16-1:0] node28798;
	wire [16-1:0] node28799;
	wire [16-1:0] node28801;
	wire [16-1:0] node28804;
	wire [16-1:0] node28805;
	wire [16-1:0] node28807;
	wire [16-1:0] node28809;
	wire [16-1:0] node28812;
	wire [16-1:0] node28813;
	wire [16-1:0] node28817;
	wire [16-1:0] node28818;
	wire [16-1:0] node28819;
	wire [16-1:0] node28820;
	wire [16-1:0] node28821;
	wire [16-1:0] node28822;
	wire [16-1:0] node28823;
	wire [16-1:0] node28826;
	wire [16-1:0] node28828;
	wire [16-1:0] node28831;
	wire [16-1:0] node28832;
	wire [16-1:0] node28833;
	wire [16-1:0] node28835;
	wire [16-1:0] node28839;
	wire [16-1:0] node28840;
	wire [16-1:0] node28844;
	wire [16-1:0] node28845;
	wire [16-1:0] node28848;
	wire [16-1:0] node28851;
	wire [16-1:0] node28852;
	wire [16-1:0] node28853;
	wire [16-1:0] node28854;
	wire [16-1:0] node28857;
	wire [16-1:0] node28860;
	wire [16-1:0] node28861;
	wire [16-1:0] node28865;
	wire [16-1:0] node28866;
	wire [16-1:0] node28868;
	wire [16-1:0] node28869;
	wire [16-1:0] node28870;
	wire [16-1:0] node28875;
	wire [16-1:0] node28877;
	wire [16-1:0] node28880;
	wire [16-1:0] node28881;
	wire [16-1:0] node28882;
	wire [16-1:0] node28883;
	wire [16-1:0] node28884;
	wire [16-1:0] node28887;
	wire [16-1:0] node28888;
	wire [16-1:0] node28890;
	wire [16-1:0] node28894;
	wire [16-1:0] node28895;
	wire [16-1:0] node28896;
	wire [16-1:0] node28901;
	wire [16-1:0] node28902;
	wire [16-1:0] node28903;
	wire [16-1:0] node28904;
	wire [16-1:0] node28906;
	wire [16-1:0] node28910;
	wire [16-1:0] node28913;
	wire [16-1:0] node28914;
	wire [16-1:0] node28917;
	wire [16-1:0] node28918;
	wire [16-1:0] node28921;
	wire [16-1:0] node28923;
	wire [16-1:0] node28926;
	wire [16-1:0] node28927;
	wire [16-1:0] node28928;
	wire [16-1:0] node28929;
	wire [16-1:0] node28932;
	wire [16-1:0] node28933;
	wire [16-1:0] node28935;
	wire [16-1:0] node28939;
	wire [16-1:0] node28940;
	wire [16-1:0] node28941;
	wire [16-1:0] node28945;
	wire [16-1:0] node28948;
	wire [16-1:0] node28950;
	wire [16-1:0] node28951;
	wire [16-1:0] node28954;
	wire [16-1:0] node28955;
	wire [16-1:0] node28958;
	wire [16-1:0] node28959;
	wire [16-1:0] node28963;
	wire [16-1:0] node28964;
	wire [16-1:0] node28965;
	wire [16-1:0] node28966;
	wire [16-1:0] node28967;
	wire [16-1:0] node28971;
	wire [16-1:0] node28972;
	wire [16-1:0] node28973;
	wire [16-1:0] node28976;
	wire [16-1:0] node28979;
	wire [16-1:0] node28981;
	wire [16-1:0] node28983;
	wire [16-1:0] node28986;
	wire [16-1:0] node28987;
	wire [16-1:0] node28988;
	wire [16-1:0] node28990;
	wire [16-1:0] node28993;
	wire [16-1:0] node28994;
	wire [16-1:0] node28997;
	wire [16-1:0] node28999;
	wire [16-1:0] node29000;
	wire [16-1:0] node29004;
	wire [16-1:0] node29006;
	wire [16-1:0] node29008;
	wire [16-1:0] node29009;
	wire [16-1:0] node29013;
	wire [16-1:0] node29014;
	wire [16-1:0] node29015;
	wire [16-1:0] node29016;
	wire [16-1:0] node29018;
	wire [16-1:0] node29019;
	wire [16-1:0] node29021;
	wire [16-1:0] node29025;
	wire [16-1:0] node29026;
	wire [16-1:0] node29027;
	wire [16-1:0] node29029;
	wire [16-1:0] node29033;
	wire [16-1:0] node29036;
	wire [16-1:0] node29037;
	wire [16-1:0] node29038;
	wire [16-1:0] node29041;
	wire [16-1:0] node29042;
	wire [16-1:0] node29046;
	wire [16-1:0] node29048;
	wire [16-1:0] node29051;
	wire [16-1:0] node29052;
	wire [16-1:0] node29054;
	wire [16-1:0] node29056;
	wire [16-1:0] node29058;
	wire [16-1:0] node29061;
	wire [16-1:0] node29062;
	wire [16-1:0] node29063;
	wire [16-1:0] node29066;
	wire [16-1:0] node29067;
	wire [16-1:0] node29069;
	wire [16-1:0] node29073;
	wire [16-1:0] node29074;
	wire [16-1:0] node29077;
	wire [16-1:0] node29079;
	wire [16-1:0] node29082;
	wire [16-1:0] node29083;
	wire [16-1:0] node29084;
	wire [16-1:0] node29085;
	wire [16-1:0] node29086;
	wire [16-1:0] node29087;
	wire [16-1:0] node29088;
	wire [16-1:0] node29089;
	wire [16-1:0] node29090;
	wire [16-1:0] node29091;
	wire [16-1:0] node29093;
	wire [16-1:0] node29094;
	wire [16-1:0] node29096;
	wire [16-1:0] node29100;
	wire [16-1:0] node29101;
	wire [16-1:0] node29102;
	wire [16-1:0] node29104;
	wire [16-1:0] node29109;
	wire [16-1:0] node29110;
	wire [16-1:0] node29111;
	wire [16-1:0] node29112;
	wire [16-1:0] node29114;
	wire [16-1:0] node29118;
	wire [16-1:0] node29120;
	wire [16-1:0] node29123;
	wire [16-1:0] node29124;
	wire [16-1:0] node29125;
	wire [16-1:0] node29126;
	wire [16-1:0] node29131;
	wire [16-1:0] node29132;
	wire [16-1:0] node29136;
	wire [16-1:0] node29137;
	wire [16-1:0] node29138;
	wire [16-1:0] node29139;
	wire [16-1:0] node29143;
	wire [16-1:0] node29144;
	wire [16-1:0] node29146;
	wire [16-1:0] node29147;
	wire [16-1:0] node29152;
	wire [16-1:0] node29153;
	wire [16-1:0] node29154;
	wire [16-1:0] node29155;
	wire [16-1:0] node29159;
	wire [16-1:0] node29161;
	wire [16-1:0] node29164;
	wire [16-1:0] node29165;
	wire [16-1:0] node29168;
	wire [16-1:0] node29171;
	wire [16-1:0] node29172;
	wire [16-1:0] node29173;
	wire [16-1:0] node29175;
	wire [16-1:0] node29176;
	wire [16-1:0] node29179;
	wire [16-1:0] node29181;
	wire [16-1:0] node29184;
	wire [16-1:0] node29185;
	wire [16-1:0] node29187;
	wire [16-1:0] node29190;
	wire [16-1:0] node29191;
	wire [16-1:0] node29195;
	wire [16-1:0] node29196;
	wire [16-1:0] node29197;
	wire [16-1:0] node29199;
	wire [16-1:0] node29202;
	wire [16-1:0] node29204;
	wire [16-1:0] node29207;
	wire [16-1:0] node29208;
	wire [16-1:0] node29209;
	wire [16-1:0] node29212;
	wire [16-1:0] node29214;
	wire [16-1:0] node29217;
	wire [16-1:0] node29218;
	wire [16-1:0] node29219;
	wire [16-1:0] node29224;
	wire [16-1:0] node29225;
	wire [16-1:0] node29226;
	wire [16-1:0] node29227;
	wire [16-1:0] node29228;
	wire [16-1:0] node29229;
	wire [16-1:0] node29233;
	wire [16-1:0] node29235;
	wire [16-1:0] node29238;
	wire [16-1:0] node29239;
	wire [16-1:0] node29241;
	wire [16-1:0] node29243;
	wire [16-1:0] node29246;
	wire [16-1:0] node29249;
	wire [16-1:0] node29250;
	wire [16-1:0] node29251;
	wire [16-1:0] node29252;
	wire [16-1:0] node29254;
	wire [16-1:0] node29257;
	wire [16-1:0] node29259;
	wire [16-1:0] node29260;
	wire [16-1:0] node29264;
	wire [16-1:0] node29265;
	wire [16-1:0] node29268;
	wire [16-1:0] node29270;
	wire [16-1:0] node29271;
	wire [16-1:0] node29275;
	wire [16-1:0] node29276;
	wire [16-1:0] node29279;
	wire [16-1:0] node29281;
	wire [16-1:0] node29282;
	wire [16-1:0] node29286;
	wire [16-1:0] node29287;
	wire [16-1:0] node29288;
	wire [16-1:0] node29289;
	wire [16-1:0] node29290;
	wire [16-1:0] node29291;
	wire [16-1:0] node29295;
	wire [16-1:0] node29298;
	wire [16-1:0] node29299;
	wire [16-1:0] node29303;
	wire [16-1:0] node29304;
	wire [16-1:0] node29305;
	wire [16-1:0] node29306;
	wire [16-1:0] node29310;
	wire [16-1:0] node29313;
	wire [16-1:0] node29316;
	wire [16-1:0] node29317;
	wire [16-1:0] node29318;
	wire [16-1:0] node29320;
	wire [16-1:0] node29323;
	wire [16-1:0] node29324;
	wire [16-1:0] node29328;
	wire [16-1:0] node29329;
	wire [16-1:0] node29330;
	wire [16-1:0] node29333;
	wire [16-1:0] node29334;
	wire [16-1:0] node29338;
	wire [16-1:0] node29340;
	wire [16-1:0] node29341;
	wire [16-1:0] node29343;
	wire [16-1:0] node29346;
	wire [16-1:0] node29349;
	wire [16-1:0] node29350;
	wire [16-1:0] node29351;
	wire [16-1:0] node29352;
	wire [16-1:0] node29353;
	wire [16-1:0] node29354;
	wire [16-1:0] node29356;
	wire [16-1:0] node29357;
	wire [16-1:0] node29358;
	wire [16-1:0] node29364;
	wire [16-1:0] node29365;
	wire [16-1:0] node29366;
	wire [16-1:0] node29368;
	wire [16-1:0] node29369;
	wire [16-1:0] node29373;
	wire [16-1:0] node29375;
	wire [16-1:0] node29376;
	wire [16-1:0] node29380;
	wire [16-1:0] node29382;
	wire [16-1:0] node29385;
	wire [16-1:0] node29386;
	wire [16-1:0] node29387;
	wire [16-1:0] node29388;
	wire [16-1:0] node29391;
	wire [16-1:0] node29394;
	wire [16-1:0] node29395;
	wire [16-1:0] node29399;
	wire [16-1:0] node29401;
	wire [16-1:0] node29402;
	wire [16-1:0] node29404;
	wire [16-1:0] node29405;
	wire [16-1:0] node29409;
	wire [16-1:0] node29411;
	wire [16-1:0] node29414;
	wire [16-1:0] node29415;
	wire [16-1:0] node29416;
	wire [16-1:0] node29417;
	wire [16-1:0] node29419;
	wire [16-1:0] node29421;
	wire [16-1:0] node29424;
	wire [16-1:0] node29425;
	wire [16-1:0] node29426;
	wire [16-1:0] node29430;
	wire [16-1:0] node29433;
	wire [16-1:0] node29434;
	wire [16-1:0] node29436;
	wire [16-1:0] node29437;
	wire [16-1:0] node29441;
	wire [16-1:0] node29443;
	wire [16-1:0] node29446;
	wire [16-1:0] node29447;
	wire [16-1:0] node29448;
	wire [16-1:0] node29450;
	wire [16-1:0] node29451;
	wire [16-1:0] node29453;
	wire [16-1:0] node29457;
	wire [16-1:0] node29458;
	wire [16-1:0] node29459;
	wire [16-1:0] node29464;
	wire [16-1:0] node29466;
	wire [16-1:0] node29467;
	wire [16-1:0] node29469;
	wire [16-1:0] node29470;
	wire [16-1:0] node29475;
	wire [16-1:0] node29476;
	wire [16-1:0] node29477;
	wire [16-1:0] node29478;
	wire [16-1:0] node29479;
	wire [16-1:0] node29480;
	wire [16-1:0] node29483;
	wire [16-1:0] node29486;
	wire [16-1:0] node29488;
	wire [16-1:0] node29489;
	wire [16-1:0] node29490;
	wire [16-1:0] node29495;
	wire [16-1:0] node29497;
	wire [16-1:0] node29498;
	wire [16-1:0] node29499;
	wire [16-1:0] node29500;
	wire [16-1:0] node29504;
	wire [16-1:0] node29507;
	wire [16-1:0] node29508;
	wire [16-1:0] node29512;
	wire [16-1:0] node29513;
	wire [16-1:0] node29514;
	wire [16-1:0] node29515;
	wire [16-1:0] node29518;
	wire [16-1:0] node29521;
	wire [16-1:0] node29522;
	wire [16-1:0] node29525;
	wire [16-1:0] node29528;
	wire [16-1:0] node29529;
	wire [16-1:0] node29530;
	wire [16-1:0] node29531;
	wire [16-1:0] node29535;
	wire [16-1:0] node29538;
	wire [16-1:0] node29539;
	wire [16-1:0] node29542;
	wire [16-1:0] node29545;
	wire [16-1:0] node29546;
	wire [16-1:0] node29547;
	wire [16-1:0] node29548;
	wire [16-1:0] node29551;
	wire [16-1:0] node29552;
	wire [16-1:0] node29553;
	wire [16-1:0] node29558;
	wire [16-1:0] node29559;
	wire [16-1:0] node29560;
	wire [16-1:0] node29563;
	wire [16-1:0] node29566;
	wire [16-1:0] node29567;
	wire [16-1:0] node29569;
	wire [16-1:0] node29570;
	wire [16-1:0] node29574;
	wire [16-1:0] node29577;
	wire [16-1:0] node29578;
	wire [16-1:0] node29579;
	wire [16-1:0] node29580;
	wire [16-1:0] node29583;
	wire [16-1:0] node29585;
	wire [16-1:0] node29586;
	wire [16-1:0] node29590;
	wire [16-1:0] node29591;
	wire [16-1:0] node29594;
	wire [16-1:0] node29595;
	wire [16-1:0] node29599;
	wire [16-1:0] node29600;
	wire [16-1:0] node29602;
	wire [16-1:0] node29604;
	wire [16-1:0] node29605;
	wire [16-1:0] node29609;
	wire [16-1:0] node29610;
	wire [16-1:0] node29611;
	wire [16-1:0] node29615;
	wire [16-1:0] node29618;
	wire [16-1:0] node29619;
	wire [16-1:0] node29620;
	wire [16-1:0] node29621;
	wire [16-1:0] node29622;
	wire [16-1:0] node29623;
	wire [16-1:0] node29624;
	wire [16-1:0] node29625;
	wire [16-1:0] node29628;
	wire [16-1:0] node29630;
	wire [16-1:0] node29631;
	wire [16-1:0] node29635;
	wire [16-1:0] node29636;
	wire [16-1:0] node29639;
	wire [16-1:0] node29641;
	wire [16-1:0] node29642;
	wire [16-1:0] node29646;
	wire [16-1:0] node29647;
	wire [16-1:0] node29648;
	wire [16-1:0] node29649;
	wire [16-1:0] node29654;
	wire [16-1:0] node29655;
	wire [16-1:0] node29658;
	wire [16-1:0] node29661;
	wire [16-1:0] node29662;
	wire [16-1:0] node29663;
	wire [16-1:0] node29664;
	wire [16-1:0] node29666;
	wire [16-1:0] node29667;
	wire [16-1:0] node29671;
	wire [16-1:0] node29673;
	wire [16-1:0] node29676;
	wire [16-1:0] node29677;
	wire [16-1:0] node29680;
	wire [16-1:0] node29682;
	wire [16-1:0] node29685;
	wire [16-1:0] node29686;
	wire [16-1:0] node29689;
	wire [16-1:0] node29690;
	wire [16-1:0] node29691;
	wire [16-1:0] node29693;
	wire [16-1:0] node29696;
	wire [16-1:0] node29699;
	wire [16-1:0] node29702;
	wire [16-1:0] node29703;
	wire [16-1:0] node29704;
	wire [16-1:0] node29705;
	wire [16-1:0] node29706;
	wire [16-1:0] node29710;
	wire [16-1:0] node29712;
	wire [16-1:0] node29713;
	wire [16-1:0] node29717;
	wire [16-1:0] node29718;
	wire [16-1:0] node29719;
	wire [16-1:0] node29722;
	wire [16-1:0] node29724;
	wire [16-1:0] node29727;
	wire [16-1:0] node29728;
	wire [16-1:0] node29732;
	wire [16-1:0] node29733;
	wire [16-1:0] node29734;
	wire [16-1:0] node29736;
	wire [16-1:0] node29739;
	wire [16-1:0] node29740;
	wire [16-1:0] node29741;
	wire [16-1:0] node29746;
	wire [16-1:0] node29747;
	wire [16-1:0] node29748;
	wire [16-1:0] node29751;
	wire [16-1:0] node29754;
	wire [16-1:0] node29755;
	wire [16-1:0] node29758;
	wire [16-1:0] node29761;
	wire [16-1:0] node29762;
	wire [16-1:0] node29763;
	wire [16-1:0] node29764;
	wire [16-1:0] node29765;
	wire [16-1:0] node29767;
	wire [16-1:0] node29768;
	wire [16-1:0] node29773;
	wire [16-1:0] node29774;
	wire [16-1:0] node29775;
	wire [16-1:0] node29776;
	wire [16-1:0] node29778;
	wire [16-1:0] node29781;
	wire [16-1:0] node29782;
	wire [16-1:0] node29786;
	wire [16-1:0] node29789;
	wire [16-1:0] node29790;
	wire [16-1:0] node29792;
	wire [16-1:0] node29795;
	wire [16-1:0] node29796;
	wire [16-1:0] node29800;
	wire [16-1:0] node29801;
	wire [16-1:0] node29802;
	wire [16-1:0] node29803;
	wire [16-1:0] node29806;
	wire [16-1:0] node29807;
	wire [16-1:0] node29809;
	wire [16-1:0] node29813;
	wire [16-1:0] node29814;
	wire [16-1:0] node29816;
	wire [16-1:0] node29820;
	wire [16-1:0] node29821;
	wire [16-1:0] node29822;
	wire [16-1:0] node29823;
	wire [16-1:0] node29828;
	wire [16-1:0] node29831;
	wire [16-1:0] node29832;
	wire [16-1:0] node29833;
	wire [16-1:0] node29834;
	wire [16-1:0] node29835;
	wire [16-1:0] node29838;
	wire [16-1:0] node29839;
	wire [16-1:0] node29841;
	wire [16-1:0] node29845;
	wire [16-1:0] node29846;
	wire [16-1:0] node29847;
	wire [16-1:0] node29849;
	wire [16-1:0] node29852;
	wire [16-1:0] node29855;
	wire [16-1:0] node29857;
	wire [16-1:0] node29860;
	wire [16-1:0] node29861;
	wire [16-1:0] node29862;
	wire [16-1:0] node29865;
	wire [16-1:0] node29866;
	wire [16-1:0] node29870;
	wire [16-1:0] node29872;
	wire [16-1:0] node29875;
	wire [16-1:0] node29876;
	wire [16-1:0] node29877;
	wire [16-1:0] node29880;
	wire [16-1:0] node29882;
	wire [16-1:0] node29884;
	wire [16-1:0] node29887;
	wire [16-1:0] node29888;
	wire [16-1:0] node29890;
	wire [16-1:0] node29893;
	wire [16-1:0] node29894;
	wire [16-1:0] node29897;
	wire [16-1:0] node29898;
	wire [16-1:0] node29900;
	wire [16-1:0] node29903;
	wire [16-1:0] node29905;
	wire [16-1:0] node29908;
	wire [16-1:0] node29909;
	wire [16-1:0] node29910;
	wire [16-1:0] node29911;
	wire [16-1:0] node29912;
	wire [16-1:0] node29913;
	wire [16-1:0] node29914;
	wire [16-1:0] node29916;
	wire [16-1:0] node29920;
	wire [16-1:0] node29922;
	wire [16-1:0] node29925;
	wire [16-1:0] node29926;
	wire [16-1:0] node29927;
	wire [16-1:0] node29930;
	wire [16-1:0] node29932;
	wire [16-1:0] node29933;
	wire [16-1:0] node29937;
	wire [16-1:0] node29939;
	wire [16-1:0] node29942;
	wire [16-1:0] node29943;
	wire [16-1:0] node29944;
	wire [16-1:0] node29946;
	wire [16-1:0] node29948;
	wire [16-1:0] node29952;
	wire [16-1:0] node29953;
	wire [16-1:0] node29955;
	wire [16-1:0] node29958;
	wire [16-1:0] node29960;
	wire [16-1:0] node29963;
	wire [16-1:0] node29964;
	wire [16-1:0] node29965;
	wire [16-1:0] node29966;
	wire [16-1:0] node29967;
	wire [16-1:0] node29971;
	wire [16-1:0] node29972;
	wire [16-1:0] node29973;
	wire [16-1:0] node29975;
	wire [16-1:0] node29979;
	wire [16-1:0] node29981;
	wire [16-1:0] node29984;
	wire [16-1:0] node29985;
	wire [16-1:0] node29986;
	wire [16-1:0] node29988;
	wire [16-1:0] node29991;
	wire [16-1:0] node29992;
	wire [16-1:0] node29994;
	wire [16-1:0] node29997;
	wire [16-1:0] node29998;
	wire [16-1:0] node30002;
	wire [16-1:0] node30003;
	wire [16-1:0] node30007;
	wire [16-1:0] node30008;
	wire [16-1:0] node30009;
	wire [16-1:0] node30012;
	wire [16-1:0] node30013;
	wire [16-1:0] node30016;
	wire [16-1:0] node30019;
	wire [16-1:0] node30020;
	wire [16-1:0] node30021;
	wire [16-1:0] node30022;
	wire [16-1:0] node30026;
	wire [16-1:0] node30029;
	wire [16-1:0] node30030;
	wire [16-1:0] node30034;
	wire [16-1:0] node30035;
	wire [16-1:0] node30036;
	wire [16-1:0] node30037;
	wire [16-1:0] node30038;
	wire [16-1:0] node30041;
	wire [16-1:0] node30043;
	wire [16-1:0] node30046;
	wire [16-1:0] node30047;
	wire [16-1:0] node30050;
	wire [16-1:0] node30051;
	wire [16-1:0] node30053;
	wire [16-1:0] node30054;
	wire [16-1:0] node30059;
	wire [16-1:0] node30060;
	wire [16-1:0] node30061;
	wire [16-1:0] node30062;
	wire [16-1:0] node30063;
	wire [16-1:0] node30067;
	wire [16-1:0] node30069;
	wire [16-1:0] node30072;
	wire [16-1:0] node30073;
	wire [16-1:0] node30077;
	wire [16-1:0] node30078;
	wire [16-1:0] node30081;
	wire [16-1:0] node30083;
	wire [16-1:0] node30086;
	wire [16-1:0] node30087;
	wire [16-1:0] node30088;
	wire [16-1:0] node30089;
	wire [16-1:0] node30090;
	wire [16-1:0] node30093;
	wire [16-1:0] node30095;
	wire [16-1:0] node30097;
	wire [16-1:0] node30100;
	wire [16-1:0] node30101;
	wire [16-1:0] node30104;
	wire [16-1:0] node30107;
	wire [16-1:0] node30108;
	wire [16-1:0] node30109;
	wire [16-1:0] node30111;
	wire [16-1:0] node30114;
	wire [16-1:0] node30117;
	wire [16-1:0] node30118;
	wire [16-1:0] node30119;
	wire [16-1:0] node30124;
	wire [16-1:0] node30125;
	wire [16-1:0] node30126;
	wire [16-1:0] node30128;
	wire [16-1:0] node30130;
	wire [16-1:0] node30131;
	wire [16-1:0] node30135;
	wire [16-1:0] node30136;
	wire [16-1:0] node30140;
	wire [16-1:0] node30141;
	wire [16-1:0] node30142;
	wire [16-1:0] node30144;
	wire [16-1:0] node30145;
	wire [16-1:0] node30149;
	wire [16-1:0] node30151;
	wire [16-1:0] node30154;
	wire [16-1:0] node30155;
	wire [16-1:0] node30158;
	wire [16-1:0] node30159;
	wire [16-1:0] node30161;
	wire [16-1:0] node30165;
	wire [16-1:0] node30166;
	wire [16-1:0] node30167;
	wire [16-1:0] node30168;
	wire [16-1:0] node30169;
	wire [16-1:0] node30170;
	wire [16-1:0] node30171;
	wire [16-1:0] node30172;
	wire [16-1:0] node30173;
	wire [16-1:0] node30175;
	wire [16-1:0] node30176;
	wire [16-1:0] node30180;
	wire [16-1:0] node30184;
	wire [16-1:0] node30186;
	wire [16-1:0] node30187;
	wire [16-1:0] node30188;
	wire [16-1:0] node30193;
	wire [16-1:0] node30194;
	wire [16-1:0] node30195;
	wire [16-1:0] node30196;
	wire [16-1:0] node30199;
	wire [16-1:0] node30201;
	wire [16-1:0] node30204;
	wire [16-1:0] node30205;
	wire [16-1:0] node30206;
	wire [16-1:0] node30208;
	wire [16-1:0] node30211;
	wire [16-1:0] node30215;
	wire [16-1:0] node30216;
	wire [16-1:0] node30217;
	wire [16-1:0] node30220;
	wire [16-1:0] node30222;
	wire [16-1:0] node30223;
	wire [16-1:0] node30227;
	wire [16-1:0] node30228;
	wire [16-1:0] node30231;
	wire [16-1:0] node30233;
	wire [16-1:0] node30234;
	wire [16-1:0] node30238;
	wire [16-1:0] node30239;
	wire [16-1:0] node30240;
	wire [16-1:0] node30241;
	wire [16-1:0] node30242;
	wire [16-1:0] node30247;
	wire [16-1:0] node30248;
	wire [16-1:0] node30249;
	wire [16-1:0] node30250;
	wire [16-1:0] node30254;
	wire [16-1:0] node30255;
	wire [16-1:0] node30257;
	wire [16-1:0] node30261;
	wire [16-1:0] node30262;
	wire [16-1:0] node30263;
	wire [16-1:0] node30268;
	wire [16-1:0] node30269;
	wire [16-1:0] node30270;
	wire [16-1:0] node30271;
	wire [16-1:0] node30273;
	wire [16-1:0] node30276;
	wire [16-1:0] node30279;
	wire [16-1:0] node30281;
	wire [16-1:0] node30284;
	wire [16-1:0] node30285;
	wire [16-1:0] node30286;
	wire [16-1:0] node30290;
	wire [16-1:0] node30291;
	wire [16-1:0] node30294;
	wire [16-1:0] node30296;
	wire [16-1:0] node30297;
	wire [16-1:0] node30301;
	wire [16-1:0] node30302;
	wire [16-1:0] node30303;
	wire [16-1:0] node30304;
	wire [16-1:0] node30305;
	wire [16-1:0] node30306;
	wire [16-1:0] node30308;
	wire [16-1:0] node30311;
	wire [16-1:0] node30314;
	wire [16-1:0] node30315;
	wire [16-1:0] node30317;
	wire [16-1:0] node30321;
	wire [16-1:0] node30322;
	wire [16-1:0] node30323;
	wire [16-1:0] node30327;
	wire [16-1:0] node30328;
	wire [16-1:0] node30331;
	wire [16-1:0] node30334;
	wire [16-1:0] node30335;
	wire [16-1:0] node30336;
	wire [16-1:0] node30338;
	wire [16-1:0] node30341;
	wire [16-1:0] node30342;
	wire [16-1:0] node30343;
	wire [16-1:0] node30348;
	wire [16-1:0] node30349;
	wire [16-1:0] node30350;
	wire [16-1:0] node30354;
	wire [16-1:0] node30356;
	wire [16-1:0] node30359;
	wire [16-1:0] node30360;
	wire [16-1:0] node30361;
	wire [16-1:0] node30362;
	wire [16-1:0] node30363;
	wire [16-1:0] node30367;
	wire [16-1:0] node30368;
	wire [16-1:0] node30371;
	wire [16-1:0] node30372;
	wire [16-1:0] node30374;
	wire [16-1:0] node30378;
	wire [16-1:0] node30379;
	wire [16-1:0] node30381;
	wire [16-1:0] node30385;
	wire [16-1:0] node30386;
	wire [16-1:0] node30388;
	wire [16-1:0] node30389;
	wire [16-1:0] node30392;
	wire [16-1:0] node30395;
	wire [16-1:0] node30396;
	wire [16-1:0] node30397;
	wire [16-1:0] node30400;
	wire [16-1:0] node30402;
	wire [16-1:0] node30404;
	wire [16-1:0] node30407;
	wire [16-1:0] node30409;
	wire [16-1:0] node30412;
	wire [16-1:0] node30413;
	wire [16-1:0] node30414;
	wire [16-1:0] node30415;
	wire [16-1:0] node30416;
	wire [16-1:0] node30417;
	wire [16-1:0] node30418;
	wire [16-1:0] node30419;
	wire [16-1:0] node30423;
	wire [16-1:0] node30426;
	wire [16-1:0] node30427;
	wire [16-1:0] node30429;
	wire [16-1:0] node30432;
	wire [16-1:0] node30433;
	wire [16-1:0] node30434;
	wire [16-1:0] node30438;
	wire [16-1:0] node30439;
	wire [16-1:0] node30443;
	wire [16-1:0] node30445;
	wire [16-1:0] node30446;
	wire [16-1:0] node30449;
	wire [16-1:0] node30452;
	wire [16-1:0] node30453;
	wire [16-1:0] node30454;
	wire [16-1:0] node30456;
	wire [16-1:0] node30458;
	wire [16-1:0] node30459;
	wire [16-1:0] node30463;
	wire [16-1:0] node30464;
	wire [16-1:0] node30467;
	wire [16-1:0] node30470;
	wire [16-1:0] node30471;
	wire [16-1:0] node30473;
	wire [16-1:0] node30476;
	wire [16-1:0] node30477;
	wire [16-1:0] node30478;
	wire [16-1:0] node30482;
	wire [16-1:0] node30485;
	wire [16-1:0] node30486;
	wire [16-1:0] node30487;
	wire [16-1:0] node30488;
	wire [16-1:0] node30489;
	wire [16-1:0] node30492;
	wire [16-1:0] node30494;
	wire [16-1:0] node30495;
	wire [16-1:0] node30499;
	wire [16-1:0] node30501;
	wire [16-1:0] node30504;
	wire [16-1:0] node30505;
	wire [16-1:0] node30506;
	wire [16-1:0] node30507;
	wire [16-1:0] node30509;
	wire [16-1:0] node30514;
	wire [16-1:0] node30515;
	wire [16-1:0] node30518;
	wire [16-1:0] node30521;
	wire [16-1:0] node30522;
	wire [16-1:0] node30523;
	wire [16-1:0] node30525;
	wire [16-1:0] node30526;
	wire [16-1:0] node30527;
	wire [16-1:0] node30530;
	wire [16-1:0] node30534;
	wire [16-1:0] node30535;
	wire [16-1:0] node30537;
	wire [16-1:0] node30538;
	wire [16-1:0] node30542;
	wire [16-1:0] node30544;
	wire [16-1:0] node30547;
	wire [16-1:0] node30548;
	wire [16-1:0] node30549;
	wire [16-1:0] node30551;
	wire [16-1:0] node30554;
	wire [16-1:0] node30556;
	wire [16-1:0] node30558;
	wire [16-1:0] node30561;
	wire [16-1:0] node30562;
	wire [16-1:0] node30563;
	wire [16-1:0] node30565;
	wire [16-1:0] node30568;
	wire [16-1:0] node30569;
	wire [16-1:0] node30574;
	wire [16-1:0] node30575;
	wire [16-1:0] node30576;
	wire [16-1:0] node30577;
	wire [16-1:0] node30578;
	wire [16-1:0] node30579;
	wire [16-1:0] node30582;
	wire [16-1:0] node30585;
	wire [16-1:0] node30587;
	wire [16-1:0] node30590;
	wire [16-1:0] node30591;
	wire [16-1:0] node30592;
	wire [16-1:0] node30595;
	wire [16-1:0] node30598;
	wire [16-1:0] node30600;
	wire [16-1:0] node30603;
	wire [16-1:0] node30604;
	wire [16-1:0] node30605;
	wire [16-1:0] node30606;
	wire [16-1:0] node30609;
	wire [16-1:0] node30612;
	wire [16-1:0] node30613;
	wire [16-1:0] node30616;
	wire [16-1:0] node30617;
	wire [16-1:0] node30621;
	wire [16-1:0] node30622;
	wire [16-1:0] node30625;
	wire [16-1:0] node30627;
	wire [16-1:0] node30630;
	wire [16-1:0] node30631;
	wire [16-1:0] node30632;
	wire [16-1:0] node30633;
	wire [16-1:0] node30634;
	wire [16-1:0] node30639;
	wire [16-1:0] node30640;
	wire [16-1:0] node30642;
	wire [16-1:0] node30645;
	wire [16-1:0] node30646;
	wire [16-1:0] node30650;
	wire [16-1:0] node30651;
	wire [16-1:0] node30652;
	wire [16-1:0] node30653;
	wire [16-1:0] node30656;
	wire [16-1:0] node30659;
	wire [16-1:0] node30660;
	wire [16-1:0] node30663;
	wire [16-1:0] node30666;
	wire [16-1:0] node30667;
	wire [16-1:0] node30669;
	wire [16-1:0] node30673;
	wire [16-1:0] node30674;
	wire [16-1:0] node30675;
	wire [16-1:0] node30676;
	wire [16-1:0] node30677;
	wire [16-1:0] node30678;
	wire [16-1:0] node30679;
	wire [16-1:0] node30682;
	wire [16-1:0] node30683;
	wire [16-1:0] node30685;
	wire [16-1:0] node30689;
	wire [16-1:0] node30690;
	wire [16-1:0] node30693;
	wire [16-1:0] node30694;
	wire [16-1:0] node30696;
	wire [16-1:0] node30700;
	wire [16-1:0] node30701;
	wire [16-1:0] node30702;
	wire [16-1:0] node30703;
	wire [16-1:0] node30706;
	wire [16-1:0] node30709;
	wire [16-1:0] node30710;
	wire [16-1:0] node30714;
	wire [16-1:0] node30715;
	wire [16-1:0] node30717;
	wire [16-1:0] node30719;
	wire [16-1:0] node30722;
	wire [16-1:0] node30723;
	wire [16-1:0] node30727;
	wire [16-1:0] node30728;
	wire [16-1:0] node30729;
	wire [16-1:0] node30730;
	wire [16-1:0] node30731;
	wire [16-1:0] node30734;
	wire [16-1:0] node30736;
	wire [16-1:0] node30739;
	wire [16-1:0] node30740;
	wire [16-1:0] node30742;
	wire [16-1:0] node30743;
	wire [16-1:0] node30747;
	wire [16-1:0] node30750;
	wire [16-1:0] node30751;
	wire [16-1:0] node30752;
	wire [16-1:0] node30755;
	wire [16-1:0] node30758;
	wire [16-1:0] node30759;
	wire [16-1:0] node30762;
	wire [16-1:0] node30765;
	wire [16-1:0] node30766;
	wire [16-1:0] node30767;
	wire [16-1:0] node30769;
	wire [16-1:0] node30770;
	wire [16-1:0] node30772;
	wire [16-1:0] node30776;
	wire [16-1:0] node30777;
	wire [16-1:0] node30778;
	wire [16-1:0] node30782;
	wire [16-1:0] node30784;
	wire [16-1:0] node30787;
	wire [16-1:0] node30788;
	wire [16-1:0] node30790;
	wire [16-1:0] node30793;
	wire [16-1:0] node30794;
	wire [16-1:0] node30797;
	wire [16-1:0] node30800;
	wire [16-1:0] node30801;
	wire [16-1:0] node30802;
	wire [16-1:0] node30803;
	wire [16-1:0] node30804;
	wire [16-1:0] node30805;
	wire [16-1:0] node30808;
	wire [16-1:0] node30809;
	wire [16-1:0] node30813;
	wire [16-1:0] node30814;
	wire [16-1:0] node30817;
	wire [16-1:0] node30819;
	wire [16-1:0] node30820;
	wire [16-1:0] node30824;
	wire [16-1:0] node30825;
	wire [16-1:0] node30826;
	wire [16-1:0] node30829;
	wire [16-1:0] node30832;
	wire [16-1:0] node30833;
	wire [16-1:0] node30836;
	wire [16-1:0] node30839;
	wire [16-1:0] node30840;
	wire [16-1:0] node30841;
	wire [16-1:0] node30842;
	wire [16-1:0] node30845;
	wire [16-1:0] node30847;
	wire [16-1:0] node30850;
	wire [16-1:0] node30851;
	wire [16-1:0] node30853;
	wire [16-1:0] node30854;
	wire [16-1:0] node30858;
	wire [16-1:0] node30861;
	wire [16-1:0] node30862;
	wire [16-1:0] node30864;
	wire [16-1:0] node30867;
	wire [16-1:0] node30868;
	wire [16-1:0] node30871;
	wire [16-1:0] node30872;
	wire [16-1:0] node30876;
	wire [16-1:0] node30877;
	wire [16-1:0] node30878;
	wire [16-1:0] node30879;
	wire [16-1:0] node30880;
	wire [16-1:0] node30884;
	wire [16-1:0] node30885;
	wire [16-1:0] node30889;
	wire [16-1:0] node30890;
	wire [16-1:0] node30893;
	wire [16-1:0] node30894;
	wire [16-1:0] node30897;
	wire [16-1:0] node30899;
	wire [16-1:0] node30902;
	wire [16-1:0] node30903;
	wire [16-1:0] node30904;
	wire [16-1:0] node30906;
	wire [16-1:0] node30909;
	wire [16-1:0] node30910;
	wire [16-1:0] node30911;
	wire [16-1:0] node30913;
	wire [16-1:0] node30916;
	wire [16-1:0] node30918;
	wire [16-1:0] node30921;
	wire [16-1:0] node30924;
	wire [16-1:0] node30926;
	wire [16-1:0] node30927;
	wire [16-1:0] node30930;
	wire [16-1:0] node30933;
	wire [16-1:0] node30934;
	wire [16-1:0] node30935;
	wire [16-1:0] node30936;
	wire [16-1:0] node30937;
	wire [16-1:0] node30938;
	wire [16-1:0] node30939;
	wire [16-1:0] node30941;
	wire [16-1:0] node30944;
	wire [16-1:0] node30947;
	wire [16-1:0] node30948;
	wire [16-1:0] node30952;
	wire [16-1:0] node30953;
	wire [16-1:0] node30954;
	wire [16-1:0] node30958;
	wire [16-1:0] node30959;
	wire [16-1:0] node30962;
	wire [16-1:0] node30963;
	wire [16-1:0] node30965;
	wire [16-1:0] node30969;
	wire [16-1:0] node30970;
	wire [16-1:0] node30971;
	wire [16-1:0] node30972;
	wire [16-1:0] node30973;
	wire [16-1:0] node30977;
	wire [16-1:0] node30980;
	wire [16-1:0] node30981;
	wire [16-1:0] node30983;
	wire [16-1:0] node30986;
	wire [16-1:0] node30987;
	wire [16-1:0] node30988;
	wire [16-1:0] node30993;
	wire [16-1:0] node30994;
	wire [16-1:0] node30995;
	wire [16-1:0] node30999;
	wire [16-1:0] node31000;
	wire [16-1:0] node31002;
	wire [16-1:0] node31005;
	wire [16-1:0] node31006;
	wire [16-1:0] node31010;
	wire [16-1:0] node31011;
	wire [16-1:0] node31012;
	wire [16-1:0] node31013;
	wire [16-1:0] node31014;
	wire [16-1:0] node31017;
	wire [16-1:0] node31019;
	wire [16-1:0] node31020;
	wire [16-1:0] node31025;
	wire [16-1:0] node31026;
	wire [16-1:0] node31027;
	wire [16-1:0] node31030;
	wire [16-1:0] node31033;
	wire [16-1:0] node31034;
	wire [16-1:0] node31037;
	wire [16-1:0] node31038;
	wire [16-1:0] node31040;
	wire [16-1:0] node31043;
	wire [16-1:0] node31046;
	wire [16-1:0] node31047;
	wire [16-1:0] node31048;
	wire [16-1:0] node31050;
	wire [16-1:0] node31053;
	wire [16-1:0] node31055;
	wire [16-1:0] node31058;
	wire [16-1:0] node31059;
	wire [16-1:0] node31062;
	wire [16-1:0] node31063;
	wire [16-1:0] node31064;
	wire [16-1:0] node31067;
	wire [16-1:0] node31069;
	wire [16-1:0] node31072;
	wire [16-1:0] node31073;
	wire [16-1:0] node31075;
	wire [16-1:0] node31078;
	wire [16-1:0] node31081;
	wire [16-1:0] node31082;
	wire [16-1:0] node31083;
	wire [16-1:0] node31084;
	wire [16-1:0] node31085;
	wire [16-1:0] node31086;
	wire [16-1:0] node31087;
	wire [16-1:0] node31091;
	wire [16-1:0] node31092;
	wire [16-1:0] node31094;
	wire [16-1:0] node31098;
	wire [16-1:0] node31101;
	wire [16-1:0] node31102;
	wire [16-1:0] node31103;
	wire [16-1:0] node31106;
	wire [16-1:0] node31109;
	wire [16-1:0] node31111;
	wire [16-1:0] node31114;
	wire [16-1:0] node31115;
	wire [16-1:0] node31116;
	wire [16-1:0] node31117;
	wire [16-1:0] node31120;
	wire [16-1:0] node31123;
	wire [16-1:0] node31125;
	wire [16-1:0] node31128;
	wire [16-1:0] node31129;
	wire [16-1:0] node31131;
	wire [16-1:0] node31132;
	wire [16-1:0] node31135;
	wire [16-1:0] node31137;
	wire [16-1:0] node31140;
	wire [16-1:0] node31142;
	wire [16-1:0] node31145;
	wire [16-1:0] node31146;
	wire [16-1:0] node31147;
	wire [16-1:0] node31148;
	wire [16-1:0] node31152;
	wire [16-1:0] node31153;
	wire [16-1:0] node31154;
	wire [16-1:0] node31155;
	wire [16-1:0] node31159;
	wire [16-1:0] node31161;
	wire [16-1:0] node31163;
	wire [16-1:0] node31166;
	wire [16-1:0] node31167;
	wire [16-1:0] node31169;
	wire [16-1:0] node31173;
	wire [16-1:0] node31174;
	wire [16-1:0] node31175;
	wire [16-1:0] node31177;
	wire [16-1:0] node31178;
	wire [16-1:0] node31182;
	wire [16-1:0] node31183;
	wire [16-1:0] node31185;
	wire [16-1:0] node31187;
	wire [16-1:0] node31190;
	wire [16-1:0] node31191;
	wire [16-1:0] node31195;
	wire [16-1:0] node31196;
	wire [16-1:0] node31197;
	wire [16-1:0] node31201;
	wire [16-1:0] node31202;
	wire [16-1:0] node31203;
	wire [16-1:0] node31206;
	wire [16-1:0] node31208;
	wire [16-1:0] node31211;
	wire [16-1:0] node31213;
	wire [16-1:0] node31215;
	wire [16-1:0] node31218;
	wire [16-1:0] node31219;
	wire [16-1:0] node31220;
	wire [16-1:0] node31221;
	wire [16-1:0] node31222;
	wire [16-1:0] node31223;
	wire [16-1:0] node31224;
	wire [16-1:0] node31225;
	wire [16-1:0] node31226;
	wire [16-1:0] node31227;
	wire [16-1:0] node31228;
	wire [16-1:0] node31231;
	wire [16-1:0] node31235;
	wire [16-1:0] node31236;
	wire [16-1:0] node31237;
	wire [16-1:0] node31240;
	wire [16-1:0] node31243;
	wire [16-1:0] node31246;
	wire [16-1:0] node31247;
	wire [16-1:0] node31248;
	wire [16-1:0] node31249;
	wire [16-1:0] node31253;
	wire [16-1:0] node31256;
	wire [16-1:0] node31258;
	wire [16-1:0] node31259;
	wire [16-1:0] node31263;
	wire [16-1:0] node31264;
	wire [16-1:0] node31265;
	wire [16-1:0] node31267;
	wire [16-1:0] node31268;
	wire [16-1:0] node31271;
	wire [16-1:0] node31272;
	wire [16-1:0] node31277;
	wire [16-1:0] node31278;
	wire [16-1:0] node31279;
	wire [16-1:0] node31281;
	wire [16-1:0] node31284;
	wire [16-1:0] node31286;
	wire [16-1:0] node31289;
	wire [16-1:0] node31291;
	wire [16-1:0] node31294;
	wire [16-1:0] node31295;
	wire [16-1:0] node31296;
	wire [16-1:0] node31297;
	wire [16-1:0] node31298;
	wire [16-1:0] node31300;
	wire [16-1:0] node31301;
	wire [16-1:0] node31305;
	wire [16-1:0] node31306;
	wire [16-1:0] node31310;
	wire [16-1:0] node31312;
	wire [16-1:0] node31313;
	wire [16-1:0] node31317;
	wire [16-1:0] node31318;
	wire [16-1:0] node31319;
	wire [16-1:0] node31322;
	wire [16-1:0] node31326;
	wire [16-1:0] node31327;
	wire [16-1:0] node31328;
	wire [16-1:0] node31331;
	wire [16-1:0] node31333;
	wire [16-1:0] node31335;
	wire [16-1:0] node31338;
	wire [16-1:0] node31339;
	wire [16-1:0] node31340;
	wire [16-1:0] node31343;
	wire [16-1:0] node31344;
	wire [16-1:0] node31346;
	wire [16-1:0] node31350;
	wire [16-1:0] node31351;
	wire [16-1:0] node31354;
	wire [16-1:0] node31356;
	wire [16-1:0] node31359;
	wire [16-1:0] node31360;
	wire [16-1:0] node31361;
	wire [16-1:0] node31362;
	wire [16-1:0] node31363;
	wire [16-1:0] node31364;
	wire [16-1:0] node31366;
	wire [16-1:0] node31367;
	wire [16-1:0] node31370;
	wire [16-1:0] node31373;
	wire [16-1:0] node31376;
	wire [16-1:0] node31377;
	wire [16-1:0] node31381;
	wire [16-1:0] node31382;
	wire [16-1:0] node31383;
	wire [16-1:0] node31384;
	wire [16-1:0] node31388;
	wire [16-1:0] node31390;
	wire [16-1:0] node31391;
	wire [16-1:0] node31395;
	wire [16-1:0] node31397;
	wire [16-1:0] node31400;
	wire [16-1:0] node31401;
	wire [16-1:0] node31402;
	wire [16-1:0] node31403;
	wire [16-1:0] node31404;
	wire [16-1:0] node31406;
	wire [16-1:0] node31409;
	wire [16-1:0] node31412;
	wire [16-1:0] node31414;
	wire [16-1:0] node31417;
	wire [16-1:0] node31419;
	wire [16-1:0] node31422;
	wire [16-1:0] node31424;
	wire [16-1:0] node31425;
	wire [16-1:0] node31428;
	wire [16-1:0] node31429;
	wire [16-1:0] node31430;
	wire [16-1:0] node31435;
	wire [16-1:0] node31436;
	wire [16-1:0] node31437;
	wire [16-1:0] node31438;
	wire [16-1:0] node31439;
	wire [16-1:0] node31443;
	wire [16-1:0] node31444;
	wire [16-1:0] node31447;
	wire [16-1:0] node31449;
	wire [16-1:0] node31452;
	wire [16-1:0] node31453;
	wire [16-1:0] node31454;
	wire [16-1:0] node31457;
	wire [16-1:0] node31459;
	wire [16-1:0] node31460;
	wire [16-1:0] node31464;
	wire [16-1:0] node31465;
	wire [16-1:0] node31467;
	wire [16-1:0] node31468;
	wire [16-1:0] node31473;
	wire [16-1:0] node31474;
	wire [16-1:0] node31475;
	wire [16-1:0] node31476;
	wire [16-1:0] node31478;
	wire [16-1:0] node31479;
	wire [16-1:0] node31484;
	wire [16-1:0] node31485;
	wire [16-1:0] node31486;
	wire [16-1:0] node31491;
	wire [16-1:0] node31492;
	wire [16-1:0] node31493;
	wire [16-1:0] node31495;
	wire [16-1:0] node31496;
	wire [16-1:0] node31501;
	wire [16-1:0] node31503;
	wire [16-1:0] node31505;
	wire [16-1:0] node31508;
	wire [16-1:0] node31509;
	wire [16-1:0] node31510;
	wire [16-1:0] node31511;
	wire [16-1:0] node31512;
	wire [16-1:0] node31513;
	wire [16-1:0] node31514;
	wire [16-1:0] node31517;
	wire [16-1:0] node31520;
	wire [16-1:0] node31522;
	wire [16-1:0] node31525;
	wire [16-1:0] node31526;
	wire [16-1:0] node31527;
	wire [16-1:0] node31530;
	wire [16-1:0] node31533;
	wire [16-1:0] node31534;
	wire [16-1:0] node31537;
	wire [16-1:0] node31540;
	wire [16-1:0] node31541;
	wire [16-1:0] node31542;
	wire [16-1:0] node31543;
	wire [16-1:0] node31546;
	wire [16-1:0] node31549;
	wire [16-1:0] node31550;
	wire [16-1:0] node31553;
	wire [16-1:0] node31556;
	wire [16-1:0] node31557;
	wire [16-1:0] node31558;
	wire [16-1:0] node31561;
	wire [16-1:0] node31564;
	wire [16-1:0] node31565;
	wire [16-1:0] node31568;
	wire [16-1:0] node31571;
	wire [16-1:0] node31572;
	wire [16-1:0] node31573;
	wire [16-1:0] node31574;
	wire [16-1:0] node31575;
	wire [16-1:0] node31579;
	wire [16-1:0] node31581;
	wire [16-1:0] node31584;
	wire [16-1:0] node31585;
	wire [16-1:0] node31586;
	wire [16-1:0] node31589;
	wire [16-1:0] node31592;
	wire [16-1:0] node31593;
	wire [16-1:0] node31596;
	wire [16-1:0] node31599;
	wire [16-1:0] node31600;
	wire [16-1:0] node31601;
	wire [16-1:0] node31603;
	wire [16-1:0] node31606;
	wire [16-1:0] node31607;
	wire [16-1:0] node31608;
	wire [16-1:0] node31612;
	wire [16-1:0] node31615;
	wire [16-1:0] node31616;
	wire [16-1:0] node31617;
	wire [16-1:0] node31620;
	wire [16-1:0] node31621;
	wire [16-1:0] node31623;
	wire [16-1:0] node31627;
	wire [16-1:0] node31628;
	wire [16-1:0] node31630;
	wire [16-1:0] node31632;
	wire [16-1:0] node31635;
	wire [16-1:0] node31637;
	wire [16-1:0] node31640;
	wire [16-1:0] node31641;
	wire [16-1:0] node31642;
	wire [16-1:0] node31643;
	wire [16-1:0] node31644;
	wire [16-1:0] node31647;
	wire [16-1:0] node31648;
	wire [16-1:0] node31651;
	wire [16-1:0] node31654;
	wire [16-1:0] node31655;
	wire [16-1:0] node31657;
	wire [16-1:0] node31660;
	wire [16-1:0] node31661;
	wire [16-1:0] node31662;
	wire [16-1:0] node31666;
	wire [16-1:0] node31668;
	wire [16-1:0] node31671;
	wire [16-1:0] node31672;
	wire [16-1:0] node31673;
	wire [16-1:0] node31675;
	wire [16-1:0] node31678;
	wire [16-1:0] node31679;
	wire [16-1:0] node31682;
	wire [16-1:0] node31684;
	wire [16-1:0] node31685;
	wire [16-1:0] node31689;
	wire [16-1:0] node31690;
	wire [16-1:0] node31692;
	wire [16-1:0] node31694;
	wire [16-1:0] node31697;
	wire [16-1:0] node31699;
	wire [16-1:0] node31702;
	wire [16-1:0] node31703;
	wire [16-1:0] node31704;
	wire [16-1:0] node31705;
	wire [16-1:0] node31708;
	wire [16-1:0] node31710;
	wire [16-1:0] node31711;
	wire [16-1:0] node31715;
	wire [16-1:0] node31716;
	wire [16-1:0] node31718;
	wire [16-1:0] node31719;
	wire [16-1:0] node31720;
	wire [16-1:0] node31724;
	wire [16-1:0] node31725;
	wire [16-1:0] node31729;
	wire [16-1:0] node31730;
	wire [16-1:0] node31731;
	wire [16-1:0] node31733;
	wire [16-1:0] node31738;
	wire [16-1:0] node31739;
	wire [16-1:0] node31740;
	wire [16-1:0] node31741;
	wire [16-1:0] node31746;
	wire [16-1:0] node31747;
	wire [16-1:0] node31749;
	wire [16-1:0] node31751;
	wire [16-1:0] node31754;
	wire [16-1:0] node31755;
	wire [16-1:0] node31756;
	wire [16-1:0] node31760;
	wire [16-1:0] node31761;
	wire [16-1:0] node31763;
	wire [16-1:0] node31767;
	wire [16-1:0] node31768;
	wire [16-1:0] node31769;
	wire [16-1:0] node31770;
	wire [16-1:0] node31771;
	wire [16-1:0] node31772;
	wire [16-1:0] node31773;
	wire [16-1:0] node31774;
	wire [16-1:0] node31775;
	wire [16-1:0] node31777;
	wire [16-1:0] node31781;
	wire [16-1:0] node31783;
	wire [16-1:0] node31786;
	wire [16-1:0] node31788;
	wire [16-1:0] node31791;
	wire [16-1:0] node31792;
	wire [16-1:0] node31793;
	wire [16-1:0] node31794;
	wire [16-1:0] node31799;
	wire [16-1:0] node31800;
	wire [16-1:0] node31801;
	wire [16-1:0] node31806;
	wire [16-1:0] node31807;
	wire [16-1:0] node31808;
	wire [16-1:0] node31811;
	wire [16-1:0] node31812;
	wire [16-1:0] node31816;
	wire [16-1:0] node31817;
	wire [16-1:0] node31819;
	wire [16-1:0] node31823;
	wire [16-1:0] node31824;
	wire [16-1:0] node31825;
	wire [16-1:0] node31826;
	wire [16-1:0] node31827;
	wire [16-1:0] node31828;
	wire [16-1:0] node31833;
	wire [16-1:0] node31836;
	wire [16-1:0] node31837;
	wire [16-1:0] node31838;
	wire [16-1:0] node31842;
	wire [16-1:0] node31843;
	wire [16-1:0] node31845;
	wire [16-1:0] node31848;
	wire [16-1:0] node31851;
	wire [16-1:0] node31852;
	wire [16-1:0] node31853;
	wire [16-1:0] node31855;
	wire [16-1:0] node31859;
	wire [16-1:0] node31860;
	wire [16-1:0] node31861;
	wire [16-1:0] node31865;
	wire [16-1:0] node31866;
	wire [16-1:0] node31867;
	wire [16-1:0] node31871;
	wire [16-1:0] node31874;
	wire [16-1:0] node31875;
	wire [16-1:0] node31876;
	wire [16-1:0] node31877;
	wire [16-1:0] node31878;
	wire [16-1:0] node31879;
	wire [16-1:0] node31882;
	wire [16-1:0] node31885;
	wire [16-1:0] node31886;
	wire [16-1:0] node31888;
	wire [16-1:0] node31889;
	wire [16-1:0] node31893;
	wire [16-1:0] node31896;
	wire [16-1:0] node31897;
	wire [16-1:0] node31898;
	wire [16-1:0] node31900;
	wire [16-1:0] node31901;
	wire [16-1:0] node31905;
	wire [16-1:0] node31906;
	wire [16-1:0] node31910;
	wire [16-1:0] node31912;
	wire [16-1:0] node31915;
	wire [16-1:0] node31916;
	wire [16-1:0] node31917;
	wire [16-1:0] node31918;
	wire [16-1:0] node31921;
	wire [16-1:0] node31924;
	wire [16-1:0] node31925;
	wire [16-1:0] node31926;
	wire [16-1:0] node31928;
	wire [16-1:0] node31933;
	wire [16-1:0] node31934;
	wire [16-1:0] node31936;
	wire [16-1:0] node31939;
	wire [16-1:0] node31940;
	wire [16-1:0] node31943;
	wire [16-1:0] node31946;
	wire [16-1:0] node31947;
	wire [16-1:0] node31948;
	wire [16-1:0] node31950;
	wire [16-1:0] node31951;
	wire [16-1:0] node31953;
	wire [16-1:0] node31954;
	wire [16-1:0] node31958;
	wire [16-1:0] node31961;
	wire [16-1:0] node31962;
	wire [16-1:0] node31963;
	wire [16-1:0] node31966;
	wire [16-1:0] node31969;
	wire [16-1:0] node31971;
	wire [16-1:0] node31972;
	wire [16-1:0] node31973;
	wire [16-1:0] node31978;
	wire [16-1:0] node31979;
	wire [16-1:0] node31980;
	wire [16-1:0] node31981;
	wire [16-1:0] node31984;
	wire [16-1:0] node31986;
	wire [16-1:0] node31987;
	wire [16-1:0] node31991;
	wire [16-1:0] node31992;
	wire [16-1:0] node31995;
	wire [16-1:0] node31997;
	wire [16-1:0] node32000;
	wire [16-1:0] node32001;
	wire [16-1:0] node32002;
	wire [16-1:0] node32003;
	wire [16-1:0] node32007;
	wire [16-1:0] node32008;
	wire [16-1:0] node32011;
	wire [16-1:0] node32012;
	wire [16-1:0] node32016;
	wire [16-1:0] node32017;
	wire [16-1:0] node32021;
	wire [16-1:0] node32022;
	wire [16-1:0] node32023;
	wire [16-1:0] node32024;
	wire [16-1:0] node32025;
	wire [16-1:0] node32026;
	wire [16-1:0] node32027;
	wire [16-1:0] node32031;
	wire [16-1:0] node32032;
	wire [16-1:0] node32035;
	wire [16-1:0] node32038;
	wire [16-1:0] node32040;
	wire [16-1:0] node32043;
	wire [16-1:0] node32044;
	wire [16-1:0] node32045;
	wire [16-1:0] node32046;
	wire [16-1:0] node32050;
	wire [16-1:0] node32051;
	wire [16-1:0] node32055;
	wire [16-1:0] node32056;
	wire [16-1:0] node32057;
	wire [16-1:0] node32059;
	wire [16-1:0] node32062;
	wire [16-1:0] node32064;
	wire [16-1:0] node32067;
	wire [16-1:0] node32068;
	wire [16-1:0] node32070;
	wire [16-1:0] node32074;
	wire [16-1:0] node32075;
	wire [16-1:0] node32076;
	wire [16-1:0] node32077;
	wire [16-1:0] node32078;
	wire [16-1:0] node32079;
	wire [16-1:0] node32083;
	wire [16-1:0] node32085;
	wire [16-1:0] node32086;
	wire [16-1:0] node32090;
	wire [16-1:0] node32092;
	wire [16-1:0] node32094;
	wire [16-1:0] node32097;
	wire [16-1:0] node32098;
	wire [16-1:0] node32099;
	wire [16-1:0] node32102;
	wire [16-1:0] node32105;
	wire [16-1:0] node32106;
	wire [16-1:0] node32108;
	wire [16-1:0] node32109;
	wire [16-1:0] node32114;
	wire [16-1:0] node32115;
	wire [16-1:0] node32116;
	wire [16-1:0] node32117;
	wire [16-1:0] node32118;
	wire [16-1:0] node32122;
	wire [16-1:0] node32123;
	wire [16-1:0] node32125;
	wire [16-1:0] node32129;
	wire [16-1:0] node32130;
	wire [16-1:0] node32134;
	wire [16-1:0] node32135;
	wire [16-1:0] node32139;
	wire [16-1:0] node32140;
	wire [16-1:0] node32141;
	wire [16-1:0] node32142;
	wire [16-1:0] node32143;
	wire [16-1:0] node32144;
	wire [16-1:0] node32145;
	wire [16-1:0] node32149;
	wire [16-1:0] node32151;
	wire [16-1:0] node32154;
	wire [16-1:0] node32155;
	wire [16-1:0] node32158;
	wire [16-1:0] node32161;
	wire [16-1:0] node32162;
	wire [16-1:0] node32163;
	wire [16-1:0] node32166;
	wire [16-1:0] node32168;
	wire [16-1:0] node32171;
	wire [16-1:0] node32172;
	wire [16-1:0] node32174;
	wire [16-1:0] node32175;
	wire [16-1:0] node32179;
	wire [16-1:0] node32182;
	wire [16-1:0] node32183;
	wire [16-1:0] node32184;
	wire [16-1:0] node32185;
	wire [16-1:0] node32189;
	wire [16-1:0] node32190;
	wire [16-1:0] node32193;
	wire [16-1:0] node32195;
	wire [16-1:0] node32198;
	wire [16-1:0] node32199;
	wire [16-1:0] node32200;
	wire [16-1:0] node32203;
	wire [16-1:0] node32206;
	wire [16-1:0] node32207;
	wire [16-1:0] node32208;
	wire [16-1:0] node32213;
	wire [16-1:0] node32214;
	wire [16-1:0] node32215;
	wire [16-1:0] node32216;
	wire [16-1:0] node32217;
	wire [16-1:0] node32218;
	wire [16-1:0] node32222;
	wire [16-1:0] node32226;
	wire [16-1:0] node32227;
	wire [16-1:0] node32228;
	wire [16-1:0] node32231;
	wire [16-1:0] node32233;
	wire [16-1:0] node32236;
	wire [16-1:0] node32237;
	wire [16-1:0] node32240;
	wire [16-1:0] node32241;
	wire [16-1:0] node32244;
	wire [16-1:0] node32245;
	wire [16-1:0] node32249;
	wire [16-1:0] node32250;
	wire [16-1:0] node32251;
	wire [16-1:0] node32253;
	wire [16-1:0] node32255;
	wire [16-1:0] node32257;
	wire [16-1:0] node32261;
	wire [16-1:0] node32262;
	wire [16-1:0] node32263;
	wire [16-1:0] node32264;
	wire [16-1:0] node32269;
	wire [16-1:0] node32270;
	wire [16-1:0] node32273;
	wire [16-1:0] node32276;
	wire [16-1:0] node32277;
	wire [16-1:0] node32278;
	wire [16-1:0] node32279;
	wire [16-1:0] node32280;
	wire [16-1:0] node32281;
	wire [16-1:0] node32282;
	wire [16-1:0] node32283;
	wire [16-1:0] node32284;
	wire [16-1:0] node32286;
	wire [16-1:0] node32289;
	wire [16-1:0] node32292;
	wire [16-1:0] node32293;
	wire [16-1:0] node32295;
	wire [16-1:0] node32298;
	wire [16-1:0] node32301;
	wire [16-1:0] node32302;
	wire [16-1:0] node32303;
	wire [16-1:0] node32304;
	wire [16-1:0] node32308;
	wire [16-1:0] node32310;
	wire [16-1:0] node32311;
	wire [16-1:0] node32315;
	wire [16-1:0] node32316;
	wire [16-1:0] node32317;
	wire [16-1:0] node32322;
	wire [16-1:0] node32323;
	wire [16-1:0] node32324;
	wire [16-1:0] node32325;
	wire [16-1:0] node32329;
	wire [16-1:0] node32330;
	wire [16-1:0] node32334;
	wire [16-1:0] node32335;
	wire [16-1:0] node32336;
	wire [16-1:0] node32337;
	wire [16-1:0] node32341;
	wire [16-1:0] node32342;
	wire [16-1:0] node32343;
	wire [16-1:0] node32348;
	wire [16-1:0] node32349;
	wire [16-1:0] node32351;
	wire [16-1:0] node32354;
	wire [16-1:0] node32357;
	wire [16-1:0] node32358;
	wire [16-1:0] node32359;
	wire [16-1:0] node32360;
	wire [16-1:0] node32362;
	wire [16-1:0] node32364;
	wire [16-1:0] node32365;
	wire [16-1:0] node32368;
	wire [16-1:0] node32371;
	wire [16-1:0] node32373;
	wire [16-1:0] node32374;
	wire [16-1:0] node32375;
	wire [16-1:0] node32380;
	wire [16-1:0] node32382;
	wire [16-1:0] node32383;
	wire [16-1:0] node32387;
	wire [16-1:0] node32388;
	wire [16-1:0] node32389;
	wire [16-1:0] node32391;
	wire [16-1:0] node32394;
	wire [16-1:0] node32395;
	wire [16-1:0] node32398;
	wire [16-1:0] node32401;
	wire [16-1:0] node32402;
	wire [16-1:0] node32403;
	wire [16-1:0] node32406;
	wire [16-1:0] node32407;
	wire [16-1:0] node32411;
	wire [16-1:0] node32413;
	wire [16-1:0] node32416;
	wire [16-1:0] node32417;
	wire [16-1:0] node32418;
	wire [16-1:0] node32419;
	wire [16-1:0] node32420;
	wire [16-1:0] node32422;
	wire [16-1:0] node32425;
	wire [16-1:0] node32426;
	wire [16-1:0] node32430;
	wire [16-1:0] node32431;
	wire [16-1:0] node32434;
	wire [16-1:0] node32435;
	wire [16-1:0] node32437;
	wire [16-1:0] node32438;
	wire [16-1:0] node32442;
	wire [16-1:0] node32445;
	wire [16-1:0] node32446;
	wire [16-1:0] node32447;
	wire [16-1:0] node32448;
	wire [16-1:0] node32451;
	wire [16-1:0] node32453;
	wire [16-1:0] node32456;
	wire [16-1:0] node32457;
	wire [16-1:0] node32461;
	wire [16-1:0] node32462;
	wire [16-1:0] node32463;
	wire [16-1:0] node32465;
	wire [16-1:0] node32466;
	wire [16-1:0] node32470;
	wire [16-1:0] node32471;
	wire [16-1:0] node32475;
	wire [16-1:0] node32476;
	wire [16-1:0] node32478;
	wire [16-1:0] node32479;
	wire [16-1:0] node32484;
	wire [16-1:0] node32485;
	wire [16-1:0] node32486;
	wire [16-1:0] node32487;
	wire [16-1:0] node32488;
	wire [16-1:0] node32490;
	wire [16-1:0] node32493;
	wire [16-1:0] node32496;
	wire [16-1:0] node32498;
	wire [16-1:0] node32499;
	wire [16-1:0] node32503;
	wire [16-1:0] node32504;
	wire [16-1:0] node32505;
	wire [16-1:0] node32508;
	wire [16-1:0] node32510;
	wire [16-1:0] node32511;
	wire [16-1:0] node32515;
	wire [16-1:0] node32516;
	wire [16-1:0] node32517;
	wire [16-1:0] node32521;
	wire [16-1:0] node32524;
	wire [16-1:0] node32525;
	wire [16-1:0] node32526;
	wire [16-1:0] node32529;
	wire [16-1:0] node32530;
	wire [16-1:0] node32533;
	wire [16-1:0] node32534;
	wire [16-1:0] node32538;
	wire [16-1:0] node32539;
	wire [16-1:0] node32541;
	wire [16-1:0] node32544;
	wire [16-1:0] node32545;
	wire [16-1:0] node32547;
	wire [16-1:0] node32550;
	wire [16-1:0] node32551;
	wire [16-1:0] node32554;
	wire [16-1:0] node32556;
	wire [16-1:0] node32559;
	wire [16-1:0] node32560;
	wire [16-1:0] node32561;
	wire [16-1:0] node32562;
	wire [16-1:0] node32563;
	wire [16-1:0] node32565;
	wire [16-1:0] node32566;
	wire [16-1:0] node32568;
	wire [16-1:0] node32572;
	wire [16-1:0] node32573;
	wire [16-1:0] node32574;
	wire [16-1:0] node32578;
	wire [16-1:0] node32579;
	wire [16-1:0] node32581;
	wire [16-1:0] node32585;
	wire [16-1:0] node32586;
	wire [16-1:0] node32587;
	wire [16-1:0] node32588;
	wire [16-1:0] node32589;
	wire [16-1:0] node32594;
	wire [16-1:0] node32595;
	wire [16-1:0] node32598;
	wire [16-1:0] node32600;
	wire [16-1:0] node32603;
	wire [16-1:0] node32604;
	wire [16-1:0] node32605;
	wire [16-1:0] node32609;
	wire [16-1:0] node32610;
	wire [16-1:0] node32611;
	wire [16-1:0] node32616;
	wire [16-1:0] node32617;
	wire [16-1:0] node32618;
	wire [16-1:0] node32620;
	wire [16-1:0] node32621;
	wire [16-1:0] node32624;
	wire [16-1:0] node32627;
	wire [16-1:0] node32628;
	wire [16-1:0] node32629;
	wire [16-1:0] node32630;
	wire [16-1:0] node32634;
	wire [16-1:0] node32636;
	wire [16-1:0] node32639;
	wire [16-1:0] node32641;
	wire [16-1:0] node32643;
	wire [16-1:0] node32646;
	wire [16-1:0] node32647;
	wire [16-1:0] node32648;
	wire [16-1:0] node32649;
	wire [16-1:0] node32652;
	wire [16-1:0] node32653;
	wire [16-1:0] node32655;
	wire [16-1:0] node32659;
	wire [16-1:0] node32660;
	wire [16-1:0] node32662;
	wire [16-1:0] node32665;
	wire [16-1:0] node32668;
	wire [16-1:0] node32669;
	wire [16-1:0] node32670;
	wire [16-1:0] node32671;
	wire [16-1:0] node32675;
	wire [16-1:0] node32678;
	wire [16-1:0] node32679;
	wire [16-1:0] node32683;
	wire [16-1:0] node32684;
	wire [16-1:0] node32685;
	wire [16-1:0] node32686;
	wire [16-1:0] node32687;
	wire [16-1:0] node32688;
	wire [16-1:0] node32692;
	wire [16-1:0] node32693;
	wire [16-1:0] node32696;
	wire [16-1:0] node32698;
	wire [16-1:0] node32701;
	wire [16-1:0] node32702;
	wire [16-1:0] node32703;
	wire [16-1:0] node32706;
	wire [16-1:0] node32708;
	wire [16-1:0] node32711;
	wire [16-1:0] node32712;
	wire [16-1:0] node32715;
	wire [16-1:0] node32716;
	wire [16-1:0] node32718;
	wire [16-1:0] node32722;
	wire [16-1:0] node32723;
	wire [16-1:0] node32724;
	wire [16-1:0] node32725;
	wire [16-1:0] node32726;
	wire [16-1:0] node32728;
	wire [16-1:0] node32731;
	wire [16-1:0] node32734;
	wire [16-1:0] node32736;
	wire [16-1:0] node32739;
	wire [16-1:0] node32740;
	wire [16-1:0] node32744;
	wire [16-1:0] node32745;
	wire [16-1:0] node32746;
	wire [16-1:0] node32747;
	wire [16-1:0] node32752;
	wire [16-1:0] node32754;
	wire [16-1:0] node32756;
	wire [16-1:0] node32758;
	wire [16-1:0] node32761;
	wire [16-1:0] node32762;
	wire [16-1:0] node32763;
	wire [16-1:0] node32764;
	wire [16-1:0] node32766;
	wire [16-1:0] node32769;
	wire [16-1:0] node32770;
	wire [16-1:0] node32773;
	wire [16-1:0] node32776;
	wire [16-1:0] node32777;
	wire [16-1:0] node32778;
	wire [16-1:0] node32782;
	wire [16-1:0] node32785;
	wire [16-1:0] node32786;
	wire [16-1:0] node32787;
	wire [16-1:0] node32788;
	wire [16-1:0] node32789;
	wire [16-1:0] node32793;
	wire [16-1:0] node32795;
	wire [16-1:0] node32796;
	wire [16-1:0] node32800;
	wire [16-1:0] node32801;
	wire [16-1:0] node32804;
	wire [16-1:0] node32806;
	wire [16-1:0] node32808;
	wire [16-1:0] node32811;
	wire [16-1:0] node32812;
	wire [16-1:0] node32814;
	wire [16-1:0] node32817;
	wire [16-1:0] node32819;
	wire [16-1:0] node32821;
	wire [16-1:0] node32823;
	wire [16-1:0] node32826;
	wire [16-1:0] node32827;
	wire [16-1:0] node32828;
	wire [16-1:0] node32829;
	wire [16-1:0] node32830;
	wire [16-1:0] node32831;
	wire [16-1:0] node32832;
	wire [16-1:0] node32834;
	wire [16-1:0] node32835;
	wire [16-1:0] node32839;
	wire [16-1:0] node32840;
	wire [16-1:0] node32843;
	wire [16-1:0] node32844;
	wire [16-1:0] node32848;
	wire [16-1:0] node32849;
	wire [16-1:0] node32851;
	wire [16-1:0] node32852;
	wire [16-1:0] node32854;
	wire [16-1:0] node32858;
	wire [16-1:0] node32859;
	wire [16-1:0] node32860;
	wire [16-1:0] node32864;
	wire [16-1:0] node32867;
	wire [16-1:0] node32868;
	wire [16-1:0] node32871;
	wire [16-1:0] node32873;
	wire [16-1:0] node32876;
	wire [16-1:0] node32877;
	wire [16-1:0] node32878;
	wire [16-1:0] node32879;
	wire [16-1:0] node32881;
	wire [16-1:0] node32882;
	wire [16-1:0] node32886;
	wire [16-1:0] node32888;
	wire [16-1:0] node32891;
	wire [16-1:0] node32892;
	wire [16-1:0] node32893;
	wire [16-1:0] node32896;
	wire [16-1:0] node32899;
	wire [16-1:0] node32901;
	wire [16-1:0] node32904;
	wire [16-1:0] node32905;
	wire [16-1:0] node32906;
	wire [16-1:0] node32907;
	wire [16-1:0] node32910;
	wire [16-1:0] node32913;
	wire [16-1:0] node32914;
	wire [16-1:0] node32915;
	wire [16-1:0] node32919;
	wire [16-1:0] node32922;
	wire [16-1:0] node32923;
	wire [16-1:0] node32924;
	wire [16-1:0] node32927;
	wire [16-1:0] node32930;
	wire [16-1:0] node32931;
	wire [16-1:0] node32933;
	wire [16-1:0] node32936;
	wire [16-1:0] node32939;
	wire [16-1:0] node32940;
	wire [16-1:0] node32941;
	wire [16-1:0] node32942;
	wire [16-1:0] node32943;
	wire [16-1:0] node32944;
	wire [16-1:0] node32947;
	wire [16-1:0] node32949;
	wire [16-1:0] node32952;
	wire [16-1:0] node32953;
	wire [16-1:0] node32955;
	wire [16-1:0] node32958;
	wire [16-1:0] node32961;
	wire [16-1:0] node32962;
	wire [16-1:0] node32963;
	wire [16-1:0] node32964;
	wire [16-1:0] node32968;
	wire [16-1:0] node32969;
	wire [16-1:0] node32970;
	wire [16-1:0] node32975;
	wire [16-1:0] node32978;
	wire [16-1:0] node32979;
	wire [16-1:0] node32980;
	wire [16-1:0] node32982;
	wire [16-1:0] node32985;
	wire [16-1:0] node32986;
	wire [16-1:0] node32988;
	wire [16-1:0] node32989;
	wire [16-1:0] node32994;
	wire [16-1:0] node32995;
	wire [16-1:0] node32996;
	wire [16-1:0] node32998;
	wire [16-1:0] node32999;
	wire [16-1:0] node33003;
	wire [16-1:0] node33006;
	wire [16-1:0] node33007;
	wire [16-1:0] node33010;
	wire [16-1:0] node33011;
	wire [16-1:0] node33013;
	wire [16-1:0] node33017;
	wire [16-1:0] node33018;
	wire [16-1:0] node33019;
	wire [16-1:0] node33020;
	wire [16-1:0] node33022;
	wire [16-1:0] node33025;
	wire [16-1:0] node33027;
	wire [16-1:0] node33030;
	wire [16-1:0] node33031;
	wire [16-1:0] node33032;
	wire [16-1:0] node33035;
	wire [16-1:0] node33036;
	wire [16-1:0] node33039;
	wire [16-1:0] node33041;
	wire [16-1:0] node33044;
	wire [16-1:0] node33046;
	wire [16-1:0] node33047;
	wire [16-1:0] node33051;
	wire [16-1:0] node33052;
	wire [16-1:0] node33054;
	wire [16-1:0] node33055;
	wire [16-1:0] node33058;
	wire [16-1:0] node33061;
	wire [16-1:0] node33062;
	wire [16-1:0] node33063;
	wire [16-1:0] node33065;
	wire [16-1:0] node33069;
	wire [16-1:0] node33071;
	wire [16-1:0] node33074;
	wire [16-1:0] node33075;
	wire [16-1:0] node33076;
	wire [16-1:0] node33077;
	wire [16-1:0] node33078;
	wire [16-1:0] node33079;
	wire [16-1:0] node33080;
	wire [16-1:0] node33083;
	wire [16-1:0] node33084;
	wire [16-1:0] node33088;
	wire [16-1:0] node33090;
	wire [16-1:0] node33093;
	wire [16-1:0] node33094;
	wire [16-1:0] node33097;
	wire [16-1:0] node33098;
	wire [16-1:0] node33099;
	wire [16-1:0] node33103;
	wire [16-1:0] node33106;
	wire [16-1:0] node33107;
	wire [16-1:0] node33108;
	wire [16-1:0] node33110;
	wire [16-1:0] node33113;
	wire [16-1:0] node33114;
	wire [16-1:0] node33116;
	wire [16-1:0] node33119;
	wire [16-1:0] node33121;
	wire [16-1:0] node33124;
	wire [16-1:0] node33125;
	wire [16-1:0] node33126;
	wire [16-1:0] node33129;
	wire [16-1:0] node33131;
	wire [16-1:0] node33132;
	wire [16-1:0] node33136;
	wire [16-1:0] node33137;
	wire [16-1:0] node33139;
	wire [16-1:0] node33140;
	wire [16-1:0] node33144;
	wire [16-1:0] node33145;
	wire [16-1:0] node33148;
	wire [16-1:0] node33151;
	wire [16-1:0] node33152;
	wire [16-1:0] node33153;
	wire [16-1:0] node33154;
	wire [16-1:0] node33157;
	wire [16-1:0] node33158;
	wire [16-1:0] node33159;
	wire [16-1:0] node33163;
	wire [16-1:0] node33165;
	wire [16-1:0] node33166;
	wire [16-1:0] node33170;
	wire [16-1:0] node33171;
	wire [16-1:0] node33173;
	wire [16-1:0] node33176;
	wire [16-1:0] node33177;
	wire [16-1:0] node33181;
	wire [16-1:0] node33182;
	wire [16-1:0] node33183;
	wire [16-1:0] node33185;
	wire [16-1:0] node33188;
	wire [16-1:0] node33191;
	wire [16-1:0] node33193;
	wire [16-1:0] node33196;
	wire [16-1:0] node33197;
	wire [16-1:0] node33198;
	wire [16-1:0] node33199;
	wire [16-1:0] node33200;
	wire [16-1:0] node33202;
	wire [16-1:0] node33206;
	wire [16-1:0] node33208;
	wire [16-1:0] node33209;
	wire [16-1:0] node33211;
	wire [16-1:0] node33214;
	wire [16-1:0] node33217;
	wire [16-1:0] node33218;
	wire [16-1:0] node33219;
	wire [16-1:0] node33221;
	wire [16-1:0] node33224;
	wire [16-1:0] node33225;
	wire [16-1:0] node33226;
	wire [16-1:0] node33230;
	wire [16-1:0] node33232;
	wire [16-1:0] node33235;
	wire [16-1:0] node33236;
	wire [16-1:0] node33237;
	wire [16-1:0] node33240;
	wire [16-1:0] node33243;
	wire [16-1:0] node33245;
	wire [16-1:0] node33247;
	wire [16-1:0] node33250;
	wire [16-1:0] node33251;
	wire [16-1:0] node33252;
	wire [16-1:0] node33253;
	wire [16-1:0] node33255;
	wire [16-1:0] node33259;
	wire [16-1:0] node33260;
	wire [16-1:0] node33261;
	wire [16-1:0] node33264;
	wire [16-1:0] node33266;
	wire [16-1:0] node33269;
	wire [16-1:0] node33270;
	wire [16-1:0] node33273;
	wire [16-1:0] node33275;
	wire [16-1:0] node33278;
	wire [16-1:0] node33279;
	wire [16-1:0] node33280;
	wire [16-1:0] node33282;
	wire [16-1:0] node33285;
	wire [16-1:0] node33286;
	wire [16-1:0] node33290;
	wire [16-1:0] node33291;
	wire [16-1:0] node33292;
	wire [16-1:0] node33294;
	wire [16-1:0] node33297;
	wire [16-1:0] node33298;
	wire [16-1:0] node33300;
	wire [16-1:0] node33304;
	wire [16-1:0] node33305;
	wire [16-1:0] node33306;
	wire [16-1:0] node33308;
	wire [16-1:0] node33311;
	wire [16-1:0] node33312;
	wire [16-1:0] node33316;

	assign outp = (inp[0]) ? node16642 : node1;
		assign node1 = (inp[4]) ? node8371 : node2;
			assign node2 = (inp[10]) ? node4156 : node3;
				assign node3 = (inp[11]) ? node2093 : node4;
					assign node4 = (inp[9]) ? node1080 : node5;
						assign node5 = (inp[15]) ? node555 : node6;
							assign node6 = (inp[6]) ? node292 : node7;
								assign node7 = (inp[2]) ? node161 : node8;
									assign node8 = (inp[7]) ? node94 : node9;
										assign node9 = (inp[12]) ? node61 : node10;
											assign node10 = (inp[8]) ? node40 : node11;
												assign node11 = (inp[14]) ? node29 : node12;
													assign node12 = (inp[13]) ? node20 : node13;
														assign node13 = (inp[5]) ? 16'b0011111111111111 : node14;
															assign node14 = (inp[3]) ? 16'b0111111111111111 : node15;
																assign node15 = (inp[1]) ? 16'b0111111111111111 : 16'b1111111111111111;
														assign node20 = (inp[1]) ? node24 : node21;
															assign node21 = (inp[3]) ? 16'b0011111111111111 : 16'b0111111111111111;
															assign node24 = (inp[5]) ? 16'b0001111111111111 : node25;
																assign node25 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node29 = (inp[3]) ? node37 : node30;
														assign node30 = (inp[13]) ? node32 : 16'b0011111111111111;
															assign node32 = (inp[1]) ? 16'b0001111111111111 : node33;
																assign node33 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node37 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node40 = (inp[13]) ? node56 : node41;
													assign node41 = (inp[5]) ? node53 : node42;
														assign node42 = (inp[1]) ? node48 : node43;
															assign node43 = (inp[14]) ? node45 : 16'b0011111111111111;
																assign node45 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node48 = (inp[14]) ? 16'b0001111111111111 : node49;
																assign node49 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node53 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node56 = (inp[14]) ? 16'b0000111111111111 : node57;
														assign node57 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node61 = (inp[3]) ? node79 : node62;
												assign node62 = (inp[5]) ? node70 : node63;
													assign node63 = (inp[13]) ? node65 : 16'b0001111111111111;
														assign node65 = (inp[8]) ? 16'b0001111111111111 : node66;
															assign node66 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node70 = (inp[14]) ? node74 : node71;
														assign node71 = (inp[1]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node74 = (inp[8]) ? node76 : 16'b0000111111111111;
															assign node76 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node79 = (inp[5]) ? node89 : node80;
													assign node80 = (inp[8]) ? node84 : node81;
														assign node81 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node84 = (inp[1]) ? 16'b0000011111111111 : node85;
															assign node85 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node89 = (inp[1]) ? node91 : 16'b0000011111111111;
														assign node91 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node94 = (inp[13]) ? node126 : node95;
											assign node95 = (inp[3]) ? node115 : node96;
												assign node96 = (inp[8]) ? node112 : node97;
													assign node97 = (inp[1]) ? node107 : node98;
														assign node98 = (inp[5]) ? node104 : node99;
															assign node99 = (inp[12]) ? 16'b0011111111111111 : node100;
																assign node100 = (inp[14]) ? 16'b0011111111111111 : 16'b0111111111111111;
															assign node104 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node107 = (inp[12]) ? 16'b0000111111111111 : node108;
															assign node108 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node112 = (inp[14]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node115 = (inp[5]) ? node117 : 16'b0000111111111111;
													assign node117 = (inp[8]) ? 16'b0000001111111111 : node118;
														assign node118 = (inp[1]) ? node120 : 16'b0000111111111111;
															assign node120 = (inp[12]) ? node122 : 16'b0000011111111111;
																assign node122 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node126 = (inp[8]) ? node142 : node127;
												assign node127 = (inp[5]) ? node139 : node128;
													assign node128 = (inp[12]) ? node136 : node129;
														assign node129 = (inp[1]) ? node131 : 16'b0000111111111111;
															assign node131 = (inp[3]) ? node133 : 16'b0000111111111111;
																assign node133 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node136 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node139 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node142 = (inp[1]) ? node150 : node143;
													assign node143 = (inp[3]) ? node147 : node144;
														assign node144 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node147 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node150 = (inp[3]) ? node156 : node151;
														assign node151 = (inp[5]) ? node153 : 16'b0000011111111111;
															assign node153 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node156 = (inp[12]) ? 16'b0000000111111111 : node157;
															assign node157 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node161 = (inp[1]) ? node241 : node162;
										assign node162 = (inp[7]) ? node210 : node163;
											assign node163 = (inp[13]) ? node183 : node164;
												assign node164 = (inp[5]) ? node176 : node165;
													assign node165 = (inp[12]) ? node167 : 16'b0011111111111111;
														assign node167 = (inp[14]) ? node171 : node168;
															assign node168 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node171 = (inp[8]) ? 16'b0000111111111111 : node172;
																assign node172 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node176 = (inp[12]) ? node180 : node177;
														assign node177 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node180 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node183 = (inp[3]) ? node191 : node184;
													assign node184 = (inp[14]) ? node188 : node185;
														assign node185 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node188 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node191 = (inp[12]) ? node203 : node192;
														assign node192 = (inp[8]) ? node198 : node193;
															assign node193 = (inp[5]) ? node195 : 16'b0000111111111111;
																assign node195 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node198 = (inp[5]) ? 16'b0000011111111111 : node199;
																assign node199 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node203 = (inp[8]) ? 16'b0000011111111111 : node204;
															assign node204 = (inp[5]) ? 16'b0000011111111111 : node205;
																assign node205 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node210 = (inp[12]) ? node222 : node211;
												assign node211 = (inp[3]) ? 16'b0000011111111111 : node212;
													assign node212 = (inp[14]) ? node216 : node213;
														assign node213 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node216 = (inp[5]) ? node218 : 16'b0000111111111111;
															assign node218 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node222 = (inp[5]) ? node234 : node223;
													assign node223 = (inp[14]) ? node227 : node224;
														assign node224 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node227 = (inp[3]) ? 16'b0000001111111111 : node228;
															assign node228 = (inp[8]) ? node230 : 16'b0000011111111111;
																assign node230 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node234 = (inp[8]) ? node238 : node235;
														assign node235 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node238 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node241 = (inp[12]) ? node267 : node242;
											assign node242 = (inp[14]) ? node256 : node243;
												assign node243 = (inp[13]) ? node247 : node244;
													assign node244 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node247 = (inp[7]) ? node249 : 16'b0000111111111111;
														assign node249 = (inp[8]) ? node253 : node250;
															assign node250 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node253 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node256 = (inp[3]) ? node262 : node257;
													assign node257 = (inp[5]) ? node259 : 16'b0000111111111111;
														assign node259 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node262 = (inp[8]) ? 16'b0000001111111111 : node263;
														assign node263 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node267 = (inp[8]) ? node279 : node268;
												assign node268 = (inp[13]) ? node270 : 16'b0000011111111111;
													assign node270 = (inp[7]) ? node274 : node271;
														assign node271 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node274 = (inp[14]) ? 16'b0000000111111111 : node275;
															assign node275 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node279 = (inp[14]) ? node289 : node280;
													assign node280 = (inp[5]) ? node286 : node281;
														assign node281 = (inp[7]) ? 16'b0000001111111111 : node282;
															assign node282 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node286 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node289 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node292 = (inp[13]) ? node452 : node293;
									assign node293 = (inp[3]) ? node365 : node294;
										assign node294 = (inp[14]) ? node326 : node295;
											assign node295 = (inp[12]) ? node317 : node296;
												assign node296 = (inp[1]) ? node310 : node297;
													assign node297 = (inp[5]) ? node305 : node298;
														assign node298 = (inp[2]) ? node300 : 16'b0111111111111111;
															assign node300 = (inp[8]) ? 16'b0001111111111111 : node301;
																assign node301 = (inp[7]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node305 = (inp[8]) ? node307 : 16'b0001111111111111;
															assign node307 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node310 = (inp[8]) ? node314 : node311;
														assign node311 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node314 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node317 = (inp[2]) ? node319 : 16'b0000111111111111;
													assign node319 = (inp[7]) ? node323 : node320;
														assign node320 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node323 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node326 = (inp[8]) ? node350 : node327;
												assign node327 = (inp[7]) ? node343 : node328;
													assign node328 = (inp[1]) ? node336 : node329;
														assign node329 = (inp[2]) ? 16'b0000111111111111 : node330;
															assign node330 = (inp[5]) ? node332 : 16'b0001111111111111;
																assign node332 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node336 = (inp[12]) ? 16'b0000011111111111 : node337;
															assign node337 = (inp[2]) ? node339 : 16'b0000111111111111;
																assign node339 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node343 = (inp[5]) ? node347 : node344;
														assign node344 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node347 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node350 = (inp[5]) ? node354 : node351;
													assign node351 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node354 = (inp[12]) ? node362 : node355;
														assign node355 = (inp[2]) ? node357 : 16'b0000011111111111;
															assign node357 = (inp[1]) ? 16'b0000001111111111 : node358;
																assign node358 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node362 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node365 = (inp[5]) ? node403 : node366;
											assign node366 = (inp[2]) ? node386 : node367;
												assign node367 = (inp[7]) ? node373 : node368;
													assign node368 = (inp[12]) ? node370 : 16'b0000111111111111;
														assign node370 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node373 = (inp[1]) ? node381 : node374;
														assign node374 = (inp[8]) ? node376 : 16'b0000111111111111;
															assign node376 = (inp[12]) ? 16'b0000011111111111 : node377;
																assign node377 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node381 = (inp[8]) ? 16'b0000001111111111 : node382;
															assign node382 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node386 = (inp[7]) ? node396 : node387;
													assign node387 = (inp[12]) ? node393 : node388;
														assign node388 = (inp[8]) ? 16'b0000011111111111 : node389;
															assign node389 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node393 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node396 = (inp[14]) ? node400 : node397;
														assign node397 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node400 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node403 = (inp[8]) ? node431 : node404;
												assign node404 = (inp[12]) ? node420 : node405;
													assign node405 = (inp[14]) ? node415 : node406;
														assign node406 = (inp[2]) ? node412 : node407;
															assign node407 = (inp[7]) ? node409 : 16'b0000111111111111;
																assign node409 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node412 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node415 = (inp[1]) ? node417 : 16'b0000011111111111;
															assign node417 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node420 = (inp[7]) ? node426 : node421;
														assign node421 = (inp[14]) ? node423 : 16'b0000011111111111;
															assign node423 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node426 = (inp[1]) ? node428 : 16'b0000000111111111;
															assign node428 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node431 = (inp[7]) ? node441 : node432;
													assign node432 = (inp[12]) ? node436 : node433;
														assign node433 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node436 = (inp[14]) ? 16'b0000000111111111 : node437;
															assign node437 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node441 = (inp[2]) ? node447 : node442;
														assign node442 = (inp[12]) ? 16'b0000000111111111 : node443;
															assign node443 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node447 = (inp[1]) ? node449 : 16'b0000000111111111;
															assign node449 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node452 = (inp[2]) ? node486 : node453;
										assign node453 = (inp[14]) ? node469 : node454;
											assign node454 = (inp[5]) ? node462 : node455;
												assign node455 = (inp[3]) ? 16'b0000011111111111 : node456;
													assign node456 = (inp[8]) ? node458 : 16'b0001111111111111;
														assign node458 = (inp[1]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node462 = (inp[1]) ? node464 : 16'b0000011111111111;
													assign node464 = (inp[7]) ? 16'b0000001111111111 : node465;
														assign node465 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node469 = (inp[12]) ? node481 : node470;
												assign node470 = (inp[3]) ? node476 : node471;
													assign node471 = (inp[7]) ? 16'b0000011111111111 : node472;
														assign node472 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node476 = (inp[1]) ? node478 : 16'b0000011111111111;
														assign node478 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node481 = (inp[8]) ? node483 : 16'b0000001111111111;
													assign node483 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node486 = (inp[1]) ? node514 : node487;
											assign node487 = (inp[5]) ? node509 : node488;
												assign node488 = (inp[7]) ? node498 : node489;
													assign node489 = (inp[3]) ? node495 : node490;
														assign node490 = (inp[12]) ? 16'b0000011111111111 : node491;
															assign node491 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node495 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node498 = (inp[8]) ? node506 : node499;
														assign node499 = (inp[12]) ? 16'b0000001111111111 : node500;
															assign node500 = (inp[3]) ? node502 : 16'b0000011111111111;
																assign node502 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node506 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node509 = (inp[12]) ? 16'b0000000111111111 : node510;
													assign node510 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node514 = (inp[8]) ? node532 : node515;
												assign node515 = (inp[3]) ? node525 : node516;
													assign node516 = (inp[7]) ? node520 : node517;
														assign node517 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node520 = (inp[12]) ? 16'b0000000111111111 : node521;
															assign node521 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node525 = (inp[7]) ? 16'b0000000011111111 : node526;
														assign node526 = (inp[5]) ? 16'b0000000111111111 : node527;
															assign node527 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node532 = (inp[14]) ? node542 : node533;
													assign node533 = (inp[5]) ? node537 : node534;
														assign node534 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node537 = (inp[7]) ? node539 : 16'b0000000111111111;
															assign node539 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node542 = (inp[3]) ? node546 : node543;
														assign node543 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node546 = (inp[12]) ? node552 : node547;
															assign node547 = (inp[5]) ? node549 : 16'b0000000011111111;
																assign node549 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node552 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node555 = (inp[8]) ? node803 : node556;
								assign node556 = (inp[2]) ? node684 : node557;
									assign node557 = (inp[6]) ? node619 : node558;
										assign node558 = (inp[13]) ? node588 : node559;
											assign node559 = (inp[12]) ? node573 : node560;
												assign node560 = (inp[7]) ? node568 : node561;
													assign node561 = (inp[14]) ? node565 : node562;
														assign node562 = (inp[1]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node565 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node568 = (inp[1]) ? node570 : 16'b0001111111111111;
														assign node570 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node573 = (inp[5]) ? node581 : node574;
													assign node574 = (inp[3]) ? 16'b0000111111111111 : node575;
														assign node575 = (inp[1]) ? node577 : 16'b0001111111111111;
															assign node577 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node581 = (inp[3]) ? 16'b0000001111111111 : node582;
														assign node582 = (inp[1]) ? node584 : 16'b0000011111111111;
															assign node584 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node588 = (inp[1]) ? node612 : node589;
												assign node589 = (inp[14]) ? node603 : node590;
													assign node590 = (inp[7]) ? node592 : 16'b0000111111111111;
														assign node592 = (inp[3]) ? node598 : node593;
															assign node593 = (inp[5]) ? node595 : 16'b0000111111111111;
																assign node595 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node598 = (inp[5]) ? node600 : 16'b0000011111111111;
																assign node600 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node603 = (inp[5]) ? node609 : node604;
														assign node604 = (inp[7]) ? 16'b0000011111111111 : node605;
															assign node605 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node609 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node612 = (inp[14]) ? node614 : 16'b0000011111111111;
													assign node614 = (inp[3]) ? 16'b0000000111111111 : node615;
														assign node615 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node619 = (inp[7]) ? node653 : node620;
											assign node620 = (inp[13]) ? node642 : node621;
												assign node621 = (inp[12]) ? node631 : node622;
													assign node622 = (inp[3]) ? 16'b0000011111111111 : node623;
														assign node623 = (inp[5]) ? node625 : 16'b0001111111111111;
															assign node625 = (inp[1]) ? 16'b0000111111111111 : node626;
																assign node626 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node631 = (inp[14]) ? node637 : node632;
														assign node632 = (inp[1]) ? 16'b0000011111111111 : node633;
															assign node633 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node637 = (inp[1]) ? node639 : 16'b0000011111111111;
															assign node639 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node642 = (inp[1]) ? node648 : node643;
													assign node643 = (inp[5]) ? node645 : 16'b0000011111111111;
														assign node645 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node648 = (inp[5]) ? node650 : 16'b0000001111111111;
														assign node650 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node653 = (inp[3]) ? node671 : node654;
												assign node654 = (inp[14]) ? node660 : node655;
													assign node655 = (inp[5]) ? node657 : 16'b0000011111111111;
														assign node657 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node660 = (inp[5]) ? node668 : node661;
														assign node661 = (inp[13]) ? 16'b0000001111111111 : node662;
															assign node662 = (inp[1]) ? node664 : 16'b0000011111111111;
																assign node664 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node668 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node671 = (inp[12]) ? node677 : node672;
													assign node672 = (inp[14]) ? node674 : 16'b0000001111111111;
														assign node674 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node677 = (inp[1]) ? node679 : 16'b0000000111111111;
														assign node679 = (inp[13]) ? node681 : 16'b0000000111111111;
															assign node681 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node684 = (inp[1]) ? node746 : node685;
										assign node685 = (inp[14]) ? node721 : node686;
											assign node686 = (inp[12]) ? node706 : node687;
												assign node687 = (inp[3]) ? node699 : node688;
													assign node688 = (inp[7]) ? node692 : node689;
														assign node689 = (inp[6]) ? 16'b0000111111111111 : 16'b0011111111111111;
														assign node692 = (inp[6]) ? node696 : node693;
															assign node693 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node696 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node699 = (inp[13]) ? node701 : 16'b0000011111111111;
														assign node701 = (inp[7]) ? node703 : 16'b0000011111111111;
															assign node703 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node706 = (inp[6]) ? node712 : node707;
													assign node707 = (inp[7]) ? node709 : 16'b0001111111111111;
														assign node709 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node712 = (inp[13]) ? node716 : node713;
														assign node713 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node716 = (inp[3]) ? 16'b0000000111111111 : node717;
															assign node717 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node721 = (inp[13]) ? node731 : node722;
												assign node722 = (inp[7]) ? node724 : 16'b0000011111111111;
													assign node724 = (inp[12]) ? 16'b0000000111111111 : node725;
														assign node725 = (inp[6]) ? 16'b0000001111111111 : node726;
															assign node726 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node731 = (inp[6]) ? node741 : node732;
													assign node732 = (inp[12]) ? node736 : node733;
														assign node733 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node736 = (inp[7]) ? node738 : 16'b0000001111111111;
															assign node738 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node741 = (inp[7]) ? 16'b0000000111111111 : node742;
														assign node742 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node746 = (inp[7]) ? node782 : node747;
											assign node747 = (inp[13]) ? node761 : node748;
												assign node748 = (inp[12]) ? 16'b0000001111111111 : node749;
													assign node749 = (inp[3]) ? node753 : node750;
														assign node750 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node753 = (inp[5]) ? 16'b0000001111111111 : node754;
															assign node754 = (inp[6]) ? node756 : 16'b0000011111111111;
																assign node756 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node761 = (inp[3]) ? node773 : node762;
													assign node762 = (inp[12]) ? node764 : 16'b0000001111111111;
														assign node764 = (inp[5]) ? 16'b0000000111111111 : node765;
															assign node765 = (inp[14]) ? node769 : node766;
																assign node766 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
																assign node769 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node773 = (inp[14]) ? node779 : node774;
														assign node774 = (inp[12]) ? node776 : 16'b0000001111111111;
															assign node776 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node779 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node782 = (inp[5]) ? node790 : node783;
												assign node783 = (inp[12]) ? node785 : 16'b0000001111111111;
													assign node785 = (inp[13]) ? 16'b0000000111111111 : node786;
														assign node786 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node790 = (inp[3]) ? node796 : node791;
													assign node791 = (inp[13]) ? node793 : 16'b0000000111111111;
														assign node793 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node796 = (inp[12]) ? 16'b0000000011111111 : node797;
														assign node797 = (inp[13]) ? 16'b0000000011111111 : node798;
															assign node798 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node803 = (inp[5]) ? node931 : node804;
									assign node804 = (inp[7]) ? node870 : node805;
										assign node805 = (inp[2]) ? node839 : node806;
											assign node806 = (inp[12]) ? node824 : node807;
												assign node807 = (inp[14]) ? 16'b0000011111111111 : node808;
													assign node808 = (inp[3]) ? node816 : node809;
														assign node809 = (inp[13]) ? node813 : node810;
															assign node810 = (inp[1]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node813 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node816 = (inp[13]) ? node820 : node817;
															assign node817 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node820 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node824 = (inp[3]) ? node836 : node825;
													assign node825 = (inp[6]) ? node833 : node826;
														assign node826 = (inp[14]) ? node828 : 16'b0000111111111111;
															assign node828 = (inp[1]) ? 16'b0000011111111111 : node829;
																assign node829 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node833 = (inp[13]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node836 = (inp[6]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node839 = (inp[13]) ? node853 : node840;
												assign node840 = (inp[6]) ? node848 : node841;
													assign node841 = (inp[14]) ? node843 : 16'b0000011111111111;
														assign node843 = (inp[1]) ? 16'b0000011111111111 : node844;
															assign node844 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node848 = (inp[14]) ? node850 : 16'b0000011111111111;
														assign node850 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node853 = (inp[6]) ? node865 : node854;
													assign node854 = (inp[12]) ? node860 : node855;
														assign node855 = (inp[3]) ? 16'b0000001111111111 : node856;
															assign node856 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node860 = (inp[1]) ? 16'b0000000111111111 : node861;
															assign node861 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node865 = (inp[12]) ? node867 : 16'b0000000111111111;
														assign node867 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node870 = (inp[3]) ? node904 : node871;
											assign node871 = (inp[6]) ? node885 : node872;
												assign node872 = (inp[2]) ? node878 : node873;
													assign node873 = (inp[12]) ? 16'b0000111111111111 : node874;
														assign node874 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node878 = (inp[1]) ? 16'b0000001111111111 : node879;
														assign node879 = (inp[14]) ? 16'b0000001111111111 : node880;
															assign node880 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node885 = (inp[14]) ? node895 : node886;
													assign node886 = (inp[2]) ? 16'b0000000011111111 : node887;
														assign node887 = (inp[12]) ? 16'b0000001111111111 : node888;
															assign node888 = (inp[1]) ? node890 : 16'b0000011111111111;
																assign node890 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node895 = (inp[13]) ? node901 : node896;
														assign node896 = (inp[12]) ? 16'b0000000111111111 : node897;
															assign node897 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node901 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node904 = (inp[6]) ? node920 : node905;
												assign node905 = (inp[14]) ? node911 : node906;
													assign node906 = (inp[13]) ? node908 : 16'b0000001111111111;
														assign node908 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node911 = (inp[12]) ? node915 : node912;
														assign node912 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node915 = (inp[1]) ? 16'b0000000001111111 : node916;
															assign node916 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node920 = (inp[1]) ? node926 : node921;
													assign node921 = (inp[14]) ? node923 : 16'b0000000111111111;
														assign node923 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node926 = (inp[12]) ? 16'b0000000011111111 : node927;
														assign node927 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node931 = (inp[13]) ? node1011 : node932;
										assign node932 = (inp[7]) ? node960 : node933;
											assign node933 = (inp[12]) ? node951 : node934;
												assign node934 = (inp[6]) ? node938 : node935;
													assign node935 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node938 = (inp[1]) ? node944 : node939;
														assign node939 = (inp[14]) ? 16'b0000001111111111 : node940;
															assign node940 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node944 = (inp[3]) ? 16'b0000000111111111 : node945;
															assign node945 = (inp[14]) ? node947 : 16'b0000001111111111;
																assign node947 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node951 = (inp[3]) ? node957 : node952;
													assign node952 = (inp[6]) ? node954 : 16'b0000001111111111;
														assign node954 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node957 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node960 = (inp[14]) ? node982 : node961;
												assign node961 = (inp[1]) ? node975 : node962;
													assign node962 = (inp[6]) ? node970 : node963;
														assign node963 = (inp[12]) ? 16'b0000001111111111 : node964;
															assign node964 = (inp[3]) ? node966 : 16'b0000011111111111;
																assign node966 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node970 = (inp[3]) ? node972 : 16'b0000001111111111;
															assign node972 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node975 = (inp[3]) ? node979 : node976;
														assign node976 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node979 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node982 = (inp[2]) ? node1004 : node983;
													assign node983 = (inp[6]) ? node993 : node984;
														assign node984 = (inp[12]) ? node988 : node985;
															assign node985 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node988 = (inp[1]) ? node990 : 16'b0000000111111111;
																assign node990 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node993 = (inp[1]) ? node999 : node994;
															assign node994 = (inp[12]) ? node996 : 16'b0000000111111111;
																assign node996 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node999 = (inp[3]) ? node1001 : 16'b0000000011111111;
																assign node1001 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1004 = (inp[12]) ? node1008 : node1005;
														assign node1005 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1008 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1011 = (inp[6]) ? node1047 : node1012;
											assign node1012 = (inp[2]) ? node1032 : node1013;
												assign node1013 = (inp[14]) ? node1029 : node1014;
													assign node1014 = (inp[12]) ? node1018 : node1015;
														assign node1015 = (inp[3]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node1018 = (inp[7]) ? node1024 : node1019;
															assign node1019 = (inp[3]) ? node1021 : 16'b0000001111111111;
																assign node1021 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node1024 = (inp[3]) ? 16'b0000000111111111 : node1025;
																assign node1025 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1029 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1032 = (inp[3]) ? node1042 : node1033;
													assign node1033 = (inp[7]) ? node1037 : node1034;
														assign node1034 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1037 = (inp[1]) ? 16'b0000000011111111 : node1038;
															assign node1038 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1042 = (inp[7]) ? node1044 : 16'b0000000011111111;
														assign node1044 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1047 = (inp[3]) ? node1063 : node1048;
												assign node1048 = (inp[1]) ? node1054 : node1049;
													assign node1049 = (inp[12]) ? 16'b0000000111111111 : node1050;
														assign node1050 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1054 = (inp[12]) ? node1056 : 16'b0000000111111111;
														assign node1056 = (inp[2]) ? node1058 : 16'b0000000011111111;
															assign node1058 = (inp[14]) ? node1060 : 16'b0000000001111111;
																assign node1060 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1063 = (inp[14]) ? node1071 : node1064;
													assign node1064 = (inp[2]) ? node1066 : 16'b0000000011111111;
														assign node1066 = (inp[12]) ? 16'b0000000001111111 : node1067;
															assign node1067 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1071 = (inp[7]) ? node1073 : 16'b0000000001111111;
														assign node1073 = (inp[12]) ? node1075 : 16'b0000000001111111;
															assign node1075 = (inp[1]) ? node1077 : 16'b0000000000111111;
																assign node1077 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1080 = (inp[5]) ? node1606 : node1081;
							assign node1081 = (inp[13]) ? node1347 : node1082;
								assign node1082 = (inp[12]) ? node1228 : node1083;
									assign node1083 = (inp[6]) ? node1159 : node1084;
										assign node1084 = (inp[2]) ? node1120 : node1085;
											assign node1085 = (inp[1]) ? node1107 : node1086;
												assign node1086 = (inp[15]) ? node1096 : node1087;
													assign node1087 = (inp[3]) ? node1093 : node1088;
														assign node1088 = (inp[7]) ? 16'b0011111111111111 : node1089;
															assign node1089 = (inp[14]) ? 16'b0011111111111111 : 16'b0111111111111111;
														assign node1093 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1096 = (inp[3]) ? node1102 : node1097;
														assign node1097 = (inp[8]) ? node1099 : 16'b0001111111111111;
															assign node1099 = (inp[14]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node1102 = (inp[7]) ? node1104 : 16'b0000111111111111;
															assign node1104 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1107 = (inp[15]) ? node1115 : node1108;
													assign node1108 = (inp[3]) ? node1112 : node1109;
														assign node1109 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1112 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1115 = (inp[8]) ? node1117 : 16'b0000011111111111;
														assign node1117 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node1120 = (inp[7]) ? node1142 : node1121;
												assign node1121 = (inp[8]) ? node1129 : node1122;
													assign node1122 = (inp[1]) ? node1126 : node1123;
														assign node1123 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1126 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1129 = (inp[15]) ? node1135 : node1130;
														assign node1130 = (inp[14]) ? 16'b0000011111111111 : node1131;
															assign node1131 = (inp[1]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node1135 = (inp[1]) ? 16'b0000001111111111 : node1136;
															assign node1136 = (inp[14]) ? node1138 : 16'b0000011111111111;
																assign node1138 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1142 = (inp[1]) ? node1154 : node1143;
													assign node1143 = (inp[8]) ? node1145 : 16'b0000011111111111;
														assign node1145 = (inp[14]) ? 16'b0000001111111111 : node1146;
															assign node1146 = (inp[3]) ? node1150 : node1147;
																assign node1147 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
																assign node1150 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1154 = (inp[15]) ? 16'b0000000111111111 : node1155;
														assign node1155 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1159 = (inp[2]) ? node1197 : node1160;
											assign node1160 = (inp[1]) ? node1178 : node1161;
												assign node1161 = (inp[8]) ? node1175 : node1162;
													assign node1162 = (inp[7]) ? node1168 : node1163;
														assign node1163 = (inp[15]) ? 16'b0000111111111111 : node1164;
															assign node1164 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1168 = (inp[15]) ? 16'b0000011111111111 : node1169;
															assign node1169 = (inp[3]) ? node1171 : 16'b0000111111111111;
																assign node1171 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1175 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1178 = (inp[3]) ? node1188 : node1179;
													assign node1179 = (inp[15]) ? 16'b0000001111111111 : node1180;
														assign node1180 = (inp[14]) ? 16'b0000011111111111 : node1181;
															assign node1181 = (inp[7]) ? node1183 : 16'b0000111111111111;
																assign node1183 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1188 = (inp[7]) ? node1192 : node1189;
														assign node1189 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1192 = (inp[8]) ? node1194 : 16'b0000001111111111;
															assign node1194 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1197 = (inp[14]) ? node1217 : node1198;
												assign node1198 = (inp[1]) ? node1210 : node1199;
													assign node1199 = (inp[15]) ? node1203 : node1200;
														assign node1200 = (inp[3]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node1203 = (inp[3]) ? 16'b0000001111111111 : node1204;
															assign node1204 = (inp[8]) ? node1206 : 16'b0000011111111111;
																assign node1206 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1210 = (inp[15]) ? node1214 : node1211;
														assign node1211 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1214 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1217 = (inp[1]) ? node1225 : node1218;
													assign node1218 = (inp[3]) ? node1222 : node1219;
														assign node1219 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1222 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1225 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1228 = (inp[8]) ? node1274 : node1229;
										assign node1229 = (inp[14]) ? node1255 : node1230;
											assign node1230 = (inp[2]) ? node1246 : node1231;
												assign node1231 = (inp[6]) ? node1241 : node1232;
													assign node1232 = (inp[15]) ? 16'b0000111111111111 : node1233;
														assign node1233 = (inp[1]) ? node1235 : 16'b0001111111111111;
															assign node1235 = (inp[7]) ? 16'b0000111111111111 : node1236;
																assign node1236 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1241 = (inp[3]) ? 16'b0000011111111111 : node1242;
														assign node1242 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1246 = (inp[15]) ? node1252 : node1247;
													assign node1247 = (inp[3]) ? node1249 : 16'b0001111111111111;
														assign node1249 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1252 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1255 = (inp[6]) ? node1269 : node1256;
												assign node1256 = (inp[15]) ? node1264 : node1257;
													assign node1257 = (inp[7]) ? node1259 : 16'b0000011111111111;
														assign node1259 = (inp[2]) ? 16'b0000001111111111 : node1260;
															assign node1260 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1264 = (inp[2]) ? node1266 : 16'b0000001111111111;
														assign node1266 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1269 = (inp[2]) ? node1271 : 16'b0000001111111111;
													assign node1271 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1274 = (inp[7]) ? node1304 : node1275;
											assign node1275 = (inp[3]) ? node1291 : node1276;
												assign node1276 = (inp[15]) ? node1286 : node1277;
													assign node1277 = (inp[2]) ? node1281 : node1278;
														assign node1278 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1281 = (inp[14]) ? node1283 : 16'b0000011111111111;
															assign node1283 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1286 = (inp[6]) ? 16'b0000000111111111 : node1287;
														assign node1287 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1291 = (inp[2]) ? node1299 : node1292;
													assign node1292 = (inp[1]) ? node1294 : 16'b0000001111111111;
														assign node1294 = (inp[14]) ? node1296 : 16'b0000001111111111;
															assign node1296 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1299 = (inp[14]) ? 16'b0000000011111111 : node1300;
														assign node1300 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1304 = (inp[1]) ? node1324 : node1305;
												assign node1305 = (inp[6]) ? node1315 : node1306;
													assign node1306 = (inp[3]) ? node1312 : node1307;
														assign node1307 = (inp[14]) ? 16'b0000001111111111 : node1308;
															assign node1308 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1312 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1315 = (inp[15]) ? 16'b0000000111111111 : node1316;
														assign node1316 = (inp[14]) ? node1318 : 16'b0000001111111111;
															assign node1318 = (inp[2]) ? 16'b0000000111111111 : node1319;
																assign node1319 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1324 = (inp[2]) ? node1336 : node1325;
													assign node1325 = (inp[6]) ? node1333 : node1326;
														assign node1326 = (inp[14]) ? 16'b0000000111111111 : node1327;
															assign node1327 = (inp[3]) ? node1329 : 16'b0000001111111111;
																assign node1329 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1333 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1336 = (inp[15]) ? node1342 : node1337;
														assign node1337 = (inp[6]) ? 16'b0000000011111111 : node1338;
															assign node1338 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1342 = (inp[3]) ? node1344 : 16'b0000000011111111;
															assign node1344 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1347 = (inp[3]) ? node1453 : node1348;
									assign node1348 = (inp[8]) ? node1398 : node1349;
										assign node1349 = (inp[6]) ? node1367 : node1350;
											assign node1350 = (inp[2]) ? node1360 : node1351;
												assign node1351 = (inp[7]) ? node1353 : 16'b0000111111111111;
													assign node1353 = (inp[14]) ? node1357 : node1354;
														assign node1354 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1357 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1360 = (inp[1]) ? node1362 : 16'b0000011111111111;
													assign node1362 = (inp[14]) ? 16'b0000001111111111 : node1363;
														assign node1363 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1367 = (inp[14]) ? node1377 : node1368;
												assign node1368 = (inp[15]) ? node1370 : 16'b0000011111111111;
													assign node1370 = (inp[7]) ? node1372 : 16'b0000011111111111;
														assign node1372 = (inp[12]) ? 16'b0000001111111111 : node1373;
															assign node1373 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1377 = (inp[1]) ? node1391 : node1378;
													assign node1378 = (inp[2]) ? 16'b0000001111111111 : node1379;
														assign node1379 = (inp[7]) ? node1385 : node1380;
															assign node1380 = (inp[15]) ? 16'b0000011111111111 : node1381;
																assign node1381 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node1385 = (inp[15]) ? 16'b0000001111111111 : node1386;
																assign node1386 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1391 = (inp[12]) ? 16'b0000001111111111 : node1392;
														assign node1392 = (inp[2]) ? 16'b0000000111111111 : node1393;
															assign node1393 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1398 = (inp[1]) ? node1426 : node1399;
											assign node1399 = (inp[15]) ? node1413 : node1400;
												assign node1400 = (inp[6]) ? node1410 : node1401;
													assign node1401 = (inp[2]) ? 16'b0000011111111111 : node1402;
														assign node1402 = (inp[14]) ? 16'b0000011111111111 : node1403;
															assign node1403 = (inp[12]) ? 16'b0000111111111111 : node1404;
																assign node1404 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1410 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1413 = (inp[7]) ? node1421 : node1414;
													assign node1414 = (inp[2]) ? node1416 : 16'b0000011111111111;
														assign node1416 = (inp[6]) ? node1418 : 16'b0000001111111111;
															assign node1418 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1421 = (inp[2]) ? 16'b0000000111111111 : node1422;
														assign node1422 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1426 = (inp[15]) ? node1448 : node1427;
												assign node1427 = (inp[6]) ? node1441 : node1428;
													assign node1428 = (inp[14]) ? node1432 : node1429;
														assign node1429 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node1432 = (inp[12]) ? node1438 : node1433;
															assign node1433 = (inp[2]) ? node1435 : 16'b0000001111111111;
																assign node1435 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node1438 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1441 = (inp[12]) ? 16'b0000000111111111 : node1442;
														assign node1442 = (inp[7]) ? node1444 : 16'b0000000111111111;
															assign node1444 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1448 = (inp[14]) ? node1450 : 16'b0000000111111111;
													assign node1450 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node1453 = (inp[15]) ? node1531 : node1454;
										assign node1454 = (inp[7]) ? node1490 : node1455;
											assign node1455 = (inp[8]) ? node1483 : node1456;
												assign node1456 = (inp[14]) ? node1472 : node1457;
													assign node1457 = (inp[6]) ? node1465 : node1458;
														assign node1458 = (inp[12]) ? 16'b0000011111111111 : node1459;
															assign node1459 = (inp[2]) ? node1461 : 16'b0000111111111111;
																assign node1461 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1465 = (inp[12]) ? 16'b0000001111111111 : node1466;
															assign node1466 = (inp[2]) ? node1468 : 16'b0000011111111111;
																assign node1468 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1472 = (inp[2]) ? node1474 : 16'b0000011111111111;
														assign node1474 = (inp[1]) ? node1478 : node1475;
															assign node1475 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node1478 = (inp[12]) ? 16'b0000000111111111 : node1479;
																assign node1479 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1483 = (inp[1]) ? node1485 : 16'b0000001111111111;
													assign node1485 = (inp[14]) ? node1487 : 16'b0000001111111111;
														assign node1487 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1490 = (inp[6]) ? node1510 : node1491;
												assign node1491 = (inp[12]) ? node1501 : node1492;
													assign node1492 = (inp[8]) ? 16'b0000001111111111 : node1493;
														assign node1493 = (inp[1]) ? node1495 : 16'b0000011111111111;
															assign node1495 = (inp[2]) ? 16'b0000001111111111 : node1496;
																assign node1496 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1501 = (inp[2]) ? node1505 : node1502;
														assign node1502 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1505 = (inp[8]) ? node1507 : 16'b0000000111111111;
															assign node1507 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1510 = (inp[1]) ? node1522 : node1511;
													assign node1511 = (inp[8]) ? node1517 : node1512;
														assign node1512 = (inp[2]) ? 16'b0000000111111111 : node1513;
															assign node1513 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1517 = (inp[2]) ? node1519 : 16'b0000000111111111;
															assign node1519 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1522 = (inp[14]) ? node1526 : node1523;
														assign node1523 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1526 = (inp[2]) ? node1528 : 16'b0000000011111111;
															assign node1528 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1531 = (inp[2]) ? node1567 : node1532;
											assign node1532 = (inp[14]) ? node1548 : node1533;
												assign node1533 = (inp[7]) ? node1539 : node1534;
													assign node1534 = (inp[8]) ? 16'b0000000111111111 : node1535;
														assign node1535 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1539 = (inp[6]) ? node1545 : node1540;
														assign node1540 = (inp[8]) ? 16'b0000000111111111 : node1541;
															assign node1541 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1545 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1548 = (inp[6]) ? node1556 : node1549;
													assign node1549 = (inp[8]) ? node1553 : node1550;
														assign node1550 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1553 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1556 = (inp[7]) ? node1560 : node1557;
														assign node1557 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1560 = (inp[8]) ? 16'b0000000001111111 : node1561;
															assign node1561 = (inp[12]) ? node1563 : 16'b0000000011111111;
																assign node1563 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1567 = (inp[6]) ? node1585 : node1568;
												assign node1568 = (inp[1]) ? node1578 : node1569;
													assign node1569 = (inp[8]) ? node1575 : node1570;
														assign node1570 = (inp[14]) ? node1572 : 16'b0000001111111111;
															assign node1572 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1575 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1578 = (inp[12]) ? node1582 : node1579;
														assign node1579 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1582 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1585 = (inp[14]) ? node1595 : node1586;
													assign node1586 = (inp[12]) ? 16'b0000000001111111 : node1587;
														assign node1587 = (inp[7]) ? node1589 : 16'b0000000111111111;
															assign node1589 = (inp[1]) ? node1591 : 16'b0000000011111111;
																assign node1591 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1595 = (inp[8]) ? node1599 : node1596;
														assign node1596 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1599 = (inp[12]) ? node1603 : node1600;
															assign node1600 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node1603 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1606 = (inp[14]) ? node1876 : node1607;
								assign node1607 = (inp[13]) ? node1737 : node1608;
									assign node1608 = (inp[7]) ? node1670 : node1609;
										assign node1609 = (inp[1]) ? node1635 : node1610;
											assign node1610 = (inp[3]) ? node1632 : node1611;
												assign node1611 = (inp[2]) ? node1621 : node1612;
													assign node1612 = (inp[6]) ? node1616 : node1613;
														assign node1613 = (inp[8]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node1616 = (inp[8]) ? 16'b0000111111111111 : node1617;
															assign node1617 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1621 = (inp[12]) ? node1627 : node1622;
														assign node1622 = (inp[15]) ? 16'b0000011111111111 : node1623;
															assign node1623 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1627 = (inp[6]) ? 16'b0000001111111111 : node1628;
															assign node1628 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1632 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1635 = (inp[6]) ? node1655 : node1636;
												assign node1636 = (inp[3]) ? node1644 : node1637;
													assign node1637 = (inp[2]) ? node1641 : node1638;
														assign node1638 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1641 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1644 = (inp[2]) ? node1650 : node1645;
														assign node1645 = (inp[15]) ? 16'b0000001111111111 : node1646;
															assign node1646 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node1650 = (inp[15]) ? node1652 : 16'b0000001111111111;
															assign node1652 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1655 = (inp[8]) ? node1661 : node1656;
													assign node1656 = (inp[3]) ? 16'b0000000111111111 : node1657;
														assign node1657 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1661 = (inp[12]) ? node1665 : node1662;
														assign node1662 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1665 = (inp[15]) ? node1667 : 16'b0000000111111111;
															assign node1667 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1670 = (inp[8]) ? node1706 : node1671;
											assign node1671 = (inp[1]) ? node1699 : node1672;
												assign node1672 = (inp[2]) ? node1684 : node1673;
													assign node1673 = (inp[15]) ? node1681 : node1674;
														assign node1674 = (inp[3]) ? 16'b0000011111111111 : node1675;
															assign node1675 = (inp[6]) ? node1677 : 16'b0000111111111111;
																assign node1677 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1681 = (inp[6]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node1684 = (inp[15]) ? node1692 : node1685;
														assign node1685 = (inp[6]) ? 16'b0000001111111111 : node1686;
															assign node1686 = (inp[12]) ? node1688 : 16'b0000011111111111;
																assign node1688 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1692 = (inp[6]) ? 16'b0000000111111111 : node1693;
															assign node1693 = (inp[12]) ? node1695 : 16'b0000001111111111;
																assign node1695 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1699 = (inp[6]) ? 16'b0000000111111111 : node1700;
													assign node1700 = (inp[2]) ? node1702 : 16'b0000001111111111;
														assign node1702 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1706 = (inp[6]) ? node1724 : node1707;
												assign node1707 = (inp[1]) ? node1715 : node1708;
													assign node1708 = (inp[3]) ? node1710 : 16'b0000001111111111;
														assign node1710 = (inp[15]) ? node1712 : 16'b0000001111111111;
															assign node1712 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1715 = (inp[3]) ? node1721 : node1716;
														assign node1716 = (inp[15]) ? 16'b0000000111111111 : node1717;
															assign node1717 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1721 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1724 = (inp[15]) ? node1732 : node1725;
													assign node1725 = (inp[3]) ? node1727 : 16'b0000001111111111;
														assign node1727 = (inp[12]) ? node1729 : 16'b0000000111111111;
															assign node1729 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1732 = (inp[12]) ? 16'b0000000001111111 : node1733;
														assign node1733 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1737 = (inp[8]) ? node1801 : node1738;
										assign node1738 = (inp[2]) ? node1768 : node1739;
											assign node1739 = (inp[6]) ? node1755 : node1740;
												assign node1740 = (inp[1]) ? node1746 : node1741;
													assign node1741 = (inp[3]) ? 16'b0000011111111111 : node1742;
														assign node1742 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1746 = (inp[3]) ? node1752 : node1747;
														assign node1747 = (inp[12]) ? node1749 : 16'b0000011111111111;
															assign node1749 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1752 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1755 = (inp[15]) ? node1765 : node1756;
													assign node1756 = (inp[3]) ? node1760 : node1757;
														assign node1757 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1760 = (inp[12]) ? 16'b0000000111111111 : node1761;
															assign node1761 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1765 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1768 = (inp[15]) ? node1782 : node1769;
												assign node1769 = (inp[12]) ? node1775 : node1770;
													assign node1770 = (inp[1]) ? 16'b0000001111111111 : node1771;
														assign node1771 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1775 = (inp[6]) ? 16'b0000000011111111 : node1776;
														assign node1776 = (inp[7]) ? 16'b0000000111111111 : node1777;
															assign node1777 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node1782 = (inp[1]) ? node1796 : node1783;
													assign node1783 = (inp[3]) ? node1791 : node1784;
														assign node1784 = (inp[12]) ? 16'b0000000111111111 : node1785;
															assign node1785 = (inp[7]) ? node1787 : 16'b0000001111111111;
																assign node1787 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1791 = (inp[12]) ? node1793 : 16'b0000000111111111;
															assign node1793 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1796 = (inp[7]) ? node1798 : 16'b0000000111111111;
														assign node1798 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1801 = (inp[7]) ? node1827 : node1802;
											assign node1802 = (inp[15]) ? node1812 : node1803;
												assign node1803 = (inp[2]) ? 16'b0000000111111111 : node1804;
													assign node1804 = (inp[1]) ? node1808 : node1805;
														assign node1805 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1808 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1812 = (inp[3]) ? node1822 : node1813;
													assign node1813 = (inp[1]) ? node1815 : 16'b0000001111111111;
														assign node1815 = (inp[2]) ? node1817 : 16'b0000000111111111;
															assign node1817 = (inp[6]) ? 16'b0000000011111111 : node1818;
																assign node1818 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1822 = (inp[2]) ? 16'b0000000011111111 : node1823;
														assign node1823 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node1827 = (inp[12]) ? node1857 : node1828;
												assign node1828 = (inp[3]) ? node1842 : node1829;
													assign node1829 = (inp[15]) ? node1839 : node1830;
														assign node1830 = (inp[6]) ? node1834 : node1831;
															assign node1831 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node1834 = (inp[1]) ? 16'b0000000111111111 : node1835;
																assign node1835 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1839 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1842 = (inp[1]) ? node1850 : node1843;
														assign node1843 = (inp[15]) ? node1845 : 16'b0000000111111111;
															assign node1845 = (inp[2]) ? 16'b0000000011111111 : node1846;
																assign node1846 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1850 = (inp[15]) ? 16'b0000000000111111 : node1851;
															assign node1851 = (inp[6]) ? node1853 : 16'b0000000011111111;
																assign node1853 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1857 = (inp[1]) ? node1869 : node1858;
													assign node1858 = (inp[15]) ? node1862 : node1859;
														assign node1859 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1862 = (inp[2]) ? 16'b0000000000111111 : node1863;
															assign node1863 = (inp[3]) ? node1865 : 16'b0000000011111111;
																assign node1865 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1869 = (inp[2]) ? 16'b0000000001111111 : node1870;
														assign node1870 = (inp[15]) ? 16'b0000000001111111 : node1871;
															assign node1871 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1876 = (inp[1]) ? node1970 : node1877;
									assign node1877 = (inp[13]) ? node1921 : node1878;
										assign node1878 = (inp[12]) ? node1890 : node1879;
											assign node1879 = (inp[2]) ? node1883 : node1880;
												assign node1880 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1883 = (inp[15]) ? node1885 : 16'b0000001111111111;
													assign node1885 = (inp[3]) ? node1887 : 16'b0000001111111111;
														assign node1887 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1890 = (inp[7]) ? node1906 : node1891;
												assign node1891 = (inp[6]) ? node1901 : node1892;
													assign node1892 = (inp[2]) ? node1898 : node1893;
														assign node1893 = (inp[15]) ? 16'b0000001111111111 : node1894;
															assign node1894 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1898 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1901 = (inp[2]) ? 16'b0000000111111111 : node1902;
														assign node1902 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1906 = (inp[15]) ? node1914 : node1907;
													assign node1907 = (inp[2]) ? node1911 : node1908;
														assign node1908 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1911 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1914 = (inp[6]) ? node1918 : node1915;
														assign node1915 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1918 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1921 = (inp[3]) ? node1949 : node1922;
											assign node1922 = (inp[6]) ? node1932 : node1923;
												assign node1923 = (inp[12]) ? node1927 : node1924;
													assign node1924 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1927 = (inp[8]) ? 16'b0000000111111111 : node1928;
														assign node1928 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1932 = (inp[2]) ? node1940 : node1933;
													assign node1933 = (inp[8]) ? node1937 : node1934;
														assign node1934 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1937 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1940 = (inp[7]) ? 16'b0000000011111111 : node1941;
														assign node1941 = (inp[8]) ? node1943 : 16'b0000000111111111;
															assign node1943 = (inp[15]) ? 16'b0000000011111111 : node1944;
																assign node1944 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1949 = (inp[6]) ? node1961 : node1950;
												assign node1950 = (inp[15]) ? node1956 : node1951;
													assign node1951 = (inp[7]) ? node1953 : 16'b0000000111111111;
														assign node1953 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1956 = (inp[12]) ? node1958 : 16'b0000000011111111;
														assign node1958 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1961 = (inp[12]) ? node1967 : node1962;
													assign node1962 = (inp[2]) ? node1964 : 16'b0000000011111111;
														assign node1964 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1967 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1970 = (inp[8]) ? node2040 : node1971;
										assign node1971 = (inp[6]) ? node2007 : node1972;
											assign node1972 = (inp[15]) ? node1990 : node1973;
												assign node1973 = (inp[13]) ? node1979 : node1974;
													assign node1974 = (inp[2]) ? node1976 : 16'b0000011111111111;
														assign node1976 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1979 = (inp[3]) ? node1983 : node1980;
														assign node1980 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1983 = (inp[12]) ? node1985 : 16'b0000000111111111;
															assign node1985 = (inp[7]) ? 16'b0000000011111111 : node1986;
																assign node1986 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1990 = (inp[13]) ? node1996 : node1991;
													assign node1991 = (inp[2]) ? node1993 : 16'b0000000111111111;
														assign node1993 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1996 = (inp[2]) ? node2000 : node1997;
														assign node1997 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2000 = (inp[3]) ? node2004 : node2001;
															assign node2001 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node2004 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2007 = (inp[13]) ? node2025 : node2008;
												assign node2008 = (inp[3]) ? node2018 : node2009;
													assign node2009 = (inp[15]) ? node2013 : node2010;
														assign node2010 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2013 = (inp[2]) ? 16'b0000000011111111 : node2014;
															assign node2014 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2018 = (inp[7]) ? node2020 : 16'b0000000011111111;
														assign node2020 = (inp[2]) ? node2022 : 16'b0000000011111111;
															assign node2022 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2025 = (inp[12]) ? node2033 : node2026;
													assign node2026 = (inp[7]) ? node2028 : 16'b0000000011111111;
														assign node2028 = (inp[2]) ? node2030 : 16'b0000000011111111;
															assign node2030 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2033 = (inp[2]) ? 16'b0000000001111111 : node2034;
														assign node2034 = (inp[15]) ? node2036 : 16'b0000000011111111;
															assign node2036 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2040 = (inp[2]) ? node2060 : node2041;
											assign node2041 = (inp[6]) ? node2049 : node2042;
												assign node2042 = (inp[7]) ? node2046 : node2043;
													assign node2043 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node2046 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node2049 = (inp[7]) ? 16'b0000000000111111 : node2050;
													assign node2050 = (inp[3]) ? node2056 : node2051;
														assign node2051 = (inp[12]) ? 16'b0000000011111111 : node2052;
															assign node2052 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2056 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2060 = (inp[12]) ? node2072 : node2061;
												assign node2061 = (inp[7]) ? node2063 : 16'b0000000011111111;
													assign node2063 = (inp[3]) ? node2069 : node2064;
														assign node2064 = (inp[13]) ? 16'b0000000001111111 : node2065;
															assign node2065 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2069 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node2072 = (inp[7]) ? node2080 : node2073;
													assign node2073 = (inp[13]) ? node2075 : 16'b0000000001111111;
														assign node2075 = (inp[3]) ? 16'b0000000000111111 : node2076;
															assign node2076 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2080 = (inp[15]) ? node2084 : node2081;
														assign node2081 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node2084 = (inp[13]) ? node2088 : node2085;
															assign node2085 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
															assign node2088 = (inp[6]) ? node2090 : 16'b0000000000011111;
																assign node2090 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node2093 = (inp[1]) ? node3161 : node2094;
						assign node2094 = (inp[14]) ? node2638 : node2095;
							assign node2095 = (inp[12]) ? node2383 : node2096;
								assign node2096 = (inp[2]) ? node2248 : node2097;
									assign node2097 = (inp[8]) ? node2165 : node2098;
										assign node2098 = (inp[15]) ? node2138 : node2099;
											assign node2099 = (inp[6]) ? node2111 : node2100;
												assign node2100 = (inp[13]) ? node2106 : node2101;
													assign node2101 = (inp[3]) ? 16'b0001111111111111 : node2102;
														assign node2102 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node2106 = (inp[5]) ? 16'b0000111111111111 : node2107;
														assign node2107 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node2111 = (inp[9]) ? node2123 : node2112;
													assign node2112 = (inp[7]) ? node2120 : node2113;
														assign node2113 = (inp[13]) ? node2115 : 16'b0001111111111111;
															assign node2115 = (inp[5]) ? 16'b0000111111111111 : node2116;
																assign node2116 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2120 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2123 = (inp[13]) ? node2131 : node2124;
														assign node2124 = (inp[5]) ? node2126 : 16'b0001111111111111;
															assign node2126 = (inp[7]) ? 16'b0000011111111111 : node2127;
																assign node2127 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2131 = (inp[3]) ? 16'b0000001111111111 : node2132;
															assign node2132 = (inp[5]) ? node2134 : 16'b0000011111111111;
																assign node2134 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2138 = (inp[5]) ? node2152 : node2139;
												assign node2139 = (inp[7]) ? node2145 : node2140;
													assign node2140 = (inp[13]) ? node2142 : 16'b0000111111111111;
														assign node2142 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2145 = (inp[6]) ? 16'b0000001111111111 : node2146;
														assign node2146 = (inp[13]) ? 16'b0000011111111111 : node2147;
															assign node2147 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2152 = (inp[13]) ? node2160 : node2153;
													assign node2153 = (inp[9]) ? node2155 : 16'b0000111111111111;
														assign node2155 = (inp[3]) ? node2157 : 16'b0000011111111111;
															assign node2157 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2160 = (inp[3]) ? 16'b0000000111111111 : node2161;
														assign node2161 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node2165 = (inp[6]) ? node2203 : node2166;
											assign node2166 = (inp[7]) ? node2186 : node2167;
												assign node2167 = (inp[13]) ? node2177 : node2168;
													assign node2168 = (inp[3]) ? 16'b0000011111111111 : node2169;
														assign node2169 = (inp[15]) ? node2171 : 16'b0000111111111111;
															assign node2171 = (inp[9]) ? node2173 : 16'b0000111111111111;
																assign node2173 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2177 = (inp[9]) ? node2181 : node2178;
														assign node2178 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2181 = (inp[15]) ? node2183 : 16'b0000011111111111;
															assign node2183 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2186 = (inp[5]) ? node2198 : node2187;
													assign node2187 = (inp[13]) ? node2191 : node2188;
														assign node2188 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2191 = (inp[9]) ? node2193 : 16'b0000011111111111;
															assign node2193 = (inp[3]) ? 16'b0000001111111111 : node2194;
																assign node2194 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2198 = (inp[9]) ? 16'b0000001111111111 : node2199;
														assign node2199 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2203 = (inp[9]) ? node2233 : node2204;
												assign node2204 = (inp[3]) ? node2226 : node2205;
													assign node2205 = (inp[5]) ? node2217 : node2206;
														assign node2206 = (inp[13]) ? node2212 : node2207;
															assign node2207 = (inp[15]) ? node2209 : 16'b0000111111111111;
																assign node2209 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node2212 = (inp[15]) ? node2214 : 16'b0000011111111111;
																assign node2214 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2217 = (inp[15]) ? node2223 : node2218;
															assign node2218 = (inp[13]) ? node2220 : 16'b0000011111111111;
																assign node2220 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node2223 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2226 = (inp[7]) ? node2230 : node2227;
														assign node2227 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2230 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2233 = (inp[7]) ? node2241 : node2234;
													assign node2234 = (inp[15]) ? 16'b0000001111111111 : node2235;
														assign node2235 = (inp[13]) ? 16'b0000001111111111 : node2236;
															assign node2236 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2241 = (inp[3]) ? node2245 : node2242;
														assign node2242 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2245 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node2248 = (inp[9]) ? node2310 : node2249;
										assign node2249 = (inp[7]) ? node2279 : node2250;
											assign node2250 = (inp[15]) ? node2268 : node2251;
												assign node2251 = (inp[13]) ? node2257 : node2252;
													assign node2252 = (inp[6]) ? node2254 : 16'b0000111111111111;
														assign node2254 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2257 = (inp[8]) ? node2261 : node2258;
														assign node2258 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2261 = (inp[3]) ? node2263 : 16'b0000011111111111;
															assign node2263 = (inp[5]) ? 16'b0000001111111111 : node2264;
																assign node2264 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2268 = (inp[5]) ? node2274 : node2269;
													assign node2269 = (inp[13]) ? node2271 : 16'b0000011111111111;
														assign node2271 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2274 = (inp[6]) ? 16'b0000001111111111 : node2275;
														assign node2275 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2279 = (inp[3]) ? node2301 : node2280;
												assign node2280 = (inp[6]) ? node2294 : node2281;
													assign node2281 = (inp[5]) ? node2289 : node2282;
														assign node2282 = (inp[15]) ? node2284 : 16'b0001111111111111;
															assign node2284 = (inp[13]) ? 16'b0000011111111111 : node2285;
																assign node2285 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2289 = (inp[8]) ? node2291 : 16'b0000011111111111;
															assign node2291 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2294 = (inp[15]) ? node2298 : node2295;
														assign node2295 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2298 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2301 = (inp[13]) ? node2303 : 16'b0000001111111111;
													assign node2303 = (inp[15]) ? node2307 : node2304;
														assign node2304 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2307 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2310 = (inp[13]) ? node2350 : node2311;
											assign node2311 = (inp[5]) ? node2335 : node2312;
												assign node2312 = (inp[3]) ? node2324 : node2313;
													assign node2313 = (inp[15]) ? node2319 : node2314;
														assign node2314 = (inp[8]) ? 16'b0000011111111111 : node2315;
															assign node2315 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2319 = (inp[6]) ? node2321 : 16'b0000011111111111;
															assign node2321 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2324 = (inp[15]) ? 16'b0000000111111111 : node2325;
														assign node2325 = (inp[8]) ? 16'b0000001111111111 : node2326;
															assign node2326 = (inp[6]) ? node2330 : node2327;
																assign node2327 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
																assign node2330 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2335 = (inp[6]) ? node2345 : node2336;
													assign node2336 = (inp[8]) ? node2340 : node2337;
														assign node2337 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2340 = (inp[15]) ? node2342 : 16'b0000001111111111;
															assign node2342 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2345 = (inp[15]) ? node2347 : 16'b0000000111111111;
														assign node2347 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2350 = (inp[6]) ? node2368 : node2351;
												assign node2351 = (inp[3]) ? node2359 : node2352;
													assign node2352 = (inp[7]) ? node2354 : 16'b0000001111111111;
														assign node2354 = (inp[5]) ? node2356 : 16'b0000001111111111;
															assign node2356 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2359 = (inp[7]) ? node2365 : node2360;
														assign node2360 = (inp[15]) ? node2362 : 16'b0000001111111111;
															assign node2362 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node2365 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node2368 = (inp[8]) ? node2378 : node2369;
													assign node2369 = (inp[3]) ? node2375 : node2370;
														assign node2370 = (inp[5]) ? node2372 : 16'b0000001111111111;
															assign node2372 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2375 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2378 = (inp[5]) ? node2380 : 16'b0000000111111111;
														assign node2380 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2383 = (inp[7]) ? node2521 : node2384;
									assign node2384 = (inp[15]) ? node2456 : node2385;
										assign node2385 = (inp[3]) ? node2417 : node2386;
											assign node2386 = (inp[5]) ? node2404 : node2387;
												assign node2387 = (inp[13]) ? node2399 : node2388;
													assign node2388 = (inp[8]) ? node2394 : node2389;
														assign node2389 = (inp[9]) ? node2391 : 16'b0001111111111111;
															assign node2391 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2394 = (inp[6]) ? node2396 : 16'b0000111111111111;
															assign node2396 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2399 = (inp[8]) ? 16'b0000011111111111 : node2400;
														assign node2400 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2404 = (inp[8]) ? node2412 : node2405;
													assign node2405 = (inp[2]) ? node2409 : node2406;
														assign node2406 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2409 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2412 = (inp[6]) ? 16'b0000001111111111 : node2413;
														assign node2413 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2417 = (inp[9]) ? node2435 : node2418;
												assign node2418 = (inp[13]) ? node2424 : node2419;
													assign node2419 = (inp[2]) ? 16'b0000011111111111 : node2420;
														assign node2420 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2424 = (inp[5]) ? node2432 : node2425;
														assign node2425 = (inp[2]) ? node2427 : 16'b0000011111111111;
															assign node2427 = (inp[8]) ? 16'b0000001111111111 : node2428;
																assign node2428 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2432 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2435 = (inp[5]) ? node2451 : node2436;
													assign node2436 = (inp[6]) ? node2444 : node2437;
														assign node2437 = (inp[13]) ? node2439 : 16'b0000011111111111;
															assign node2439 = (inp[2]) ? node2441 : 16'b0000001111111111;
																assign node2441 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2444 = (inp[13]) ? 16'b0000000111111111 : node2445;
															assign node2445 = (inp[2]) ? node2447 : 16'b0000001111111111;
																assign node2447 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2451 = (inp[2]) ? 16'b0000000001111111 : node2452;
														assign node2452 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2456 = (inp[6]) ? node2488 : node2457;
											assign node2457 = (inp[5]) ? node2471 : node2458;
												assign node2458 = (inp[2]) ? node2468 : node2459;
													assign node2459 = (inp[13]) ? node2461 : 16'b0000011111111111;
														assign node2461 = (inp[9]) ? node2463 : 16'b0000011111111111;
															assign node2463 = (inp[8]) ? 16'b0000001111111111 : node2464;
																assign node2464 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2468 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2471 = (inp[9]) ? node2479 : node2472;
													assign node2472 = (inp[3]) ? 16'b0000000111111111 : node2473;
														assign node2473 = (inp[8]) ? 16'b0000001111111111 : node2474;
															assign node2474 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node2479 = (inp[13]) ? node2485 : node2480;
														assign node2480 = (inp[8]) ? node2482 : 16'b0000001111111111;
															assign node2482 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2485 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2488 = (inp[3]) ? node2500 : node2489;
												assign node2489 = (inp[5]) ? node2493 : node2490;
													assign node2490 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2493 = (inp[2]) ? node2497 : node2494;
														assign node2494 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2497 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2500 = (inp[8]) ? node2510 : node2501;
													assign node2501 = (inp[5]) ? node2503 : 16'b0000000111111111;
														assign node2503 = (inp[2]) ? node2505 : 16'b0000000111111111;
															assign node2505 = (inp[9]) ? 16'b0000000011111111 : node2506;
																assign node2506 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2510 = (inp[13]) ? node2512 : 16'b0000000111111111;
														assign node2512 = (inp[9]) ? node2516 : node2513;
															assign node2513 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node2516 = (inp[2]) ? node2518 : 16'b0000000001111111;
																assign node2518 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2521 = (inp[9]) ? node2571 : node2522;
										assign node2522 = (inp[3]) ? node2548 : node2523;
											assign node2523 = (inp[2]) ? node2539 : node2524;
												assign node2524 = (inp[8]) ? node2530 : node2525;
													assign node2525 = (inp[5]) ? node2527 : 16'b0000011111111111;
														assign node2527 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2530 = (inp[5]) ? node2534 : node2531;
														assign node2531 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2534 = (inp[6]) ? 16'b0000000111111111 : node2535;
															assign node2535 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2539 = (inp[15]) ? node2543 : node2540;
													assign node2540 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2543 = (inp[8]) ? 16'b0000000111111111 : node2544;
														assign node2544 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2548 = (inp[13]) ? node2562 : node2549;
												assign node2549 = (inp[2]) ? node2557 : node2550;
													assign node2550 = (inp[6]) ? 16'b0000001111111111 : node2551;
														assign node2551 = (inp[5]) ? node2553 : 16'b0000001111111111;
															assign node2553 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2557 = (inp[15]) ? 16'b0000000011111111 : node2558;
														assign node2558 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2562 = (inp[6]) ? node2564 : 16'b0000000111111111;
													assign node2564 = (inp[15]) ? node2568 : node2565;
														assign node2565 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2568 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2571 = (inp[8]) ? node2607 : node2572;
											assign node2572 = (inp[3]) ? node2586 : node2573;
												assign node2573 = (inp[5]) ? node2581 : node2574;
													assign node2574 = (inp[2]) ? node2578 : node2575;
														assign node2575 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2578 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2581 = (inp[13]) ? 16'b0000000011111111 : node2582;
														assign node2582 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2586 = (inp[15]) ? node2596 : node2587;
													assign node2587 = (inp[6]) ? node2593 : node2588;
														assign node2588 = (inp[13]) ? 16'b0000000111111111 : node2589;
															assign node2589 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2593 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2596 = (inp[13]) ? node2604 : node2597;
														assign node2597 = (inp[5]) ? 16'b0000000011111111 : node2598;
															assign node2598 = (inp[6]) ? node2600 : 16'b0000000111111111;
																assign node2600 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2604 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2607 = (inp[15]) ? node2623 : node2608;
												assign node2608 = (inp[6]) ? node2612 : node2609;
													assign node2609 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2612 = (inp[13]) ? node2618 : node2613;
														assign node2613 = (inp[3]) ? 16'b0000000011111111 : node2614;
															assign node2614 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2618 = (inp[3]) ? node2620 : 16'b0000000011111111;
															assign node2620 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2623 = (inp[6]) ? node2629 : node2624;
													assign node2624 = (inp[13]) ? 16'b0000000011111111 : node2625;
														assign node2625 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2629 = (inp[13]) ? node2631 : 16'b0000000001111111;
														assign node2631 = (inp[5]) ? node2635 : node2632;
															assign node2632 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node2635 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node2638 = (inp[9]) ? node2904 : node2639;
								assign node2639 = (inp[2]) ? node2759 : node2640;
									assign node2640 = (inp[5]) ? node2698 : node2641;
										assign node2641 = (inp[7]) ? node2671 : node2642;
											assign node2642 = (inp[13]) ? node2660 : node2643;
												assign node2643 = (inp[6]) ? node2655 : node2644;
													assign node2644 = (inp[15]) ? node2648 : node2645;
														assign node2645 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2648 = (inp[3]) ? node2652 : node2649;
															assign node2649 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node2652 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2655 = (inp[8]) ? node2657 : 16'b0000111111111111;
														assign node2657 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2660 = (inp[3]) ? node2664 : node2661;
													assign node2661 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2664 = (inp[8]) ? node2666 : 16'b0000011111111111;
														assign node2666 = (inp[15]) ? 16'b0000001111111111 : node2667;
															assign node2667 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2671 = (inp[13]) ? node2687 : node2672;
												assign node2672 = (inp[3]) ? node2682 : node2673;
													assign node2673 = (inp[6]) ? 16'b0000011111111111 : node2674;
														assign node2674 = (inp[8]) ? node2676 : 16'b0000111111111111;
															assign node2676 = (inp[12]) ? 16'b0000011111111111 : node2677;
																assign node2677 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2682 = (inp[15]) ? 16'b0000000111111111 : node2683;
														assign node2683 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2687 = (inp[15]) ? node2691 : node2688;
													assign node2688 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node2691 = (inp[8]) ? 16'b0000000111111111 : node2692;
														assign node2692 = (inp[3]) ? node2694 : 16'b0000000111111111;
															assign node2694 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2698 = (inp[15]) ? node2722 : node2699;
											assign node2699 = (inp[12]) ? node2711 : node2700;
												assign node2700 = (inp[8]) ? node2706 : node2701;
													assign node2701 = (inp[3]) ? node2703 : 16'b0000011111111111;
														assign node2703 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node2706 = (inp[6]) ? 16'b0000001111111111 : node2707;
														assign node2707 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2711 = (inp[8]) ? 16'b0000000111111111 : node2712;
													assign node2712 = (inp[6]) ? node2716 : node2713;
														assign node2713 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2716 = (inp[3]) ? node2718 : 16'b0000001111111111;
															assign node2718 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2722 = (inp[7]) ? node2740 : node2723;
												assign node2723 = (inp[13]) ? node2733 : node2724;
													assign node2724 = (inp[12]) ? node2730 : node2725;
														assign node2725 = (inp[3]) ? 16'b0000001111111111 : node2726;
															assign node2726 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2730 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2733 = (inp[8]) ? node2737 : node2734;
														assign node2734 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2737 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2740 = (inp[3]) ? node2752 : node2741;
													assign node2741 = (inp[12]) ? node2749 : node2742;
														assign node2742 = (inp[6]) ? 16'b0000000111111111 : node2743;
															assign node2743 = (inp[13]) ? node2745 : 16'b0000001111111111;
																assign node2745 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2749 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2752 = (inp[13]) ? node2754 : 16'b0000000011111111;
														assign node2754 = (inp[8]) ? node2756 : 16'b0000000011111111;
															assign node2756 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2759 = (inp[6]) ? node2839 : node2760;
										assign node2760 = (inp[13]) ? node2804 : node2761;
											assign node2761 = (inp[8]) ? node2787 : node2762;
												assign node2762 = (inp[12]) ? node2774 : node2763;
													assign node2763 = (inp[3]) ? node2769 : node2764;
														assign node2764 = (inp[15]) ? 16'b0000011111111111 : node2765;
															assign node2765 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2769 = (inp[7]) ? node2771 : 16'b0000011111111111;
															assign node2771 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node2774 = (inp[7]) ? node2782 : node2775;
														assign node2775 = (inp[5]) ? node2777 : 16'b0000001111111111;
															assign node2777 = (inp[15]) ? node2779 : 16'b0000001111111111;
																assign node2779 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2782 = (inp[5]) ? 16'b0000000111111111 : node2783;
															assign node2783 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2787 = (inp[3]) ? node2795 : node2788;
													assign node2788 = (inp[5]) ? node2792 : node2789;
														assign node2789 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2792 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2795 = (inp[5]) ? node2799 : node2796;
														assign node2796 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2799 = (inp[15]) ? node2801 : 16'b0000000111111111;
															assign node2801 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2804 = (inp[5]) ? node2832 : node2805;
												assign node2805 = (inp[12]) ? node2817 : node2806;
													assign node2806 = (inp[3]) ? node2812 : node2807;
														assign node2807 = (inp[8]) ? node2809 : 16'b0000011111111111;
															assign node2809 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2812 = (inp[7]) ? 16'b0000000111111111 : node2813;
															assign node2813 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2817 = (inp[7]) ? node2827 : node2818;
														assign node2818 = (inp[8]) ? node2824 : node2819;
															assign node2819 = (inp[15]) ? node2821 : 16'b0000001111111111;
																assign node2821 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node2824 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2827 = (inp[15]) ? 16'b0000000011111111 : node2828;
															assign node2828 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2832 = (inp[8]) ? 16'b0000000011111111 : node2833;
													assign node2833 = (inp[15]) ? node2835 : 16'b0000000111111111;
														assign node2835 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2839 = (inp[12]) ? node2875 : node2840;
											assign node2840 = (inp[7]) ? node2854 : node2841;
												assign node2841 = (inp[3]) ? node2849 : node2842;
													assign node2842 = (inp[8]) ? 16'b0000000111111111 : node2843;
														assign node2843 = (inp[13]) ? node2845 : 16'b0000011111111111;
															assign node2845 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2849 = (inp[13]) ? node2851 : 16'b0000000111111111;
														assign node2851 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2854 = (inp[8]) ? node2864 : node2855;
													assign node2855 = (inp[5]) ? node2859 : node2856;
														assign node2856 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node2859 = (inp[13]) ? node2861 : 16'b0000000111111111;
															assign node2861 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2864 = (inp[15]) ? node2872 : node2865;
														assign node2865 = (inp[13]) ? 16'b0000000011111111 : node2866;
															assign node2866 = (inp[3]) ? node2868 : 16'b0000000111111111;
																assign node2868 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2872 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node2875 = (inp[5]) ? node2887 : node2876;
												assign node2876 = (inp[3]) ? node2882 : node2877;
													assign node2877 = (inp[8]) ? node2879 : 16'b0000001111111111;
														assign node2879 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2882 = (inp[13]) ? 16'b0000000001111111 : node2883;
														assign node2883 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2887 = (inp[15]) ? node2897 : node2888;
													assign node2888 = (inp[8]) ? node2892 : node2889;
														assign node2889 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2892 = (inp[3]) ? node2894 : 16'b0000000011111111;
															assign node2894 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2897 = (inp[13]) ? node2901 : node2898;
														assign node2898 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2901 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2904 = (inp[8]) ? node3040 : node2905;
									assign node2905 = (inp[7]) ? node2975 : node2906;
										assign node2906 = (inp[13]) ? node2938 : node2907;
											assign node2907 = (inp[15]) ? node2915 : node2908;
												assign node2908 = (inp[12]) ? node2910 : 16'b0000011111111111;
													assign node2910 = (inp[2]) ? 16'b0000001111111111 : node2911;
														assign node2911 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2915 = (inp[3]) ? node2927 : node2916;
													assign node2916 = (inp[12]) ? node2924 : node2917;
														assign node2917 = (inp[6]) ? 16'b0000001111111111 : node2918;
															assign node2918 = (inp[5]) ? 16'b0000011111111111 : node2919;
																assign node2919 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2924 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2927 = (inp[2]) ? node2933 : node2928;
														assign node2928 = (inp[12]) ? node2930 : 16'b0000001111111111;
															assign node2930 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2933 = (inp[6]) ? node2935 : 16'b0000000011111111;
															assign node2935 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2938 = (inp[3]) ? node2958 : node2939;
												assign node2939 = (inp[15]) ? node2951 : node2940;
													assign node2940 = (inp[6]) ? node2942 : 16'b0000011111111111;
														assign node2942 = (inp[2]) ? node2946 : node2943;
															assign node2943 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node2946 = (inp[12]) ? 16'b0000000111111111 : node2947;
																assign node2947 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2951 = (inp[6]) ? node2955 : node2952;
														assign node2952 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2955 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2958 = (inp[6]) ? node2964 : node2959;
													assign node2959 = (inp[2]) ? 16'b0000000011111111 : node2960;
														assign node2960 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2964 = (inp[12]) ? node2968 : node2965;
														assign node2965 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2968 = (inp[2]) ? 16'b0000000001111111 : node2969;
															assign node2969 = (inp[5]) ? node2971 : 16'b0000000011111111;
																assign node2971 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2975 = (inp[13]) ? node3015 : node2976;
											assign node2976 = (inp[5]) ? node2996 : node2977;
												assign node2977 = (inp[15]) ? node2985 : node2978;
													assign node2978 = (inp[3]) ? node2980 : 16'b0000001111111111;
														assign node2980 = (inp[2]) ? 16'b0000000111111111 : node2981;
															assign node2981 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2985 = (inp[6]) ? node2989 : node2986;
														assign node2986 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2989 = (inp[3]) ? 16'b0000000011111111 : node2990;
															assign node2990 = (inp[12]) ? node2992 : 16'b0000000111111111;
																assign node2992 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2996 = (inp[12]) ? node3004 : node2997;
													assign node2997 = (inp[6]) ? 16'b0000000001111111 : node2998;
														assign node2998 = (inp[15]) ? 16'b0000000111111111 : node2999;
															assign node2999 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3004 = (inp[15]) ? node3012 : node3005;
														assign node3005 = (inp[2]) ? 16'b0000000011111111 : node3006;
															assign node3006 = (inp[6]) ? node3008 : 16'b0000000111111111;
																assign node3008 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3012 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3015 = (inp[15]) ? node3027 : node3016;
												assign node3016 = (inp[6]) ? node3022 : node3017;
													assign node3017 = (inp[12]) ? node3019 : 16'b0000001111111111;
														assign node3019 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3022 = (inp[3]) ? node3024 : 16'b0000000011111111;
														assign node3024 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3027 = (inp[6]) ? node3035 : node3028;
													assign node3028 = (inp[3]) ? node3030 : 16'b0000000011111111;
														assign node3030 = (inp[2]) ? 16'b0000000001111111 : node3031;
															assign node3031 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3035 = (inp[12]) ? 16'b0000000000111111 : node3036;
														assign node3036 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3040 = (inp[7]) ? node3112 : node3041;
										assign node3041 = (inp[3]) ? node3077 : node3042;
											assign node3042 = (inp[15]) ? node3062 : node3043;
												assign node3043 = (inp[5]) ? node3053 : node3044;
													assign node3044 = (inp[6]) ? node3050 : node3045;
														assign node3045 = (inp[13]) ? 16'b0000001111111111 : node3046;
															assign node3046 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3050 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3053 = (inp[12]) ? node3059 : node3054;
														assign node3054 = (inp[13]) ? 16'b0000000111111111 : node3055;
															assign node3055 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3059 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3062 = (inp[6]) ? node3064 : 16'b0000000111111111;
													assign node3064 = (inp[12]) ? node3074 : node3065;
														assign node3065 = (inp[13]) ? node3069 : node3066;
															assign node3066 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3069 = (inp[2]) ? 16'b0000000011111111 : node3070;
																assign node3070 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3074 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3077 = (inp[12]) ? node3097 : node3078;
												assign node3078 = (inp[2]) ? node3088 : node3079;
													assign node3079 = (inp[5]) ? node3081 : 16'b0000001111111111;
														assign node3081 = (inp[6]) ? node3083 : 16'b0000001111111111;
															assign node3083 = (inp[15]) ? 16'b0000000011111111 : node3084;
																assign node3084 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3088 = (inp[5]) ? node3090 : 16'b0000000011111111;
														assign node3090 = (inp[15]) ? 16'b0000000001111111 : node3091;
															assign node3091 = (inp[13]) ? 16'b0000000001111111 : node3092;
																assign node3092 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3097 = (inp[5]) ? node3105 : node3098;
													assign node3098 = (inp[2]) ? 16'b0000000001111111 : node3099;
														assign node3099 = (inp[15]) ? 16'b0000000011111111 : node3100;
															assign node3100 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3105 = (inp[6]) ? node3107 : 16'b0000000001111111;
														assign node3107 = (inp[15]) ? node3109 : 16'b0000000001111111;
															assign node3109 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node3112 = (inp[15]) ? node3132 : node3113;
											assign node3113 = (inp[3]) ? node3125 : node3114;
												assign node3114 = (inp[13]) ? node3118 : node3115;
													assign node3115 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3118 = (inp[2]) ? node3122 : node3119;
														assign node3119 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3122 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node3125 = (inp[12]) ? 16'b0000000001111111 : node3126;
													assign node3126 = (inp[5]) ? node3128 : 16'b0000000011111111;
														assign node3128 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3132 = (inp[2]) ? node3144 : node3133;
												assign node3133 = (inp[3]) ? 16'b0000000001111111 : node3134;
													assign node3134 = (inp[6]) ? node3136 : 16'b0000000011111111;
														assign node3136 = (inp[5]) ? node3138 : 16'b0000000011111111;
															assign node3138 = (inp[13]) ? 16'b0000000001111111 : node3139;
																assign node3139 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3144 = (inp[13]) ? node3154 : node3145;
													assign node3145 = (inp[6]) ? node3147 : 16'b0000000001111111;
														assign node3147 = (inp[5]) ? node3149 : 16'b0000000001111111;
															assign node3149 = (inp[12]) ? 16'b0000000000111111 : node3150;
																assign node3150 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3154 = (inp[3]) ? node3158 : node3155;
														assign node3155 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3158 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node3161 = (inp[8]) ? node3627 : node3162;
							assign node3162 = (inp[12]) ? node3384 : node3163;
								assign node3163 = (inp[15]) ? node3273 : node3164;
									assign node3164 = (inp[13]) ? node3234 : node3165;
										assign node3165 = (inp[5]) ? node3203 : node3166;
											assign node3166 = (inp[9]) ? node3184 : node3167;
												assign node3167 = (inp[14]) ? node3177 : node3168;
													assign node3168 = (inp[6]) ? node3172 : node3169;
														assign node3169 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3172 = (inp[2]) ? 16'b0000011111111111 : node3173;
															assign node3173 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3177 = (inp[7]) ? node3181 : node3178;
														assign node3178 = (inp[3]) ? 16'b0000111111111111 : 16'b0000011111111111;
														assign node3181 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3184 = (inp[2]) ? node3196 : node3185;
													assign node3185 = (inp[7]) ? node3189 : node3186;
														assign node3186 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3189 = (inp[14]) ? node3191 : 16'b0000011111111111;
															assign node3191 = (inp[3]) ? 16'b0000001111111111 : node3192;
																assign node3192 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3196 = (inp[7]) ? node3200 : node3197;
														assign node3197 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3200 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3203 = (inp[6]) ? node3217 : node3204;
												assign node3204 = (inp[2]) ? node3210 : node3205;
													assign node3205 = (inp[14]) ? node3207 : 16'b0000011111111111;
														assign node3207 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3210 = (inp[7]) ? node3214 : node3211;
														assign node3211 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3214 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3217 = (inp[2]) ? node3229 : node3218;
													assign node3218 = (inp[9]) ? node3224 : node3219;
														assign node3219 = (inp[7]) ? 16'b0000001111111111 : node3220;
															assign node3220 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3224 = (inp[14]) ? node3226 : 16'b0000001111111111;
															assign node3226 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3229 = (inp[9]) ? 16'b0000000111111111 : node3230;
														assign node3230 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3234 = (inp[7]) ? node3248 : node3235;
											assign node3235 = (inp[14]) ? node3245 : node3236;
												assign node3236 = (inp[5]) ? node3242 : node3237;
													assign node3237 = (inp[3]) ? node3239 : 16'b0000111111111111;
														assign node3239 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3242 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3245 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3248 = (inp[5]) ? node3262 : node3249;
												assign node3249 = (inp[2]) ? node3257 : node3250;
													assign node3250 = (inp[3]) ? node3254 : node3251;
														assign node3251 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3254 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3257 = (inp[3]) ? node3259 : 16'b0000000111111111;
														assign node3259 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3262 = (inp[6]) ? node3268 : node3263;
													assign node3263 = (inp[9]) ? node3265 : 16'b0000000111111111;
														assign node3265 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3268 = (inp[2]) ? node3270 : 16'b0000000011111111;
														assign node3270 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node3273 = (inp[3]) ? node3317 : node3274;
										assign node3274 = (inp[6]) ? node3296 : node3275;
											assign node3275 = (inp[9]) ? node3285 : node3276;
												assign node3276 = (inp[5]) ? node3280 : node3277;
													assign node3277 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3280 = (inp[2]) ? 16'b0000001111111111 : node3281;
														assign node3281 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3285 = (inp[14]) ? node3291 : node3286;
													assign node3286 = (inp[5]) ? 16'b0000001111111111 : node3287;
														assign node3287 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3291 = (inp[7]) ? node3293 : 16'b0000001111111111;
														assign node3293 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3296 = (inp[7]) ? node3308 : node3297;
												assign node3297 = (inp[5]) ? 16'b0000000111111111 : node3298;
													assign node3298 = (inp[9]) ? node3302 : node3299;
														assign node3299 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node3302 = (inp[14]) ? node3304 : 16'b0000001111111111;
															assign node3304 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3308 = (inp[5]) ? node3314 : node3309;
													assign node3309 = (inp[14]) ? node3311 : 16'b0000000111111111;
														assign node3311 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3314 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3317 = (inp[2]) ? node3357 : node3318;
											assign node3318 = (inp[9]) ? node3332 : node3319;
												assign node3319 = (inp[13]) ? 16'b0000000111111111 : node3320;
													assign node3320 = (inp[14]) ? node3326 : node3321;
														assign node3321 = (inp[6]) ? 16'b0000001111111111 : node3322;
															assign node3322 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3326 = (inp[5]) ? 16'b0000000111111111 : node3327;
															assign node3327 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3332 = (inp[5]) ? node3342 : node3333;
													assign node3333 = (inp[14]) ? node3339 : node3334;
														assign node3334 = (inp[7]) ? 16'b0000001111111111 : node3335;
															assign node3335 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3339 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3342 = (inp[6]) ? node3346 : node3343;
														assign node3343 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3346 = (inp[7]) ? node3352 : node3347;
															assign node3347 = (inp[14]) ? node3349 : 16'b0000000011111111;
																assign node3349 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node3352 = (inp[13]) ? 16'b0000000001111111 : node3353;
																assign node3353 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3357 = (inp[14]) ? node3367 : node3358;
												assign node3358 = (inp[7]) ? node3364 : node3359;
													assign node3359 = (inp[6]) ? 16'b0000000111111111 : node3360;
														assign node3360 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3364 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3367 = (inp[5]) ? node3377 : node3368;
													assign node3368 = (inp[6]) ? node3372 : node3369;
														assign node3369 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3372 = (inp[13]) ? node3374 : 16'b0000000001111111;
															assign node3374 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3377 = (inp[13]) ? node3379 : 16'b0000000001111111;
														assign node3379 = (inp[7]) ? 16'b0000000000111111 : node3380;
															assign node3380 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3384 = (inp[6]) ? node3496 : node3385;
									assign node3385 = (inp[7]) ? node3437 : node3386;
										assign node3386 = (inp[3]) ? node3410 : node3387;
											assign node3387 = (inp[5]) ? node3399 : node3388;
												assign node3388 = (inp[2]) ? node3394 : node3389;
													assign node3389 = (inp[13]) ? 16'b0000011111111111 : node3390;
														assign node3390 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3394 = (inp[13]) ? node3396 : 16'b0000001111111111;
														assign node3396 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3399 = (inp[14]) ? node3401 : 16'b0000001111111111;
													assign node3401 = (inp[13]) ? node3407 : node3402;
														assign node3402 = (inp[2]) ? 16'b0000000111111111 : node3403;
															assign node3403 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3407 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3410 = (inp[14]) ? node3430 : node3411;
												assign node3411 = (inp[13]) ? node3421 : node3412;
													assign node3412 = (inp[2]) ? 16'b0000000111111111 : node3413;
														assign node3413 = (inp[9]) ? 16'b0000001111111111 : node3414;
															assign node3414 = (inp[15]) ? node3416 : 16'b0000011111111111;
																assign node3416 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3421 = (inp[15]) ? node3427 : node3422;
														assign node3422 = (inp[2]) ? node3424 : 16'b0000001111111111;
															assign node3424 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3427 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3430 = (inp[13]) ? 16'b0000000011111111 : node3431;
													assign node3431 = (inp[9]) ? node3433 : 16'b0000000111111111;
														assign node3433 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node3437 = (inp[13]) ? node3469 : node3438;
											assign node3438 = (inp[5]) ? node3448 : node3439;
												assign node3439 = (inp[14]) ? node3441 : 16'b0000001111111111;
													assign node3441 = (inp[2]) ? 16'b0000000111111111 : node3442;
														assign node3442 = (inp[9]) ? node3444 : 16'b0000001111111111;
															assign node3444 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3448 = (inp[14]) ? node3464 : node3449;
													assign node3449 = (inp[3]) ? node3455 : node3450;
														assign node3450 = (inp[9]) ? 16'b0000000111111111 : node3451;
															assign node3451 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3455 = (inp[2]) ? node3459 : node3456;
															assign node3456 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3459 = (inp[15]) ? 16'b0000000011111111 : node3460;
																assign node3460 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3464 = (inp[9]) ? node3466 : 16'b0000000011111111;
														assign node3466 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3469 = (inp[3]) ? node3485 : node3470;
												assign node3470 = (inp[5]) ? node3480 : node3471;
													assign node3471 = (inp[14]) ? node3475 : node3472;
														assign node3472 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3475 = (inp[9]) ? 16'b0000000011111111 : node3476;
															assign node3476 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3480 = (inp[14]) ? node3482 : 16'b0000000011111111;
														assign node3482 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3485 = (inp[2]) ? node3493 : node3486;
													assign node3486 = (inp[9]) ? node3488 : 16'b0000000111111111;
														assign node3488 = (inp[15]) ? 16'b0000000001111111 : node3489;
															assign node3489 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3493 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3496 = (inp[15]) ? node3560 : node3497;
										assign node3497 = (inp[14]) ? node3523 : node3498;
											assign node3498 = (inp[5]) ? node3512 : node3499;
												assign node3499 = (inp[7]) ? node3507 : node3500;
													assign node3500 = (inp[2]) ? 16'b0000001111111111 : node3501;
														assign node3501 = (inp[13]) ? 16'b0000001111111111 : node3502;
															assign node3502 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3507 = (inp[9]) ? 16'b0000000111111111 : node3508;
														assign node3508 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3512 = (inp[9]) ? node3514 : 16'b0000000111111111;
													assign node3514 = (inp[13]) ? node3520 : node3515;
														assign node3515 = (inp[7]) ? node3517 : 16'b0000001111111111;
															assign node3517 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3520 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3523 = (inp[7]) ? node3537 : node3524;
												assign node3524 = (inp[5]) ? node3526 : 16'b0000001111111111;
													assign node3526 = (inp[9]) ? node3534 : node3527;
														assign node3527 = (inp[2]) ? 16'b0000000011111111 : node3528;
															assign node3528 = (inp[3]) ? node3530 : 16'b0000000111111111;
																assign node3530 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3534 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3537 = (inp[5]) ? node3547 : node3538;
													assign node3538 = (inp[13]) ? node3540 : 16'b0000000111111111;
														assign node3540 = (inp[9]) ? 16'b0000000001111111 : node3541;
															assign node3541 = (inp[2]) ? node3543 : 16'b0000000011111111;
																assign node3543 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3547 = (inp[3]) ? node3555 : node3548;
														assign node3548 = (inp[2]) ? node3550 : 16'b0000000011111111;
															assign node3550 = (inp[13]) ? 16'b0000000001111111 : node3551;
																assign node3551 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3555 = (inp[13]) ? node3557 : 16'b0000000001111111;
															assign node3557 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3560 = (inp[13]) ? node3598 : node3561;
											assign node3561 = (inp[7]) ? node3585 : node3562;
												assign node3562 = (inp[5]) ? node3572 : node3563;
													assign node3563 = (inp[2]) ? node3569 : node3564;
														assign node3564 = (inp[14]) ? 16'b0000000111111111 : node3565;
															assign node3565 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node3569 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3572 = (inp[14]) ? node3576 : node3573;
														assign node3573 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3576 = (inp[9]) ? node3580 : node3577;
															assign node3577 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node3580 = (inp[3]) ? node3582 : 16'b0000000001111111;
																assign node3582 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3585 = (inp[2]) ? node3591 : node3586;
													assign node3586 = (inp[3]) ? node3588 : 16'b0000000011111111;
														assign node3588 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3591 = (inp[9]) ? node3595 : node3592;
														assign node3592 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3595 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3598 = (inp[14]) ? node3610 : node3599;
												assign node3599 = (inp[2]) ? 16'b0000000001111111 : node3600;
													assign node3600 = (inp[3]) ? node3602 : 16'b0000000011111111;
														assign node3602 = (inp[9]) ? node3604 : 16'b0000000011111111;
															assign node3604 = (inp[7]) ? 16'b0000000001111111 : node3605;
																assign node3605 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3610 = (inp[9]) ? node3620 : node3611;
													assign node3611 = (inp[7]) ? node3617 : node3612;
														assign node3612 = (inp[2]) ? 16'b0000000001111111 : node3613;
															assign node3613 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3617 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node3620 = (inp[3]) ? node3624 : node3621;
														assign node3621 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3624 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node3627 = (inp[3]) ? node3891 : node3628;
								assign node3628 = (inp[7]) ? node3762 : node3629;
									assign node3629 = (inp[14]) ? node3701 : node3630;
										assign node3630 = (inp[5]) ? node3668 : node3631;
											assign node3631 = (inp[9]) ? node3653 : node3632;
												assign node3632 = (inp[15]) ? node3642 : node3633;
													assign node3633 = (inp[12]) ? node3639 : node3634;
														assign node3634 = (inp[13]) ? 16'b0000011111111111 : node3635;
															assign node3635 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3639 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3642 = (inp[6]) ? node3648 : node3643;
														assign node3643 = (inp[12]) ? node3645 : 16'b0000011111111111;
															assign node3645 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3648 = (inp[13]) ? node3650 : 16'b0000001111111111;
															assign node3650 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3653 = (inp[12]) ? node3659 : node3654;
													assign node3654 = (inp[13]) ? node3656 : 16'b0000011111111111;
														assign node3656 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3659 = (inp[15]) ? 16'b0000000011111111 : node3660;
														assign node3660 = (inp[6]) ? 16'b0000000111111111 : node3661;
															assign node3661 = (inp[2]) ? node3663 : 16'b0000001111111111;
																assign node3663 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3668 = (inp[12]) ? node3686 : node3669;
												assign node3669 = (inp[2]) ? node3673 : node3670;
													assign node3670 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3673 = (inp[9]) ? node3681 : node3674;
														assign node3674 = (inp[13]) ? node3676 : 16'b0000001111111111;
															assign node3676 = (inp[6]) ? 16'b0000000111111111 : node3677;
																assign node3677 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3681 = (inp[6]) ? node3683 : 16'b0000000111111111;
															assign node3683 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3686 = (inp[13]) ? node3694 : node3687;
													assign node3687 = (inp[2]) ? 16'b0000000111111111 : node3688;
														assign node3688 = (inp[6]) ? 16'b0000000111111111 : node3689;
															assign node3689 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3694 = (inp[15]) ? 16'b0000000001111111 : node3695;
														assign node3695 = (inp[9]) ? node3697 : 16'b0000000111111111;
															assign node3697 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3701 = (inp[12]) ? node3729 : node3702;
											assign node3702 = (inp[6]) ? node3718 : node3703;
												assign node3703 = (inp[13]) ? node3709 : node3704;
													assign node3704 = (inp[9]) ? node3706 : 16'b0000011111111111;
														assign node3706 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3709 = (inp[9]) ? node3715 : node3710;
														assign node3710 = (inp[2]) ? 16'b0000000111111111 : node3711;
															assign node3711 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3715 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3718 = (inp[2]) ? node3724 : node3719;
													assign node3719 = (inp[9]) ? 16'b0000000111111111 : node3720;
														assign node3720 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3724 = (inp[9]) ? 16'b0000000001111111 : node3725;
														assign node3725 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3729 = (inp[9]) ? node3749 : node3730;
												assign node3730 = (inp[2]) ? node3740 : node3731;
													assign node3731 = (inp[6]) ? node3735 : node3732;
														assign node3732 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3735 = (inp[15]) ? node3737 : 16'b0000000111111111;
															assign node3737 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3740 = (inp[13]) ? node3744 : node3741;
														assign node3741 = (inp[6]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node3744 = (inp[15]) ? 16'b0000000001111111 : node3745;
															assign node3745 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3749 = (inp[5]) ? node3753 : node3750;
													assign node3750 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3753 = (inp[13]) ? node3759 : node3754;
														assign node3754 = (inp[2]) ? 16'b0000000001111111 : node3755;
															assign node3755 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3759 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3762 = (inp[15]) ? node3836 : node3763;
										assign node3763 = (inp[2]) ? node3793 : node3764;
											assign node3764 = (inp[6]) ? node3776 : node3765;
												assign node3765 = (inp[14]) ? node3769 : node3766;
													assign node3766 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3769 = (inp[13]) ? node3773 : node3770;
														assign node3770 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3773 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3776 = (inp[14]) ? node3784 : node3777;
													assign node3777 = (inp[13]) ? node3781 : node3778;
														assign node3778 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node3781 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3784 = (inp[9]) ? node3790 : node3785;
														assign node3785 = (inp[5]) ? node3787 : 16'b0000000111111111;
															assign node3787 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3790 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3793 = (inp[14]) ? node3819 : node3794;
												assign node3794 = (inp[13]) ? node3808 : node3795;
													assign node3795 = (inp[5]) ? node3805 : node3796;
														assign node3796 = (inp[9]) ? node3802 : node3797;
															assign node3797 = (inp[6]) ? 16'b0000001111111111 : node3798;
																assign node3798 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node3802 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3805 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3808 = (inp[12]) ? node3812 : node3809;
														assign node3809 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3812 = (inp[6]) ? 16'b0000000001111111 : node3813;
															assign node3813 = (inp[5]) ? node3815 : 16'b0000000011111111;
																assign node3815 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3819 = (inp[13]) ? node3831 : node3820;
													assign node3820 = (inp[5]) ? node3826 : node3821;
														assign node3821 = (inp[12]) ? 16'b0000000011111111 : node3822;
															assign node3822 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3826 = (inp[12]) ? 16'b0000000001111111 : node3827;
															assign node3827 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3831 = (inp[9]) ? node3833 : 16'b0000000001111111;
														assign node3833 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3836 = (inp[6]) ? node3858 : node3837;
											assign node3837 = (inp[2]) ? node3853 : node3838;
												assign node3838 = (inp[5]) ? node3842 : node3839;
													assign node3839 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node3842 = (inp[12]) ? node3848 : node3843;
														assign node3843 = (inp[13]) ? 16'b0000000011111111 : node3844;
															assign node3844 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3848 = (inp[9]) ? 16'b0000000001111111 : node3849;
															assign node3849 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3853 = (inp[5]) ? 16'b0000000001111111 : node3854;
													assign node3854 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3858 = (inp[13]) ? node3882 : node3859;
												assign node3859 = (inp[9]) ? node3871 : node3860;
													assign node3860 = (inp[14]) ? 16'b0000000000111111 : node3861;
														assign node3861 = (inp[5]) ? node3865 : node3862;
															assign node3862 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3865 = (inp[12]) ? 16'b0000000011111111 : node3866;
																assign node3866 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3871 = (inp[12]) ? node3875 : node3872;
														assign node3872 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3875 = (inp[14]) ? 16'b0000000000111111 : node3876;
															assign node3876 = (inp[2]) ? node3878 : 16'b0000000001111111;
																assign node3878 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3882 = (inp[5]) ? node3884 : 16'b0000000001111111;
													assign node3884 = (inp[9]) ? node3888 : node3885;
														assign node3885 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3888 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3891 = (inp[6]) ? node4013 : node3892;
									assign node3892 = (inp[12]) ? node3962 : node3893;
										assign node3893 = (inp[13]) ? node3929 : node3894;
											assign node3894 = (inp[2]) ? node3908 : node3895;
												assign node3895 = (inp[14]) ? node3901 : node3896;
													assign node3896 = (inp[9]) ? node3898 : 16'b0000011111111111;
														assign node3898 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node3901 = (inp[15]) ? node3905 : node3902;
														assign node3902 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3905 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3908 = (inp[7]) ? node3920 : node3909;
													assign node3909 = (inp[15]) ? node3913 : node3910;
														assign node3910 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3913 = (inp[9]) ? 16'b0000000011111111 : node3914;
															assign node3914 = (inp[5]) ? node3916 : 16'b0000000111111111;
																assign node3916 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3920 = (inp[15]) ? node3926 : node3921;
														assign node3921 = (inp[14]) ? 16'b0000000011111111 : node3922;
															assign node3922 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3926 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node3929 = (inp[5]) ? node3943 : node3930;
												assign node3930 = (inp[15]) ? node3934 : node3931;
													assign node3931 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3934 = (inp[14]) ? node3938 : node3935;
														assign node3935 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3938 = (inp[2]) ? node3940 : 16'b0000000011111111;
															assign node3940 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3943 = (inp[2]) ? node3953 : node3944;
													assign node3944 = (inp[7]) ? node3948 : node3945;
														assign node3945 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3948 = (inp[14]) ? 16'b0000000000111111 : node3949;
															assign node3949 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3953 = (inp[15]) ? node3957 : node3954;
														assign node3954 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3957 = (inp[14]) ? node3959 : 16'b0000000001111111;
															assign node3959 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3962 = (inp[14]) ? node3984 : node3963;
											assign node3963 = (inp[7]) ? node3971 : node3964;
												assign node3964 = (inp[15]) ? node3966 : 16'b0000000111111111;
													assign node3966 = (inp[9]) ? 16'b0000000011111111 : node3967;
														assign node3967 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3971 = (inp[15]) ? node3973 : 16'b0000000011111111;
													assign node3973 = (inp[2]) ? node3979 : node3974;
														assign node3974 = (inp[5]) ? 16'b0000000001111111 : node3975;
															assign node3975 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3979 = (inp[5]) ? node3981 : 16'b0000000000111111;
															assign node3981 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3984 = (inp[13]) ? node4002 : node3985;
												assign node3985 = (inp[9]) ? node3991 : node3986;
													assign node3986 = (inp[15]) ? 16'b0000000011111111 : node3987;
														assign node3987 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3991 = (inp[15]) ? node3999 : node3992;
														assign node3992 = (inp[7]) ? 16'b0000000001111111 : node3993;
															assign node3993 = (inp[5]) ? node3995 : 16'b0000000011111111;
																assign node3995 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3999 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4002 = (inp[9]) ? node4010 : node4003;
													assign node4003 = (inp[5]) ? 16'b0000000000111111 : node4004;
														assign node4004 = (inp[15]) ? node4006 : 16'b0000000011111111;
															assign node4006 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4010 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4013 = (inp[7]) ? node4097 : node4014;
										assign node4014 = (inp[5]) ? node4060 : node4015;
											assign node4015 = (inp[15]) ? node4037 : node4016;
												assign node4016 = (inp[12]) ? node4034 : node4017;
													assign node4017 = (inp[14]) ? node4025 : node4018;
														assign node4018 = (inp[13]) ? 16'b0000001111111111 : node4019;
															assign node4019 = (inp[2]) ? 16'b0000001111111111 : node4020;
																assign node4020 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4025 = (inp[2]) ? node4029 : node4026;
															assign node4026 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node4029 = (inp[9]) ? 16'b0000000011111111 : node4030;
																assign node4030 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4034 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4037 = (inp[14]) ? node4049 : node4038;
													assign node4038 = (inp[12]) ? node4044 : node4039;
														assign node4039 = (inp[13]) ? node4041 : 16'b0000000011111111;
															assign node4041 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4044 = (inp[2]) ? 16'b0000000011111111 : node4045;
															assign node4045 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4049 = (inp[2]) ? node4055 : node4050;
														assign node4050 = (inp[9]) ? 16'b0000000001111111 : node4051;
															assign node4051 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4055 = (inp[13]) ? node4057 : 16'b0000000001111111;
															assign node4057 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4060 = (inp[14]) ? node4080 : node4061;
												assign node4061 = (inp[13]) ? node4069 : node4062;
													assign node4062 = (inp[2]) ? node4064 : 16'b0000000011111111;
														assign node4064 = (inp[12]) ? 16'b0000000001111111 : node4065;
															assign node4065 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4069 = (inp[12]) ? node4073 : node4070;
														assign node4070 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4073 = (inp[9]) ? node4075 : 16'b0000000001111111;
															assign node4075 = (inp[15]) ? 16'b0000000000111111 : node4076;
																assign node4076 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4080 = (inp[9]) ? node4090 : node4081;
													assign node4081 = (inp[12]) ? node4087 : node4082;
														assign node4082 = (inp[2]) ? 16'b0000000001111111 : node4083;
															assign node4083 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4087 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4090 = (inp[15]) ? 16'b0000000000011111 : node4091;
														assign node4091 = (inp[2]) ? node4093 : 16'b0000000001111111;
															assign node4093 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4097 = (inp[2]) ? node4123 : node4098;
											assign node4098 = (inp[13]) ? node4112 : node4099;
												assign node4099 = (inp[14]) ? node4109 : node4100;
													assign node4100 = (inp[5]) ? node4102 : 16'b0000000111111111;
														assign node4102 = (inp[15]) ? node4104 : 16'b0000000011111111;
															assign node4104 = (inp[12]) ? 16'b0000000001111111 : node4105;
																assign node4105 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4109 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4112 = (inp[12]) ? node4118 : node4113;
													assign node4113 = (inp[9]) ? node4115 : 16'b0000000001111111;
														assign node4115 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4118 = (inp[14]) ? 16'b0000000000011111 : node4119;
														assign node4119 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4123 = (inp[15]) ? node4135 : node4124;
												assign node4124 = (inp[5]) ? node4126 : 16'b0000000001111111;
													assign node4126 = (inp[12]) ? node4132 : node4127;
														assign node4127 = (inp[9]) ? node4129 : 16'b0000000001111111;
															assign node4129 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node4132 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node4135 = (inp[9]) ? node4143 : node4136;
													assign node4136 = (inp[13]) ? node4140 : node4137;
														assign node4137 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node4140 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node4143 = (inp[12]) ? node4151 : node4144;
														assign node4144 = (inp[13]) ? 16'b0000000000011111 : node4145;
															assign node4145 = (inp[5]) ? node4147 : 16'b0000000000111111;
																assign node4147 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node4151 = (inp[13]) ? 16'b0000000000001111 : node4152;
															assign node4152 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
				assign node4156 = (inp[14]) ? node6282 : node4157;
					assign node4157 = (inp[13]) ? node5209 : node4158;
						assign node4158 = (inp[2]) ? node4684 : node4159;
							assign node4159 = (inp[3]) ? node4423 : node4160;
								assign node4160 = (inp[9]) ? node4288 : node4161;
									assign node4161 = (inp[1]) ? node4219 : node4162;
										assign node4162 = (inp[5]) ? node4198 : node4163;
											assign node4163 = (inp[6]) ? node4183 : node4164;
												assign node4164 = (inp[12]) ? node4174 : node4165;
													assign node4165 = (inp[8]) ? node4171 : node4166;
														assign node4166 = (inp[11]) ? 16'b0001111111111111 : node4167;
															assign node4167 = (inp[7]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node4171 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node4174 = (inp[15]) ? node4180 : node4175;
														assign node4175 = (inp[7]) ? 16'b0000111111111111 : node4176;
															assign node4176 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4180 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4183 = (inp[11]) ? node4187 : node4184;
													assign node4184 = (inp[8]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node4187 = (inp[15]) ? node4191 : node4188;
														assign node4188 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4191 = (inp[12]) ? node4193 : 16'b0000011111111111;
															assign node4193 = (inp[8]) ? 16'b0000001111111111 : node4194;
																assign node4194 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4198 = (inp[15]) ? node4208 : node4199;
												assign node4199 = (inp[11]) ? 16'b0000011111111111 : node4200;
													assign node4200 = (inp[12]) ? node4202 : 16'b0000011111111111;
														assign node4202 = (inp[7]) ? 16'b0000111111111111 : node4203;
															assign node4203 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node4208 = (inp[7]) ? node4210 : 16'b0000011111111111;
													assign node4210 = (inp[11]) ? node4214 : node4211;
														assign node4211 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4214 = (inp[12]) ? node4216 : 16'b0000001111111111;
															assign node4216 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4219 = (inp[11]) ? node4253 : node4220;
											assign node4220 = (inp[15]) ? node4234 : node4221;
												assign node4221 = (inp[12]) ? node4229 : node4222;
													assign node4222 = (inp[6]) ? node4224 : 16'b0001111111111111;
														assign node4224 = (inp[7]) ? node4226 : 16'b0000111111111111;
															assign node4226 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4229 = (inp[7]) ? 16'b0000011111111111 : node4230;
														assign node4230 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4234 = (inp[12]) ? node4246 : node4235;
													assign node4235 = (inp[6]) ? node4241 : node4236;
														assign node4236 = (inp[8]) ? node4238 : 16'b0001111111111111;
															assign node4238 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4241 = (inp[8]) ? 16'b0000001111111111 : node4242;
															assign node4242 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4246 = (inp[7]) ? node4250 : node4247;
														assign node4247 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4250 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node4253 = (inp[12]) ? node4277 : node4254;
												assign node4254 = (inp[15]) ? node4266 : node4255;
													assign node4255 = (inp[6]) ? node4263 : node4256;
														assign node4256 = (inp[7]) ? node4260 : node4257;
															assign node4257 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node4260 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4263 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4266 = (inp[8]) ? node4270 : node4267;
														assign node4267 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4270 = (inp[5]) ? 16'b0000000111111111 : node4271;
															assign node4271 = (inp[6]) ? node4273 : 16'b0000001111111111;
																assign node4273 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4277 = (inp[5]) ? node4285 : node4278;
													assign node4278 = (inp[15]) ? 16'b0000000111111111 : node4279;
														assign node4279 = (inp[8]) ? 16'b0000001111111111 : node4280;
															assign node4280 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4285 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4288 = (inp[1]) ? node4354 : node4289;
										assign node4289 = (inp[6]) ? node4325 : node4290;
											assign node4290 = (inp[8]) ? node4306 : node4291;
												assign node4291 = (inp[12]) ? node4297 : node4292;
													assign node4292 = (inp[5]) ? node4294 : 16'b0001111111111111;
														assign node4294 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4297 = (inp[7]) ? 16'b0000011111111111 : node4298;
														assign node4298 = (inp[5]) ? node4300 : 16'b0000111111111111;
															assign node4300 = (inp[11]) ? 16'b0000011111111111 : node4301;
																assign node4301 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4306 = (inp[11]) ? node4318 : node4307;
													assign node4307 = (inp[7]) ? node4311 : node4308;
														assign node4308 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4311 = (inp[15]) ? 16'b0000001111111111 : node4312;
															assign node4312 = (inp[5]) ? node4314 : 16'b0000011111111111;
																assign node4314 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4318 = (inp[12]) ? 16'b0000001111111111 : node4319;
														assign node4319 = (inp[15]) ? 16'b0000001111111111 : node4320;
															assign node4320 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4325 = (inp[12]) ? node4343 : node4326;
												assign node4326 = (inp[7]) ? node4332 : node4327;
													assign node4327 = (inp[11]) ? node4329 : 16'b0000111111111111;
														assign node4329 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4332 = (inp[11]) ? node4336 : node4333;
														assign node4333 = (inp[5]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node4336 = (inp[5]) ? 16'b0000000111111111 : node4337;
															assign node4337 = (inp[8]) ? node4339 : 16'b0000001111111111;
																assign node4339 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4343 = (inp[8]) ? node4349 : node4344;
													assign node4344 = (inp[11]) ? node4346 : 16'b0000001111111111;
														assign node4346 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4349 = (inp[7]) ? node4351 : 16'b0000001111111111;
														assign node4351 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4354 = (inp[7]) ? node4388 : node4355;
											assign node4355 = (inp[11]) ? node4377 : node4356;
												assign node4356 = (inp[8]) ? node4366 : node4357;
													assign node4357 = (inp[15]) ? node4359 : 16'b0000111111111111;
														assign node4359 = (inp[5]) ? node4361 : 16'b0000011111111111;
															assign node4361 = (inp[12]) ? 16'b0000001111111111 : node4362;
																assign node4362 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4366 = (inp[15]) ? node4372 : node4367;
														assign node4367 = (inp[6]) ? 16'b0000001111111111 : node4368;
															assign node4368 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4372 = (inp[12]) ? 16'b0000000111111111 : node4373;
															assign node4373 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4377 = (inp[5]) ? node4379 : 16'b0000001111111111;
													assign node4379 = (inp[15]) ? 16'b0000000111111111 : node4380;
														assign node4380 = (inp[6]) ? 16'b0000000111111111 : node4381;
															assign node4381 = (inp[12]) ? node4383 : 16'b0000001111111111;
																assign node4383 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4388 = (inp[5]) ? node4406 : node4389;
												assign node4389 = (inp[8]) ? node4401 : node4390;
													assign node4390 = (inp[6]) ? node4398 : node4391;
														assign node4391 = (inp[12]) ? 16'b0000000111111111 : node4392;
															assign node4392 = (inp[11]) ? node4394 : 16'b0000011111111111;
																assign node4394 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4398 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4401 = (inp[11]) ? 16'b0000000011111111 : node4402;
														assign node4402 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4406 = (inp[15]) ? node4412 : node4407;
													assign node4407 = (inp[12]) ? 16'b0000000111111111 : node4408;
														assign node4408 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4412 = (inp[8]) ? node4420 : node4413;
														assign node4413 = (inp[6]) ? 16'b0000000001111111 : node4414;
															assign node4414 = (inp[11]) ? node4416 : 16'b0000000111111111;
																assign node4416 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4420 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node4423 = (inp[12]) ? node4555 : node4424;
									assign node4424 = (inp[8]) ? node4490 : node4425;
										assign node4425 = (inp[15]) ? node4473 : node4426;
											assign node4426 = (inp[6]) ? node4456 : node4427;
												assign node4427 = (inp[7]) ? node4443 : node4428;
													assign node4428 = (inp[5]) ? node4434 : node4429;
														assign node4429 = (inp[1]) ? node4431 : 16'b0001111111111111;
															assign node4431 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4434 = (inp[11]) ? node4438 : node4435;
															assign node4435 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node4438 = (inp[9]) ? 16'b0000011111111111 : node4439;
																assign node4439 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4443 = (inp[11]) ? node4449 : node4444;
														assign node4444 = (inp[5]) ? node4446 : 16'b0000111111111111;
															assign node4446 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4449 = (inp[5]) ? 16'b0000011111111111 : node4450;
															assign node4450 = (inp[9]) ? 16'b0000011111111111 : node4451;
																assign node4451 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4456 = (inp[1]) ? node4466 : node4457;
													assign node4457 = (inp[7]) ? node4461 : node4458;
														assign node4458 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4461 = (inp[5]) ? node4463 : 16'b0000011111111111;
															assign node4463 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4466 = (inp[9]) ? node4468 : 16'b0000001111111111;
														assign node4468 = (inp[11]) ? node4470 : 16'b0000001111111111;
															assign node4470 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4473 = (inp[1]) ? node4483 : node4474;
												assign node4474 = (inp[6]) ? 16'b0000001111111111 : node4475;
													assign node4475 = (inp[11]) ? 16'b0000001111111111 : node4476;
														assign node4476 = (inp[9]) ? 16'b0000011111111111 : node4477;
															assign node4477 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node4483 = (inp[5]) ? 16'b0000000111111111 : node4484;
													assign node4484 = (inp[11]) ? 16'b0000000111111111 : node4485;
														assign node4485 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node4490 = (inp[7]) ? node4528 : node4491;
											assign node4491 = (inp[5]) ? node4505 : node4492;
												assign node4492 = (inp[15]) ? node4500 : node4493;
													assign node4493 = (inp[11]) ? node4497 : node4494;
														assign node4494 = (inp[9]) ? 16'b0000111111111111 : 16'b0000011111111111;
														assign node4497 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4500 = (inp[1]) ? 16'b0000001111111111 : node4501;
														assign node4501 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4505 = (inp[11]) ? node4515 : node4506;
													assign node4506 = (inp[6]) ? node4510 : node4507;
														assign node4507 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4510 = (inp[15]) ? node4512 : 16'b0000001111111111;
															assign node4512 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4515 = (inp[15]) ? node4523 : node4516;
														assign node4516 = (inp[6]) ? 16'b0000000111111111 : node4517;
															assign node4517 = (inp[1]) ? node4519 : 16'b0000001111111111;
																assign node4519 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4523 = (inp[6]) ? node4525 : 16'b0000000111111111;
															assign node4525 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4528 = (inp[9]) ? node4540 : node4529;
												assign node4529 = (inp[1]) ? 16'b0000000111111111 : node4530;
													assign node4530 = (inp[6]) ? node4536 : node4531;
														assign node4531 = (inp[11]) ? 16'b0000001111111111 : node4532;
															assign node4532 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node4536 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4540 = (inp[6]) ? node4550 : node4541;
													assign node4541 = (inp[5]) ? 16'b0000000011111111 : node4542;
														assign node4542 = (inp[11]) ? node4544 : 16'b0000001111111111;
															assign node4544 = (inp[15]) ? 16'b0000000111111111 : node4545;
																assign node4545 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4550 = (inp[11]) ? 16'b0000000011111111 : node4551;
														assign node4551 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4555 = (inp[5]) ? node4619 : node4556;
										assign node4556 = (inp[1]) ? node4582 : node4557;
											assign node4557 = (inp[6]) ? node4567 : node4558;
												assign node4558 = (inp[9]) ? 16'b0000001111111111 : node4559;
													assign node4559 = (inp[8]) ? node4563 : node4560;
														assign node4560 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4563 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4567 = (inp[7]) ? node4575 : node4568;
													assign node4568 = (inp[11]) ? node4572 : node4569;
														assign node4569 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4572 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4575 = (inp[9]) ? node4579 : node4576;
														assign node4576 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4579 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4582 = (inp[8]) ? node4602 : node4583;
												assign node4583 = (inp[6]) ? node4591 : node4584;
													assign node4584 = (inp[15]) ? node4586 : 16'b0000011111111111;
														assign node4586 = (inp[9]) ? node4588 : 16'b0000001111111111;
															assign node4588 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4591 = (inp[15]) ? node4597 : node4592;
														assign node4592 = (inp[7]) ? node4594 : 16'b0000001111111111;
															assign node4594 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4597 = (inp[11]) ? node4599 : 16'b0000000111111111;
															assign node4599 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4602 = (inp[6]) ? node4612 : node4603;
													assign node4603 = (inp[11]) ? node4607 : node4604;
														assign node4604 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4607 = (inp[15]) ? node4609 : 16'b0000000111111111;
															assign node4609 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4612 = (inp[7]) ? node4616 : node4613;
														assign node4613 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4616 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4619 = (inp[15]) ? node4645 : node4620;
											assign node4620 = (inp[9]) ? node4636 : node4621;
												assign node4621 = (inp[1]) ? node4629 : node4622;
													assign node4622 = (inp[6]) ? node4626 : node4623;
														assign node4623 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4626 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4629 = (inp[11]) ? 16'b0000000001111111 : node4630;
														assign node4630 = (inp[7]) ? 16'b0000000111111111 : node4631;
															assign node4631 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4636 = (inp[7]) ? node4638 : 16'b0000000111111111;
													assign node4638 = (inp[6]) ? node4640 : 16'b0000000111111111;
														assign node4640 = (inp[1]) ? node4642 : 16'b0000000011111111;
															assign node4642 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4645 = (inp[8]) ? node4661 : node4646;
												assign node4646 = (inp[11]) ? node4652 : node4647;
													assign node4647 = (inp[9]) ? node4649 : 16'b0000000111111111;
														assign node4649 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4652 = (inp[7]) ? node4654 : 16'b0000001111111111;
														assign node4654 = (inp[6]) ? 16'b0000000001111111 : node4655;
															assign node4655 = (inp[9]) ? 16'b0000000011111111 : node4656;
																assign node4656 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4661 = (inp[1]) ? node4675 : node4662;
													assign node4662 = (inp[7]) ? node4668 : node4663;
														assign node4663 = (inp[6]) ? node4665 : 16'b0000000111111111;
															assign node4665 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4668 = (inp[11]) ? node4670 : 16'b0000000011111111;
															assign node4670 = (inp[9]) ? 16'b0000000001111111 : node4671;
																assign node4671 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4675 = (inp[7]) ? node4677 : 16'b0000000001111111;
														assign node4677 = (inp[9]) ? node4679 : 16'b0000000001111111;
															assign node4679 = (inp[11]) ? 16'b0000000000111111 : node4680;
																assign node4680 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4684 = (inp[9]) ? node4950 : node4685;
								assign node4685 = (inp[15]) ? node4819 : node4686;
									assign node4686 = (inp[5]) ? node4752 : node4687;
										assign node4687 = (inp[3]) ? node4715 : node4688;
											assign node4688 = (inp[7]) ? node4702 : node4689;
												assign node4689 = (inp[1]) ? node4697 : node4690;
													assign node4690 = (inp[12]) ? 16'b0000111111111111 : node4691;
														assign node4691 = (inp[6]) ? 16'b0001111111111111 : node4692;
															assign node4692 = (inp[8]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node4697 = (inp[12]) ? 16'b0000001111111111 : node4698;
														assign node4698 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4702 = (inp[6]) ? node4708 : node4703;
													assign node4703 = (inp[8]) ? 16'b0000011111111111 : node4704;
														assign node4704 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4708 = (inp[12]) ? 16'b0000001111111111 : node4709;
														assign node4709 = (inp[11]) ? node4711 : 16'b0000111111111111;
															assign node4711 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node4715 = (inp[1]) ? node4745 : node4716;
												assign node4716 = (inp[12]) ? node4732 : node4717;
													assign node4717 = (inp[11]) ? node4723 : node4718;
														assign node4718 = (inp[8]) ? 16'b0000011111111111 : node4719;
															assign node4719 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4723 = (inp[8]) ? 16'b0000001111111111 : node4724;
															assign node4724 = (inp[7]) ? node4728 : node4725;
																assign node4725 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
																assign node4728 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4732 = (inp[6]) ? node4740 : node4733;
														assign node4733 = (inp[11]) ? node4735 : 16'b0000011111111111;
															assign node4735 = (inp[7]) ? 16'b0000001111111111 : node4736;
																assign node4736 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4740 = (inp[11]) ? node4742 : 16'b0000001111111111;
															assign node4742 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4745 = (inp[11]) ? 16'b0000000111111111 : node4746;
													assign node4746 = (inp[7]) ? node4748 : 16'b0000011111111111;
														assign node4748 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node4752 = (inp[7]) ? node4790 : node4753;
											assign node4753 = (inp[1]) ? node4777 : node4754;
												assign node4754 = (inp[6]) ? node4770 : node4755;
													assign node4755 = (inp[3]) ? node4761 : node4756;
														assign node4756 = (inp[8]) ? node4758 : 16'b0000111111111111;
															assign node4758 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4761 = (inp[11]) ? node4765 : node4762;
															assign node4762 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node4765 = (inp[12]) ? 16'b0000001111111111 : node4766;
																assign node4766 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4770 = (inp[8]) ? node4772 : 16'b0000011111111111;
														assign node4772 = (inp[11]) ? node4774 : 16'b0000001111111111;
															assign node4774 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4777 = (inp[8]) ? node4783 : node4778;
													assign node4778 = (inp[11]) ? 16'b0000001111111111 : node4779;
														assign node4779 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4783 = (inp[11]) ? node4785 : 16'b0000001111111111;
														assign node4785 = (inp[6]) ? 16'b0000000111111111 : node4786;
															assign node4786 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4790 = (inp[3]) ? node4806 : node4791;
												assign node4791 = (inp[8]) ? node4799 : node4792;
													assign node4792 = (inp[11]) ? node4796 : node4793;
														assign node4793 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4796 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4799 = (inp[12]) ? node4801 : 16'b0000000011111111;
														assign node4801 = (inp[6]) ? node4803 : 16'b0000000111111111;
															assign node4803 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4806 = (inp[11]) ? node4814 : node4807;
													assign node4807 = (inp[12]) ? node4809 : 16'b0000000111111111;
														assign node4809 = (inp[6]) ? 16'b0000000011111111 : node4810;
															assign node4810 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4814 = (inp[1]) ? node4816 : 16'b0000000011111111;
														assign node4816 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4819 = (inp[11]) ? node4873 : node4820;
										assign node4820 = (inp[3]) ? node4844 : node4821;
											assign node4821 = (inp[1]) ? node4837 : node4822;
												assign node4822 = (inp[6]) ? node4826 : node4823;
													assign node4823 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4826 = (inp[12]) ? node4830 : node4827;
														assign node4827 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4830 = (inp[5]) ? node4832 : 16'b0000001111111111;
															assign node4832 = (inp[7]) ? 16'b0000000111111111 : node4833;
																assign node4833 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4837 = (inp[7]) ? node4839 : 16'b0000001111111111;
													assign node4839 = (inp[6]) ? 16'b0000000111111111 : node4840;
														assign node4840 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4844 = (inp[12]) ? node4862 : node4845;
												assign node4845 = (inp[6]) ? node4857 : node4846;
													assign node4846 = (inp[8]) ? node4850 : node4847;
														assign node4847 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4850 = (inp[5]) ? node4852 : 16'b0000001111111111;
															assign node4852 = (inp[7]) ? 16'b0000000111111111 : node4853;
																assign node4853 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4857 = (inp[8]) ? 16'b0000000111111111 : node4858;
														assign node4858 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4862 = (inp[8]) ? node4868 : node4863;
													assign node4863 = (inp[5]) ? 16'b0000000111111111 : node4864;
														assign node4864 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4868 = (inp[1]) ? node4870 : 16'b0000000011111111;
														assign node4870 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4873 = (inp[8]) ? node4921 : node4874;
											assign node4874 = (inp[12]) ? node4896 : node4875;
												assign node4875 = (inp[1]) ? node4885 : node4876;
													assign node4876 = (inp[6]) ? node4882 : node4877;
														assign node4877 = (inp[3]) ? 16'b0000001111111111 : node4878;
															assign node4878 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4882 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4885 = (inp[7]) ? node4889 : node4886;
														assign node4886 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4889 = (inp[5]) ? 16'b0000000011111111 : node4890;
															assign node4890 = (inp[3]) ? node4892 : 16'b0000000111111111;
																assign node4892 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4896 = (inp[7]) ? node4912 : node4897;
													assign node4897 = (inp[6]) ? node4901 : node4898;
														assign node4898 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4901 = (inp[1]) ? node4907 : node4902;
															assign node4902 = (inp[5]) ? node4904 : 16'b0000000111111111;
																assign node4904 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node4907 = (inp[5]) ? 16'b0000000011111111 : node4908;
																assign node4908 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4912 = (inp[5]) ? node4916 : node4913;
														assign node4913 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4916 = (inp[6]) ? 16'b0000000001111111 : node4917;
															assign node4917 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4921 = (inp[7]) ? node4935 : node4922;
												assign node4922 = (inp[3]) ? node4926 : node4923;
													assign node4923 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4926 = (inp[6]) ? node4928 : 16'b0000000011111111;
														assign node4928 = (inp[1]) ? 16'b0000000001111111 : node4929;
															assign node4929 = (inp[12]) ? node4931 : 16'b0000000111111111;
																assign node4931 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4935 = (inp[12]) ? node4941 : node4936;
													assign node4936 = (inp[3]) ? 16'b0000000011111111 : node4937;
														assign node4937 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4941 = (inp[5]) ? node4945 : node4942;
														assign node4942 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node4945 = (inp[6]) ? node4947 : 16'b0000000000111111;
															assign node4947 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node4950 = (inp[8]) ? node5094 : node4951;
									assign node4951 = (inp[5]) ? node5011 : node4952;
										assign node4952 = (inp[1]) ? node4984 : node4953;
											assign node4953 = (inp[3]) ? node4965 : node4954;
												assign node4954 = (inp[6]) ? 16'b0000001111111111 : node4955;
													assign node4955 = (inp[15]) ? node4957 : 16'b0000111111111111;
														assign node4957 = (inp[11]) ? 16'b0000011111111111 : node4958;
															assign node4958 = (inp[7]) ? 16'b0000011111111111 : node4959;
																assign node4959 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4965 = (inp[12]) ? node4975 : node4966;
													assign node4966 = (inp[6]) ? node4970 : node4967;
														assign node4967 = (inp[7]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node4970 = (inp[15]) ? node4972 : 16'b0000001111111111;
															assign node4972 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4975 = (inp[15]) ? node4981 : node4976;
														assign node4976 = (inp[11]) ? node4978 : 16'b0000001111111111;
															assign node4978 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4981 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4984 = (inp[7]) ? node4998 : node4985;
												assign node4985 = (inp[6]) ? node4989 : node4986;
													assign node4986 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node4989 = (inp[12]) ? 16'b0000000011111111 : node4990;
														assign node4990 = (inp[11]) ? node4992 : 16'b0000001111111111;
															assign node4992 = (inp[15]) ? 16'b0000000111111111 : node4993;
																assign node4993 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4998 = (inp[6]) ? 16'b0000000011111111 : node4999;
													assign node4999 = (inp[12]) ? node5005 : node5000;
														assign node5000 = (inp[11]) ? 16'b0000000111111111 : node5001;
															assign node5001 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5005 = (inp[11]) ? 16'b0000000011111111 : node5006;
															assign node5006 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5011 = (inp[6]) ? node5043 : node5012;
											assign node5012 = (inp[3]) ? node5022 : node5013;
												assign node5013 = (inp[11]) ? node5017 : node5014;
													assign node5014 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5017 = (inp[12]) ? 16'b0000000011111111 : node5018;
														assign node5018 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5022 = (inp[7]) ? node5030 : node5023;
													assign node5023 = (inp[12]) ? 16'b0000000111111111 : node5024;
														assign node5024 = (inp[1]) ? 16'b0000000111111111 : node5025;
															assign node5025 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5030 = (inp[1]) ? node5036 : node5031;
														assign node5031 = (inp[15]) ? node5033 : 16'b0000000111111111;
															assign node5033 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5036 = (inp[11]) ? 16'b0000000001111111 : node5037;
															assign node5037 = (inp[12]) ? 16'b0000000011111111 : node5038;
																assign node5038 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5043 = (inp[3]) ? node5073 : node5044;
												assign node5044 = (inp[1]) ? node5056 : node5045;
													assign node5045 = (inp[15]) ? node5049 : node5046;
														assign node5046 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5049 = (inp[11]) ? node5051 : 16'b0000000111111111;
															assign node5051 = (inp[7]) ? 16'b0000000011111111 : node5052;
																assign node5052 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5056 = (inp[7]) ? node5066 : node5057;
														assign node5057 = (inp[15]) ? node5061 : node5058;
															assign node5058 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node5061 = (inp[12]) ? 16'b0000000011111111 : node5062;
																assign node5062 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5066 = (inp[12]) ? 16'b0000000001111111 : node5067;
															assign node5067 = (inp[11]) ? node5069 : 16'b0000000111111111;
																assign node5069 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5073 = (inp[15]) ? node5085 : node5074;
													assign node5074 = (inp[1]) ? node5082 : node5075;
														assign node5075 = (inp[11]) ? node5077 : 16'b0000000111111111;
															assign node5077 = (inp[12]) ? 16'b0000000011111111 : node5078;
																assign node5078 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5082 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5085 = (inp[11]) ? node5087 : 16'b0000000011111111;
														assign node5087 = (inp[7]) ? 16'b0000000001111111 : node5088;
															assign node5088 = (inp[12]) ? 16'b0000000001111111 : node5089;
																assign node5089 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5094 = (inp[15]) ? node5158 : node5095;
										assign node5095 = (inp[6]) ? node5123 : node5096;
											assign node5096 = (inp[3]) ? node5118 : node5097;
												assign node5097 = (inp[1]) ? node5109 : node5098;
													assign node5098 = (inp[12]) ? node5106 : node5099;
														assign node5099 = (inp[11]) ? 16'b0000001111111111 : node5100;
															assign node5100 = (inp[5]) ? node5102 : 16'b0000011111111111;
																assign node5102 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5106 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5109 = (inp[11]) ? node5115 : node5110;
														assign node5110 = (inp[7]) ? 16'b0000000111111111 : node5111;
															assign node5111 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5115 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5118 = (inp[5]) ? 16'b0000000011111111 : node5119;
													assign node5119 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5123 = (inp[11]) ? node5135 : node5124;
												assign node5124 = (inp[12]) ? 16'b0000000011111111 : node5125;
													assign node5125 = (inp[7]) ? node5131 : node5126;
														assign node5126 = (inp[5]) ? 16'b0000000111111111 : node5127;
															assign node5127 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5131 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node5135 = (inp[3]) ? node5145 : node5136;
													assign node5136 = (inp[1]) ? node5140 : node5137;
														assign node5137 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5140 = (inp[12]) ? node5142 : 16'b0000000011111111;
															assign node5142 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5145 = (inp[12]) ? node5153 : node5146;
														assign node5146 = (inp[5]) ? 16'b0000000001111111 : node5147;
															assign node5147 = (inp[7]) ? node5149 : 16'b0000000011111111;
																assign node5149 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5153 = (inp[7]) ? node5155 : 16'b0000000001111111;
															assign node5155 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5158 = (inp[7]) ? node5186 : node5159;
											assign node5159 = (inp[6]) ? node5177 : node5160;
												assign node5160 = (inp[1]) ? node5172 : node5161;
													assign node5161 = (inp[11]) ? node5163 : 16'b0000000111111111;
														assign node5163 = (inp[12]) ? node5169 : node5164;
															assign node5164 = (inp[3]) ? node5166 : 16'b0000000111111111;
																assign node5166 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node5169 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5172 = (inp[12]) ? node5174 : 16'b0000000011111111;
														assign node5174 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5177 = (inp[12]) ? node5181 : node5178;
													assign node5178 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5181 = (inp[3]) ? node5183 : 16'b0000000001111111;
														assign node5183 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5186 = (inp[5]) ? node5196 : node5187;
												assign node5187 = (inp[12]) ? node5191 : node5188;
													assign node5188 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5191 = (inp[1]) ? node5193 : 16'b0000000001111111;
														assign node5193 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5196 = (inp[3]) ? node5202 : node5197;
													assign node5197 = (inp[1]) ? 16'b0000000001111111 : node5198;
														assign node5198 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5202 = (inp[12]) ? 16'b0000000000011111 : node5203;
														assign node5203 = (inp[1]) ? node5205 : 16'b0000000000111111;
															assign node5205 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node5209 = (inp[7]) ? node5743 : node5210;
							assign node5210 = (inp[11]) ? node5482 : node5211;
								assign node5211 = (inp[5]) ? node5369 : node5212;
									assign node5212 = (inp[6]) ? node5290 : node5213;
										assign node5213 = (inp[8]) ? node5265 : node5214;
											assign node5214 = (inp[15]) ? node5238 : node5215;
												assign node5215 = (inp[9]) ? node5229 : node5216;
													assign node5216 = (inp[12]) ? node5224 : node5217;
														assign node5217 = (inp[3]) ? 16'b0000111111111111 : node5218;
															assign node5218 = (inp[1]) ? node5220 : 16'b0001111111111111;
																assign node5220 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node5224 = (inp[1]) ? 16'b0000011111111111 : node5225;
															assign node5225 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5229 = (inp[2]) ? node5231 : 16'b0000111111111111;
														assign node5231 = (inp[12]) ? node5233 : 16'b0000011111111111;
															assign node5233 = (inp[1]) ? 16'b0000000111111111 : node5234;
																assign node5234 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5238 = (inp[1]) ? node5252 : node5239;
													assign node5239 = (inp[9]) ? node5245 : node5240;
														assign node5240 = (inp[12]) ? node5242 : 16'b0000011111111111;
															assign node5242 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5245 = (inp[2]) ? 16'b0000011111111111 : node5246;
															assign node5246 = (inp[3]) ? 16'b0000011111111111 : node5247;
																assign node5247 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5252 = (inp[9]) ? node5260 : node5253;
														assign node5253 = (inp[12]) ? 16'b0000001111111111 : node5254;
															assign node5254 = (inp[3]) ? node5256 : 16'b0000011111111111;
																assign node5256 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5260 = (inp[3]) ? node5262 : 16'b0000001111111111;
															assign node5262 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5265 = (inp[9]) ? node5283 : node5266;
												assign node5266 = (inp[1]) ? node5278 : node5267;
													assign node5267 = (inp[2]) ? node5271 : node5268;
														assign node5268 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5271 = (inp[15]) ? node5273 : 16'b0000011111111111;
															assign node5273 = (inp[12]) ? 16'b0000001111111111 : node5274;
																assign node5274 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5278 = (inp[2]) ? 16'b0000001111111111 : node5279;
														assign node5279 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5283 = (inp[2]) ? node5285 : 16'b0000001111111111;
													assign node5285 = (inp[15]) ? node5287 : 16'b0000000111111111;
														assign node5287 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node5290 = (inp[15]) ? node5324 : node5291;
											assign node5291 = (inp[1]) ? node5313 : node5292;
												assign node5292 = (inp[3]) ? node5302 : node5293;
													assign node5293 = (inp[9]) ? 16'b0000011111111111 : node5294;
														assign node5294 = (inp[8]) ? node5296 : 16'b0000111111111111;
															assign node5296 = (inp[2]) ? 16'b0000011111111111 : node5297;
																assign node5297 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5302 = (inp[12]) ? node5310 : node5303;
														assign node5303 = (inp[2]) ? 16'b0000001111111111 : node5304;
															assign node5304 = (inp[9]) ? node5306 : 16'b0000011111111111;
																assign node5306 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5310 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5313 = (inp[8]) ? node5319 : node5314;
													assign node5314 = (inp[3]) ? 16'b0000001111111111 : node5315;
														assign node5315 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5319 = (inp[12]) ? 16'b0000000111111111 : node5320;
														assign node5320 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5324 = (inp[12]) ? node5346 : node5325;
												assign node5325 = (inp[2]) ? node5337 : node5326;
													assign node5326 = (inp[3]) ? node5332 : node5327;
														assign node5327 = (inp[8]) ? node5329 : 16'b0000111111111111;
															assign node5329 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5332 = (inp[8]) ? 16'b0000000111111111 : node5333;
															assign node5333 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5337 = (inp[8]) ? node5343 : node5338;
														assign node5338 = (inp[1]) ? 16'b0000000111111111 : node5339;
															assign node5339 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5343 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5346 = (inp[1]) ? node5358 : node5347;
													assign node5347 = (inp[2]) ? node5355 : node5348;
														assign node5348 = (inp[8]) ? node5350 : 16'b0000001111111111;
															assign node5350 = (inp[3]) ? node5352 : 16'b0000001111111111;
																assign node5352 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5355 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5358 = (inp[2]) ? node5364 : node5359;
														assign node5359 = (inp[8]) ? node5361 : 16'b0000000011111111;
															assign node5361 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5364 = (inp[8]) ? 16'b0000000001111111 : node5365;
															assign node5365 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5369 = (inp[15]) ? node5427 : node5370;
										assign node5370 = (inp[8]) ? node5388 : node5371;
											assign node5371 = (inp[9]) ? node5383 : node5372;
												assign node5372 = (inp[3]) ? node5378 : node5373;
													assign node5373 = (inp[2]) ? 16'b0000011111111111 : node5374;
														assign node5374 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5378 = (inp[2]) ? 16'b0000000111111111 : node5379;
														assign node5379 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5383 = (inp[6]) ? node5385 : 16'b0000001111111111;
													assign node5385 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5388 = (inp[12]) ? node5414 : node5389;
												assign node5389 = (inp[9]) ? node5403 : node5390;
													assign node5390 = (inp[6]) ? node5396 : node5391;
														assign node5391 = (inp[2]) ? 16'b0000001111111111 : node5392;
															assign node5392 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5396 = (inp[1]) ? 16'b0000000111111111 : node5397;
															assign node5397 = (inp[2]) ? node5399 : 16'b0000001111111111;
																assign node5399 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5403 = (inp[3]) ? node5411 : node5404;
														assign node5404 = (inp[2]) ? 16'b0000000111111111 : node5405;
															assign node5405 = (inp[1]) ? node5407 : 16'b0000001111111111;
																assign node5407 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5411 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5414 = (inp[9]) ? node5416 : 16'b0000000111111111;
													assign node5416 = (inp[1]) ? node5422 : node5417;
														assign node5417 = (inp[3]) ? node5419 : 16'b0000000111111111;
															assign node5419 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5422 = (inp[3]) ? node5424 : 16'b0000000001111111;
															assign node5424 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5427 = (inp[6]) ? node5457 : node5428;
											assign node5428 = (inp[1]) ? node5438 : node5429;
												assign node5429 = (inp[2]) ? node5431 : 16'b0000001111111111;
													assign node5431 = (inp[3]) ? 16'b0000000111111111 : node5432;
														assign node5432 = (inp[12]) ? node5434 : 16'b0000001111111111;
															assign node5434 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5438 = (inp[2]) ? node5448 : node5439;
													assign node5439 = (inp[9]) ? node5445 : node5440;
														assign node5440 = (inp[8]) ? 16'b0000000111111111 : node5441;
															assign node5441 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5445 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5448 = (inp[3]) ? node5452 : node5449;
														assign node5449 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5452 = (inp[9]) ? 16'b0000000001111111 : node5453;
															assign node5453 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5457 = (inp[8]) ? node5471 : node5458;
												assign node5458 = (inp[2]) ? node5464 : node5459;
													assign node5459 = (inp[9]) ? node5461 : 16'b0000001111111111;
														assign node5461 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node5464 = (inp[9]) ? node5468 : node5465;
														assign node5465 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5468 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5471 = (inp[2]) ? node5473 : 16'b0000000011111111;
													assign node5473 = (inp[3]) ? node5477 : node5474;
														assign node5474 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5477 = (inp[1]) ? node5479 : 16'b0000000001111111;
															assign node5479 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5482 = (inp[1]) ? node5624 : node5483;
									assign node5483 = (inp[6]) ? node5569 : node5484;
										assign node5484 = (inp[9]) ? node5544 : node5485;
											assign node5485 = (inp[5]) ? node5509 : node5486;
												assign node5486 = (inp[3]) ? node5496 : node5487;
													assign node5487 = (inp[8]) ? 16'b0000011111111111 : node5488;
														assign node5488 = (inp[2]) ? node5490 : 16'b0000111111111111;
															assign node5490 = (inp[12]) ? 16'b0000011111111111 : node5491;
																assign node5491 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5496 = (inp[8]) ? node5504 : node5497;
														assign node5497 = (inp[15]) ? 16'b0000001111111111 : node5498;
															assign node5498 = (inp[12]) ? node5500 : 16'b0000011111111111;
																assign node5500 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5504 = (inp[15]) ? node5506 : 16'b0000001111111111;
															assign node5506 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5509 = (inp[12]) ? node5525 : node5510;
													assign node5510 = (inp[2]) ? node5518 : node5511;
														assign node5511 = (inp[15]) ? node5513 : 16'b0000011111111111;
															assign node5513 = (inp[8]) ? 16'b0000001111111111 : node5514;
																assign node5514 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5518 = (inp[15]) ? 16'b0000000111111111 : node5519;
															assign node5519 = (inp[3]) ? node5521 : 16'b0000001111111111;
																assign node5521 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5525 = (inp[8]) ? node5537 : node5526;
														assign node5526 = (inp[2]) ? node5532 : node5527;
															assign node5527 = (inp[3]) ? node5529 : 16'b0000001111111111;
																assign node5529 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node5532 = (inp[15]) ? node5534 : 16'b0000000111111111;
																assign node5534 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5537 = (inp[3]) ? 16'b0000000011111111 : node5538;
															assign node5538 = (inp[15]) ? node5540 : 16'b0000000111111111;
																assign node5540 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5544 = (inp[15]) ? node5556 : node5545;
												assign node5545 = (inp[2]) ? node5547 : 16'b0000001111111111;
													assign node5547 = (inp[12]) ? node5553 : node5548;
														assign node5548 = (inp[5]) ? 16'b0000000111111111 : node5549;
															assign node5549 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5553 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5556 = (inp[8]) ? node5566 : node5557;
													assign node5557 = (inp[12]) ? node5561 : node5558;
														assign node5558 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5561 = (inp[3]) ? node5563 : 16'b0000000111111111;
															assign node5563 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5566 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5569 = (inp[8]) ? node5601 : node5570;
											assign node5570 = (inp[15]) ? node5588 : node5571;
												assign node5571 = (inp[5]) ? node5583 : node5572;
													assign node5572 = (inp[9]) ? node5580 : node5573;
														assign node5573 = (inp[3]) ? node5575 : 16'b0000011111111111;
															assign node5575 = (inp[2]) ? 16'b0000001111111111 : node5576;
																assign node5576 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5580 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5583 = (inp[3]) ? 16'b0000000011111111 : node5584;
														assign node5584 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5588 = (inp[5]) ? node5594 : node5589;
													assign node5589 = (inp[3]) ? node5591 : 16'b0000000111111111;
														assign node5591 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5594 = (inp[9]) ? node5598 : node5595;
														assign node5595 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5598 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node5601 = (inp[2]) ? node5607 : node5602;
												assign node5602 = (inp[3]) ? 16'b0000000011111111 : node5603;
													assign node5603 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node5607 = (inp[5]) ? node5617 : node5608;
													assign node5608 = (inp[3]) ? node5610 : 16'b0000000011111111;
														assign node5610 = (inp[9]) ? node5612 : 16'b0000000011111111;
															assign node5612 = (inp[15]) ? 16'b0000000001111111 : node5613;
																assign node5613 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5617 = (inp[12]) ? node5619 : 16'b0000000011111111;
														assign node5619 = (inp[9]) ? 16'b0000000000111111 : node5620;
															assign node5620 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5624 = (inp[2]) ? node5682 : node5625;
										assign node5625 = (inp[6]) ? node5655 : node5626;
											assign node5626 = (inp[5]) ? node5638 : node5627;
												assign node5627 = (inp[8]) ? node5629 : 16'b0000001111111111;
													assign node5629 = (inp[12]) ? node5635 : node5630;
														assign node5630 = (inp[15]) ? node5632 : 16'b0000001111111111;
															assign node5632 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5635 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5638 = (inp[15]) ? node5646 : node5639;
													assign node5639 = (inp[9]) ? node5641 : 16'b0000001111111111;
														assign node5641 = (inp[12]) ? node5643 : 16'b0000000111111111;
															assign node5643 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node5646 = (inp[12]) ? node5650 : node5647;
														assign node5647 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5650 = (inp[9]) ? node5652 : 16'b0000000011111111;
															assign node5652 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5655 = (inp[12]) ? node5673 : node5656;
												assign node5656 = (inp[5]) ? node5664 : node5657;
													assign node5657 = (inp[9]) ? node5661 : node5658;
														assign node5658 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5661 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5664 = (inp[8]) ? 16'b0000000011111111 : node5665;
														assign node5665 = (inp[3]) ? node5667 : 16'b0000000111111111;
															assign node5667 = (inp[9]) ? 16'b0000000011111111 : node5668;
																assign node5668 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5673 = (inp[9]) ? node5677 : node5674;
													assign node5674 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5677 = (inp[3]) ? 16'b0000000001111111 : node5678;
														assign node5678 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5682 = (inp[9]) ? node5708 : node5683;
											assign node5683 = (inp[15]) ? node5697 : node5684;
												assign node5684 = (inp[12]) ? node5690 : node5685;
													assign node5685 = (inp[3]) ? node5687 : 16'b0000000111111111;
														assign node5687 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node5690 = (inp[6]) ? node5694 : node5691;
														assign node5691 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5694 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node5697 = (inp[6]) ? node5703 : node5698;
													assign node5698 = (inp[12]) ? node5700 : 16'b0000000011111111;
														assign node5700 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5703 = (inp[3]) ? 16'b0000000001111111 : node5704;
														assign node5704 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5708 = (inp[15]) ? node5732 : node5709;
												assign node5709 = (inp[5]) ? node5719 : node5710;
													assign node5710 = (inp[12]) ? node5714 : node5711;
														assign node5711 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5714 = (inp[3]) ? node5716 : 16'b0000000011111111;
															assign node5716 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5719 = (inp[3]) ? node5723 : node5720;
														assign node5720 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5723 = (inp[8]) ? node5727 : node5724;
															assign node5724 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node5727 = (inp[12]) ? 16'b0000000000111111 : node5728;
																assign node5728 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5732 = (inp[3]) ? node5738 : node5733;
													assign node5733 = (inp[5]) ? node5735 : 16'b0000000011111111;
														assign node5735 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5738 = (inp[5]) ? node5740 : 16'b0000000000111111;
														assign node5740 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node5743 = (inp[6]) ? node6025 : node5744;
								assign node5744 = (inp[11]) ? node5864 : node5745;
									assign node5745 = (inp[2]) ? node5815 : node5746;
										assign node5746 = (inp[1]) ? node5770 : node5747;
											assign node5747 = (inp[12]) ? node5761 : node5748;
												assign node5748 = (inp[15]) ? 16'b0000001111111111 : node5749;
													assign node5749 = (inp[5]) ? node5753 : node5750;
														assign node5750 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5753 = (inp[3]) ? 16'b0000001111111111 : node5754;
															assign node5754 = (inp[8]) ? node5756 : 16'b0000011111111111;
																assign node5756 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5761 = (inp[8]) ? node5765 : node5762;
													assign node5762 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5765 = (inp[5]) ? 16'b0000000111111111 : node5766;
														assign node5766 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5770 = (inp[8]) ? node5794 : node5771;
												assign node5771 = (inp[15]) ? node5789 : node5772;
													assign node5772 = (inp[3]) ? node5780 : node5773;
														assign node5773 = (inp[9]) ? node5775 : 16'b0000011111111111;
															assign node5775 = (inp[12]) ? 16'b0000001111111111 : node5776;
																assign node5776 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5780 = (inp[5]) ? node5786 : node5781;
															assign node5781 = (inp[12]) ? 16'b0000001111111111 : node5782;
																assign node5782 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node5786 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node5789 = (inp[12]) ? 16'b0000000011111111 : node5790;
														assign node5790 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5794 = (inp[9]) ? node5806 : node5795;
													assign node5795 = (inp[5]) ? node5799 : node5796;
														assign node5796 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5799 = (inp[12]) ? 16'b0000000011111111 : node5800;
															assign node5800 = (inp[3]) ? node5802 : 16'b0000000111111111;
																assign node5802 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5806 = (inp[15]) ? node5810 : node5807;
														assign node5807 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5810 = (inp[5]) ? node5812 : 16'b0000000011111111;
															assign node5812 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5815 = (inp[15]) ? node5839 : node5816;
											assign node5816 = (inp[1]) ? node5830 : node5817;
												assign node5817 = (inp[12]) ? node5823 : node5818;
													assign node5818 = (inp[5]) ? node5820 : 16'b0000001111111111;
														assign node5820 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5823 = (inp[3]) ? node5825 : 16'b0000000111111111;
														assign node5825 = (inp[5]) ? 16'b0000000011111111 : node5826;
															assign node5826 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node5830 = (inp[3]) ? node5834 : node5831;
													assign node5831 = (inp[8]) ? 16'b0000000011111111 : 16'b0000011111111111;
													assign node5834 = (inp[8]) ? 16'b0000000011111111 : node5835;
														assign node5835 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5839 = (inp[8]) ? node5853 : node5840;
												assign node5840 = (inp[12]) ? node5848 : node5841;
													assign node5841 = (inp[1]) ? node5843 : 16'b0000000111111111;
														assign node5843 = (inp[3]) ? 16'b0000000011111111 : node5844;
															assign node5844 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5848 = (inp[1]) ? node5850 : 16'b0000000011111111;
														assign node5850 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5853 = (inp[9]) ? node5855 : 16'b0000000011111111;
													assign node5855 = (inp[12]) ? node5861 : node5856;
														assign node5856 = (inp[1]) ? 16'b0000000001111111 : node5857;
															assign node5857 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5861 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
									assign node5864 = (inp[9]) ? node5938 : node5865;
										assign node5865 = (inp[5]) ? node5893 : node5866;
											assign node5866 = (inp[1]) ? node5882 : node5867;
												assign node5867 = (inp[15]) ? node5875 : node5868;
													assign node5868 = (inp[2]) ? node5872 : node5869;
														assign node5869 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5872 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5875 = (inp[12]) ? node5877 : 16'b0000001111111111;
														assign node5877 = (inp[2]) ? node5879 : 16'b0000000111111111;
															assign node5879 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5882 = (inp[3]) ? node5888 : node5883;
													assign node5883 = (inp[15]) ? node5885 : 16'b0000000111111111;
														assign node5885 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5888 = (inp[2]) ? 16'b0000000011111111 : node5889;
														assign node5889 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5893 = (inp[2]) ? node5917 : node5894;
												assign node5894 = (inp[3]) ? node5902 : node5895;
													assign node5895 = (inp[12]) ? node5899 : node5896;
														assign node5896 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5899 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node5902 = (inp[15]) ? 16'b0000000011111111 : node5903;
														assign node5903 = (inp[12]) ? node5909 : node5904;
															assign node5904 = (inp[1]) ? node5906 : 16'b0000000111111111;
																assign node5906 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node5909 = (inp[1]) ? node5913 : node5910;
																assign node5910 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node5913 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5917 = (inp[8]) ? node5923 : node5918;
													assign node5918 = (inp[3]) ? 16'b0000000011111111 : node5919;
														assign node5919 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5923 = (inp[3]) ? node5933 : node5924;
														assign node5924 = (inp[15]) ? node5928 : node5925;
															assign node5925 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node5928 = (inp[12]) ? 16'b0000000001111111 : node5929;
																assign node5929 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5933 = (inp[12]) ? node5935 : 16'b0000000001111111;
															assign node5935 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5938 = (inp[3]) ? node5978 : node5939;
											assign node5939 = (inp[1]) ? node5959 : node5940;
												assign node5940 = (inp[8]) ? node5952 : node5941;
													assign node5941 = (inp[5]) ? node5947 : node5942;
														assign node5942 = (inp[2]) ? 16'b0000000111111111 : node5943;
															assign node5943 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5947 = (inp[15]) ? node5949 : 16'b0000000111111111;
															assign node5949 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5952 = (inp[15]) ? node5956 : node5953;
														assign node5953 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5956 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5959 = (inp[12]) ? node5971 : node5960;
													assign node5960 = (inp[8]) ? node5964 : node5961;
														assign node5961 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5964 = (inp[15]) ? node5966 : 16'b0000000011111111;
															assign node5966 = (inp[5]) ? 16'b0000000001111111 : node5967;
																assign node5967 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5971 = (inp[5]) ? 16'b0000000000111111 : node5972;
														assign node5972 = (inp[15]) ? node5974 : 16'b0000000001111111;
															assign node5974 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5978 = (inp[2]) ? node6002 : node5979;
												assign node5979 = (inp[12]) ? node5995 : node5980;
													assign node5980 = (inp[5]) ? node5988 : node5981;
														assign node5981 = (inp[1]) ? node5983 : 16'b0000000011111111;
															assign node5983 = (inp[8]) ? node5985 : 16'b0000000011111111;
																assign node5985 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5988 = (inp[8]) ? 16'b0000000001111111 : node5989;
															assign node5989 = (inp[15]) ? node5991 : 16'b0000000011111111;
																assign node5991 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5995 = (inp[8]) ? 16'b0000000000111111 : node5996;
														assign node5996 = (inp[5]) ? 16'b0000000001111111 : node5997;
															assign node5997 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6002 = (inp[1]) ? node6014 : node6003;
													assign node6003 = (inp[15]) ? node6009 : node6004;
														assign node6004 = (inp[5]) ? node6006 : 16'b0000000011111111;
															assign node6006 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6009 = (inp[8]) ? node6011 : 16'b0000000000111111;
															assign node6011 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node6014 = (inp[12]) ? node6020 : node6015;
														assign node6015 = (inp[5]) ? node6017 : 16'b0000000000111111;
															assign node6017 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node6020 = (inp[15]) ? node6022 : 16'b0000000000011111;
															assign node6022 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node6025 = (inp[5]) ? node6129 : node6026;
									assign node6026 = (inp[8]) ? node6074 : node6027;
										assign node6027 = (inp[11]) ? node6043 : node6028;
											assign node6028 = (inp[15]) ? node6034 : node6029;
												assign node6029 = (inp[12]) ? node6031 : 16'b0000001111111111;
													assign node6031 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6034 = (inp[12]) ? node6036 : 16'b0000000111111111;
													assign node6036 = (inp[9]) ? 16'b0000000011111111 : node6037;
														assign node6037 = (inp[2]) ? node6039 : 16'b0000000111111111;
															assign node6039 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6043 = (inp[15]) ? node6055 : node6044;
												assign node6044 = (inp[12]) ? node6050 : node6045;
													assign node6045 = (inp[3]) ? 16'b0000000111111111 : node6046;
														assign node6046 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6050 = (inp[3]) ? node6052 : 16'b0000000111111111;
														assign node6052 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node6055 = (inp[9]) ? node6063 : node6056;
													assign node6056 = (inp[12]) ? 16'b0000000011111111 : node6057;
														assign node6057 = (inp[3]) ? node6059 : 16'b0000001111111111;
															assign node6059 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6063 = (inp[2]) ? 16'b0000000000111111 : node6064;
														assign node6064 = (inp[3]) ? 16'b0000000001111111 : node6065;
															assign node6065 = (inp[1]) ? node6069 : node6066;
																assign node6066 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node6069 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6074 = (inp[12]) ? node6094 : node6075;
											assign node6075 = (inp[11]) ? node6091 : node6076;
												assign node6076 = (inp[9]) ? node6082 : node6077;
													assign node6077 = (inp[3]) ? node6079 : 16'b0000000111111111;
														assign node6079 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6082 = (inp[15]) ? node6088 : node6083;
														assign node6083 = (inp[2]) ? 16'b0000000011111111 : node6084;
															assign node6084 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6088 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node6091 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6094 = (inp[15]) ? node6116 : node6095;
												assign node6095 = (inp[3]) ? node6105 : node6096;
													assign node6096 = (inp[2]) ? node6102 : node6097;
														assign node6097 = (inp[1]) ? node6099 : 16'b0000000111111111;
															assign node6099 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6102 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6105 = (inp[9]) ? node6111 : node6106;
														assign node6106 = (inp[1]) ? 16'b0000000001111111 : node6107;
															assign node6107 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node6111 = (inp[11]) ? 16'b0000000000111111 : node6112;
															assign node6112 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6116 = (inp[9]) ? node6122 : node6117;
													assign node6117 = (inp[11]) ? node6119 : 16'b0000000001111111;
														assign node6119 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6122 = (inp[3]) ? node6126 : node6123;
														assign node6123 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6126 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node6129 = (inp[15]) ? node6211 : node6130;
										assign node6130 = (inp[1]) ? node6184 : node6131;
											assign node6131 = (inp[9]) ? node6155 : node6132;
												assign node6132 = (inp[11]) ? node6144 : node6133;
													assign node6133 = (inp[12]) ? node6137 : node6134;
														assign node6134 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6137 = (inp[2]) ? 16'b0000000011111111 : node6138;
															assign node6138 = (inp[8]) ? node6140 : 16'b0000000111111111;
																assign node6140 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6144 = (inp[12]) ? node6152 : node6145;
														assign node6145 = (inp[2]) ? 16'b0000000011111111 : node6146;
															assign node6146 = (inp[3]) ? node6148 : 16'b0000000111111111;
																assign node6148 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6152 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6155 = (inp[11]) ? node6169 : node6156;
													assign node6156 = (inp[12]) ? node6164 : node6157;
														assign node6157 = (inp[3]) ? 16'b0000000011111111 : node6158;
															assign node6158 = (inp[2]) ? node6160 : 16'b0000000111111111;
																assign node6160 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6164 = (inp[2]) ? 16'b0000000001111111 : node6165;
															assign node6165 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6169 = (inp[8]) ? node6175 : node6170;
														assign node6170 = (inp[2]) ? node6172 : 16'b0000000011111111;
															assign node6172 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6175 = (inp[3]) ? node6177 : 16'b0000000001111111;
															assign node6177 = (inp[2]) ? node6181 : node6178;
																assign node6178 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
																assign node6181 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node6184 = (inp[12]) ? node6196 : node6185;
												assign node6185 = (inp[3]) ? node6191 : node6186;
													assign node6186 = (inp[11]) ? node6188 : 16'b0000000111111111;
														assign node6188 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6191 = (inp[8]) ? 16'b0000000001111111 : node6192;
														assign node6192 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6196 = (inp[3]) ? node6206 : node6197;
													assign node6197 = (inp[9]) ? node6203 : node6198;
														assign node6198 = (inp[8]) ? node6200 : 16'b0000000011111111;
															assign node6200 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6203 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node6206 = (inp[9]) ? node6208 : 16'b0000000000111111;
														assign node6208 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node6211 = (inp[8]) ? node6253 : node6212;
											assign node6212 = (inp[12]) ? node6234 : node6213;
												assign node6213 = (inp[11]) ? node6225 : node6214;
													assign node6214 = (inp[2]) ? node6218 : node6215;
														assign node6215 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6218 = (inp[9]) ? 16'b0000000001111111 : node6219;
															assign node6219 = (inp[3]) ? 16'b0000000011111111 : node6220;
																assign node6220 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6225 = (inp[2]) ? node6229 : node6226;
														assign node6226 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6229 = (inp[9]) ? node6231 : 16'b0000000001111111;
															assign node6231 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node6234 = (inp[2]) ? node6244 : node6235;
													assign node6235 = (inp[1]) ? node6237 : 16'b0000000001111111;
														assign node6237 = (inp[3]) ? node6239 : 16'b0000000001111111;
															assign node6239 = (inp[9]) ? 16'b0000000000111111 : node6240;
																assign node6240 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6244 = (inp[9]) ? node6248 : node6245;
														assign node6245 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6248 = (inp[1]) ? node6250 : 16'b0000000000011111;
															assign node6250 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node6253 = (inp[2]) ? node6265 : node6254;
												assign node6254 = (inp[9]) ? 16'b0000000000111111 : node6255;
													assign node6255 = (inp[11]) ? node6257 : 16'b0000000001111111;
														assign node6257 = (inp[12]) ? 16'b0000000000111111 : node6258;
															assign node6258 = (inp[1]) ? node6260 : 16'b0000000001111111;
																assign node6260 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6265 = (inp[3]) ? node6273 : node6266;
													assign node6266 = (inp[1]) ? node6268 : 16'b0000000000111111;
														assign node6268 = (inp[11]) ? 16'b0000000000011111 : node6269;
															assign node6269 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6273 = (inp[11]) ? 16'b0000000000001111 : node6274;
														assign node6274 = (inp[9]) ? 16'b0000000000011111 : node6275;
															assign node6275 = (inp[1]) ? node6277 : 16'b0000000000111111;
																assign node6277 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node6282 = (inp[2]) ? node7282 : node6283;
						assign node6283 = (inp[3]) ? node6749 : node6284;
							assign node6284 = (inp[9]) ? node6508 : node6285;
								assign node6285 = (inp[15]) ? node6395 : node6286;
									assign node6286 = (inp[6]) ? node6336 : node6287;
										assign node6287 = (inp[13]) ? node6319 : node6288;
											assign node6288 = (inp[7]) ? node6304 : node6289;
												assign node6289 = (inp[8]) ? node6297 : node6290;
													assign node6290 = (inp[5]) ? 16'b0000111111111111 : node6291;
														assign node6291 = (inp[12]) ? 16'b0000111111111111 : node6292;
															assign node6292 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node6297 = (inp[1]) ? node6301 : node6298;
														assign node6298 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6301 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6304 = (inp[12]) ? node6310 : node6305;
													assign node6305 = (inp[8]) ? 16'b0000011111111111 : node6306;
														assign node6306 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6310 = (inp[8]) ? 16'b0000000011111111 : node6311;
														assign node6311 = (inp[5]) ? node6313 : 16'b0000011111111111;
															assign node6313 = (inp[11]) ? node6315 : 16'b0000001111111111;
																assign node6315 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6319 = (inp[12]) ? node6323 : node6320;
												assign node6320 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6323 = (inp[5]) ? node6329 : node6324;
													assign node6324 = (inp[8]) ? 16'b0000001111111111 : node6325;
														assign node6325 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6329 = (inp[1]) ? node6333 : node6330;
														assign node6330 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6333 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6336 = (inp[1]) ? node6364 : node6337;
											assign node6337 = (inp[11]) ? node6359 : node6338;
												assign node6338 = (inp[12]) ? node6346 : node6339;
													assign node6339 = (inp[5]) ? 16'b0000011111111111 : node6340;
														assign node6340 = (inp[13]) ? 16'b0000011111111111 : node6341;
															assign node6341 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6346 = (inp[13]) ? node6352 : node6347;
														assign node6347 = (inp[8]) ? node6349 : 16'b0000011111111111;
															assign node6349 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6352 = (inp[5]) ? node6354 : 16'b0000001111111111;
															assign node6354 = (inp[8]) ? 16'b0000000111111111 : node6355;
																assign node6355 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6359 = (inp[8]) ? 16'b0000000111111111 : node6360;
													assign node6360 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node6364 = (inp[8]) ? node6376 : node6365;
												assign node6365 = (inp[5]) ? node6371 : node6366;
													assign node6366 = (inp[7]) ? node6368 : 16'b0000001111111111;
														assign node6368 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6371 = (inp[11]) ? 16'b0000000111111111 : node6372;
														assign node6372 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6376 = (inp[13]) ? node6392 : node6377;
													assign node6377 = (inp[5]) ? node6389 : node6378;
														assign node6378 = (inp[12]) ? node6384 : node6379;
															assign node6379 = (inp[11]) ? node6381 : 16'b0000001111111111;
																assign node6381 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node6384 = (inp[7]) ? 16'b0000000111111111 : node6385;
																assign node6385 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6389 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6392 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node6395 = (inp[11]) ? node6459 : node6396;
										assign node6396 = (inp[13]) ? node6432 : node6397;
											assign node6397 = (inp[12]) ? node6415 : node6398;
												assign node6398 = (inp[6]) ? node6408 : node6399;
													assign node6399 = (inp[7]) ? 16'b0000011111111111 : node6400;
														assign node6400 = (inp[5]) ? node6404 : node6401;
															assign node6401 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node6404 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6408 = (inp[8]) ? 16'b0000000111111111 : node6409;
														assign node6409 = (inp[5]) ? node6411 : 16'b0000011111111111;
															assign node6411 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6415 = (inp[6]) ? node6425 : node6416;
													assign node6416 = (inp[7]) ? node6422 : node6417;
														assign node6417 = (inp[5]) ? 16'b0000001111111111 : node6418;
															assign node6418 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6422 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6425 = (inp[5]) ? node6429 : node6426;
														assign node6426 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node6429 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6432 = (inp[1]) ? node6450 : node6433;
												assign node6433 = (inp[6]) ? node6441 : node6434;
													assign node6434 = (inp[12]) ? 16'b0000000111111111 : node6435;
														assign node6435 = (inp[7]) ? 16'b0000001111111111 : node6436;
															assign node6436 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node6441 = (inp[7]) ? node6447 : node6442;
														assign node6442 = (inp[5]) ? 16'b0000000111111111 : node6443;
															assign node6443 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6447 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6450 = (inp[5]) ? node6452 : 16'b0000000111111111;
													assign node6452 = (inp[7]) ? node6456 : node6453;
														assign node6453 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6456 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node6459 = (inp[1]) ? node6481 : node6460;
											assign node6460 = (inp[6]) ? node6470 : node6461;
												assign node6461 = (inp[8]) ? 16'b0000000111111111 : node6462;
													assign node6462 = (inp[7]) ? node6466 : node6463;
														assign node6463 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6466 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6470 = (inp[12]) ? node6474 : node6471;
													assign node6471 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6474 = (inp[5]) ? 16'b0000000011111111 : node6475;
														assign node6475 = (inp[8]) ? node6477 : 16'b0000000111111111;
															assign node6477 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6481 = (inp[8]) ? node6495 : node6482;
												assign node6482 = (inp[5]) ? node6488 : node6483;
													assign node6483 = (inp[12]) ? node6485 : 16'b0000001111111111;
														assign node6485 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6488 = (inp[13]) ? node6492 : node6489;
														assign node6489 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6492 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6495 = (inp[13]) ? node6501 : node6496;
													assign node6496 = (inp[12]) ? 16'b0000000001111111 : node6497;
														assign node6497 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6501 = (inp[7]) ? node6503 : 16'b0000000001111111;
														assign node6503 = (inp[6]) ? node6505 : 16'b0000000001111111;
															assign node6505 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node6508 = (inp[15]) ? node6632 : node6509;
									assign node6509 = (inp[5]) ? node6585 : node6510;
										assign node6510 = (inp[1]) ? node6548 : node6511;
											assign node6511 = (inp[13]) ? node6533 : node6512;
												assign node6512 = (inp[11]) ? node6524 : node6513;
													assign node6513 = (inp[8]) ? node6517 : node6514;
														assign node6514 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6517 = (inp[7]) ? node6519 : 16'b0000011111111111;
															assign node6519 = (inp[12]) ? 16'b0000001111111111 : node6520;
																assign node6520 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6524 = (inp[7]) ? node6530 : node6525;
														assign node6525 = (inp[12]) ? 16'b0000001111111111 : node6526;
															assign node6526 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6530 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6533 = (inp[8]) ? node6543 : node6534;
													assign node6534 = (inp[11]) ? node6540 : node6535;
														assign node6535 = (inp[12]) ? node6537 : 16'b0000011111111111;
															assign node6537 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6540 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6543 = (inp[7]) ? node6545 : 16'b0000000111111111;
														assign node6545 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6548 = (inp[8]) ? node6562 : node6549;
												assign node6549 = (inp[7]) ? node6551 : 16'b0000001111111111;
													assign node6551 = (inp[13]) ? node6559 : node6552;
														assign node6552 = (inp[11]) ? node6554 : 16'b0000001111111111;
															assign node6554 = (inp[12]) ? 16'b0000000011111111 : node6555;
																assign node6555 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6559 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6562 = (inp[11]) ? node6572 : node6563;
													assign node6563 = (inp[13]) ? node6567 : node6564;
														assign node6564 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6567 = (inp[7]) ? node6569 : 16'b0000000111111111;
															assign node6569 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6572 = (inp[13]) ? node6582 : node6573;
														assign node6573 = (inp[7]) ? node6577 : node6574;
															assign node6574 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node6577 = (inp[6]) ? 16'b0000000011111111 : node6578;
																assign node6578 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6582 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6585 = (inp[1]) ? node6617 : node6586;
											assign node6586 = (inp[12]) ? node6606 : node6587;
												assign node6587 = (inp[11]) ? node6599 : node6588;
													assign node6588 = (inp[6]) ? node6590 : 16'b0000001111111111;
														assign node6590 = (inp[13]) ? 16'b0000000111111111 : node6591;
															assign node6591 = (inp[8]) ? node6595 : node6592;
																assign node6592 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
																assign node6595 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6599 = (inp[6]) ? node6601 : 16'b0000000111111111;
														assign node6601 = (inp[8]) ? 16'b0000000011111111 : node6602;
															assign node6602 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6606 = (inp[6]) ? node6608 : 16'b0000000111111111;
													assign node6608 = (inp[7]) ? node6614 : node6609;
														assign node6609 = (inp[11]) ? 16'b0000000011111111 : node6610;
															assign node6610 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6614 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6617 = (inp[6]) ? node6625 : node6618;
												assign node6618 = (inp[13]) ? 16'b0000000011111111 : node6619;
													assign node6619 = (inp[11]) ? 16'b0000000011111111 : node6620;
														assign node6620 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6625 = (inp[8]) ? 16'b0000000001111111 : node6626;
													assign node6626 = (inp[7]) ? 16'b0000000001111111 : node6627;
														assign node6627 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node6632 = (inp[6]) ? node6704 : node6633;
										assign node6633 = (inp[8]) ? node6673 : node6634;
											assign node6634 = (inp[5]) ? node6646 : node6635;
												assign node6635 = (inp[7]) ? node6641 : node6636;
													assign node6636 = (inp[11]) ? 16'b0000001111111111 : node6637;
														assign node6637 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6641 = (inp[11]) ? 16'b0000000111111111 : node6642;
														assign node6642 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6646 = (inp[13]) ? node6668 : node6647;
													assign node6647 = (inp[7]) ? node6655 : node6648;
														assign node6648 = (inp[11]) ? 16'b0000000111111111 : node6649;
															assign node6649 = (inp[12]) ? node6651 : 16'b0000001111111111;
																assign node6651 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6655 = (inp[1]) ? node6663 : node6656;
															assign node6656 = (inp[12]) ? node6660 : node6657;
																assign node6657 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
																assign node6660 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node6663 = (inp[11]) ? 16'b0000000011111111 : node6664;
																assign node6664 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6668 = (inp[11]) ? 16'b0000000001111111 : node6669;
														assign node6669 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node6673 = (inp[11]) ? node6687 : node6674;
												assign node6674 = (inp[5]) ? node6678 : node6675;
													assign node6675 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6678 = (inp[1]) ? node6684 : node6679;
														assign node6679 = (inp[12]) ? node6681 : 16'b0000000111111111;
															assign node6681 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6684 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6687 = (inp[12]) ? node6697 : node6688;
													assign node6688 = (inp[1]) ? node6692 : node6689;
														assign node6689 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node6692 = (inp[5]) ? 16'b0000000001111111 : node6693;
															assign node6693 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6697 = (inp[5]) ? node6701 : node6698;
														assign node6698 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6701 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6704 = (inp[12]) ? node6720 : node6705;
											assign node6705 = (inp[5]) ? node6717 : node6706;
												assign node6706 = (inp[13]) ? node6712 : node6707;
													assign node6707 = (inp[1]) ? node6709 : 16'b0000000111111111;
														assign node6709 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6712 = (inp[7]) ? 16'b0000000011111111 : node6713;
														assign node6713 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6717 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6720 = (inp[11]) ? node6738 : node6721;
												assign node6721 = (inp[7]) ? node6729 : node6722;
													assign node6722 = (inp[5]) ? node6724 : 16'b0000000111111111;
														assign node6724 = (inp[1]) ? node6726 : 16'b0000000011111111;
															assign node6726 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6729 = (inp[5]) ? node6733 : node6730;
														assign node6730 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6733 = (inp[1]) ? node6735 : 16'b0000000001111111;
															assign node6735 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6738 = (inp[8]) ? 16'b0000000000111111 : node6739;
													assign node6739 = (inp[13]) ? node6745 : node6740;
														assign node6740 = (inp[5]) ? 16'b0000000001111111 : node6741;
															assign node6741 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6745 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node6749 = (inp[1]) ? node7019 : node6750;
								assign node6750 = (inp[5]) ? node6878 : node6751;
									assign node6751 = (inp[7]) ? node6825 : node6752;
										assign node6752 = (inp[8]) ? node6790 : node6753;
											assign node6753 = (inp[11]) ? node6777 : node6754;
												assign node6754 = (inp[9]) ? node6768 : node6755;
													assign node6755 = (inp[13]) ? node6761 : node6756;
														assign node6756 = (inp[12]) ? node6758 : 16'b0000111111111111;
															assign node6758 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6761 = (inp[12]) ? 16'b0000001111111111 : node6762;
															assign node6762 = (inp[15]) ? 16'b0000011111111111 : node6763;
																assign node6763 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6768 = (inp[6]) ? node6774 : node6769;
														assign node6769 = (inp[15]) ? 16'b0000001111111111 : node6770;
															assign node6770 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6774 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6777 = (inp[12]) ? node6783 : node6778;
													assign node6778 = (inp[13]) ? node6780 : 16'b0000011111111111;
														assign node6780 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6783 = (inp[15]) ? node6787 : node6784;
														assign node6784 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6787 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6790 = (inp[6]) ? node6810 : node6791;
												assign node6791 = (inp[11]) ? node6803 : node6792;
													assign node6792 = (inp[13]) ? node6796 : node6793;
														assign node6793 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6796 = (inp[12]) ? node6798 : 16'b0000001111111111;
															assign node6798 = (inp[9]) ? 16'b0000000111111111 : node6799;
																assign node6799 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6803 = (inp[13]) ? node6807 : node6804;
														assign node6804 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6807 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6810 = (inp[13]) ? node6818 : node6811;
													assign node6811 = (inp[15]) ? 16'b0000000111111111 : node6812;
														assign node6812 = (inp[9]) ? 16'b0000000111111111 : node6813;
															assign node6813 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6818 = (inp[11]) ? node6822 : node6819;
														assign node6819 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6822 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6825 = (inp[6]) ? node6853 : node6826;
											assign node6826 = (inp[11]) ? node6844 : node6827;
												assign node6827 = (inp[8]) ? node6837 : node6828;
													assign node6828 = (inp[12]) ? node6830 : 16'b0000011111111111;
														assign node6830 = (inp[15]) ? 16'b0000000111111111 : node6831;
															assign node6831 = (inp[9]) ? 16'b0000001111111111 : node6832;
																assign node6832 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6837 = (inp[15]) ? node6841 : node6838;
														assign node6838 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6841 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6844 = (inp[9]) ? node6846 : 16'b0000000111111111;
													assign node6846 = (inp[13]) ? 16'b0000000001111111 : node6847;
														assign node6847 = (inp[15]) ? 16'b0000000011111111 : node6848;
															assign node6848 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node6853 = (inp[12]) ? node6871 : node6854;
												assign node6854 = (inp[15]) ? node6858 : node6855;
													assign node6855 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6858 = (inp[9]) ? node6866 : node6859;
														assign node6859 = (inp[13]) ? node6861 : 16'b0000000111111111;
															assign node6861 = (inp[8]) ? 16'b0000000011111111 : node6862;
																assign node6862 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6866 = (inp[13]) ? node6868 : 16'b0000000011111111;
															assign node6868 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6871 = (inp[9]) ? 16'b0000000000111111 : node6872;
													assign node6872 = (inp[13]) ? node6874 : 16'b0000000111111111;
														assign node6874 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node6878 = (inp[15]) ? node6948 : node6879;
										assign node6879 = (inp[9]) ? node6917 : node6880;
											assign node6880 = (inp[12]) ? node6894 : node6881;
												assign node6881 = (inp[11]) ? node6887 : node6882;
													assign node6882 = (inp[7]) ? 16'b0000000111111111 : node6883;
														assign node6883 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6887 = (inp[6]) ? node6891 : node6888;
														assign node6888 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6891 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6894 = (inp[6]) ? node6910 : node6895;
													assign node6895 = (inp[11]) ? node6899 : node6896;
														assign node6896 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6899 = (inp[13]) ? node6905 : node6900;
															assign node6900 = (inp[8]) ? node6902 : 16'b0000000111111111;
																assign node6902 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node6905 = (inp[8]) ? 16'b0000000011111111 : node6906;
																assign node6906 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6910 = (inp[7]) ? node6914 : node6911;
														assign node6911 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6914 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6917 = (inp[11]) ? node6941 : node6918;
												assign node6918 = (inp[8]) ? node6930 : node6919;
													assign node6919 = (inp[13]) ? node6927 : node6920;
														assign node6920 = (inp[7]) ? node6922 : 16'b0000001111111111;
															assign node6922 = (inp[6]) ? 16'b0000000111111111 : node6923;
																assign node6923 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6927 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6930 = (inp[6]) ? node6934 : node6931;
														assign node6931 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node6934 = (inp[7]) ? node6936 : 16'b0000000011111111;
															assign node6936 = (inp[12]) ? 16'b0000000001111111 : node6937;
																assign node6937 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6941 = (inp[12]) ? 16'b0000000001111111 : node6942;
													assign node6942 = (inp[8]) ? 16'b0000000001111111 : node6943;
														assign node6943 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6948 = (inp[7]) ? node6982 : node6949;
											assign node6949 = (inp[8]) ? node6973 : node6950;
												assign node6950 = (inp[11]) ? node6960 : node6951;
													assign node6951 = (inp[13]) ? node6955 : node6952;
														assign node6952 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node6955 = (inp[12]) ? node6957 : 16'b0000000111111111;
															assign node6957 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6960 = (inp[6]) ? node6968 : node6961;
														assign node6961 = (inp[12]) ? node6963 : 16'b0000000111111111;
															assign node6963 = (inp[9]) ? 16'b0000000011111111 : node6964;
																assign node6964 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6968 = (inp[12]) ? node6970 : 16'b0000000001111111;
															assign node6970 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6973 = (inp[12]) ? 16'b0000000001111111 : node6974;
													assign node6974 = (inp[11]) ? node6976 : 16'b0000000011111111;
														assign node6976 = (inp[9]) ? 16'b0000000001111111 : node6977;
															assign node6977 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6982 = (inp[12]) ? node6998 : node6983;
												assign node6983 = (inp[6]) ? node6991 : node6984;
													assign node6984 = (inp[11]) ? 16'b0000000001111111 : node6985;
														assign node6985 = (inp[9]) ? 16'b0000000011111111 : node6986;
															assign node6986 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6991 = (inp[13]) ? 16'b0000000001111111 : node6992;
														assign node6992 = (inp[8]) ? node6994 : 16'b0000000011111111;
															assign node6994 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6998 = (inp[11]) ? node7014 : node6999;
													assign node6999 = (inp[6]) ? node7007 : node7000;
														assign node7000 = (inp[9]) ? node7002 : 16'b0000000011111111;
															assign node7002 = (inp[8]) ? 16'b0000000001111111 : node7003;
																assign node7003 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7007 = (inp[13]) ? node7009 : 16'b0000000001111111;
															assign node7009 = (inp[8]) ? 16'b0000000000111111 : node7010;
																assign node7010 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7014 = (inp[13]) ? node7016 : 16'b0000000000111111;
														assign node7016 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7019 = (inp[13]) ? node7161 : node7020;
									assign node7020 = (inp[7]) ? node7090 : node7021;
										assign node7021 = (inp[11]) ? node7059 : node7022;
											assign node7022 = (inp[9]) ? node7042 : node7023;
												assign node7023 = (inp[12]) ? node7037 : node7024;
													assign node7024 = (inp[5]) ? node7032 : node7025;
														assign node7025 = (inp[6]) ? node7027 : 16'b0000011111111111;
															assign node7027 = (inp[15]) ? 16'b0000001111111111 : node7028;
																assign node7028 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7032 = (inp[15]) ? node7034 : 16'b0000001111111111;
															assign node7034 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7037 = (inp[6]) ? node7039 : 16'b0000001111111111;
														assign node7039 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7042 = (inp[6]) ? node7046 : node7043;
													assign node7043 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7046 = (inp[15]) ? node7056 : node7047;
														assign node7047 = (inp[8]) ? node7051 : node7048;
															assign node7048 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node7051 = (inp[12]) ? 16'b0000000011111111 : node7052;
																assign node7052 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7056 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7059 = (inp[8]) ? node7079 : node7060;
												assign node7060 = (inp[6]) ? node7068 : node7061;
													assign node7061 = (inp[15]) ? node7063 : 16'b0000000111111111;
														assign node7063 = (inp[12]) ? 16'b0000000011111111 : node7064;
															assign node7064 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7068 = (inp[12]) ? node7076 : node7069;
														assign node7069 = (inp[9]) ? node7071 : 16'b0000000111111111;
															assign node7071 = (inp[5]) ? 16'b0000000011111111 : node7072;
																assign node7072 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7076 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7079 = (inp[6]) ? node7081 : 16'b0000000111111111;
													assign node7081 = (inp[5]) ? 16'b0000000000111111 : node7082;
														assign node7082 = (inp[15]) ? node7086 : node7083;
															assign node7083 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node7086 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7090 = (inp[15]) ? node7118 : node7091;
											assign node7091 = (inp[6]) ? node7099 : node7092;
												assign node7092 = (inp[9]) ? node7094 : 16'b0000000111111111;
													assign node7094 = (inp[8]) ? node7096 : 16'b0000000111111111;
														assign node7096 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7099 = (inp[11]) ? node7109 : node7100;
													assign node7100 = (inp[12]) ? 16'b0000000001111111 : node7101;
														assign node7101 = (inp[5]) ? node7103 : 16'b0000000111111111;
															assign node7103 = (inp[8]) ? 16'b0000000011111111 : node7104;
																assign node7104 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7109 = (inp[8]) ? node7113 : node7110;
														assign node7110 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7113 = (inp[5]) ? 16'b0000000001111111 : node7114;
															assign node7114 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7118 = (inp[8]) ? node7144 : node7119;
												assign node7119 = (inp[9]) ? node7131 : node7120;
													assign node7120 = (inp[5]) ? node7128 : node7121;
														assign node7121 = (inp[11]) ? 16'b0000000011111111 : node7122;
															assign node7122 = (inp[12]) ? node7124 : 16'b0000000111111111;
																assign node7124 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7128 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7131 = (inp[12]) ? node7133 : 16'b0000000011111111;
														assign node7133 = (inp[5]) ? node7139 : node7134;
															assign node7134 = (inp[6]) ? 16'b0000000001111111 : node7135;
																assign node7135 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node7139 = (inp[6]) ? 16'b0000000000111111 : node7140;
																assign node7140 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7144 = (inp[9]) ? node7154 : node7145;
													assign node7145 = (inp[5]) ? node7147 : 16'b0000000001111111;
														assign node7147 = (inp[12]) ? node7149 : 16'b0000000001111111;
															assign node7149 = (inp[11]) ? 16'b0000000000111111 : node7150;
																assign node7150 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7154 = (inp[11]) ? node7156 : 16'b0000000001111111;
														assign node7156 = (inp[5]) ? node7158 : 16'b0000000000111111;
															assign node7158 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node7161 = (inp[12]) ? node7227 : node7162;
										assign node7162 = (inp[15]) ? node7194 : node7163;
											assign node7163 = (inp[7]) ? node7187 : node7164;
												assign node7164 = (inp[11]) ? node7180 : node7165;
													assign node7165 = (inp[9]) ? node7173 : node7166;
														assign node7166 = (inp[8]) ? node7168 : 16'b0000001111111111;
															assign node7168 = (inp[6]) ? node7170 : 16'b0000000111111111;
																assign node7170 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7173 = (inp[5]) ? 16'b0000000011111111 : node7174;
															assign node7174 = (inp[6]) ? node7176 : 16'b0000000111111111;
																assign node7176 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7180 = (inp[5]) ? node7184 : node7181;
														assign node7181 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node7184 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7187 = (inp[8]) ? 16'b0000000001111111 : node7188;
													assign node7188 = (inp[11]) ? 16'b0000000001111111 : node7189;
														assign node7189 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7194 = (inp[8]) ? node7210 : node7195;
												assign node7195 = (inp[9]) ? node7207 : node7196;
													assign node7196 = (inp[11]) ? node7202 : node7197;
														assign node7197 = (inp[5]) ? node7199 : 16'b0000000111111111;
															assign node7199 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7202 = (inp[6]) ? node7204 : 16'b0000000011111111;
															assign node7204 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7207 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7210 = (inp[7]) ? node7218 : node7211;
													assign node7211 = (inp[6]) ? node7213 : 16'b0000000001111111;
														assign node7213 = (inp[9]) ? 16'b0000000000111111 : node7214;
															assign node7214 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7218 = (inp[5]) ? node7220 : 16'b0000000000111111;
														assign node7220 = (inp[6]) ? node7222 : 16'b0000000000111111;
															assign node7222 = (inp[11]) ? 16'b0000000000011111 : node7223;
																assign node7223 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7227 = (inp[9]) ? node7249 : node7228;
											assign node7228 = (inp[15]) ? node7238 : node7229;
												assign node7229 = (inp[6]) ? node7235 : node7230;
													assign node7230 = (inp[8]) ? node7232 : 16'b0000000011111111;
														assign node7232 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7235 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7238 = (inp[5]) ? node7244 : node7239;
													assign node7239 = (inp[7]) ? node7241 : 16'b0000000001111111;
														assign node7241 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7244 = (inp[6]) ? node7246 : 16'b0000000000111111;
														assign node7246 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7249 = (inp[5]) ? node7263 : node7250;
												assign node7250 = (inp[11]) ? node7260 : node7251;
													assign node7251 = (inp[15]) ? 16'b0000000000111111 : node7252;
														assign node7252 = (inp[8]) ? node7254 : 16'b0000000011111111;
															assign node7254 = (inp[6]) ? node7256 : 16'b0000000001111111;
																assign node7256 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7260 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7263 = (inp[7]) ? node7267 : node7264;
													assign node7264 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node7267 = (inp[8]) ? node7275 : node7268;
														assign node7268 = (inp[15]) ? node7270 : 16'b0000000000111111;
															assign node7270 = (inp[6]) ? node7272 : 16'b0000000000011111;
																assign node7272 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node7275 = (inp[6]) ? 16'b0000000000001111 : node7276;
															assign node7276 = (inp[11]) ? node7278 : 16'b0000000000011111;
																assign node7278 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node7282 = (inp[3]) ? node7790 : node7283;
							assign node7283 = (inp[5]) ? node7523 : node7284;
								assign node7284 = (inp[12]) ? node7396 : node7285;
									assign node7285 = (inp[6]) ? node7337 : node7286;
										assign node7286 = (inp[7]) ? node7312 : node7287;
											assign node7287 = (inp[1]) ? node7301 : node7288;
												assign node7288 = (inp[11]) ? node7298 : node7289;
													assign node7289 = (inp[15]) ? 16'b0000011111111111 : node7290;
														assign node7290 = (inp[9]) ? 16'b0000011111111111 : node7291;
															assign node7291 = (inp[8]) ? node7293 : 16'b0000111111111111;
																assign node7293 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7298 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7301 = (inp[11]) ? node7305 : node7302;
													assign node7302 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7305 = (inp[8]) ? node7309 : node7306;
														assign node7306 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7309 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7312 = (inp[15]) ? node7330 : node7313;
												assign node7313 = (inp[9]) ? node7323 : node7314;
													assign node7314 = (inp[1]) ? node7318 : node7315;
														assign node7315 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7318 = (inp[8]) ? node7320 : 16'b0000001111111111;
															assign node7320 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7323 = (inp[13]) ? node7327 : node7324;
														assign node7324 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7327 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7330 = (inp[1]) ? 16'b0000000011111111 : node7331;
													assign node7331 = (inp[13]) ? node7333 : 16'b0000000111111111;
														assign node7333 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7337 = (inp[8]) ? node7371 : node7338;
											assign node7338 = (inp[7]) ? node7356 : node7339;
												assign node7339 = (inp[9]) ? node7351 : node7340;
													assign node7340 = (inp[11]) ? node7344 : node7341;
														assign node7341 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7344 = (inp[13]) ? 16'b0000000111111111 : node7345;
															assign node7345 = (inp[1]) ? node7347 : 16'b0000001111111111;
																assign node7347 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7351 = (inp[1]) ? node7353 : 16'b0000000111111111;
														assign node7353 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7356 = (inp[11]) ? 16'b0000000011111111 : node7357;
													assign node7357 = (inp[13]) ? node7365 : node7358;
														assign node7358 = (inp[1]) ? node7360 : 16'b0000001111111111;
															assign node7360 = (inp[9]) ? node7362 : 16'b0000000111111111;
																assign node7362 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7365 = (inp[9]) ? 16'b0000000011111111 : node7366;
															assign node7366 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7371 = (inp[11]) ? node7387 : node7372;
												assign node7372 = (inp[15]) ? node7380 : node7373;
													assign node7373 = (inp[1]) ? node7377 : node7374;
														assign node7374 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7377 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7380 = (inp[1]) ? node7384 : node7381;
														assign node7381 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7384 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7387 = (inp[9]) ? node7393 : node7388;
													assign node7388 = (inp[1]) ? node7390 : 16'b0000000011111111;
														assign node7390 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7393 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7396 = (inp[11]) ? node7466 : node7397;
										assign node7397 = (inp[8]) ? node7433 : node7398;
											assign node7398 = (inp[1]) ? node7412 : node7399;
												assign node7399 = (inp[9]) ? node7405 : node7400;
													assign node7400 = (inp[15]) ? node7402 : 16'b0000011111111111;
														assign node7402 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7405 = (inp[15]) ? 16'b0000000111111111 : node7406;
														assign node7406 = (inp[13]) ? node7408 : 16'b0000001111111111;
															assign node7408 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7412 = (inp[13]) ? node7424 : node7413;
													assign node7413 = (inp[15]) ? node7421 : node7414;
														assign node7414 = (inp[9]) ? node7416 : 16'b0000001111111111;
															assign node7416 = (inp[7]) ? 16'b0000000111111111 : node7417;
																assign node7417 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7421 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7424 = (inp[7]) ? node7430 : node7425;
														assign node7425 = (inp[9]) ? node7427 : 16'b0000000111111111;
															assign node7427 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7430 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7433 = (inp[9]) ? node7453 : node7434;
												assign node7434 = (inp[13]) ? node7442 : node7435;
													assign node7435 = (inp[1]) ? node7439 : node7436;
														assign node7436 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7439 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node7442 = (inp[7]) ? 16'b0000000011111111 : node7443;
														assign node7443 = (inp[6]) ? node7445 : 16'b0000000111111111;
															assign node7445 = (inp[15]) ? node7449 : node7446;
																assign node7446 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node7449 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7453 = (inp[1]) ? node7461 : node7454;
													assign node7454 = (inp[7]) ? node7458 : node7455;
														assign node7455 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7458 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7461 = (inp[15]) ? node7463 : 16'b0000000001111111;
														assign node7463 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7466 = (inp[13]) ? node7498 : node7467;
											assign node7467 = (inp[9]) ? node7483 : node7468;
												assign node7468 = (inp[7]) ? node7476 : node7469;
													assign node7469 = (inp[8]) ? node7473 : node7470;
														assign node7470 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7473 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7476 = (inp[8]) ? node7478 : 16'b0000000011111111;
														assign node7478 = (inp[1]) ? node7480 : 16'b0000000011111111;
															assign node7480 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7483 = (inp[8]) ? node7493 : node7484;
													assign node7484 = (inp[15]) ? node7490 : node7485;
														assign node7485 = (inp[1]) ? 16'b0000000011111111 : node7486;
															assign node7486 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7490 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7493 = (inp[7]) ? 16'b0000000001111111 : node7494;
														assign node7494 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7498 = (inp[1]) ? node7508 : node7499;
												assign node7499 = (inp[15]) ? node7503 : node7500;
													assign node7500 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7503 = (inp[9]) ? 16'b0000000001111111 : node7504;
														assign node7504 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7508 = (inp[6]) ? node7514 : node7509;
													assign node7509 = (inp[15]) ? 16'b0000000001111111 : node7510;
														assign node7510 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7514 = (inp[7]) ? 16'b0000000000111111 : node7515;
														assign node7515 = (inp[8]) ? node7517 : 16'b0000000001111111;
															assign node7517 = (inp[9]) ? 16'b0000000000011111 : node7518;
																assign node7518 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node7523 = (inp[12]) ? node7659 : node7524;
									assign node7524 = (inp[7]) ? node7594 : node7525;
										assign node7525 = (inp[6]) ? node7559 : node7526;
											assign node7526 = (inp[8]) ? node7538 : node7527;
												assign node7527 = (inp[11]) ? node7533 : node7528;
													assign node7528 = (inp[13]) ? node7530 : 16'b0000011111111111;
														assign node7530 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7533 = (inp[15]) ? 16'b0000000111111111 : node7534;
														assign node7534 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7538 = (inp[1]) ? node7550 : node7539;
													assign node7539 = (inp[9]) ? node7547 : node7540;
														assign node7540 = (inp[15]) ? 16'b0000000011111111 : node7541;
															assign node7541 = (inp[13]) ? 16'b0000001111111111 : node7542;
																assign node7542 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7547 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7550 = (inp[13]) ? 16'b0000000011111111 : node7551;
														assign node7551 = (inp[9]) ? 16'b0000000011111111 : node7552;
															assign node7552 = (inp[15]) ? node7554 : 16'b0000000111111111;
																assign node7554 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7559 = (inp[11]) ? node7583 : node7560;
												assign node7560 = (inp[1]) ? node7570 : node7561;
													assign node7561 = (inp[9]) ? node7567 : node7562;
														assign node7562 = (inp[8]) ? 16'b0000000111111111 : node7563;
															assign node7563 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7567 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7570 = (inp[13]) ? node7578 : node7571;
														assign node7571 = (inp[15]) ? node7573 : 16'b0000001111111111;
															assign node7573 = (inp[8]) ? 16'b0000000011111111 : node7574;
																assign node7574 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7578 = (inp[8]) ? 16'b0000000001111111 : node7579;
															assign node7579 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7583 = (inp[13]) ? node7585 : 16'b0000000011111111;
													assign node7585 = (inp[9]) ? node7591 : node7586;
														assign node7586 = (inp[1]) ? node7588 : 16'b0000000011111111;
															assign node7588 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7591 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7594 = (inp[8]) ? node7626 : node7595;
											assign node7595 = (inp[11]) ? node7607 : node7596;
												assign node7596 = (inp[15]) ? 16'b0000000001111111 : node7597;
													assign node7597 = (inp[13]) ? 16'b0000000111111111 : node7598;
														assign node7598 = (inp[9]) ? node7600 : 16'b0000001111111111;
															assign node7600 = (inp[1]) ? 16'b0000000111111111 : node7601;
																assign node7601 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7607 = (inp[13]) ? node7617 : node7608;
													assign node7608 = (inp[9]) ? node7614 : node7609;
														assign node7609 = (inp[15]) ? node7611 : 16'b0000000111111111;
															assign node7611 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7614 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node7617 = (inp[1]) ? node7621 : node7618;
														assign node7618 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7621 = (inp[9]) ? 16'b0000000000111111 : node7622;
															assign node7622 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node7626 = (inp[1]) ? node7644 : node7627;
												assign node7627 = (inp[9]) ? 16'b0000000001111111 : node7628;
													assign node7628 = (inp[6]) ? node7632 : node7629;
														assign node7629 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7632 = (inp[15]) ? node7638 : node7633;
															assign node7633 = (inp[11]) ? node7635 : 16'b0000000011111111;
																assign node7635 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node7638 = (inp[11]) ? node7640 : 16'b0000000001111111;
																assign node7640 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7644 = (inp[13]) ? node7654 : node7645;
													assign node7645 = (inp[9]) ? node7649 : node7646;
														assign node7646 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7649 = (inp[6]) ? node7651 : 16'b0000000001111111;
															assign node7651 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7654 = (inp[6]) ? 16'b0000000000111111 : node7655;
														assign node7655 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7659 = (inp[13]) ? node7723 : node7660;
										assign node7660 = (inp[15]) ? node7700 : node7661;
											assign node7661 = (inp[9]) ? node7679 : node7662;
												assign node7662 = (inp[7]) ? node7670 : node7663;
													assign node7663 = (inp[8]) ? 16'b0000000111111111 : node7664;
														assign node7664 = (inp[11]) ? node7666 : 16'b0000011111111111;
															assign node7666 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7670 = (inp[1]) ? node7674 : node7671;
														assign node7671 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7674 = (inp[8]) ? node7676 : 16'b0000000011111111;
															assign node7676 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7679 = (inp[8]) ? node7689 : node7680;
													assign node7680 = (inp[1]) ? node7684 : node7681;
														assign node7681 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7684 = (inp[6]) ? node7686 : 16'b0000000011111111;
															assign node7686 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7689 = (inp[1]) ? node7697 : node7690;
														assign node7690 = (inp[7]) ? node7692 : 16'b0000000011111111;
															assign node7692 = (inp[11]) ? 16'b0000000001111111 : node7693;
																assign node7693 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7697 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node7700 = (inp[11]) ? node7710 : node7701;
												assign node7701 = (inp[1]) ? node7703 : 16'b0000000011111111;
													assign node7703 = (inp[7]) ? node7707 : node7704;
														assign node7704 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7707 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7710 = (inp[7]) ? node7718 : node7711;
													assign node7711 = (inp[8]) ? node7713 : 16'b0000000001111111;
														assign node7713 = (inp[9]) ? node7715 : 16'b0000000001111111;
															assign node7715 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7718 = (inp[8]) ? node7720 : 16'b0000000001111111;
														assign node7720 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node7723 = (inp[1]) ? node7755 : node7724;
											assign node7724 = (inp[11]) ? node7748 : node7725;
												assign node7725 = (inp[6]) ? node7743 : node7726;
													assign node7726 = (inp[15]) ? node7732 : node7727;
														assign node7727 = (inp[8]) ? 16'b0000000011111111 : node7728;
															assign node7728 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7732 = (inp[7]) ? node7738 : node7733;
															assign node7733 = (inp[9]) ? node7735 : 16'b0000000011111111;
																assign node7735 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node7738 = (inp[8]) ? node7740 : 16'b0000000001111111;
																assign node7740 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7743 = (inp[7]) ? node7745 : 16'b0000000001111111;
														assign node7745 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node7748 = (inp[15]) ? node7752 : node7749;
													assign node7749 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7752 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node7755 = (inp[15]) ? node7775 : node7756;
												assign node7756 = (inp[7]) ? node7766 : node7757;
													assign node7757 = (inp[6]) ? node7759 : 16'b0000000001111111;
														assign node7759 = (inp[9]) ? node7761 : 16'b0000000001111111;
															assign node7761 = (inp[11]) ? 16'b0000000000111111 : node7762;
																assign node7762 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7766 = (inp[6]) ? node7770 : node7767;
														assign node7767 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7770 = (inp[8]) ? node7772 : 16'b0000000000111111;
															assign node7772 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7775 = (inp[8]) ? node7781 : node7776;
													assign node7776 = (inp[9]) ? 16'b0000000000111111 : node7777;
														assign node7777 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7781 = (inp[6]) ? node7787 : node7782;
														assign node7782 = (inp[11]) ? node7784 : 16'b0000000000111111;
															assign node7784 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node7787 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7790 = (inp[11]) ? node8094 : node7791;
								assign node7791 = (inp[13]) ? node7949 : node7792;
									assign node7792 = (inp[8]) ? node7870 : node7793;
										assign node7793 = (inp[12]) ? node7833 : node7794;
											assign node7794 = (inp[5]) ? node7806 : node7795;
												assign node7795 = (inp[9]) ? 16'b0000000111111111 : node7796;
													assign node7796 = (inp[7]) ? node7800 : node7797;
														assign node7797 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7800 = (inp[15]) ? 16'b0000000111111111 : node7801;
															assign node7801 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7806 = (inp[15]) ? node7818 : node7807;
													assign node7807 = (inp[9]) ? node7813 : node7808;
														assign node7808 = (inp[1]) ? 16'b0000000111111111 : node7809;
															assign node7809 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7813 = (inp[6]) ? node7815 : 16'b0000000111111111;
															assign node7815 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7818 = (inp[6]) ? node7826 : node7819;
														assign node7819 = (inp[9]) ? node7821 : 16'b0000000111111111;
															assign node7821 = (inp[1]) ? 16'b0000000011111111 : node7822;
																assign node7822 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7826 = (inp[9]) ? 16'b0000000000111111 : node7827;
															assign node7827 = (inp[1]) ? node7829 : 16'b0000000011111111;
																assign node7829 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7833 = (inp[1]) ? node7853 : node7834;
												assign node7834 = (inp[15]) ? node7844 : node7835;
													assign node7835 = (inp[9]) ? node7839 : node7836;
														assign node7836 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7839 = (inp[5]) ? node7841 : 16'b0000000111111111;
															assign node7841 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7844 = (inp[5]) ? 16'b0000000011111111 : node7845;
														assign node7845 = (inp[9]) ? 16'b0000000011111111 : node7846;
															assign node7846 = (inp[7]) ? node7848 : 16'b0000000111111111;
																assign node7848 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7853 = (inp[6]) ? node7865 : node7854;
													assign node7854 = (inp[5]) ? node7862 : node7855;
														assign node7855 = (inp[15]) ? 16'b0000000011111111 : node7856;
															assign node7856 = (inp[9]) ? node7858 : 16'b0000000111111111;
																assign node7858 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7862 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7865 = (inp[9]) ? node7867 : 16'b0000000011111111;
														assign node7867 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7870 = (inp[6]) ? node7906 : node7871;
											assign node7871 = (inp[15]) ? node7891 : node7872;
												assign node7872 = (inp[7]) ? node7882 : node7873;
													assign node7873 = (inp[5]) ? 16'b0000000111111111 : node7874;
														assign node7874 = (inp[1]) ? 16'b0000000111111111 : node7875;
															assign node7875 = (inp[12]) ? 16'b0000001111111111 : node7876;
																assign node7876 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7882 = (inp[5]) ? node7888 : node7883;
														assign node7883 = (inp[9]) ? 16'b0000000011111111 : node7884;
															assign node7884 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7888 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7891 = (inp[1]) ? node7899 : node7892;
													assign node7892 = (inp[7]) ? node7894 : 16'b0000000011111111;
														assign node7894 = (inp[5]) ? node7896 : 16'b0000000011111111;
															assign node7896 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7899 = (inp[5]) ? 16'b0000000001111111 : node7900;
														assign node7900 = (inp[9]) ? 16'b0000000001111111 : node7901;
															assign node7901 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7906 = (inp[1]) ? node7930 : node7907;
												assign node7907 = (inp[7]) ? node7915 : node7908;
													assign node7908 = (inp[9]) ? node7912 : node7909;
														assign node7909 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7912 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7915 = (inp[12]) ? node7927 : node7916;
														assign node7916 = (inp[9]) ? node7922 : node7917;
															assign node7917 = (inp[5]) ? node7919 : 16'b0000000011111111;
																assign node7919 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node7922 = (inp[15]) ? 16'b0000000001111111 : node7923;
																assign node7923 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7927 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7930 = (inp[9]) ? node7936 : node7931;
													assign node7931 = (inp[5]) ? 16'b0000000001111111 : node7932;
														assign node7932 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7936 = (inp[5]) ? node7944 : node7937;
														assign node7937 = (inp[12]) ? 16'b0000000000111111 : node7938;
															assign node7938 = (inp[7]) ? 16'b0000000000111111 : node7939;
																assign node7939 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7944 = (inp[12]) ? node7946 : 16'b0000000000011111;
															assign node7946 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7949 = (inp[15]) ? node8019 : node7950;
										assign node7950 = (inp[7]) ? node7978 : node7951;
											assign node7951 = (inp[6]) ? node7967 : node7952;
												assign node7952 = (inp[9]) ? node7958 : node7953;
													assign node7953 = (inp[8]) ? node7955 : 16'b0000001111111111;
														assign node7955 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7958 = (inp[12]) ? 16'b0000000011111111 : node7959;
														assign node7959 = (inp[5]) ? 16'b0000000011111111 : node7960;
															assign node7960 = (inp[1]) ? node7962 : 16'b0000000111111111;
																assign node7962 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7967 = (inp[5]) ? node7969 : 16'b0000000011111111;
													assign node7969 = (inp[1]) ? node7975 : node7970;
														assign node7970 = (inp[12]) ? 16'b0000000001111111 : node7971;
															assign node7971 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7975 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7978 = (inp[1]) ? node7998 : node7979;
												assign node7979 = (inp[6]) ? node7987 : node7980;
													assign node7980 = (inp[8]) ? node7982 : 16'b0000000011111111;
														assign node7982 = (inp[9]) ? 16'b0000000001111111 : node7983;
															assign node7983 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7987 = (inp[8]) ? node7995 : node7988;
														assign node7988 = (inp[12]) ? node7990 : 16'b0000000011111111;
															assign node7990 = (inp[5]) ? 16'b0000000001111111 : node7991;
																assign node7991 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7995 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node7998 = (inp[5]) ? node8010 : node7999;
													assign node7999 = (inp[6]) ? node8005 : node8000;
														assign node8000 = (inp[12]) ? node8002 : 16'b0000000111111111;
															assign node8002 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8005 = (inp[9]) ? 16'b0000000000111111 : node8006;
															assign node8006 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8010 = (inp[12]) ? node8012 : 16'b0000000001111111;
														assign node8012 = (inp[8]) ? 16'b0000000000011111 : node8013;
															assign node8013 = (inp[9]) ? node8015 : 16'b0000000000111111;
																assign node8015 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8019 = (inp[5]) ? node8065 : node8020;
											assign node8020 = (inp[12]) ? node8044 : node8021;
												assign node8021 = (inp[6]) ? node8033 : node8022;
													assign node8022 = (inp[7]) ? node8028 : node8023;
														assign node8023 = (inp[1]) ? 16'b0000000011111111 : node8024;
															assign node8024 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8028 = (inp[9]) ? 16'b0000000001111111 : node8029;
															assign node8029 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8033 = (inp[1]) ? node8037 : node8034;
														assign node8034 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8037 = (inp[9]) ? node8039 : 16'b0000000001111111;
															assign node8039 = (inp[8]) ? 16'b0000000000111111 : node8040;
																assign node8040 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8044 = (inp[1]) ? node8056 : node8045;
													assign node8045 = (inp[8]) ? node8049 : node8046;
														assign node8046 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node8049 = (inp[9]) ? 16'b0000000000111111 : node8050;
															assign node8050 = (inp[6]) ? node8052 : 16'b0000000001111111;
																assign node8052 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8056 = (inp[6]) ? node8062 : node8057;
														assign node8057 = (inp[7]) ? 16'b0000000000111111 : node8058;
															assign node8058 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8062 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8065 = (inp[9]) ? node8081 : node8066;
												assign node8066 = (inp[8]) ? node8074 : node8067;
													assign node8067 = (inp[7]) ? 16'b0000000000111111 : node8068;
														assign node8068 = (inp[12]) ? 16'b0000000001111111 : node8069;
															assign node8069 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8074 = (inp[6]) ? node8076 : 16'b0000000001111111;
														assign node8076 = (inp[1]) ? node8078 : 16'b0000000000111111;
															assign node8078 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8081 = (inp[8]) ? node8091 : node8082;
													assign node8082 = (inp[6]) ? node8086 : node8083;
														assign node8083 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8086 = (inp[7]) ? node8088 : 16'b0000000000111111;
															assign node8088 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8091 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
								assign node8094 = (inp[12]) ? node8244 : node8095;
									assign node8095 = (inp[8]) ? node8163 : node8096;
										assign node8096 = (inp[13]) ? node8122 : node8097;
											assign node8097 = (inp[1]) ? node8113 : node8098;
												assign node8098 = (inp[7]) ? node8110 : node8099;
													assign node8099 = (inp[5]) ? node8107 : node8100;
														assign node8100 = (inp[9]) ? 16'b0000000111111111 : node8101;
															assign node8101 = (inp[15]) ? 16'b0000001111111111 : node8102;
																assign node8102 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8107 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8110 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node8113 = (inp[5]) ? node8115 : 16'b0000000011111111;
													assign node8115 = (inp[15]) ? 16'b0000000001111111 : node8116;
														assign node8116 = (inp[9]) ? node8118 : 16'b0000000011111111;
															assign node8118 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8122 = (inp[6]) ? node8142 : node8123;
												assign node8123 = (inp[1]) ? node8131 : node8124;
													assign node8124 = (inp[5]) ? node8126 : 16'b0000000111111111;
														assign node8126 = (inp[7]) ? 16'b0000000011111111 : node8127;
															assign node8127 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8131 = (inp[15]) ? node8139 : node8132;
														assign node8132 = (inp[5]) ? 16'b0000000001111111 : node8133;
															assign node8133 = (inp[7]) ? node8135 : 16'b0000000011111111;
																assign node8135 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8139 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8142 = (inp[15]) ? node8154 : node8143;
													assign node8143 = (inp[5]) ? node8151 : node8144;
														assign node8144 = (inp[1]) ? 16'b0000000001111111 : node8145;
															assign node8145 = (inp[7]) ? node8147 : 16'b0000000011111111;
																assign node8147 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8151 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8154 = (inp[9]) ? node8158 : node8155;
														assign node8155 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8158 = (inp[7]) ? node8160 : 16'b0000000000111111;
															assign node8160 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8163 = (inp[6]) ? node8211 : node8164;
											assign node8164 = (inp[15]) ? node8196 : node8165;
												assign node8165 = (inp[13]) ? node8179 : node8166;
													assign node8166 = (inp[7]) ? node8174 : node8167;
														assign node8167 = (inp[5]) ? 16'b0000000001111111 : node8168;
															assign node8168 = (inp[1]) ? node8170 : 16'b0000000111111111;
																assign node8170 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8174 = (inp[1]) ? node8176 : 16'b0000000011111111;
															assign node8176 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8179 = (inp[9]) ? node8187 : node8180;
														assign node8180 = (inp[5]) ? node8182 : 16'b0000000011111111;
															assign node8182 = (inp[1]) ? 16'b0000000001111111 : node8183;
																assign node8183 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8187 = (inp[5]) ? node8193 : node8188;
															assign node8188 = (inp[1]) ? node8190 : 16'b0000000001111111;
																assign node8190 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node8193 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8196 = (inp[9]) ? node8206 : node8197;
													assign node8197 = (inp[1]) ? node8201 : node8198;
														assign node8198 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8201 = (inp[7]) ? 16'b0000000000111111 : node8202;
															assign node8202 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8206 = (inp[5]) ? 16'b0000000000011111 : node8207;
														assign node8207 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8211 = (inp[5]) ? node8233 : node8212;
												assign node8212 = (inp[1]) ? node8218 : node8213;
													assign node8213 = (inp[7]) ? 16'b0000000001111111 : node8214;
														assign node8214 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8218 = (inp[15]) ? node8230 : node8219;
														assign node8219 = (inp[9]) ? node8225 : node8220;
															assign node8220 = (inp[7]) ? node8222 : 16'b0000000001111111;
																assign node8222 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node8225 = (inp[7]) ? node8227 : 16'b0000000000111111;
																assign node8227 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node8230 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8233 = (inp[13]) ? node8239 : node8234;
													assign node8234 = (inp[9]) ? node8236 : 16'b0000000000111111;
														assign node8236 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8239 = (inp[15]) ? 16'b0000000000001111 : node8240;
														assign node8240 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node8244 = (inp[13]) ? node8306 : node8245;
										assign node8245 = (inp[6]) ? node8275 : node8246;
											assign node8246 = (inp[15]) ? node8262 : node8247;
												assign node8247 = (inp[8]) ? node8255 : node8248;
													assign node8248 = (inp[5]) ? 16'b0000000011111111 : node8249;
														assign node8249 = (inp[7]) ? node8251 : 16'b0000000111111111;
															assign node8251 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8255 = (inp[7]) ? node8259 : node8256;
														assign node8256 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8259 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8262 = (inp[9]) ? node8272 : node8263;
													assign node8263 = (inp[7]) ? node8265 : 16'b0000000001111111;
														assign node8265 = (inp[5]) ? 16'b0000000000111111 : node8266;
															assign node8266 = (inp[1]) ? node8268 : 16'b0000000001111111;
																assign node8268 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8272 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node8275 = (inp[9]) ? node8291 : node8276;
												assign node8276 = (inp[1]) ? node8282 : node8277;
													assign node8277 = (inp[7]) ? 16'b0000000001111111 : node8278;
														assign node8278 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8282 = (inp[7]) ? node8284 : 16'b0000000001111111;
														assign node8284 = (inp[8]) ? 16'b0000000000011111 : node8285;
															assign node8285 = (inp[5]) ? node8287 : 16'b0000000000111111;
																assign node8287 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8291 = (inp[15]) ? node8297 : node8292;
													assign node8292 = (inp[7]) ? node8294 : 16'b0000000001111111;
														assign node8294 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8297 = (inp[5]) ? node8301 : node8298;
														assign node8298 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node8301 = (inp[8]) ? node8303 : 16'b0000000000011111;
															assign node8303 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node8306 = (inp[1]) ? node8338 : node8307;
											assign node8307 = (inp[8]) ? node8317 : node8308;
												assign node8308 = (inp[9]) ? node8312 : node8309;
													assign node8309 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8312 = (inp[5]) ? 16'b0000000000111111 : node8313;
														assign node8313 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8317 = (inp[6]) ? node8327 : node8318;
													assign node8318 = (inp[5]) ? node8320 : 16'b0000000000111111;
														assign node8320 = (inp[9]) ? 16'b0000000000011111 : node8321;
															assign node8321 = (inp[15]) ? node8323 : 16'b0000000000111111;
																assign node8323 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8327 = (inp[7]) ? node8335 : node8328;
														assign node8328 = (inp[9]) ? 16'b0000000000011111 : node8329;
															assign node8329 = (inp[5]) ? node8331 : 16'b0000000000111111;
																assign node8331 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node8335 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8338 = (inp[15]) ? node8360 : node8339;
												assign node8339 = (inp[9]) ? node8351 : node8340;
													assign node8340 = (inp[7]) ? node8344 : node8341;
														assign node8341 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8344 = (inp[6]) ? 16'b0000000000011111 : node8345;
															assign node8345 = (inp[8]) ? node8347 : 16'b0000000000111111;
																assign node8347 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8351 = (inp[8]) ? 16'b0000000000001111 : node8352;
														assign node8352 = (inp[7]) ? node8354 : 16'b0000000000111111;
															assign node8354 = (inp[6]) ? node8356 : 16'b0000000000011111;
																assign node8356 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node8360 = (inp[7]) ? node8366 : node8361;
													assign node8361 = (inp[6]) ? node8363 : 16'b0000000000011111;
														assign node8363 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node8366 = (inp[9]) ? node8368 : 16'b0000000000001111;
														assign node8368 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
			assign node8371 = (inp[8]) ? node12489 : node8372;
				assign node8372 = (inp[5]) ? node10488 : node8373;
					assign node8373 = (inp[1]) ? node9405 : node8374;
						assign node8374 = (inp[6]) ? node8884 : node8375;
							assign node8375 = (inp[3]) ? node8647 : node8376;
								assign node8376 = (inp[9]) ? node8530 : node8377;
									assign node8377 = (inp[7]) ? node8461 : node8378;
										assign node8378 = (inp[12]) ? node8420 : node8379;
											assign node8379 = (inp[15]) ? node8407 : node8380;
												assign node8380 = (inp[11]) ? node8400 : node8381;
													assign node8381 = (inp[10]) ? node8391 : node8382;
														assign node8382 = (inp[14]) ? node8388 : node8383;
															assign node8383 = (inp[2]) ? 16'b0011111111111111 : node8384;
																assign node8384 = (inp[13]) ? 16'b0011111111111111 : 16'b0111111111111111;
															assign node8388 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node8391 = (inp[14]) ? node8397 : node8392;
															assign node8392 = (inp[2]) ? 16'b0001111111111111 : node8393;
																assign node8393 = (inp[13]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node8397 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node8400 = (inp[14]) ? 16'b0000111111111111 : node8401;
														assign node8401 = (inp[2]) ? 16'b0000111111111111 : node8402;
															assign node8402 = (inp[13]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node8407 = (inp[2]) ? 16'b0000011111111111 : node8408;
													assign node8408 = (inp[13]) ? node8416 : node8409;
														assign node8409 = (inp[11]) ? node8411 : 16'b0001111111111111;
															assign node8411 = (inp[10]) ? 16'b0000111111111111 : node8412;
																assign node8412 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8416 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node8420 = (inp[10]) ? node8438 : node8421;
												assign node8421 = (inp[14]) ? node8433 : node8422;
													assign node8422 = (inp[11]) ? node8426 : node8423;
														assign node8423 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8426 = (inp[13]) ? node8428 : 16'b0000111111111111;
															assign node8428 = (inp[2]) ? 16'b0000011111111111 : node8429;
																assign node8429 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8433 = (inp[11]) ? 16'b0000011111111111 : node8434;
														assign node8434 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8438 = (inp[13]) ? node8452 : node8439;
													assign node8439 = (inp[14]) ? node8447 : node8440;
														assign node8440 = (inp[11]) ? 16'b0000011111111111 : node8441;
															assign node8441 = (inp[15]) ? node8443 : 16'b0000111111111111;
																assign node8443 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8447 = (inp[2]) ? node8449 : 16'b0000011111111111;
															assign node8449 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8452 = (inp[14]) ? node8458 : node8453;
														assign node8453 = (inp[15]) ? node8455 : 16'b0000011111111111;
															assign node8455 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8458 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8461 = (inp[13]) ? node8495 : node8462;
											assign node8462 = (inp[14]) ? node8478 : node8463;
												assign node8463 = (inp[10]) ? node8473 : node8464;
													assign node8464 = (inp[2]) ? node8470 : node8465;
														assign node8465 = (inp[12]) ? node8467 : 16'b0001111111111111;
															assign node8467 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8470 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8473 = (inp[2]) ? 16'b0000011111111111 : node8474;
														assign node8474 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8478 = (inp[2]) ? node8488 : node8479;
													assign node8479 = (inp[12]) ? node8485 : node8480;
														assign node8480 = (inp[10]) ? node8482 : 16'b0001111111111111;
															assign node8482 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8485 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8488 = (inp[12]) ? 16'b0000000111111111 : node8489;
														assign node8489 = (inp[11]) ? 16'b0000001111111111 : node8490;
															assign node8490 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8495 = (inp[14]) ? node8507 : node8496;
												assign node8496 = (inp[2]) ? node8502 : node8497;
													assign node8497 = (inp[10]) ? node8499 : 16'b0000011111111111;
														assign node8499 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8502 = (inp[11]) ? 16'b0000001111111111 : node8503;
														assign node8503 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8507 = (inp[2]) ? node8521 : node8508;
													assign node8508 = (inp[15]) ? node8516 : node8509;
														assign node8509 = (inp[10]) ? 16'b0000001111111111 : node8510;
															assign node8510 = (inp[12]) ? node8512 : 16'b0000011111111111;
																assign node8512 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8516 = (inp[12]) ? 16'b0000000111111111 : node8517;
															assign node8517 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8521 = (inp[11]) ? node8523 : 16'b0000000111111111;
														assign node8523 = (inp[15]) ? 16'b0000000011111111 : node8524;
															assign node8524 = (inp[10]) ? 16'b0000000011111111 : node8525;
																assign node8525 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node8530 = (inp[15]) ? node8578 : node8531;
										assign node8531 = (inp[7]) ? node8551 : node8532;
											assign node8532 = (inp[10]) ? node8540 : node8533;
												assign node8533 = (inp[11]) ? node8535 : 16'b0000111111111111;
													assign node8535 = (inp[12]) ? 16'b0000011111111111 : node8536;
														assign node8536 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8540 = (inp[12]) ? node8548 : node8541;
													assign node8541 = (inp[11]) ? node8545 : node8542;
														assign node8542 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8545 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8548 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8551 = (inp[10]) ? node8569 : node8552;
												assign node8552 = (inp[13]) ? node8556 : node8553;
													assign node8553 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8556 = (inp[11]) ? node8564 : node8557;
														assign node8557 = (inp[14]) ? node8559 : 16'b0000011111111111;
															assign node8559 = (inp[2]) ? 16'b0000001111111111 : node8560;
																assign node8560 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8564 = (inp[14]) ? node8566 : 16'b0000000111111111;
															assign node8566 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8569 = (inp[2]) ? node8571 : 16'b0000001111111111;
													assign node8571 = (inp[13]) ? 16'b0000000111111111 : node8572;
														assign node8572 = (inp[14]) ? node8574 : 16'b0000001111111111;
															assign node8574 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node8578 = (inp[14]) ? node8620 : node8579;
											assign node8579 = (inp[2]) ? node8607 : node8580;
												assign node8580 = (inp[11]) ? node8600 : node8581;
													assign node8581 = (inp[13]) ? node8591 : node8582;
														assign node8582 = (inp[7]) ? node8586 : node8583;
															assign node8583 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node8586 = (inp[12]) ? 16'b0000011111111111 : node8587;
																assign node8587 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8591 = (inp[7]) ? node8593 : 16'b0000011111111111;
															assign node8593 = (inp[10]) ? node8597 : node8594;
																assign node8594 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
																assign node8597 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8600 = (inp[13]) ? 16'b0000001111111111 : node8601;
														assign node8601 = (inp[10]) ? 16'b0000001111111111 : node8602;
															assign node8602 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8607 = (inp[12]) ? node8617 : node8608;
													assign node8608 = (inp[11]) ? node8610 : 16'b0000011111111111;
														assign node8610 = (inp[10]) ? 16'b0000000111111111 : node8611;
															assign node8611 = (inp[7]) ? node8613 : 16'b0000001111111111;
																assign node8613 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8617 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8620 = (inp[7]) ? node8632 : node8621;
												assign node8621 = (inp[11]) ? 16'b0000000111111111 : node8622;
													assign node8622 = (inp[12]) ? node8626 : node8623;
														assign node8623 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node8626 = (inp[2]) ? 16'b0000000111111111 : node8627;
															assign node8627 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8632 = (inp[10]) ? node8638 : node8633;
													assign node8633 = (inp[11]) ? node8635 : 16'b0000001111111111;
														assign node8635 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8638 = (inp[11]) ? node8642 : node8639;
														assign node8639 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8642 = (inp[2]) ? 16'b0000000000111111 : node8643;
															assign node8643 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node8647 = (inp[13]) ? node8773 : node8648;
									assign node8648 = (inp[14]) ? node8712 : node8649;
										assign node8649 = (inp[15]) ? node8679 : node8650;
											assign node8650 = (inp[11]) ? node8664 : node8651;
												assign node8651 = (inp[7]) ? node8657 : node8652;
													assign node8652 = (inp[9]) ? 16'b0000111111111111 : node8653;
														assign node8653 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node8657 = (inp[12]) ? node8661 : node8658;
														assign node8658 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8661 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8664 = (inp[2]) ? node8670 : node8665;
													assign node8665 = (inp[12]) ? node8667 : 16'b0000011111111111;
														assign node8667 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8670 = (inp[9]) ? node8676 : node8671;
														assign node8671 = (inp[10]) ? node8673 : 16'b0000001111111111;
															assign node8673 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8676 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8679 = (inp[9]) ? node8695 : node8680;
												assign node8680 = (inp[7]) ? node8688 : node8681;
													assign node8681 = (inp[11]) ? 16'b0000011111111111 : node8682;
														assign node8682 = (inp[2]) ? 16'b0000011111111111 : node8683;
															assign node8683 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8688 = (inp[12]) ? node8692 : node8689;
														assign node8689 = (inp[10]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node8692 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8695 = (inp[11]) ? node8705 : node8696;
													assign node8696 = (inp[12]) ? node8700 : node8697;
														assign node8697 = (inp[7]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node8700 = (inp[2]) ? node8702 : 16'b0000001111111111;
															assign node8702 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8705 = (inp[12]) ? node8709 : node8706;
														assign node8706 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8709 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8712 = (inp[2]) ? node8746 : node8713;
											assign node8713 = (inp[7]) ? node8735 : node8714;
												assign node8714 = (inp[9]) ? node8726 : node8715;
													assign node8715 = (inp[10]) ? node8719 : node8716;
														assign node8716 = (inp[15]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node8719 = (inp[15]) ? node8721 : 16'b0000011111111111;
															assign node8721 = (inp[12]) ? 16'b0000001111111111 : node8722;
																assign node8722 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8726 = (inp[15]) ? node8732 : node8727;
														assign node8727 = (inp[10]) ? 16'b0000001111111111 : node8728;
															assign node8728 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8732 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8735 = (inp[9]) ? node8743 : node8736;
													assign node8736 = (inp[15]) ? node8738 : 16'b0000001111111111;
														assign node8738 = (inp[10]) ? node8740 : 16'b0000001111111111;
															assign node8740 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8743 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8746 = (inp[9]) ? node8764 : node8747;
												assign node8747 = (inp[10]) ? node8755 : node8748;
													assign node8748 = (inp[7]) ? node8750 : 16'b0000001111111111;
														assign node8750 = (inp[12]) ? 16'b0000000111111111 : node8751;
															assign node8751 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8755 = (inp[11]) ? node8759 : node8756;
														assign node8756 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8759 = (inp[15]) ? node8761 : 16'b0000000111111111;
															assign node8761 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8764 = (inp[10]) ? node8770 : node8765;
													assign node8765 = (inp[11]) ? 16'b0000000011111111 : node8766;
														assign node8766 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8770 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node8773 = (inp[15]) ? node8837 : node8774;
										assign node8774 = (inp[14]) ? node8808 : node8775;
											assign node8775 = (inp[12]) ? node8795 : node8776;
												assign node8776 = (inp[7]) ? node8788 : node8777;
													assign node8777 = (inp[11]) ? node8783 : node8778;
														assign node8778 = (inp[2]) ? 16'b0000011111111111 : node8779;
															assign node8779 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8783 = (inp[9]) ? node8785 : 16'b0000011111111111;
															assign node8785 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8788 = (inp[9]) ? node8792 : node8789;
														assign node8789 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8792 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8795 = (inp[9]) ? node8801 : node8796;
													assign node8796 = (inp[2]) ? node8798 : 16'b0000001111111111;
														assign node8798 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8801 = (inp[10]) ? 16'b0000000011111111 : node8802;
														assign node8802 = (inp[7]) ? node8804 : 16'b0000001111111111;
															assign node8804 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8808 = (inp[11]) ? node8820 : node8809;
												assign node8809 = (inp[10]) ? node8817 : node8810;
													assign node8810 = (inp[2]) ? 16'b0000000111111111 : node8811;
														assign node8811 = (inp[9]) ? 16'b0000001111111111 : node8812;
															assign node8812 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8817 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8820 = (inp[7]) ? node8830 : node8821;
													assign node8821 = (inp[10]) ? node8827 : node8822;
														assign node8822 = (inp[12]) ? 16'b0000000111111111 : node8823;
															assign node8823 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8827 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8830 = (inp[2]) ? 16'b0000000001111111 : node8831;
														assign node8831 = (inp[12]) ? 16'b0000000001111111 : node8832;
															assign node8832 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8837 = (inp[11]) ? node8861 : node8838;
											assign node8838 = (inp[2]) ? node8846 : node8839;
												assign node8839 = (inp[7]) ? node8841 : 16'b0000001111111111;
													assign node8841 = (inp[12]) ? 16'b0000000111111111 : node8842;
														assign node8842 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8846 = (inp[10]) ? node8852 : node8847;
													assign node8847 = (inp[14]) ? 16'b0000000111111111 : node8848;
														assign node8848 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8852 = (inp[7]) ? 16'b0000000011111111 : node8853;
														assign node8853 = (inp[14]) ? node8855 : 16'b0000000111111111;
															assign node8855 = (inp[12]) ? 16'b0000000011111111 : node8856;
																assign node8856 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8861 = (inp[2]) ? node8873 : node8862;
												assign node8862 = (inp[12]) ? node8868 : node8863;
													assign node8863 = (inp[9]) ? node8865 : 16'b0000001111111111;
														assign node8865 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8868 = (inp[7]) ? 16'b0000000011111111 : node8869;
														assign node8869 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8873 = (inp[10]) ? node8875 : 16'b0000000011111111;
													assign node8875 = (inp[14]) ? 16'b0000000000111111 : node8876;
														assign node8876 = (inp[12]) ? 16'b0000000001111111 : node8877;
															assign node8877 = (inp[7]) ? node8879 : 16'b0000000011111111;
																assign node8879 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node8884 = (inp[9]) ? node9150 : node8885;
								assign node8885 = (inp[2]) ? node9021 : node8886;
									assign node8886 = (inp[14]) ? node8960 : node8887;
										assign node8887 = (inp[13]) ? node8919 : node8888;
											assign node8888 = (inp[10]) ? node8906 : node8889;
												assign node8889 = (inp[15]) ? node8897 : node8890;
													assign node8890 = (inp[7]) ? 16'b0000111111111111 : node8891;
														assign node8891 = (inp[12]) ? 16'b0000111111111111 : node8892;
															assign node8892 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node8897 = (inp[3]) ? node8901 : node8898;
														assign node8898 = (inp[11]) ? 16'b0000111111111111 : 16'b0000011111111111;
														assign node8901 = (inp[11]) ? node8903 : 16'b0000011111111111;
															assign node8903 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8906 = (inp[12]) ? node8916 : node8907;
													assign node8907 = (inp[3]) ? node8913 : node8908;
														assign node8908 = (inp[11]) ? 16'b0000011111111111 : node8909;
															assign node8909 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8913 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8916 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8919 = (inp[7]) ? node8933 : node8920;
												assign node8920 = (inp[10]) ? 16'b0000001111111111 : node8921;
													assign node8921 = (inp[3]) ? node8927 : node8922;
														assign node8922 = (inp[11]) ? 16'b0000011111111111 : node8923;
															assign node8923 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8927 = (inp[15]) ? node8929 : 16'b0000011111111111;
															assign node8929 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8933 = (inp[11]) ? node8949 : node8934;
													assign node8934 = (inp[3]) ? node8942 : node8935;
														assign node8935 = (inp[15]) ? 16'b0000011111111111 : node8936;
															assign node8936 = (inp[12]) ? 16'b0000011111111111 : node8937;
																assign node8937 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8942 = (inp[12]) ? 16'b0000000111111111 : node8943;
															assign node8943 = (inp[15]) ? 16'b0000000111111111 : node8944;
																assign node8944 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8949 = (inp[3]) ? node8957 : node8950;
														assign node8950 = (inp[12]) ? node8952 : 16'b0000001111111111;
															assign node8952 = (inp[15]) ? 16'b0000000111111111 : node8953;
																assign node8953 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8957 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8960 = (inp[13]) ? node8998 : node8961;
											assign node8961 = (inp[11]) ? node8975 : node8962;
												assign node8962 = (inp[3]) ? node8972 : node8963;
													assign node8963 = (inp[12]) ? node8967 : node8964;
														assign node8964 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8967 = (inp[15]) ? node8969 : 16'b0000011111111111;
															assign node8969 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8972 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node8975 = (inp[10]) ? node8987 : node8976;
													assign node8976 = (inp[15]) ? node8984 : node8977;
														assign node8977 = (inp[7]) ? node8979 : 16'b0000011111111111;
															assign node8979 = (inp[12]) ? 16'b0000000111111111 : node8980;
																assign node8980 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8984 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8987 = (inp[7]) ? node8993 : node8988;
														assign node8988 = (inp[3]) ? 16'b0000000111111111 : node8989;
															assign node8989 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8993 = (inp[15]) ? node8995 : 16'b0000000111111111;
															assign node8995 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8998 = (inp[15]) ? node9010 : node8999;
												assign node8999 = (inp[11]) ? 16'b0000000111111111 : node9000;
													assign node9000 = (inp[12]) ? node9002 : 16'b0000001111111111;
														assign node9002 = (inp[10]) ? 16'b0000000111111111 : node9003;
															assign node9003 = (inp[3]) ? node9005 : 16'b0000001111111111;
																assign node9005 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9010 = (inp[12]) ? 16'b0000000011111111 : node9011;
													assign node9011 = (inp[10]) ? node9015 : node9012;
														assign node9012 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9015 = (inp[11]) ? node9017 : 16'b0000000111111111;
															assign node9017 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node9021 = (inp[10]) ? node9089 : node9022;
										assign node9022 = (inp[3]) ? node9054 : node9023;
											assign node9023 = (inp[7]) ? node9035 : node9024;
												assign node9024 = (inp[14]) ? node9030 : node9025;
													assign node9025 = (inp[13]) ? 16'b0000011111111111 : node9026;
														assign node9026 = (inp[12]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node9030 = (inp[15]) ? 16'b0000001111111111 : node9031;
														assign node9031 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9035 = (inp[11]) ? node9045 : node9036;
													assign node9036 = (inp[14]) ? node9038 : 16'b0000001111111111;
														assign node9038 = (inp[15]) ? 16'b0000000111111111 : node9039;
															assign node9039 = (inp[13]) ? node9041 : 16'b0000001111111111;
																assign node9041 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9045 = (inp[12]) ? node9049 : node9046;
														assign node9046 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9049 = (inp[14]) ? 16'b0000000011111111 : node9050;
															assign node9050 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9054 = (inp[15]) ? node9076 : node9055;
												assign node9055 = (inp[14]) ? node9063 : node9056;
													assign node9056 = (inp[11]) ? node9060 : node9057;
														assign node9057 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9060 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9063 = (inp[13]) ? node9069 : node9064;
														assign node9064 = (inp[7]) ? node9066 : 16'b0000001111111111;
															assign node9066 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9069 = (inp[7]) ? 16'b0000000111111111 : node9070;
															assign node9070 = (inp[11]) ? 16'b0000000111111111 : node9071;
																assign node9071 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9076 = (inp[13]) ? node9082 : node9077;
													assign node9077 = (inp[12]) ? 16'b0000000111111111 : node9078;
														assign node9078 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9082 = (inp[14]) ? node9084 : 16'b0000000011111111;
														assign node9084 = (inp[12]) ? node9086 : 16'b0000000011111111;
															assign node9086 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9089 = (inp[3]) ? node9131 : node9090;
											assign node9090 = (inp[13]) ? node9106 : node9091;
												assign node9091 = (inp[7]) ? node9101 : node9092;
													assign node9092 = (inp[15]) ? node9096 : node9093;
														assign node9093 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9096 = (inp[14]) ? 16'b0000000111111111 : node9097;
															assign node9097 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9101 = (inp[11]) ? 16'b0000000111111111 : node9102;
														assign node9102 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9106 = (inp[7]) ? node9122 : node9107;
													assign node9107 = (inp[15]) ? node9115 : node9108;
														assign node9108 = (inp[12]) ? 16'b0000000111111111 : node9109;
															assign node9109 = (inp[11]) ? node9111 : 16'b0000001111111111;
																assign node9111 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9115 = (inp[11]) ? node9117 : 16'b0000000111111111;
															assign node9117 = (inp[14]) ? 16'b0000000011111111 : node9118;
																assign node9118 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9122 = (inp[12]) ? node9128 : node9123;
														assign node9123 = (inp[11]) ? 16'b0000000011111111 : node9124;
															assign node9124 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9128 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node9131 = (inp[11]) ? node9139 : node9132;
												assign node9132 = (inp[12]) ? 16'b0000000011111111 : node9133;
													assign node9133 = (inp[13]) ? node9135 : 16'b0000001111111111;
														assign node9135 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9139 = (inp[13]) ? node9143 : node9140;
													assign node9140 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node9143 = (inp[14]) ? node9145 : 16'b0000000011111111;
														assign node9145 = (inp[12]) ? 16'b0000000000111111 : node9146;
															assign node9146 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node9150 = (inp[11]) ? node9274 : node9151;
									assign node9151 = (inp[2]) ? node9213 : node9152;
										assign node9152 = (inp[13]) ? node9190 : node9153;
											assign node9153 = (inp[3]) ? node9169 : node9154;
												assign node9154 = (inp[7]) ? node9166 : node9155;
													assign node9155 = (inp[14]) ? node9163 : node9156;
														assign node9156 = (inp[10]) ? node9158 : 16'b0000111111111111;
															assign node9158 = (inp[12]) ? 16'b0000011111111111 : node9159;
																assign node9159 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9163 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9166 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9169 = (inp[14]) ? node9179 : node9170;
													assign node9170 = (inp[15]) ? node9174 : node9171;
														assign node9171 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9174 = (inp[10]) ? node9176 : 16'b0000001111111111;
															assign node9176 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9179 = (inp[7]) ? node9185 : node9180;
														assign node9180 = (inp[15]) ? 16'b0000000111111111 : node9181;
															assign node9181 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9185 = (inp[12]) ? 16'b0000000011111111 : node9186;
															assign node9186 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9190 = (inp[14]) ? node9202 : node9191;
												assign node9191 = (inp[12]) ? node9195 : node9192;
													assign node9192 = (inp[7]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node9195 = (inp[3]) ? node9199 : node9196;
														assign node9196 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9199 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9202 = (inp[15]) ? node9204 : 16'b0000000111111111;
													assign node9204 = (inp[12]) ? node9210 : node9205;
														assign node9205 = (inp[10]) ? 16'b0000000011111111 : node9206;
															assign node9206 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9210 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node9213 = (inp[15]) ? node9251 : node9214;
											assign node9214 = (inp[10]) ? node9230 : node9215;
												assign node9215 = (inp[13]) ? node9225 : node9216;
													assign node9216 = (inp[7]) ? node9220 : node9217;
														assign node9217 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9220 = (inp[3]) ? 16'b0000000111111111 : node9221;
															assign node9221 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9225 = (inp[14]) ? node9227 : 16'b0000000111111111;
														assign node9227 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9230 = (inp[3]) ? node9242 : node9231;
													assign node9231 = (inp[14]) ? node9239 : node9232;
														assign node9232 = (inp[12]) ? 16'b0000000111111111 : node9233;
															assign node9233 = (inp[13]) ? node9235 : 16'b0000001111111111;
																assign node9235 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9239 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9242 = (inp[7]) ? 16'b0000000011111111 : node9243;
														assign node9243 = (inp[14]) ? node9245 : 16'b0000000111111111;
															assign node9245 = (inp[12]) ? 16'b0000000011111111 : node9246;
																assign node9246 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9251 = (inp[7]) ? node9263 : node9252;
												assign node9252 = (inp[3]) ? node9254 : 16'b0000000111111111;
													assign node9254 = (inp[13]) ? 16'b0000000011111111 : node9255;
														assign node9255 = (inp[12]) ? node9257 : 16'b0000000111111111;
															assign node9257 = (inp[14]) ? node9259 : 16'b0000000111111111;
																assign node9259 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9263 = (inp[10]) ? 16'b0000000001111111 : node9264;
													assign node9264 = (inp[3]) ? node9270 : node9265;
														assign node9265 = (inp[13]) ? node9267 : 16'b0000000111111111;
															assign node9267 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9270 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node9274 = (inp[12]) ? node9334 : node9275;
										assign node9275 = (inp[14]) ? node9309 : node9276;
											assign node9276 = (inp[13]) ? node9292 : node9277;
												assign node9277 = (inp[15]) ? node9287 : node9278;
													assign node9278 = (inp[3]) ? node9284 : node9279;
														assign node9279 = (inp[10]) ? node9281 : 16'b0000011111111111;
															assign node9281 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9284 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9287 = (inp[10]) ? 16'b0000000111111111 : node9288;
														assign node9288 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9292 = (inp[10]) ? node9298 : node9293;
													assign node9293 = (inp[2]) ? 16'b0000000111111111 : node9294;
														assign node9294 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9298 = (inp[3]) ? node9300 : 16'b0000000111111111;
														assign node9300 = (inp[7]) ? node9306 : node9301;
															assign node9301 = (inp[15]) ? 16'b0000000011111111 : node9302;
																assign node9302 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node9306 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9309 = (inp[13]) ? node9325 : node9310;
												assign node9310 = (inp[7]) ? node9322 : node9311;
													assign node9311 = (inp[15]) ? node9317 : node9312;
														assign node9312 = (inp[3]) ? 16'b0000000111111111 : node9313;
															assign node9313 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9317 = (inp[3]) ? 16'b0000000001111111 : node9318;
															assign node9318 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9322 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9325 = (inp[2]) ? node9331 : node9326;
													assign node9326 = (inp[3]) ? node9328 : 16'b0000000011111111;
														assign node9328 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node9331 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9334 = (inp[3]) ? node9370 : node9335;
											assign node9335 = (inp[2]) ? node9355 : node9336;
												assign node9336 = (inp[7]) ? node9346 : node9337;
													assign node9337 = (inp[15]) ? node9341 : node9338;
														assign node9338 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9341 = (inp[13]) ? node9343 : 16'b0000000111111111;
															assign node9343 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9346 = (inp[15]) ? node9348 : 16'b0000000111111111;
														assign node9348 = (inp[14]) ? 16'b0000000001111111 : node9349;
															assign node9349 = (inp[13]) ? node9351 : 16'b0000000011111111;
																assign node9351 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9355 = (inp[10]) ? node9363 : node9356;
													assign node9356 = (inp[13]) ? node9360 : node9357;
														assign node9357 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9360 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9363 = (inp[15]) ? 16'b0000000000111111 : node9364;
														assign node9364 = (inp[14]) ? 16'b0000000001111111 : node9365;
															assign node9365 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9370 = (inp[14]) ? node9384 : node9371;
												assign node9371 = (inp[10]) ? node9379 : node9372;
													assign node9372 = (inp[2]) ? node9374 : 16'b0000000111111111;
														assign node9374 = (inp[13]) ? node9376 : 16'b0000000011111111;
															assign node9376 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9379 = (inp[15]) ? node9381 : 16'b0000000001111111;
														assign node9381 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9384 = (inp[2]) ? node9392 : node9385;
													assign node9385 = (inp[13]) ? node9387 : 16'b0000000001111111;
														assign node9387 = (inp[10]) ? node9389 : 16'b0000000000111111;
															assign node9389 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node9392 = (inp[15]) ? node9398 : node9393;
														assign node9393 = (inp[7]) ? 16'b0000000000011111 : node9394;
															assign node9394 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9398 = (inp[7]) ? node9400 : 16'b0000000000011111;
															assign node9400 = (inp[13]) ? node9402 : 16'b0000000000011111;
																assign node9402 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node9405 = (inp[6]) ? node9961 : node9406;
							assign node9406 = (inp[10]) ? node9702 : node9407;
								assign node9407 = (inp[3]) ? node9557 : node9408;
									assign node9408 = (inp[2]) ? node9480 : node9409;
										assign node9409 = (inp[12]) ? node9447 : node9410;
											assign node9410 = (inp[11]) ? node9426 : node9411;
												assign node9411 = (inp[9]) ? node9419 : node9412;
													assign node9412 = (inp[15]) ? node9414 : 16'b0000111111111111;
														assign node9414 = (inp[13]) ? node9416 : 16'b0000111111111111;
															assign node9416 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9419 = (inp[15]) ? 16'b0000000111111111 : node9420;
														assign node9420 = (inp[14]) ? 16'b0000011111111111 : node9421;
															assign node9421 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node9426 = (inp[15]) ? node9436 : node9427;
													assign node9427 = (inp[14]) ? node9429 : 16'b0000111111111111;
														assign node9429 = (inp[13]) ? node9431 : 16'b0000011111111111;
															assign node9431 = (inp[9]) ? 16'b0000001111111111 : node9432;
																assign node9432 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9436 = (inp[14]) ? node9444 : node9437;
														assign node9437 = (inp[13]) ? 16'b0000001111111111 : node9438;
															assign node9438 = (inp[7]) ? node9440 : 16'b0000011111111111;
																assign node9440 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9444 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9447 = (inp[11]) ? node9461 : node9448;
												assign node9448 = (inp[14]) ? node9456 : node9449;
													assign node9449 = (inp[15]) ? 16'b0000001111111111 : node9450;
														assign node9450 = (inp[13]) ? 16'b0000011111111111 : node9451;
															assign node9451 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9456 = (inp[13]) ? 16'b0000001111111111 : node9457;
														assign node9457 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9461 = (inp[9]) ? node9469 : node9462;
													assign node9462 = (inp[13]) ? node9464 : 16'b0000011111111111;
														assign node9464 = (inp[15]) ? 16'b0000000111111111 : node9465;
															assign node9465 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9469 = (inp[13]) ? node9473 : node9470;
														assign node9470 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9473 = (inp[7]) ? node9475 : 16'b0000000111111111;
															assign node9475 = (inp[15]) ? 16'b0000000011111111 : node9476;
																assign node9476 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9480 = (inp[11]) ? node9520 : node9481;
											assign node9481 = (inp[15]) ? node9499 : node9482;
												assign node9482 = (inp[7]) ? node9490 : node9483;
													assign node9483 = (inp[14]) ? 16'b0000011111111111 : node9484;
														assign node9484 = (inp[12]) ? 16'b0000011111111111 : node9485;
															assign node9485 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9490 = (inp[9]) ? node9496 : node9491;
														assign node9491 = (inp[13]) ? 16'b0000001111111111 : node9492;
															assign node9492 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9496 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9499 = (inp[12]) ? node9509 : node9500;
													assign node9500 = (inp[14]) ? node9502 : 16'b0000001111111111;
														assign node9502 = (inp[7]) ? node9504 : 16'b0000001111111111;
															assign node9504 = (inp[9]) ? 16'b0000000111111111 : node9505;
																assign node9505 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9509 = (inp[14]) ? node9513 : node9510;
														assign node9510 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node9513 = (inp[13]) ? 16'b0000000111111111 : node9514;
															assign node9514 = (inp[9]) ? 16'b0000000111111111 : node9515;
																assign node9515 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9520 = (inp[14]) ? node9540 : node9521;
												assign node9521 = (inp[7]) ? node9527 : node9522;
													assign node9522 = (inp[12]) ? 16'b0000011111111111 : node9523;
														assign node9523 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9527 = (inp[9]) ? node9535 : node9528;
														assign node9528 = (inp[15]) ? 16'b0000000111111111 : node9529;
															assign node9529 = (inp[13]) ? node9531 : 16'b0000001111111111;
																assign node9531 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9535 = (inp[13]) ? 16'b0000000011111111 : node9536;
															assign node9536 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9540 = (inp[9]) ? node9550 : node9541;
													assign node9541 = (inp[13]) ? node9543 : 16'b0000000111111111;
														assign node9543 = (inp[15]) ? node9545 : 16'b0000000111111111;
															assign node9545 = (inp[12]) ? 16'b0000000011111111 : node9546;
																assign node9546 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9550 = (inp[7]) ? node9554 : node9551;
														assign node9551 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9554 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9557 = (inp[14]) ? node9633 : node9558;
										assign node9558 = (inp[9]) ? node9596 : node9559;
											assign node9559 = (inp[2]) ? node9573 : node9560;
												assign node9560 = (inp[7]) ? node9568 : node9561;
													assign node9561 = (inp[11]) ? node9565 : node9562;
														assign node9562 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9565 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9568 = (inp[15]) ? 16'b0000001111111111 : node9569;
														assign node9569 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9573 = (inp[12]) ? node9583 : node9574;
													assign node9574 = (inp[15]) ? node9578 : node9575;
														assign node9575 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9578 = (inp[13]) ? node9580 : 16'b0000001111111111;
															assign node9580 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9583 = (inp[13]) ? node9591 : node9584;
														assign node9584 = (inp[7]) ? node9586 : 16'b0000001111111111;
															assign node9586 = (inp[11]) ? node9588 : 16'b0000001111111111;
																assign node9588 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9591 = (inp[11]) ? node9593 : 16'b0000000111111111;
															assign node9593 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9596 = (inp[2]) ? node9618 : node9597;
												assign node9597 = (inp[7]) ? node9609 : node9598;
													assign node9598 = (inp[12]) ? node9602 : node9599;
														assign node9599 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9602 = (inp[13]) ? 16'b0000000111111111 : node9603;
															assign node9603 = (inp[15]) ? node9605 : 16'b0000001111111111;
																assign node9605 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9609 = (inp[12]) ? node9615 : node9610;
														assign node9610 = (inp[11]) ? 16'b0000000111111111 : node9611;
															assign node9611 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9615 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9618 = (inp[15]) ? node9628 : node9619;
													assign node9619 = (inp[13]) ? node9623 : node9620;
														assign node9620 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9623 = (inp[12]) ? node9625 : 16'b0000000111111111;
															assign node9625 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9628 = (inp[13]) ? 16'b0000000011111111 : node9629;
														assign node9629 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9633 = (inp[7]) ? node9669 : node9634;
											assign node9634 = (inp[11]) ? node9654 : node9635;
												assign node9635 = (inp[2]) ? node9645 : node9636;
													assign node9636 = (inp[13]) ? node9638 : 16'b0000001111111111;
														assign node9638 = (inp[9]) ? node9640 : 16'b0000001111111111;
															assign node9640 = (inp[15]) ? 16'b0000000111111111 : node9641;
																assign node9641 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9645 = (inp[13]) ? node9651 : node9646;
														assign node9646 = (inp[12]) ? 16'b0000000111111111 : node9647;
															assign node9647 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9651 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9654 = (inp[9]) ? node9662 : node9655;
													assign node9655 = (inp[15]) ? node9659 : node9656;
														assign node9656 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9659 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9662 = (inp[13]) ? node9666 : node9663;
														assign node9663 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9666 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9669 = (inp[11]) ? node9695 : node9670;
												assign node9670 = (inp[2]) ? node9678 : node9671;
													assign node9671 = (inp[9]) ? node9675 : node9672;
														assign node9672 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9675 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9678 = (inp[15]) ? node9688 : node9679;
														assign node9679 = (inp[9]) ? node9685 : node9680;
															assign node9680 = (inp[13]) ? node9682 : 16'b0000000111111111;
																assign node9682 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node9685 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9688 = (inp[12]) ? 16'b0000000001111111 : node9689;
															assign node9689 = (inp[13]) ? node9691 : 16'b0000000011111111;
																assign node9691 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9695 = (inp[2]) ? node9699 : node9696;
													assign node9696 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9699 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node9702 = (inp[11]) ? node9844 : node9703;
									assign node9703 = (inp[7]) ? node9781 : node9704;
										assign node9704 = (inp[13]) ? node9742 : node9705;
											assign node9705 = (inp[12]) ? node9729 : node9706;
												assign node9706 = (inp[3]) ? node9720 : node9707;
													assign node9707 = (inp[14]) ? node9715 : node9708;
														assign node9708 = (inp[9]) ? 16'b0000111111111111 : node9709;
															assign node9709 = (inp[2]) ? 16'b0000111111111111 : node9710;
																assign node9710 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node9715 = (inp[2]) ? node9717 : 16'b0000011111111111;
															assign node9717 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9720 = (inp[15]) ? node9724 : node9721;
														assign node9721 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9724 = (inp[2]) ? node9726 : 16'b0000001111111111;
															assign node9726 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node9729 = (inp[15]) ? node9737 : node9730;
													assign node9730 = (inp[14]) ? node9734 : node9731;
														assign node9731 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9734 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9737 = (inp[9]) ? node9739 : 16'b0000000111111111;
														assign node9739 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9742 = (inp[9]) ? node9768 : node9743;
												assign node9743 = (inp[3]) ? node9757 : node9744;
													assign node9744 = (inp[12]) ? 16'b0000000011111111 : node9745;
														assign node9745 = (inp[2]) ? node9751 : node9746;
															assign node9746 = (inp[14]) ? node9748 : 16'b0000011111111111;
																assign node9748 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node9751 = (inp[14]) ? node9753 : 16'b0000001111111111;
																assign node9753 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9757 = (inp[14]) ? node9761 : node9758;
														assign node9758 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9761 = (inp[15]) ? node9763 : 16'b0000000111111111;
															assign node9763 = (inp[12]) ? 16'b0000000011111111 : node9764;
																assign node9764 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9768 = (inp[14]) ? node9776 : node9769;
													assign node9769 = (inp[15]) ? node9773 : node9770;
														assign node9770 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9773 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9776 = (inp[15]) ? node9778 : 16'b0000000011111111;
														assign node9778 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9781 = (inp[14]) ? node9809 : node9782;
											assign node9782 = (inp[13]) ? node9792 : node9783;
												assign node9783 = (inp[9]) ? node9787 : node9784;
													assign node9784 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9787 = (inp[3]) ? 16'b0000000011111111 : node9788;
														assign node9788 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9792 = (inp[3]) ? node9806 : node9793;
													assign node9793 = (inp[15]) ? node9799 : node9794;
														assign node9794 = (inp[12]) ? 16'b0000000111111111 : node9795;
															assign node9795 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9799 = (inp[2]) ? node9801 : 16'b0000001111111111;
															assign node9801 = (inp[12]) ? 16'b0000000011111111 : node9802;
																assign node9802 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9806 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9809 = (inp[2]) ? node9829 : node9810;
												assign node9810 = (inp[12]) ? node9820 : node9811;
													assign node9811 = (inp[9]) ? node9815 : node9812;
														assign node9812 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9815 = (inp[13]) ? node9817 : 16'b0000000111111111;
															assign node9817 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9820 = (inp[3]) ? 16'b0000000011111111 : node9821;
														assign node9821 = (inp[15]) ? 16'b0000000011111111 : node9822;
															assign node9822 = (inp[9]) ? node9824 : 16'b0000001111111111;
																assign node9824 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9829 = (inp[13]) ? node9835 : node9830;
													assign node9830 = (inp[12]) ? node9832 : 16'b0000000111111111;
														assign node9832 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9835 = (inp[9]) ? node9841 : node9836;
														assign node9836 = (inp[3]) ? 16'b0000000001111111 : node9837;
															assign node9837 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9841 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node9844 = (inp[15]) ? node9916 : node9845;
										assign node9845 = (inp[2]) ? node9873 : node9846;
											assign node9846 = (inp[14]) ? node9862 : node9847;
												assign node9847 = (inp[9]) ? node9853 : node9848;
													assign node9848 = (inp[7]) ? 16'b0000000111111111 : node9849;
														assign node9849 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9853 = (inp[12]) ? 16'b0000000111111111 : node9854;
														assign node9854 = (inp[13]) ? 16'b0000000111111111 : node9855;
															assign node9855 = (inp[7]) ? node9857 : 16'b0000001111111111;
																assign node9857 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9862 = (inp[12]) ? node9866 : node9863;
													assign node9863 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node9866 = (inp[9]) ? node9870 : node9867;
														assign node9867 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9870 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9873 = (inp[3]) ? node9893 : node9874;
												assign node9874 = (inp[12]) ? node9884 : node9875;
													assign node9875 = (inp[14]) ? node9881 : node9876;
														assign node9876 = (inp[7]) ? node9878 : 16'b0000001111111111;
															assign node9878 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9881 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node9884 = (inp[13]) ? 16'b0000000001111111 : node9885;
														assign node9885 = (inp[9]) ? node9887 : 16'b0000000111111111;
															assign node9887 = (inp[7]) ? 16'b0000000011111111 : node9888;
																assign node9888 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9893 = (inp[12]) ? node9905 : node9894;
													assign node9894 = (inp[13]) ? node9900 : node9895;
														assign node9895 = (inp[14]) ? 16'b0000000011111111 : node9896;
															assign node9896 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9900 = (inp[9]) ? node9902 : 16'b0000000011111111;
															assign node9902 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9905 = (inp[14]) ? node9913 : node9906;
														assign node9906 = (inp[7]) ? 16'b0000000001111111 : node9907;
															assign node9907 = (inp[13]) ? node9909 : 16'b0000000011111111;
																assign node9909 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9913 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9916 = (inp[7]) ? node9938 : node9917;
											assign node9917 = (inp[3]) ? node9929 : node9918;
												assign node9918 = (inp[12]) ? 16'b0000000011111111 : node9919;
													assign node9919 = (inp[13]) ? 16'b0000000011111111 : node9920;
														assign node9920 = (inp[9]) ? node9922 : 16'b0000000111111111;
															assign node9922 = (inp[2]) ? node9924 : 16'b0000000111111111;
																assign node9924 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9929 = (inp[14]) ? node9931 : 16'b0000000011111111;
													assign node9931 = (inp[13]) ? node9935 : node9932;
														assign node9932 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9935 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9938 = (inp[14]) ? node9948 : node9939;
												assign node9939 = (inp[9]) ? 16'b0000000001111111 : node9940;
													assign node9940 = (inp[13]) ? node9944 : node9941;
														assign node9941 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9944 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9948 = (inp[12]) ? node9956 : node9949;
													assign node9949 = (inp[3]) ? node9953 : node9950;
														assign node9950 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node9953 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9956 = (inp[2]) ? node9958 : 16'b0000000000111111;
														assign node9958 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node9961 = (inp[13]) ? node10211 : node9962;
								assign node9962 = (inp[2]) ? node10090 : node9963;
									assign node9963 = (inp[9]) ? node10029 : node9964;
										assign node9964 = (inp[15]) ? node9998 : node9965;
											assign node9965 = (inp[14]) ? node9983 : node9966;
												assign node9966 = (inp[11]) ? node9974 : node9967;
													assign node9967 = (inp[7]) ? node9971 : node9968;
														assign node9968 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9971 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9974 = (inp[12]) ? node9978 : node9975;
														assign node9975 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9978 = (inp[3]) ? node9980 : 16'b0000001111111111;
															assign node9980 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9983 = (inp[7]) ? node9985 : 16'b0000001111111111;
													assign node9985 = (inp[3]) ? node9993 : node9986;
														assign node9986 = (inp[11]) ? 16'b0000000111111111 : node9987;
															assign node9987 = (inp[12]) ? 16'b0000001111111111 : node9988;
																assign node9988 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9993 = (inp[12]) ? 16'b0000000111111111 : node9994;
															assign node9994 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9998 = (inp[3]) ? node10016 : node9999;
												assign node9999 = (inp[12]) ? node10009 : node10000;
													assign node10000 = (inp[7]) ? node10006 : node10001;
														assign node10001 = (inp[11]) ? node10003 : 16'b0000011111111111;
															assign node10003 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10006 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10009 = (inp[7]) ? node10013 : node10010;
														assign node10010 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10013 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10016 = (inp[14]) ? node10024 : node10017;
													assign node10017 = (inp[11]) ? node10019 : 16'b0000000111111111;
														assign node10019 = (inp[12]) ? 16'b0000000011111111 : node10020;
															assign node10020 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10024 = (inp[10]) ? node10026 : 16'b0000000011111111;
														assign node10026 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10029 = (inp[11]) ? node10063 : node10030;
											assign node10030 = (inp[10]) ? node10044 : node10031;
												assign node10031 = (inp[12]) ? node10041 : node10032;
													assign node10032 = (inp[15]) ? node10038 : node10033;
														assign node10033 = (inp[3]) ? 16'b0000001111111111 : node10034;
															assign node10034 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10038 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10041 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10044 = (inp[7]) ? node10056 : node10045;
													assign node10045 = (inp[3]) ? node10053 : node10046;
														assign node10046 = (inp[15]) ? 16'b0000000111111111 : node10047;
															assign node10047 = (inp[12]) ? node10049 : 16'b0000011111111111;
																assign node10049 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10053 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10056 = (inp[12]) ? node10060 : node10057;
														assign node10057 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10060 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10063 = (inp[3]) ? node10077 : node10064;
												assign node10064 = (inp[7]) ? node10070 : node10065;
													assign node10065 = (inp[15]) ? node10067 : 16'b0000000111111111;
														assign node10067 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10070 = (inp[14]) ? node10074 : node10071;
														assign node10071 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10074 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10077 = (inp[15]) ? node10087 : node10078;
													assign node10078 = (inp[10]) ? node10084 : node10079;
														assign node10079 = (inp[14]) ? 16'b0000000011111111 : node10080;
															assign node10080 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10084 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node10087 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10090 = (inp[14]) ? node10150 : node10091;
										assign node10091 = (inp[12]) ? node10123 : node10092;
											assign node10092 = (inp[15]) ? node10108 : node10093;
												assign node10093 = (inp[9]) ? node10097 : node10094;
													assign node10094 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10097 = (inp[11]) ? node10105 : node10098;
														assign node10098 = (inp[10]) ? 16'b0000000111111111 : node10099;
															assign node10099 = (inp[7]) ? node10101 : 16'b0000001111111111;
																assign node10101 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10105 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10108 = (inp[10]) ? node10120 : node10109;
													assign node10109 = (inp[9]) ? node10115 : node10110;
														assign node10110 = (inp[11]) ? node10112 : 16'b0000001111111111;
															assign node10112 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10115 = (inp[3]) ? 16'b0000000011111111 : node10116;
															assign node10116 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10120 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node10123 = (inp[9]) ? node10141 : node10124;
												assign node10124 = (inp[15]) ? node10130 : node10125;
													assign node10125 = (inp[3]) ? node10127 : 16'b0000000111111111;
														assign node10127 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10130 = (inp[3]) ? node10136 : node10131;
														assign node10131 = (inp[7]) ? 16'b0000000011111111 : node10132;
															assign node10132 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10136 = (inp[7]) ? node10138 : 16'b0000000011111111;
															assign node10138 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10141 = (inp[3]) ? node10147 : node10142;
													assign node10142 = (inp[10]) ? node10144 : 16'b0000000111111111;
														assign node10144 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node10147 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10150 = (inp[3]) ? node10176 : node10151;
											assign node10151 = (inp[15]) ? node10161 : node10152;
												assign node10152 = (inp[10]) ? node10158 : node10153;
													assign node10153 = (inp[7]) ? node10155 : 16'b0000000111111111;
														assign node10155 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10158 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10161 = (inp[10]) ? node10167 : node10162;
													assign node10162 = (inp[9]) ? 16'b0000000011111111 : node10163;
														assign node10163 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10167 = (inp[11]) ? node10171 : node10168;
														assign node10168 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10171 = (inp[9]) ? node10173 : 16'b0000000001111111;
															assign node10173 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10176 = (inp[15]) ? node10188 : node10177;
												assign node10177 = (inp[11]) ? node10181 : node10178;
													assign node10178 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10181 = (inp[9]) ? node10183 : 16'b0000000001111111;
														assign node10183 = (inp[12]) ? 16'b0000000000111111 : node10184;
															assign node10184 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10188 = (inp[12]) ? node10198 : node10189;
													assign node10189 = (inp[9]) ? node10191 : 16'b0000000001111111;
														assign node10191 = (inp[10]) ? node10193 : 16'b0000000001111111;
															assign node10193 = (inp[7]) ? node10195 : 16'b0000000000111111;
																assign node10195 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10198 = (inp[7]) ? node10200 : 16'b0000000000111111;
														assign node10200 = (inp[11]) ? node10206 : node10201;
															assign node10201 = (inp[10]) ? node10203 : 16'b0000000000111111;
																assign node10203 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node10206 = (inp[9]) ? node10208 : 16'b0000000000011111;
																assign node10208 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node10211 = (inp[10]) ? node10329 : node10212;
									assign node10212 = (inp[12]) ? node10268 : node10213;
										assign node10213 = (inp[3]) ? node10243 : node10214;
											assign node10214 = (inp[9]) ? node10226 : node10215;
												assign node10215 = (inp[7]) ? node10219 : node10216;
													assign node10216 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10219 = (inp[14]) ? node10221 : 16'b0000001111111111;
														assign node10221 = (inp[11]) ? 16'b0000000111111111 : node10222;
															assign node10222 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10226 = (inp[14]) ? node10240 : node10227;
													assign node10227 = (inp[11]) ? node10235 : node10228;
														assign node10228 = (inp[7]) ? 16'b0000000111111111 : node10229;
															assign node10229 = (inp[2]) ? node10231 : 16'b0000001111111111;
																assign node10231 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10235 = (inp[15]) ? node10237 : 16'b0000000111111111;
															assign node10237 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10240 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10243 = (inp[7]) ? node10255 : node10244;
												assign node10244 = (inp[11]) ? node10250 : node10245;
													assign node10245 = (inp[9]) ? node10247 : 16'b0000000111111111;
														assign node10247 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10250 = (inp[2]) ? 16'b0000000011111111 : node10251;
														assign node10251 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node10255 = (inp[14]) ? node10261 : node10256;
													assign node10256 = (inp[11]) ? 16'b0000000001111111 : node10257;
														assign node10257 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10261 = (inp[9]) ? node10265 : node10262;
														assign node10262 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10265 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10268 = (inp[3]) ? node10306 : node10269;
											assign node10269 = (inp[15]) ? node10287 : node10270;
												assign node10270 = (inp[2]) ? node10278 : node10271;
													assign node10271 = (inp[11]) ? node10275 : node10272;
														assign node10272 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10275 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10278 = (inp[11]) ? node10282 : node10279;
														assign node10279 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node10282 = (inp[7]) ? node10284 : 16'b0000000011111111;
															assign node10284 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10287 = (inp[14]) ? node10299 : node10288;
													assign node10288 = (inp[9]) ? node10290 : 16'b0000001111111111;
														assign node10290 = (inp[11]) ? 16'b0000000001111111 : node10291;
															assign node10291 = (inp[2]) ? node10295 : node10292;
																assign node10292 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node10295 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10299 = (inp[9]) ? node10301 : 16'b0000000001111111;
														assign node10301 = (inp[2]) ? 16'b0000000000111111 : node10302;
															assign node10302 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10306 = (inp[14]) ? node10322 : node10307;
												assign node10307 = (inp[2]) ? node10313 : node10308;
													assign node10308 = (inp[7]) ? node10310 : 16'b0000000011111111;
														assign node10310 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10313 = (inp[7]) ? node10315 : 16'b0000000001111111;
														assign node10315 = (inp[15]) ? 16'b0000000000011111 : node10316;
															assign node10316 = (inp[11]) ? node10318 : 16'b0000000001111111;
																assign node10318 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10322 = (inp[11]) ? node10324 : 16'b0000000000011111;
													assign node10324 = (inp[15]) ? 16'b0000000000111111 : node10325;
														assign node10325 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10329 = (inp[7]) ? node10405 : node10330;
										assign node10330 = (inp[12]) ? node10358 : node10331;
											assign node10331 = (inp[15]) ? node10349 : node10332;
												assign node10332 = (inp[3]) ? node10342 : node10333;
													assign node10333 = (inp[9]) ? node10339 : node10334;
														assign node10334 = (inp[2]) ? node10336 : 16'b0000011111111111;
															assign node10336 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10339 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10342 = (inp[11]) ? node10346 : node10343;
														assign node10343 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10346 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10349 = (inp[2]) ? node10353 : node10350;
													assign node10350 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10353 = (inp[9]) ? node10355 : 16'b0000000011111111;
														assign node10355 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10358 = (inp[15]) ? node10378 : node10359;
												assign node10359 = (inp[2]) ? node10369 : node10360;
													assign node10360 = (inp[3]) ? node10366 : node10361;
														assign node10361 = (inp[11]) ? node10363 : 16'b0000000111111111;
															assign node10363 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10366 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node10369 = (inp[14]) ? node10375 : node10370;
														assign node10370 = (inp[11]) ? 16'b0000000001111111 : node10371;
															assign node10371 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10375 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10378 = (inp[11]) ? node10392 : node10379;
													assign node10379 = (inp[3]) ? node10385 : node10380;
														assign node10380 = (inp[9]) ? node10382 : 16'b0000000011111111;
															assign node10382 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10385 = (inp[9]) ? 16'b0000000000111111 : node10386;
															assign node10386 = (inp[14]) ? node10388 : 16'b0000000001111111;
																assign node10388 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10392 = (inp[9]) ? node10398 : node10393;
														assign node10393 = (inp[2]) ? 16'b0000000000111111 : node10394;
															assign node10394 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10398 = (inp[3]) ? 16'b0000000000001111 : node10399;
															assign node10399 = (inp[14]) ? node10401 : 16'b0000000000111111;
																assign node10401 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10405 = (inp[3]) ? node10441 : node10406;
											assign node10406 = (inp[9]) ? node10420 : node10407;
												assign node10407 = (inp[15]) ? node10409 : 16'b0000000011111111;
													assign node10409 = (inp[14]) ? node10415 : node10410;
														assign node10410 = (inp[2]) ? node10412 : 16'b0000000011111111;
															assign node10412 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10415 = (inp[2]) ? 16'b0000000001111111 : node10416;
															assign node10416 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10420 = (inp[15]) ? node10426 : node10421;
													assign node10421 = (inp[14]) ? node10423 : 16'b0000000001111111;
														assign node10423 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10426 = (inp[2]) ? node10434 : node10427;
														assign node10427 = (inp[12]) ? 16'b0000000000111111 : node10428;
															assign node10428 = (inp[11]) ? node10430 : 16'b0000000001111111;
																assign node10430 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10434 = (inp[14]) ? 16'b0000000000011111 : node10435;
															assign node10435 = (inp[11]) ? node10437 : 16'b0000000000111111;
																assign node10437 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10441 = (inp[12]) ? node10461 : node10442;
												assign node10442 = (inp[15]) ? node10452 : node10443;
													assign node10443 = (inp[11]) ? node10445 : 16'b0000000001111111;
														assign node10445 = (inp[14]) ? node10447 : 16'b0000000001111111;
															assign node10447 = (inp[2]) ? 16'b0000000000111111 : node10448;
																assign node10448 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10452 = (inp[11]) ? node10456 : node10453;
														assign node10453 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10456 = (inp[14]) ? 16'b0000000000011111 : node10457;
															assign node10457 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10461 = (inp[2]) ? node10479 : node10462;
													assign node10462 = (inp[11]) ? node10472 : node10463;
														assign node10463 = (inp[9]) ? node10469 : node10464;
															assign node10464 = (inp[14]) ? node10466 : 16'b0000000001111111;
																assign node10466 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node10469 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node10472 = (inp[14]) ? 16'b0000000000011111 : node10473;
															assign node10473 = (inp[15]) ? node10475 : 16'b0000000000111111;
																assign node10475 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10479 = (inp[15]) ? node10481 : 16'b0000000000011111;
														assign node10481 = (inp[14]) ? 16'b0000000000001111 : node10482;
															assign node10482 = (inp[11]) ? node10484 : 16'b0000000000011111;
																assign node10484 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node10488 = (inp[11]) ? node11526 : node10489;
						assign node10489 = (inp[15]) ? node11037 : node10490;
							assign node10490 = (inp[6]) ? node10754 : node10491;
								assign node10491 = (inp[13]) ? node10631 : node10492;
									assign node10492 = (inp[2]) ? node10558 : node10493;
										assign node10493 = (inp[10]) ? node10515 : node10494;
											assign node10494 = (inp[14]) ? node10506 : node10495;
												assign node10495 = (inp[12]) ? node10501 : node10496;
													assign node10496 = (inp[3]) ? 16'b0000111111111111 : node10497;
														assign node10497 = (inp[7]) ? 16'b0000111111111111 : 16'b0011111111111111;
													assign node10501 = (inp[7]) ? 16'b0000011111111111 : node10502;
														assign node10502 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node10506 = (inp[9]) ? node10510 : node10507;
													assign node10507 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node10510 = (inp[12]) ? 16'b0000001111111111 : node10511;
														assign node10511 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node10515 = (inp[9]) ? node10535 : node10516;
												assign node10516 = (inp[7]) ? node10528 : node10517;
													assign node10517 = (inp[1]) ? node10521 : node10518;
														assign node10518 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node10521 = (inp[14]) ? node10523 : 16'b0000011111111111;
															assign node10523 = (inp[3]) ? 16'b0000001111111111 : node10524;
																assign node10524 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10528 = (inp[1]) ? 16'b0000001111111111 : node10529;
														assign node10529 = (inp[14]) ? 16'b0000001111111111 : node10530;
															assign node10530 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node10535 = (inp[3]) ? node10547 : node10536;
													assign node10536 = (inp[1]) ? node10544 : node10537;
														assign node10537 = (inp[12]) ? node10539 : 16'b0000011111111111;
															assign node10539 = (inp[7]) ? 16'b0000001111111111 : node10540;
																assign node10540 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10544 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10547 = (inp[14]) ? node10553 : node10548;
														assign node10548 = (inp[1]) ? 16'b0000000111111111 : node10549;
															assign node10549 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10553 = (inp[12]) ? node10555 : 16'b0000000111111111;
															assign node10555 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node10558 = (inp[12]) ? node10598 : node10559;
											assign node10559 = (inp[14]) ? node10573 : node10560;
												assign node10560 = (inp[3]) ? node10566 : node10561;
													assign node10561 = (inp[1]) ? 16'b0000011111111111 : node10562;
														assign node10562 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node10566 = (inp[1]) ? node10570 : node10567;
														assign node10567 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10570 = (inp[7]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node10573 = (inp[9]) ? node10587 : node10574;
													assign node10574 = (inp[7]) ? node10580 : node10575;
														assign node10575 = (inp[3]) ? 16'b0000001111111111 : node10576;
															assign node10576 = (inp[1]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node10580 = (inp[3]) ? 16'b0000000111111111 : node10581;
															assign node10581 = (inp[10]) ? node10583 : 16'b0000001111111111;
																assign node10583 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10587 = (inp[10]) ? node10595 : node10588;
														assign node10588 = (inp[3]) ? 16'b0000000111111111 : node10589;
															assign node10589 = (inp[1]) ? node10591 : 16'b0000001111111111;
																assign node10591 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10595 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10598 = (inp[1]) ? node10612 : node10599;
												assign node10599 = (inp[3]) ? node10605 : node10600;
													assign node10600 = (inp[7]) ? 16'b0000001111111111 : node10601;
														assign node10601 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node10605 = (inp[10]) ? node10609 : node10606;
														assign node10606 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10609 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10612 = (inp[10]) ? node10618 : node10613;
													assign node10613 = (inp[9]) ? node10615 : 16'b0000001111111111;
														assign node10615 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node10618 = (inp[3]) ? node10626 : node10619;
														assign node10619 = (inp[9]) ? 16'b0000000001111111 : node10620;
															assign node10620 = (inp[14]) ? node10622 : 16'b0000000111111111;
																assign node10622 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10626 = (inp[14]) ? node10628 : 16'b0000000011111111;
															assign node10628 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node10631 = (inp[9]) ? node10693 : node10632;
										assign node10632 = (inp[3]) ? node10668 : node10633;
											assign node10633 = (inp[14]) ? node10653 : node10634;
												assign node10634 = (inp[7]) ? node10646 : node10635;
													assign node10635 = (inp[1]) ? node10643 : node10636;
														assign node10636 = (inp[10]) ? 16'b0000011111111111 : node10637;
															assign node10637 = (inp[2]) ? 16'b0000111111111111 : node10638;
																assign node10638 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node10643 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10646 = (inp[12]) ? node10650 : node10647;
														assign node10647 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10650 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10653 = (inp[1]) ? node10663 : node10654;
													assign node10654 = (inp[7]) ? node10658 : node10655;
														assign node10655 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10658 = (inp[12]) ? node10660 : 16'b0000001111111111;
															assign node10660 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10663 = (inp[12]) ? node10665 : 16'b0000001111111111;
														assign node10665 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node10668 = (inp[7]) ? node10678 : node10669;
												assign node10669 = (inp[14]) ? node10673 : node10670;
													assign node10670 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10673 = (inp[1]) ? node10675 : 16'b0000000111111111;
														assign node10675 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10678 = (inp[12]) ? node10684 : node10679;
													assign node10679 = (inp[2]) ? node10681 : 16'b0000000111111111;
														assign node10681 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10684 = (inp[2]) ? node10688 : node10685;
														assign node10685 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10688 = (inp[1]) ? node10690 : 16'b0000000011111111;
															assign node10690 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10693 = (inp[10]) ? node10723 : node10694;
											assign node10694 = (inp[7]) ? node10710 : node10695;
												assign node10695 = (inp[1]) ? node10703 : node10696;
													assign node10696 = (inp[3]) ? node10698 : 16'b0000001111111111;
														assign node10698 = (inp[2]) ? node10700 : 16'b0000001111111111;
															assign node10700 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10703 = (inp[12]) ? 16'b0000000011111111 : node10704;
														assign node10704 = (inp[14]) ? node10706 : 16'b0000001111111111;
															assign node10706 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10710 = (inp[2]) ? node10714 : node10711;
													assign node10711 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10714 = (inp[3]) ? node10720 : node10715;
														assign node10715 = (inp[12]) ? node10717 : 16'b0000000111111111;
															assign node10717 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10720 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10723 = (inp[14]) ? node10739 : node10724;
												assign node10724 = (inp[3]) ? node10734 : node10725;
													assign node10725 = (inp[7]) ? node10729 : node10726;
														assign node10726 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10729 = (inp[12]) ? 16'b0000000011111111 : node10730;
															assign node10730 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10734 = (inp[1]) ? node10736 : 16'b0000000011111111;
														assign node10736 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node10739 = (inp[1]) ? node10747 : node10740;
													assign node10740 = (inp[12]) ? node10742 : 16'b0000000011111111;
														assign node10742 = (inp[7]) ? node10744 : 16'b0000000011111111;
															assign node10744 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10747 = (inp[7]) ? node10751 : node10748;
														assign node10748 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10751 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node10754 = (inp[14]) ? node10888 : node10755;
									assign node10755 = (inp[7]) ? node10837 : node10756;
										assign node10756 = (inp[12]) ? node10804 : node10757;
											assign node10757 = (inp[2]) ? node10779 : node10758;
												assign node10758 = (inp[1]) ? node10770 : node10759;
													assign node10759 = (inp[9]) ? node10767 : node10760;
														assign node10760 = (inp[3]) ? node10762 : 16'b0000111111111111;
															assign node10762 = (inp[13]) ? 16'b0000011111111111 : node10763;
																assign node10763 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node10767 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10770 = (inp[3]) ? node10776 : node10771;
														assign node10771 = (inp[13]) ? 16'b0000001111111111 : node10772;
															assign node10772 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10776 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node10779 = (inp[10]) ? node10791 : node10780;
													assign node10780 = (inp[3]) ? node10784 : node10781;
														assign node10781 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10784 = (inp[1]) ? node10786 : 16'b0000001111111111;
															assign node10786 = (inp[9]) ? 16'b0000000111111111 : node10787;
																assign node10787 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10791 = (inp[1]) ? node10799 : node10792;
														assign node10792 = (inp[3]) ? node10794 : 16'b0000001111111111;
															assign node10794 = (inp[9]) ? 16'b0000000111111111 : node10795;
																assign node10795 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10799 = (inp[3]) ? node10801 : 16'b0000000111111111;
															assign node10801 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10804 = (inp[13]) ? node10820 : node10805;
												assign node10805 = (inp[9]) ? node10811 : node10806;
													assign node10806 = (inp[10]) ? node10808 : 16'b0000011111111111;
														assign node10808 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10811 = (inp[1]) ? node10815 : node10812;
														assign node10812 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10815 = (inp[10]) ? node10817 : 16'b0000000111111111;
															assign node10817 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10820 = (inp[2]) ? node10832 : node10821;
													assign node10821 = (inp[1]) ? node10829 : node10822;
														assign node10822 = (inp[10]) ? 16'b0000000011111111 : node10823;
															assign node10823 = (inp[9]) ? node10825 : 16'b0000001111111111;
																assign node10825 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10829 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10832 = (inp[10]) ? 16'b0000000011111111 : node10833;
														assign node10833 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node10837 = (inp[3]) ? node10865 : node10838;
											assign node10838 = (inp[9]) ? node10856 : node10839;
												assign node10839 = (inp[2]) ? node10847 : node10840;
													assign node10840 = (inp[10]) ? node10842 : 16'b0000001111111111;
														assign node10842 = (inp[12]) ? 16'b0000000111111111 : node10843;
															assign node10843 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10847 = (inp[12]) ? node10851 : node10848;
														assign node10848 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10851 = (inp[13]) ? node10853 : 16'b0000000111111111;
															assign node10853 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10856 = (inp[1]) ? node10858 : 16'b0000000111111111;
													assign node10858 = (inp[2]) ? 16'b0000000011111111 : node10859;
														assign node10859 = (inp[12]) ? 16'b0000000011111111 : node10860;
															assign node10860 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10865 = (inp[12]) ? node10885 : node10866;
												assign node10866 = (inp[10]) ? node10878 : node10867;
													assign node10867 = (inp[9]) ? node10871 : node10868;
														assign node10868 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10871 = (inp[2]) ? 16'b0000000001111111 : node10872;
															assign node10872 = (inp[13]) ? node10874 : 16'b0000000111111111;
																assign node10874 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10878 = (inp[13]) ? 16'b0000000011111111 : node10879;
														assign node10879 = (inp[2]) ? 16'b0000000011111111 : node10880;
															assign node10880 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10885 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node10888 = (inp[12]) ? node10968 : node10889;
										assign node10889 = (inp[2]) ? node10925 : node10890;
											assign node10890 = (inp[1]) ? node10910 : node10891;
												assign node10891 = (inp[3]) ? node10903 : node10892;
													assign node10892 = (inp[10]) ? node10896 : node10893;
														assign node10893 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10896 = (inp[9]) ? 16'b0000000111111111 : node10897;
															assign node10897 = (inp[13]) ? node10899 : 16'b0000001111111111;
																assign node10899 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10903 = (inp[13]) ? node10907 : node10904;
														assign node10904 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10907 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10910 = (inp[3]) ? node10920 : node10911;
													assign node10911 = (inp[10]) ? node10915 : node10912;
														assign node10912 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10915 = (inp[9]) ? node10917 : 16'b0000000111111111;
															assign node10917 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10920 = (inp[7]) ? 16'b0000000001111111 : node10921;
														assign node10921 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10925 = (inp[13]) ? node10953 : node10926;
												assign node10926 = (inp[1]) ? node10938 : node10927;
													assign node10927 = (inp[7]) ? node10935 : node10928;
														assign node10928 = (inp[9]) ? node10930 : 16'b0000001111111111;
															assign node10930 = (inp[10]) ? 16'b0000000111111111 : node10931;
																assign node10931 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10935 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node10938 = (inp[3]) ? node10948 : node10939;
														assign node10939 = (inp[7]) ? node10941 : 16'b0000000111111111;
															assign node10941 = (inp[10]) ? node10945 : node10942;
																assign node10942 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node10945 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10948 = (inp[9]) ? node10950 : 16'b0000000011111111;
															assign node10950 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10953 = (inp[10]) ? node10963 : node10954;
													assign node10954 = (inp[1]) ? node10958 : node10955;
														assign node10955 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10958 = (inp[3]) ? node10960 : 16'b0000000011111111;
															assign node10960 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10963 = (inp[1]) ? 16'b0000000001111111 : node10964;
														assign node10964 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10968 = (inp[3]) ? node11002 : node10969;
											assign node10969 = (inp[1]) ? node10987 : node10970;
												assign node10970 = (inp[7]) ? node10980 : node10971;
													assign node10971 = (inp[13]) ? node10977 : node10972;
														assign node10972 = (inp[2]) ? node10974 : 16'b0000001111111111;
															assign node10974 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10977 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10980 = (inp[10]) ? node10984 : node10981;
														assign node10981 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10984 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10987 = (inp[13]) ? node10997 : node10988;
													assign node10988 = (inp[2]) ? node10992 : node10989;
														assign node10989 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10992 = (inp[7]) ? node10994 : 16'b0000000011111111;
															assign node10994 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10997 = (inp[9]) ? 16'b0000000001111111 : node10998;
														assign node10998 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11002 = (inp[13]) ? node11020 : node11003;
												assign node11003 = (inp[10]) ? node11011 : node11004;
													assign node11004 = (inp[1]) ? node11006 : 16'b0000000111111111;
														assign node11006 = (inp[7]) ? node11008 : 16'b0000000011111111;
															assign node11008 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node11011 = (inp[1]) ? node11017 : node11012;
														assign node11012 = (inp[9]) ? node11014 : 16'b0000000001111111;
															assign node11014 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11017 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11020 = (inp[1]) ? node11026 : node11021;
													assign node11021 = (inp[9]) ? node11023 : 16'b0000000011111111;
														assign node11023 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11026 = (inp[10]) ? node11034 : node11027;
														assign node11027 = (inp[9]) ? 16'b0000000000011111 : node11028;
															assign node11028 = (inp[7]) ? node11030 : 16'b0000000001111111;
																assign node11030 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11034 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node11037 = (inp[2]) ? node11283 : node11038;
								assign node11038 = (inp[3]) ? node11154 : node11039;
									assign node11039 = (inp[12]) ? node11099 : node11040;
										assign node11040 = (inp[10]) ? node11074 : node11041;
											assign node11041 = (inp[6]) ? node11059 : node11042;
												assign node11042 = (inp[1]) ? node11054 : node11043;
													assign node11043 = (inp[7]) ? node11051 : node11044;
														assign node11044 = (inp[14]) ? 16'b0000011111111111 : node11045;
															assign node11045 = (inp[13]) ? 16'b0000111111111111 : node11046;
																assign node11046 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node11051 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11054 = (inp[9]) ? 16'b0000000111111111 : node11055;
														assign node11055 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node11059 = (inp[7]) ? node11069 : node11060;
													assign node11060 = (inp[1]) ? node11064 : node11061;
														assign node11061 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11064 = (inp[14]) ? node11066 : 16'b0000001111111111;
															assign node11066 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11069 = (inp[14]) ? 16'b0000000011111111 : node11070;
														assign node11070 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node11074 = (inp[9]) ? node11088 : node11075;
												assign node11075 = (inp[6]) ? node11083 : node11076;
													assign node11076 = (inp[13]) ? node11080 : node11077;
														assign node11077 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node11080 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11083 = (inp[13]) ? 16'b0000000111111111 : node11084;
														assign node11084 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11088 = (inp[14]) ? node11090 : 16'b0000000111111111;
													assign node11090 = (inp[13]) ? node11094 : node11091;
														assign node11091 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11094 = (inp[7]) ? node11096 : 16'b0000000011111111;
															assign node11096 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11099 = (inp[6]) ? node11119 : node11100;
											assign node11100 = (inp[10]) ? node11104 : node11101;
												assign node11101 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node11104 = (inp[7]) ? node11114 : node11105;
													assign node11105 = (inp[1]) ? node11109 : node11106;
														assign node11106 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11109 = (inp[14]) ? 16'b0000000011111111 : node11110;
															assign node11110 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11114 = (inp[9]) ? 16'b0000000011111111 : node11115;
														assign node11115 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11119 = (inp[9]) ? node11141 : node11120;
												assign node11120 = (inp[13]) ? node11130 : node11121;
													assign node11121 = (inp[1]) ? 16'b0000000011111111 : node11122;
														assign node11122 = (inp[14]) ? node11124 : 16'b0000001111111111;
															assign node11124 = (inp[10]) ? 16'b0000000111111111 : node11125;
																assign node11125 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11130 = (inp[14]) ? node11134 : node11131;
														assign node11131 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11134 = (inp[10]) ? 16'b0000000001111111 : node11135;
															assign node11135 = (inp[1]) ? node11137 : 16'b0000000011111111;
																assign node11137 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11141 = (inp[7]) ? node11147 : node11142;
													assign node11142 = (inp[10]) ? node11144 : 16'b0000000011111111;
														assign node11144 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11147 = (inp[13]) ? node11149 : 16'b0000000011111111;
														assign node11149 = (inp[1]) ? node11151 : 16'b0000000001111111;
															assign node11151 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node11154 = (inp[13]) ? node11222 : node11155;
										assign node11155 = (inp[9]) ? node11183 : node11156;
											assign node11156 = (inp[14]) ? node11176 : node11157;
												assign node11157 = (inp[7]) ? node11167 : node11158;
													assign node11158 = (inp[1]) ? node11160 : 16'b0000011111111111;
														assign node11160 = (inp[6]) ? node11164 : node11161;
															assign node11161 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node11164 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11167 = (inp[12]) ? node11169 : 16'b0000001111111111;
														assign node11169 = (inp[10]) ? node11171 : 16'b0000000111111111;
															assign node11171 = (inp[1]) ? 16'b0000000011111111 : node11172;
																assign node11172 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11176 = (inp[10]) ? 16'b0000000011111111 : node11177;
													assign node11177 = (inp[1]) ? node11179 : 16'b0000000111111111;
														assign node11179 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11183 = (inp[6]) ? node11207 : node11184;
												assign node11184 = (inp[1]) ? node11192 : node11185;
													assign node11185 = (inp[10]) ? node11189 : node11186;
														assign node11186 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11189 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node11192 = (inp[7]) ? node11200 : node11193;
														assign node11193 = (inp[12]) ? 16'b0000000011111111 : node11194;
															assign node11194 = (inp[14]) ? node11196 : 16'b0000000111111111;
																assign node11196 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11200 = (inp[10]) ? 16'b0000000001111111 : node11201;
															assign node11201 = (inp[12]) ? node11203 : 16'b0000000011111111;
																assign node11203 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11207 = (inp[1]) ? node11215 : node11208;
													assign node11208 = (inp[12]) ? node11212 : node11209;
														assign node11209 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11212 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11215 = (inp[7]) ? node11219 : node11216;
														assign node11216 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11219 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11222 = (inp[6]) ? node11252 : node11223;
											assign node11223 = (inp[10]) ? node11235 : node11224;
												assign node11224 = (inp[14]) ? 16'b0000000011111111 : node11225;
													assign node11225 = (inp[1]) ? node11227 : 16'b0000001111111111;
														assign node11227 = (inp[12]) ? node11229 : 16'b0000000111111111;
															assign node11229 = (inp[7]) ? 16'b0000000011111111 : node11230;
																assign node11230 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11235 = (inp[9]) ? node11245 : node11236;
													assign node11236 = (inp[1]) ? node11240 : node11237;
														assign node11237 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11240 = (inp[14]) ? node11242 : 16'b0000000011111111;
															assign node11242 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11245 = (inp[1]) ? node11249 : node11246;
														assign node11246 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11249 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11252 = (inp[12]) ? node11270 : node11253;
												assign node11253 = (inp[1]) ? node11263 : node11254;
													assign node11254 = (inp[10]) ? node11256 : 16'b0000000111111111;
														assign node11256 = (inp[14]) ? node11258 : 16'b0000000011111111;
															assign node11258 = (inp[9]) ? 16'b0000000001111111 : node11259;
																assign node11259 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11263 = (inp[10]) ? node11267 : node11264;
														assign node11264 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11267 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11270 = (inp[1]) ? 16'b0000000000111111 : node11271;
													assign node11271 = (inp[14]) ? node11275 : node11272;
														assign node11272 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11275 = (inp[9]) ? node11277 : 16'b0000000001111111;
															assign node11277 = (inp[10]) ? 16'b0000000000111111 : node11278;
																assign node11278 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node11283 = (inp[9]) ? node11413 : node11284;
									assign node11284 = (inp[12]) ? node11344 : node11285;
										assign node11285 = (inp[7]) ? node11313 : node11286;
											assign node11286 = (inp[3]) ? node11298 : node11287;
												assign node11287 = (inp[14]) ? node11293 : node11288;
													assign node11288 = (inp[6]) ? node11290 : 16'b0000001111111111;
														assign node11290 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11293 = (inp[1]) ? node11295 : 16'b0000000111111111;
														assign node11295 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11298 = (inp[6]) ? node11304 : node11299;
													assign node11299 = (inp[10]) ? 16'b0000000111111111 : node11300;
														assign node11300 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11304 = (inp[10]) ? node11308 : node11305;
														assign node11305 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11308 = (inp[1]) ? node11310 : 16'b0000000011111111;
															assign node11310 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11313 = (inp[13]) ? node11329 : node11314;
												assign node11314 = (inp[14]) ? node11320 : node11315;
													assign node11315 = (inp[1]) ? node11317 : 16'b0000000111111111;
														assign node11317 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11320 = (inp[3]) ? node11324 : node11321;
														assign node11321 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11324 = (inp[10]) ? node11326 : 16'b0000000011111111;
															assign node11326 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11329 = (inp[6]) ? node11337 : node11330;
													assign node11330 = (inp[3]) ? node11334 : node11331;
														assign node11331 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11334 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11337 = (inp[10]) ? 16'b0000000011111111 : node11338;
														assign node11338 = (inp[1]) ? node11340 : 16'b0000000001111111;
															assign node11340 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11344 = (inp[14]) ? node11376 : node11345;
											assign node11345 = (inp[3]) ? node11365 : node11346;
												assign node11346 = (inp[6]) ? node11356 : node11347;
													assign node11347 = (inp[7]) ? node11353 : node11348;
														assign node11348 = (inp[1]) ? 16'b0000000111111111 : node11349;
															assign node11349 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11353 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11356 = (inp[1]) ? node11360 : node11357;
														assign node11357 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11360 = (inp[7]) ? node11362 : 16'b0000000011111111;
															assign node11362 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11365 = (inp[6]) ? 16'b0000000001111111 : node11366;
													assign node11366 = (inp[10]) ? node11370 : node11367;
														assign node11367 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11370 = (inp[7]) ? 16'b0000000001111111 : node11371;
															assign node11371 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11376 = (inp[7]) ? node11396 : node11377;
												assign node11377 = (inp[1]) ? node11383 : node11378;
													assign node11378 = (inp[3]) ? node11380 : 16'b0000000011111111;
														assign node11380 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11383 = (inp[13]) ? node11389 : node11384;
														assign node11384 = (inp[6]) ? 16'b0000000001111111 : node11385;
															assign node11385 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11389 = (inp[6]) ? 16'b0000000000111111 : node11390;
															assign node11390 = (inp[3]) ? node11392 : 16'b0000000001111111;
																assign node11392 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11396 = (inp[6]) ? node11406 : node11397;
													assign node11397 = (inp[10]) ? node11401 : node11398;
														assign node11398 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11401 = (inp[1]) ? node11403 : 16'b0000000001111111;
															assign node11403 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11406 = (inp[1]) ? node11410 : node11407;
														assign node11407 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11410 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node11413 = (inp[12]) ? node11469 : node11414;
										assign node11414 = (inp[13]) ? node11436 : node11415;
											assign node11415 = (inp[1]) ? node11429 : node11416;
												assign node11416 = (inp[14]) ? node11426 : node11417;
													assign node11417 = (inp[7]) ? node11419 : 16'b0000000111111111;
														assign node11419 = (inp[3]) ? node11421 : 16'b0000000111111111;
															assign node11421 = (inp[6]) ? 16'b0000000011111111 : node11422;
																assign node11422 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11426 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11429 = (inp[10]) ? 16'b0000000001111111 : node11430;
													assign node11430 = (inp[3]) ? 16'b0000000001111111 : node11431;
														assign node11431 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11436 = (inp[7]) ? node11460 : node11437;
												assign node11437 = (inp[3]) ? node11447 : node11438;
													assign node11438 = (inp[6]) ? node11440 : 16'b0000000011111111;
														assign node11440 = (inp[1]) ? node11444 : node11441;
															assign node11441 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node11444 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11447 = (inp[10]) ? node11453 : node11448;
														assign node11448 = (inp[6]) ? 16'b0000000001111111 : node11449;
															assign node11449 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11453 = (inp[6]) ? 16'b0000000000111111 : node11454;
															assign node11454 = (inp[1]) ? node11456 : 16'b0000000001111111;
																assign node11456 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11460 = (inp[1]) ? node11464 : node11461;
													assign node11461 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11464 = (inp[10]) ? node11466 : 16'b0000000000111111;
														assign node11466 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11469 = (inp[1]) ? node11499 : node11470;
											assign node11470 = (inp[14]) ? node11484 : node11471;
												assign node11471 = (inp[7]) ? node11475 : node11472;
													assign node11472 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node11475 = (inp[3]) ? node11479 : node11476;
														assign node11476 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11479 = (inp[10]) ? node11481 : 16'b0000000001111111;
															assign node11481 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11484 = (inp[7]) ? node11492 : node11485;
													assign node11485 = (inp[13]) ? node11489 : node11486;
														assign node11486 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11489 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11492 = (inp[3]) ? 16'b0000000000111111 : node11493;
														assign node11493 = (inp[13]) ? 16'b0000000000111111 : node11494;
															assign node11494 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11499 = (inp[14]) ? node11513 : node11500;
												assign node11500 = (inp[7]) ? node11506 : node11501;
													assign node11501 = (inp[3]) ? node11503 : 16'b0000000001111111;
														assign node11503 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11506 = (inp[10]) ? node11510 : node11507;
														assign node11507 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11510 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11513 = (inp[3]) ? node11519 : node11514;
													assign node11514 = (inp[10]) ? node11516 : 16'b0000000001111111;
														assign node11516 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11519 = (inp[13]) ? node11523 : node11520;
														assign node11520 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11523 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node11526 = (inp[13]) ? node12016 : node11527;
							assign node11527 = (inp[14]) ? node11781 : node11528;
								assign node11528 = (inp[3]) ? node11636 : node11529;
									assign node11529 = (inp[10]) ? node11577 : node11530;
										assign node11530 = (inp[12]) ? node11550 : node11531;
											assign node11531 = (inp[7]) ? node11543 : node11532;
												assign node11532 = (inp[9]) ? node11538 : node11533;
													assign node11533 = (inp[2]) ? 16'b0000011111111111 : node11534;
														assign node11534 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node11538 = (inp[15]) ? 16'b0000001111111111 : node11539;
														assign node11539 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node11543 = (inp[2]) ? node11547 : node11544;
													assign node11544 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11547 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node11550 = (inp[15]) ? node11560 : node11551;
												assign node11551 = (inp[9]) ? node11555 : node11552;
													assign node11552 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11555 = (inp[1]) ? 16'b0000000111111111 : node11556;
														assign node11556 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11560 = (inp[9]) ? node11570 : node11561;
													assign node11561 = (inp[6]) ? node11567 : node11562;
														assign node11562 = (inp[1]) ? node11564 : 16'b0000001111111111;
															assign node11564 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11567 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11570 = (inp[6]) ? 16'b0000000000111111 : node11571;
														assign node11571 = (inp[2]) ? node11573 : 16'b0000000011111111;
															assign node11573 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node11577 = (inp[9]) ? node11617 : node11578;
											assign node11578 = (inp[2]) ? node11590 : node11579;
												assign node11579 = (inp[12]) ? node11585 : node11580;
													assign node11580 = (inp[6]) ? node11582 : 16'b0000001111111111;
														assign node11582 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11585 = (inp[6]) ? 16'b0000000011111111 : node11586;
														assign node11586 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11590 = (inp[6]) ? node11606 : node11591;
													assign node11591 = (inp[7]) ? node11601 : node11592;
														assign node11592 = (inp[12]) ? node11598 : node11593;
															assign node11593 = (inp[15]) ? node11595 : 16'b0000001111111111;
																assign node11595 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node11598 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11601 = (inp[15]) ? node11603 : 16'b0000000111111111;
															assign node11603 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11606 = (inp[1]) ? node11614 : node11607;
														assign node11607 = (inp[7]) ? node11609 : 16'b0000000111111111;
															assign node11609 = (inp[15]) ? 16'b0000000011111111 : node11610;
																assign node11610 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11614 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11617 = (inp[15]) ? node11623 : node11618;
												assign node11618 = (inp[12]) ? node11620 : 16'b0000001111111111;
													assign node11620 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11623 = (inp[6]) ? node11631 : node11624;
													assign node11624 = (inp[7]) ? node11628 : node11625;
														assign node11625 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11628 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11631 = (inp[12]) ? node11633 : 16'b0000000001111111;
														assign node11633 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node11636 = (inp[6]) ? node11722 : node11637;
										assign node11637 = (inp[15]) ? node11679 : node11638;
											assign node11638 = (inp[10]) ? node11654 : node11639;
												assign node11639 = (inp[9]) ? node11649 : node11640;
													assign node11640 = (inp[1]) ? 16'b0000001111111111 : node11641;
														assign node11641 = (inp[12]) ? 16'b0000001111111111 : node11642;
															assign node11642 = (inp[2]) ? 16'b0000011111111111 : node11643;
																assign node11643 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node11649 = (inp[7]) ? node11651 : 16'b0000000111111111;
														assign node11651 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11654 = (inp[7]) ? node11668 : node11655;
													assign node11655 = (inp[1]) ? node11661 : node11656;
														assign node11656 = (inp[2]) ? 16'b0000000111111111 : node11657;
															assign node11657 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11661 = (inp[12]) ? node11663 : 16'b0000000111111111;
															assign node11663 = (inp[2]) ? 16'b0000000011111111 : node11664;
																assign node11664 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11668 = (inp[1]) ? node11676 : node11669;
														assign node11669 = (inp[2]) ? 16'b0000000011111111 : node11670;
															assign node11670 = (inp[9]) ? node11672 : 16'b0000000111111111;
																assign node11672 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11676 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node11679 = (inp[1]) ? node11703 : node11680;
												assign node11680 = (inp[10]) ? node11692 : node11681;
													assign node11681 = (inp[7]) ? node11685 : node11682;
														assign node11682 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11685 = (inp[9]) ? node11687 : 16'b0000000111111111;
															assign node11687 = (inp[12]) ? 16'b0000000011111111 : node11688;
																assign node11688 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11692 = (inp[2]) ? node11698 : node11693;
														assign node11693 = (inp[9]) ? 16'b0000000011111111 : node11694;
															assign node11694 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11698 = (inp[9]) ? node11700 : 16'b0000000011111111;
															assign node11700 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11703 = (inp[9]) ? node11713 : node11704;
													assign node11704 = (inp[10]) ? 16'b0000000001111111 : node11705;
														assign node11705 = (inp[7]) ? 16'b0000000011111111 : node11706;
															assign node11706 = (inp[12]) ? node11708 : 16'b0000000111111111;
																assign node11708 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11713 = (inp[12]) ? node11719 : node11714;
														assign node11714 = (inp[7]) ? 16'b0000000001111111 : node11715;
															assign node11715 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11719 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11722 = (inp[15]) ? node11756 : node11723;
											assign node11723 = (inp[9]) ? node11733 : node11724;
												assign node11724 = (inp[12]) ? node11726 : 16'b0000000111111111;
													assign node11726 = (inp[2]) ? node11730 : node11727;
														assign node11727 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11730 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11733 = (inp[1]) ? node11745 : node11734;
													assign node11734 = (inp[7]) ? node11740 : node11735;
														assign node11735 = (inp[2]) ? 16'b0000000011111111 : node11736;
															assign node11736 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11740 = (inp[2]) ? node11742 : 16'b0000000011111111;
															assign node11742 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node11745 = (inp[12]) ? node11753 : node11746;
														assign node11746 = (inp[2]) ? node11748 : 16'b0000000011111111;
															assign node11748 = (inp[10]) ? 16'b0000000001111111 : node11749;
																assign node11749 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11753 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11756 = (inp[1]) ? node11770 : node11757;
												assign node11757 = (inp[12]) ? node11767 : node11758;
													assign node11758 = (inp[2]) ? node11764 : node11759;
														assign node11759 = (inp[10]) ? node11761 : 16'b0000000111111111;
															assign node11761 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11764 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11767 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node11770 = (inp[9]) ? node11776 : node11771;
													assign node11771 = (inp[12]) ? node11773 : 16'b0000000001111111;
														assign node11773 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11776 = (inp[7]) ? node11778 : 16'b0000000000111111;
														assign node11778 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node11781 = (inp[3]) ? node11893 : node11782;
									assign node11782 = (inp[10]) ? node11828 : node11783;
										assign node11783 = (inp[9]) ? node11799 : node11784;
											assign node11784 = (inp[7]) ? node11788 : node11785;
												assign node11785 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11788 = (inp[15]) ? node11794 : node11789;
													assign node11789 = (inp[6]) ? node11791 : 16'b0000000111111111;
														assign node11791 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11794 = (inp[2]) ? 16'b0000000011111111 : node11795;
														assign node11795 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11799 = (inp[12]) ? node11819 : node11800;
												assign node11800 = (inp[15]) ? node11810 : node11801;
													assign node11801 = (inp[7]) ? 16'b0000000011111111 : node11802;
														assign node11802 = (inp[2]) ? node11806 : node11803;
															assign node11803 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node11806 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11810 = (inp[7]) ? node11816 : node11811;
														assign node11811 = (inp[6]) ? 16'b0000000011111111 : node11812;
															assign node11812 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11816 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11819 = (inp[1]) ? node11823 : node11820;
													assign node11820 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11823 = (inp[6]) ? node11825 : 16'b0000000001111111;
														assign node11825 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node11828 = (inp[12]) ? node11874 : node11829;
											assign node11829 = (inp[1]) ? node11845 : node11830;
												assign node11830 = (inp[15]) ? node11836 : node11831;
													assign node11831 = (inp[6]) ? node11833 : 16'b0000000111111111;
														assign node11833 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11836 = (inp[2]) ? node11842 : node11837;
														assign node11837 = (inp[7]) ? 16'b0000000011111111 : node11838;
															assign node11838 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11842 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11845 = (inp[7]) ? node11859 : node11846;
													assign node11846 = (inp[6]) ? node11854 : node11847;
														assign node11847 = (inp[15]) ? node11849 : 16'b0000000111111111;
															assign node11849 = (inp[9]) ? node11851 : 16'b0000000111111111;
																assign node11851 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11854 = (inp[2]) ? node11856 : 16'b0000000011111111;
															assign node11856 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11859 = (inp[2]) ? node11871 : node11860;
														assign node11860 = (inp[6]) ? node11866 : node11861;
															assign node11861 = (inp[9]) ? node11863 : 16'b0000000011111111;
																assign node11863 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node11866 = (inp[9]) ? 16'b0000000001111111 : node11867;
																assign node11867 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11871 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node11874 = (inp[2]) ? node11884 : node11875;
												assign node11875 = (inp[7]) ? node11877 : 16'b0000000011111111;
													assign node11877 = (inp[9]) ? node11881 : node11878;
														assign node11878 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11881 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11884 = (inp[7]) ? node11890 : node11885;
													assign node11885 = (inp[15]) ? 16'b0000000000111111 : node11886;
														assign node11886 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11890 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node11893 = (inp[7]) ? node11955 : node11894;
										assign node11894 = (inp[12]) ? node11922 : node11895;
											assign node11895 = (inp[9]) ? node11905 : node11896;
												assign node11896 = (inp[15]) ? node11898 : 16'b0000000111111111;
													assign node11898 = (inp[1]) ? 16'b0000000001111111 : node11899;
														assign node11899 = (inp[2]) ? 16'b0000000011111111 : node11900;
															assign node11900 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11905 = (inp[10]) ? node11917 : node11906;
													assign node11906 = (inp[6]) ? node11912 : node11907;
														assign node11907 = (inp[2]) ? node11909 : 16'b0000000111111111;
															assign node11909 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11912 = (inp[15]) ? node11914 : 16'b0000000011111111;
															assign node11914 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11917 = (inp[15]) ? 16'b0000000000111111 : node11918;
														assign node11918 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11922 = (inp[1]) ? node11940 : node11923;
												assign node11923 = (inp[2]) ? node11929 : node11924;
													assign node11924 = (inp[6]) ? 16'b0000000001111111 : node11925;
														assign node11925 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11929 = (inp[9]) ? node11937 : node11930;
														assign node11930 = (inp[6]) ? node11932 : 16'b0000000011111111;
															assign node11932 = (inp[10]) ? 16'b0000000001111111 : node11933;
																assign node11933 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11937 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11940 = (inp[2]) ? node11948 : node11941;
													assign node11941 = (inp[9]) ? node11945 : node11942;
														assign node11942 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11945 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11948 = (inp[15]) ? node11952 : node11949;
														assign node11949 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11952 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11955 = (inp[6]) ? node11979 : node11956;
											assign node11956 = (inp[2]) ? node11962 : node11957;
												assign node11957 = (inp[10]) ? node11959 : 16'b0000000011111111;
													assign node11959 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11962 = (inp[12]) ? node11970 : node11963;
													assign node11963 = (inp[10]) ? node11965 : 16'b0000000011111111;
														assign node11965 = (inp[1]) ? node11967 : 16'b0000000001111111;
															assign node11967 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11970 = (inp[15]) ? node11974 : node11971;
														assign node11971 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11974 = (inp[9]) ? node11976 : 16'b0000000000011111;
															assign node11976 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11979 = (inp[2]) ? node11995 : node11980;
												assign node11980 = (inp[10]) ? node11982 : 16'b0000000001111111;
													assign node11982 = (inp[9]) ? node11988 : node11983;
														assign node11983 = (inp[12]) ? node11985 : 16'b0000000001111111;
															assign node11985 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11988 = (inp[1]) ? 16'b0000000000011111 : node11989;
															assign node11989 = (inp[12]) ? node11991 : 16'b0000000000111111;
																assign node11991 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11995 = (inp[10]) ? node12005 : node11996;
													assign node11996 = (inp[15]) ? node11998 : 16'b0000000000111111;
														assign node11998 = (inp[1]) ? node12000 : 16'b0000000000111111;
															assign node12000 = (inp[9]) ? 16'b0000000000011111 : node12001;
																assign node12001 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node12005 = (inp[9]) ? node12013 : node12006;
														assign node12006 = (inp[12]) ? node12008 : 16'b0000000000111111;
															assign node12008 = (inp[1]) ? 16'b0000000000011111 : node12009;
																assign node12009 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node12013 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node12016 = (inp[15]) ? node12248 : node12017;
								assign node12017 = (inp[10]) ? node12131 : node12018;
									assign node12018 = (inp[7]) ? node12064 : node12019;
										assign node12019 = (inp[3]) ? node12047 : node12020;
											assign node12020 = (inp[9]) ? node12038 : node12021;
												assign node12021 = (inp[12]) ? node12029 : node12022;
													assign node12022 = (inp[2]) ? 16'b0000001111111111 : node12023;
														assign node12023 = (inp[1]) ? 16'b0000001111111111 : node12024;
															assign node12024 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12029 = (inp[6]) ? node12035 : node12030;
														assign node12030 = (inp[14]) ? 16'b0000000111111111 : node12031;
															assign node12031 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12035 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12038 = (inp[14]) ? node12042 : node12039;
													assign node12039 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node12042 = (inp[12]) ? node12044 : 16'b0000000011111111;
														assign node12044 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node12047 = (inp[6]) ? node12055 : node12048;
												assign node12048 = (inp[9]) ? 16'b0000000011111111 : node12049;
													assign node12049 = (inp[2]) ? node12051 : 16'b0000000111111111;
														assign node12051 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12055 = (inp[2]) ? node12061 : node12056;
													assign node12056 = (inp[12]) ? 16'b0000000011111111 : node12057;
														assign node12057 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12061 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node12064 = (inp[6]) ? node12092 : node12065;
											assign node12065 = (inp[2]) ? node12077 : node12066;
												assign node12066 = (inp[1]) ? node12068 : 16'b0000000111111111;
													assign node12068 = (inp[12]) ? node12074 : node12069;
														assign node12069 = (inp[9]) ? node12071 : 16'b0000000111111111;
															assign node12071 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12074 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12077 = (inp[14]) ? node12085 : node12078;
													assign node12078 = (inp[12]) ? node12080 : 16'b0000000011111111;
														assign node12080 = (inp[3]) ? 16'b0000000011111111 : node12081;
															assign node12081 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12085 = (inp[1]) ? node12089 : node12086;
														assign node12086 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12089 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12092 = (inp[3]) ? node12116 : node12093;
												assign node12093 = (inp[9]) ? node12107 : node12094;
													assign node12094 = (inp[12]) ? node12100 : node12095;
														assign node12095 = (inp[14]) ? node12097 : 16'b0000000111111111;
															assign node12097 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12100 = (inp[2]) ? node12102 : 16'b0000000011111111;
															assign node12102 = (inp[1]) ? 16'b0000000001111111 : node12103;
																assign node12103 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12107 = (inp[12]) ? node12111 : node12108;
														assign node12108 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12111 = (inp[1]) ? 16'b0000000000111111 : node12112;
															assign node12112 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12116 = (inp[14]) ? node12126 : node12117;
													assign node12117 = (inp[1]) ? node12119 : 16'b0000000001111111;
														assign node12119 = (inp[12]) ? 16'b0000000000111111 : node12120;
															assign node12120 = (inp[9]) ? node12122 : 16'b0000000001111111;
																assign node12122 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12126 = (inp[12]) ? 16'b0000000000011111 : node12127;
														assign node12127 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12131 = (inp[14]) ? node12181 : node12132;
										assign node12132 = (inp[1]) ? node12152 : node12133;
											assign node12133 = (inp[6]) ? node12141 : node12134;
												assign node12134 = (inp[12]) ? node12136 : 16'b0000000111111111;
													assign node12136 = (inp[9]) ? node12138 : 16'b0000000011111111;
														assign node12138 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12141 = (inp[7]) ? node12147 : node12142;
													assign node12142 = (inp[9]) ? node12144 : 16'b0000000111111111;
														assign node12144 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12147 = (inp[9]) ? node12149 : 16'b0000000001111111;
														assign node12149 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node12152 = (inp[3]) ? node12168 : node12153;
												assign node12153 = (inp[9]) ? node12161 : node12154;
													assign node12154 = (inp[2]) ? node12158 : node12155;
														assign node12155 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node12158 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12161 = (inp[7]) ? node12165 : node12162;
														assign node12162 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12165 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12168 = (inp[7]) ? node12176 : node12169;
													assign node12169 = (inp[2]) ? node12171 : 16'b0000000001111111;
														assign node12171 = (inp[12]) ? 16'b0000000000111111 : node12172;
															assign node12172 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12176 = (inp[12]) ? node12178 : 16'b0000000000111111;
														assign node12178 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node12181 = (inp[2]) ? node12221 : node12182;
											assign node12182 = (inp[6]) ? node12196 : node12183;
												assign node12183 = (inp[3]) ? node12189 : node12184;
													assign node12184 = (inp[9]) ? node12186 : 16'b0000000011111111;
														assign node12186 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12189 = (inp[1]) ? node12191 : 16'b0000000001111111;
														assign node12191 = (inp[9]) ? node12193 : 16'b0000000001111111;
															assign node12193 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12196 = (inp[1]) ? node12212 : node12197;
													assign node12197 = (inp[12]) ? node12205 : node12198;
														assign node12198 = (inp[9]) ? node12200 : 16'b0000000011111111;
															assign node12200 = (inp[7]) ? 16'b0000000001111111 : node12201;
																assign node12201 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12205 = (inp[7]) ? node12207 : 16'b0000000001111111;
															assign node12207 = (inp[3]) ? 16'b0000000000111111 : node12208;
																assign node12208 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12212 = (inp[9]) ? 16'b0000000000111111 : node12213;
														assign node12213 = (inp[7]) ? 16'b0000000000111111 : node12214;
															assign node12214 = (inp[3]) ? node12216 : 16'b0000000001111111;
																assign node12216 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12221 = (inp[6]) ? node12235 : node12222;
												assign node12222 = (inp[7]) ? node12228 : node12223;
													assign node12223 = (inp[12]) ? node12225 : 16'b0000000001111111;
														assign node12225 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12228 = (inp[12]) ? node12230 : 16'b0000000000111111;
														assign node12230 = (inp[3]) ? 16'b0000000000111111 : node12231;
															assign node12231 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12235 = (inp[9]) ? node12239 : node12236;
													assign node12236 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12239 = (inp[7]) ? node12241 : 16'b0000000000111111;
														assign node12241 = (inp[3]) ? node12243 : 16'b0000000000011111;
															assign node12243 = (inp[12]) ? node12245 : 16'b0000000000001111;
																assign node12245 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node12248 = (inp[12]) ? node12362 : node12249;
									assign node12249 = (inp[2]) ? node12291 : node12250;
										assign node12250 = (inp[10]) ? node12268 : node12251;
											assign node12251 = (inp[7]) ? node12263 : node12252;
												assign node12252 = (inp[14]) ? node12258 : node12253;
													assign node12253 = (inp[1]) ? 16'b0000000111111111 : node12254;
														assign node12254 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12258 = (inp[1]) ? 16'b0000000001111111 : node12259;
														assign node12259 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12263 = (inp[14]) ? node12265 : 16'b0000000011111111;
													assign node12265 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12268 = (inp[3]) ? node12280 : node12269;
												assign node12269 = (inp[6]) ? node12275 : node12270;
													assign node12270 = (inp[14]) ? 16'b0000000011111111 : node12271;
														assign node12271 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12275 = (inp[14]) ? 16'b0000000000111111 : node12276;
														assign node12276 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12280 = (inp[9]) ? node12286 : node12281;
													assign node12281 = (inp[7]) ? node12283 : 16'b0000000111111111;
														assign node12283 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12286 = (inp[6]) ? 16'b0000000000111111 : node12287;
														assign node12287 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node12291 = (inp[9]) ? node12325 : node12292;
											assign node12292 = (inp[6]) ? node12312 : node12293;
												assign node12293 = (inp[14]) ? node12305 : node12294;
													assign node12294 = (inp[3]) ? node12302 : node12295;
														assign node12295 = (inp[7]) ? 16'b0000000001111111 : node12296;
															assign node12296 = (inp[10]) ? 16'b0000000111111111 : node12297;
																assign node12297 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12302 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12305 = (inp[1]) ? node12307 : 16'b0000000001111111;
														assign node12307 = (inp[3]) ? node12309 : 16'b0000000001111111;
															assign node12309 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12312 = (inp[7]) ? node12320 : node12313;
													assign node12313 = (inp[3]) ? node12317 : node12314;
														assign node12314 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12317 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12320 = (inp[3]) ? node12322 : 16'b0000000000111111;
														assign node12322 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node12325 = (inp[7]) ? node12347 : node12326;
												assign node12326 = (inp[6]) ? node12338 : node12327;
													assign node12327 = (inp[10]) ? 16'b0000000000111111 : node12328;
														assign node12328 = (inp[1]) ? node12332 : node12329;
															assign node12329 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node12332 = (inp[3]) ? node12334 : 16'b0000000001111111;
																assign node12334 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12338 = (inp[1]) ? node12342 : node12339;
														assign node12339 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12342 = (inp[14]) ? node12344 : 16'b0000000000111111;
															assign node12344 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node12347 = (inp[1]) ? node12357 : node12348;
													assign node12348 = (inp[6]) ? node12352 : node12349;
														assign node12349 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12352 = (inp[10]) ? node12354 : 16'b0000000000111111;
															assign node12354 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node12357 = (inp[10]) ? 16'b0000000000011111 : node12358;
														assign node12358 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node12362 = (inp[3]) ? node12418 : node12363;
										assign node12363 = (inp[14]) ? node12389 : node12364;
											assign node12364 = (inp[1]) ? node12376 : node12365;
												assign node12365 = (inp[6]) ? 16'b0000000001111111 : node12366;
													assign node12366 = (inp[2]) ? node12372 : node12367;
														assign node12367 = (inp[10]) ? 16'b0000000011111111 : node12368;
															assign node12368 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12372 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12376 = (inp[7]) ? node12382 : node12377;
													assign node12377 = (inp[10]) ? node12379 : 16'b0000000011111111;
														assign node12379 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12382 = (inp[9]) ? node12386 : node12383;
														assign node12383 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12386 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node12389 = (inp[1]) ? node12399 : node12390;
												assign node12390 = (inp[6]) ? node12394 : node12391;
													assign node12391 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12394 = (inp[9]) ? 16'b0000000000011111 : node12395;
														assign node12395 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node12399 = (inp[10]) ? node12407 : node12400;
													assign node12400 = (inp[7]) ? node12404 : node12401;
														assign node12401 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12404 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node12407 = (inp[9]) ? node12411 : node12408;
														assign node12408 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node12411 = (inp[6]) ? 16'b0000000000001111 : node12412;
															assign node12412 = (inp[7]) ? node12414 : 16'b0000000000011111;
																assign node12414 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node12418 = (inp[1]) ? node12452 : node12419;
											assign node12419 = (inp[2]) ? node12431 : node12420;
												assign node12420 = (inp[10]) ? node12422 : 16'b0000000001111111;
													assign node12422 = (inp[9]) ? node12424 : 16'b0000000000011111;
														assign node12424 = (inp[14]) ? 16'b0000000000111111 : node12425;
															assign node12425 = (inp[6]) ? 16'b0000000000111111 : node12426;
																assign node12426 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12431 = (inp[9]) ? node12445 : node12432;
													assign node12432 = (inp[7]) ? 16'b0000000000011111 : node12433;
														assign node12433 = (inp[6]) ? node12439 : node12434;
															assign node12434 = (inp[10]) ? node12436 : 16'b0000000001111111;
																assign node12436 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node12439 = (inp[10]) ? node12441 : 16'b0000000000111111;
																assign node12441 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node12445 = (inp[6]) ? node12449 : node12446;
														assign node12446 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node12449 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node12452 = (inp[9]) ? node12470 : node12453;
												assign node12453 = (inp[10]) ? node12459 : node12454;
													assign node12454 = (inp[14]) ? node12456 : 16'b0000000001111111;
														assign node12456 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node12459 = (inp[14]) ? node12463 : node12460;
														assign node12460 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node12463 = (inp[7]) ? 16'b0000000000001111 : node12464;
															assign node12464 = (inp[2]) ? node12466 : 16'b0000000000011111;
																assign node12466 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node12470 = (inp[2]) ? node12480 : node12471;
													assign node12471 = (inp[10]) ? node12473 : 16'b0000000000111111;
														assign node12473 = (inp[7]) ? node12475 : 16'b0000000000011111;
															assign node12475 = (inp[6]) ? 16'b0000000000001111 : node12476;
																assign node12476 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node12480 = (inp[14]) ? node12484 : node12481;
														assign node12481 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node12484 = (inp[6]) ? node12486 : 16'b0000000000001111;
															assign node12486 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node12489 = (inp[12]) ? node14511 : node12490;
					assign node12490 = (inp[11]) ? node13486 : node12491;
						assign node12491 = (inp[15]) ? node12983 : node12492;
							assign node12492 = (inp[3]) ? node12736 : node12493;
								assign node12493 = (inp[9]) ? node12617 : node12494;
									assign node12494 = (inp[5]) ? node12568 : node12495;
										assign node12495 = (inp[7]) ? node12539 : node12496;
											assign node12496 = (inp[1]) ? node12518 : node12497;
												assign node12497 = (inp[6]) ? node12511 : node12498;
													assign node12498 = (inp[2]) ? node12506 : node12499;
														assign node12499 = (inp[14]) ? node12501 : 16'b0001111111111111;
															assign node12501 = (inp[10]) ? 16'b0000111111111111 : node12502;
																assign node12502 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node12506 = (inp[13]) ? node12508 : 16'b0000111111111111;
															assign node12508 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12511 = (inp[13]) ? 16'b0000011111111111 : node12512;
														assign node12512 = (inp[14]) ? node12514 : 16'b0000111111111111;
															assign node12514 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node12518 = (inp[2]) ? node12532 : node12519;
													assign node12519 = (inp[6]) ? node12527 : node12520;
														assign node12520 = (inp[10]) ? 16'b0000011111111111 : node12521;
															assign node12521 = (inp[13]) ? 16'b0000111111111111 : node12522;
																assign node12522 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node12527 = (inp[13]) ? node12529 : 16'b0000011111111111;
															assign node12529 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12532 = (inp[14]) ? 16'b0000000111111111 : node12533;
														assign node12533 = (inp[6]) ? 16'b0000001111111111 : node12534;
															assign node12534 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node12539 = (inp[1]) ? node12555 : node12540;
												assign node12540 = (inp[10]) ? node12550 : node12541;
													assign node12541 = (inp[6]) ? node12543 : 16'b0000111111111111;
														assign node12543 = (inp[14]) ? 16'b0000001111111111 : node12544;
															assign node12544 = (inp[13]) ? 16'b0000011111111111 : node12545;
																assign node12545 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12550 = (inp[13]) ? node12552 : 16'b0000011111111111;
														assign node12552 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12555 = (inp[14]) ? node12563 : node12556;
													assign node12556 = (inp[2]) ? node12560 : node12557;
														assign node12557 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12560 = (inp[10]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node12563 = (inp[13]) ? node12565 : 16'b0000000111111111;
														assign node12565 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12568 = (inp[2]) ? node12590 : node12569;
											assign node12569 = (inp[13]) ? node12579 : node12570;
												assign node12570 = (inp[1]) ? node12576 : node12571;
													assign node12571 = (inp[14]) ? node12573 : 16'b0000111111111111;
														assign node12573 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12576 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12579 = (inp[10]) ? node12587 : node12580;
													assign node12580 = (inp[6]) ? 16'b0000001111111111 : node12581;
														assign node12581 = (inp[14]) ? 16'b0000001111111111 : node12582;
															assign node12582 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12587 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node12590 = (inp[13]) ? node12602 : node12591;
												assign node12591 = (inp[14]) ? node12595 : node12592;
													assign node12592 = (inp[6]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node12595 = (inp[7]) ? 16'b0000000111111111 : node12596;
														assign node12596 = (inp[6]) ? node12598 : 16'b0000001111111111;
															assign node12598 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12602 = (inp[14]) ? node12612 : node12603;
													assign node12603 = (inp[10]) ? node12609 : node12604;
														assign node12604 = (inp[6]) ? 16'b0000000111111111 : node12605;
															assign node12605 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12609 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12612 = (inp[10]) ? node12614 : 16'b0000000011111111;
														assign node12614 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node12617 = (inp[14]) ? node12675 : node12618;
										assign node12618 = (inp[1]) ? node12648 : node12619;
											assign node12619 = (inp[6]) ? node12637 : node12620;
												assign node12620 = (inp[2]) ? node12628 : node12621;
													assign node12621 = (inp[10]) ? node12625 : node12622;
														assign node12622 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12625 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12628 = (inp[13]) ? 16'b0000001111111111 : node12629;
														assign node12629 = (inp[7]) ? 16'b0000001111111111 : node12630;
															assign node12630 = (inp[10]) ? node12632 : 16'b0000011111111111;
																assign node12632 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node12637 = (inp[5]) ? node12641 : node12638;
													assign node12638 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node12641 = (inp[13]) ? 16'b0000000111111111 : node12642;
														assign node12642 = (inp[10]) ? 16'b0000000111111111 : node12643;
															assign node12643 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node12648 = (inp[10]) ? node12660 : node12649;
												assign node12649 = (inp[6]) ? node12655 : node12650;
													assign node12650 = (inp[13]) ? node12652 : 16'b0000011111111111;
														assign node12652 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12655 = (inp[7]) ? 16'b0000000111111111 : node12656;
														assign node12656 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12660 = (inp[13]) ? node12662 : 16'b0000000111111111;
													assign node12662 = (inp[2]) ? 16'b0000000011111111 : node12663;
														assign node12663 = (inp[7]) ? node12669 : node12664;
															assign node12664 = (inp[6]) ? 16'b0000000111111111 : node12665;
																assign node12665 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node12669 = (inp[6]) ? 16'b0000000011111111 : node12670;
																assign node12670 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node12675 = (inp[2]) ? node12699 : node12676;
											assign node12676 = (inp[6]) ? node12688 : node12677;
												assign node12677 = (inp[5]) ? node12683 : node12678;
													assign node12678 = (inp[13]) ? 16'b0000001111111111 : node12679;
														assign node12679 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12683 = (inp[10]) ? node12685 : 16'b0000001111111111;
														assign node12685 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node12688 = (inp[7]) ? node12694 : node12689;
													assign node12689 = (inp[1]) ? 16'b0000000111111111 : node12690;
														assign node12690 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12694 = (inp[1]) ? node12696 : 16'b0000000111111111;
														assign node12696 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12699 = (inp[6]) ? node12719 : node12700;
												assign node12700 = (inp[13]) ? node12706 : node12701;
													assign node12701 = (inp[1]) ? 16'b0000000111111111 : node12702;
														assign node12702 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12706 = (inp[10]) ? node12710 : node12707;
														assign node12707 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12710 = (inp[5]) ? node12716 : node12711;
															assign node12711 = (inp[7]) ? 16'b0000000011111111 : node12712;
																assign node12712 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node12716 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12719 = (inp[13]) ? node12731 : node12720;
													assign node12720 = (inp[10]) ? node12726 : node12721;
														assign node12721 = (inp[1]) ? node12723 : 16'b0000000111111111;
															assign node12723 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12726 = (inp[5]) ? node12728 : 16'b0000000011111111;
															assign node12728 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12731 = (inp[5]) ? 16'b0000000001111111 : node12732;
														assign node12732 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node12736 = (inp[2]) ? node12864 : node12737;
									assign node12737 = (inp[6]) ? node12801 : node12738;
										assign node12738 = (inp[14]) ? node12770 : node12739;
											assign node12739 = (inp[10]) ? node12755 : node12740;
												assign node12740 = (inp[5]) ? node12746 : node12741;
													assign node12741 = (inp[9]) ? 16'b0000011111111111 : node12742;
														assign node12742 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12746 = (inp[1]) ? 16'b0000001111111111 : node12747;
														assign node12747 = (inp[13]) ? 16'b0000001111111111 : node12748;
															assign node12748 = (inp[9]) ? 16'b0000011111111111 : node12749;
																assign node12749 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node12755 = (inp[13]) ? node12767 : node12756;
													assign node12756 = (inp[1]) ? node12764 : node12757;
														assign node12757 = (inp[7]) ? node12759 : 16'b0000011111111111;
															assign node12759 = (inp[5]) ? node12761 : 16'b0000011111111111;
																assign node12761 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12764 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12767 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node12770 = (inp[9]) ? node12782 : node12771;
												assign node12771 = (inp[13]) ? node12777 : node12772;
													assign node12772 = (inp[1]) ? node12774 : 16'b0000001111111111;
														assign node12774 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12777 = (inp[10]) ? 16'b0000000011111111 : node12778;
														assign node12778 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node12782 = (inp[5]) ? node12790 : node12783;
													assign node12783 = (inp[1]) ? node12787 : node12784;
														assign node12784 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12787 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node12790 = (inp[13]) ? node12794 : node12791;
														assign node12791 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12794 = (inp[7]) ? 16'b0000000001111111 : node12795;
															assign node12795 = (inp[10]) ? node12797 : 16'b0000000011111111;
																assign node12797 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node12801 = (inp[5]) ? node12827 : node12802;
											assign node12802 = (inp[7]) ? node12812 : node12803;
												assign node12803 = (inp[1]) ? 16'b0000000111111111 : node12804;
													assign node12804 = (inp[13]) ? node12808 : node12805;
														assign node12805 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12808 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12812 = (inp[9]) ? node12818 : node12813;
													assign node12813 = (inp[10]) ? 16'b0000000111111111 : node12814;
														assign node12814 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12818 = (inp[13]) ? node12824 : node12819;
														assign node12819 = (inp[1]) ? 16'b0000000011111111 : node12820;
															assign node12820 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12824 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12827 = (inp[13]) ? node12843 : node12828;
												assign node12828 = (inp[1]) ? node12836 : node12829;
													assign node12829 = (inp[10]) ? node12831 : 16'b0000000111111111;
														assign node12831 = (inp[14]) ? 16'b0000000011111111 : node12832;
															assign node12832 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12836 = (inp[9]) ? node12840 : node12837;
														assign node12837 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node12840 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12843 = (inp[7]) ? node12853 : node12844;
													assign node12844 = (inp[10]) ? node12850 : node12845;
														assign node12845 = (inp[9]) ? node12847 : 16'b0000001111111111;
															assign node12847 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12850 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12853 = (inp[1]) ? node12861 : node12854;
														assign node12854 = (inp[10]) ? 16'b0000000001111111 : node12855;
															assign node12855 = (inp[14]) ? node12857 : 16'b0000000011111111;
																assign node12857 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12861 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12864 = (inp[13]) ? node12932 : node12865;
										assign node12865 = (inp[7]) ? node12903 : node12866;
											assign node12866 = (inp[6]) ? node12888 : node12867;
												assign node12867 = (inp[14]) ? node12873 : node12868;
													assign node12868 = (inp[1]) ? node12870 : 16'b0000001111111111;
														assign node12870 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12873 = (inp[1]) ? node12883 : node12874;
														assign node12874 = (inp[9]) ? node12880 : node12875;
															assign node12875 = (inp[10]) ? node12877 : 16'b0000001111111111;
																assign node12877 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node12880 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12883 = (inp[10]) ? node12885 : 16'b0000000111111111;
															assign node12885 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12888 = (inp[5]) ? node12894 : node12889;
													assign node12889 = (inp[1]) ? node12891 : 16'b0000001111111111;
														assign node12891 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12894 = (inp[14]) ? node12898 : node12895;
														assign node12895 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12898 = (inp[9]) ? 16'b0000000001111111 : node12899;
															assign node12899 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12903 = (inp[9]) ? node12919 : node12904;
												assign node12904 = (inp[5]) ? node12910 : node12905;
													assign node12905 = (inp[1]) ? 16'b0000000111111111 : node12906;
														assign node12906 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12910 = (inp[6]) ? node12914 : node12911;
														assign node12911 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12914 = (inp[1]) ? 16'b0000000001111111 : node12915;
															assign node12915 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12919 = (inp[1]) ? node12921 : 16'b0000000011111111;
													assign node12921 = (inp[10]) ? node12925 : node12922;
														assign node12922 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12925 = (inp[5]) ? node12927 : 16'b0000000001111111;
															assign node12927 = (inp[14]) ? 16'b0000000000111111 : node12928;
																assign node12928 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node12932 = (inp[5]) ? node12958 : node12933;
											assign node12933 = (inp[1]) ? node12943 : node12934;
												assign node12934 = (inp[6]) ? node12936 : 16'b0000000111111111;
													assign node12936 = (inp[9]) ? 16'b0000000011111111 : node12937;
														assign node12937 = (inp[7]) ? 16'b0000000011111111 : node12938;
															assign node12938 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12943 = (inp[10]) ? node12951 : node12944;
													assign node12944 = (inp[9]) ? node12948 : node12945;
														assign node12945 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12948 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12951 = (inp[6]) ? node12955 : node12952;
														assign node12952 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12955 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12958 = (inp[14]) ? node12970 : node12959;
												assign node12959 = (inp[10]) ? node12965 : node12960;
													assign node12960 = (inp[6]) ? 16'b0000000011111111 : node12961;
														assign node12961 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12965 = (inp[7]) ? node12967 : 16'b0000000011111111;
														assign node12967 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12970 = (inp[6]) ? node12978 : node12971;
													assign node12971 = (inp[1]) ? 16'b0000000001111111 : node12972;
														assign node12972 = (inp[10]) ? node12974 : 16'b0000000001111111;
															assign node12974 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12978 = (inp[9]) ? 16'b0000000000111111 : node12979;
														assign node12979 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node12983 = (inp[10]) ? node13211 : node12984;
								assign node12984 = (inp[14]) ? node13100 : node12985;
									assign node12985 = (inp[7]) ? node13039 : node12986;
										assign node12986 = (inp[9]) ? node13016 : node12987;
											assign node12987 = (inp[6]) ? node13003 : node12988;
												assign node12988 = (inp[5]) ? node12996 : node12989;
													assign node12989 = (inp[2]) ? node12991 : 16'b0000111111111111;
														assign node12991 = (inp[13]) ? 16'b0000011111111111 : node12992;
															assign node12992 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node12996 = (inp[13]) ? node12998 : 16'b0000011111111111;
														assign node12998 = (inp[3]) ? 16'b0000001111111111 : node12999;
															assign node12999 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13003 = (inp[1]) ? 16'b0000000111111111 : node13004;
													assign node13004 = (inp[13]) ? node13010 : node13005;
														assign node13005 = (inp[3]) ? 16'b0000001111111111 : node13006;
															assign node13006 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13010 = (inp[2]) ? node13012 : 16'b0000001111111111;
															assign node13012 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13016 = (inp[13]) ? node13026 : node13017;
												assign node13017 = (inp[6]) ? node13021 : node13018;
													assign node13018 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13021 = (inp[1]) ? node13023 : 16'b0000001111111111;
														assign node13023 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13026 = (inp[6]) ? node13034 : node13027;
													assign node13027 = (inp[1]) ? node13031 : node13028;
														assign node13028 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13031 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13034 = (inp[2]) ? 16'b0000000011111111 : node13035;
														assign node13035 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node13039 = (inp[6]) ? node13073 : node13040;
											assign node13040 = (inp[5]) ? node13058 : node13041;
												assign node13041 = (inp[2]) ? node13047 : node13042;
													assign node13042 = (inp[3]) ? node13044 : 16'b0000011111111111;
														assign node13044 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13047 = (inp[3]) ? node13055 : node13048;
														assign node13048 = (inp[1]) ? node13050 : 16'b0000001111111111;
															assign node13050 = (inp[9]) ? 16'b0000000111111111 : node13051;
																assign node13051 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13055 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13058 = (inp[3]) ? node13070 : node13059;
													assign node13059 = (inp[9]) ? node13065 : node13060;
														assign node13060 = (inp[2]) ? 16'b0000000111111111 : node13061;
															assign node13061 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13065 = (inp[2]) ? 16'b0000000011111111 : node13066;
															assign node13066 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13070 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node13073 = (inp[1]) ? node13085 : node13074;
												assign node13074 = (inp[13]) ? node13076 : 16'b0000000111111111;
													assign node13076 = (inp[5]) ? 16'b0000000011111111 : node13077;
														assign node13077 = (inp[2]) ? 16'b0000000011111111 : node13078;
															assign node13078 = (inp[3]) ? node13080 : 16'b0000000111111111;
																assign node13080 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13085 = (inp[3]) ? node13091 : node13086;
													assign node13086 = (inp[5]) ? node13088 : 16'b0000000111111111;
														assign node13088 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13091 = (inp[9]) ? node13095 : node13092;
														assign node13092 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13095 = (inp[13]) ? 16'b0000000000111111 : node13096;
															assign node13096 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node13100 = (inp[2]) ? node13152 : node13101;
										assign node13101 = (inp[9]) ? node13127 : node13102;
											assign node13102 = (inp[13]) ? node13120 : node13103;
												assign node13103 = (inp[7]) ? node13111 : node13104;
													assign node13104 = (inp[1]) ? node13106 : 16'b0000001111111111;
														assign node13106 = (inp[6]) ? node13108 : 16'b0000001111111111;
															assign node13108 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13111 = (inp[1]) ? 16'b0000000111111111 : node13112;
														assign node13112 = (inp[3]) ? 16'b0000000111111111 : node13113;
															assign node13113 = (inp[5]) ? 16'b0000001111111111 : node13114;
																assign node13114 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13120 = (inp[6]) ? node13124 : node13121;
													assign node13121 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13124 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13127 = (inp[6]) ? node13141 : node13128;
												assign node13128 = (inp[3]) ? node13132 : node13129;
													assign node13129 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13132 = (inp[1]) ? node13134 : 16'b0000000111111111;
														assign node13134 = (inp[7]) ? node13136 : 16'b0000000011111111;
															assign node13136 = (inp[13]) ? 16'b0000000001111111 : node13137;
																assign node13137 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13141 = (inp[1]) ? 16'b0000000001111111 : node13142;
													assign node13142 = (inp[7]) ? node13146 : node13143;
														assign node13143 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13146 = (inp[3]) ? 16'b0000000001111111 : node13147;
															assign node13147 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13152 = (inp[3]) ? node13178 : node13153;
											assign node13153 = (inp[1]) ? node13169 : node13154;
												assign node13154 = (inp[9]) ? 16'b0000000011111111 : node13155;
													assign node13155 = (inp[13]) ? node13159 : node13156;
														assign node13156 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13159 = (inp[5]) ? node13165 : node13160;
															assign node13160 = (inp[6]) ? node13162 : 16'b0000000111111111;
																assign node13162 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node13165 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13169 = (inp[6]) ? node13173 : node13170;
													assign node13170 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13173 = (inp[9]) ? node13175 : 16'b0000000001111111;
														assign node13175 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13178 = (inp[5]) ? node13196 : node13179;
												assign node13179 = (inp[13]) ? node13189 : node13180;
													assign node13180 = (inp[7]) ? 16'b0000000011111111 : node13181;
														assign node13181 = (inp[6]) ? node13183 : 16'b0000000111111111;
															assign node13183 = (inp[9]) ? 16'b0000000011111111 : node13184;
																assign node13184 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13189 = (inp[9]) ? 16'b0000000000111111 : node13190;
														assign node13190 = (inp[7]) ? 16'b0000000001111111 : node13191;
															assign node13191 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13196 = (inp[13]) ? node13206 : node13197;
													assign node13197 = (inp[6]) ? node13199 : 16'b0000000001111111;
														assign node13199 = (inp[9]) ? 16'b0000000000111111 : node13200;
															assign node13200 = (inp[1]) ? node13202 : 16'b0000000001111111;
																assign node13202 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13206 = (inp[9]) ? node13208 : 16'b0000000000111111;
														assign node13208 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node13211 = (inp[1]) ? node13347 : node13212;
									assign node13212 = (inp[2]) ? node13276 : node13213;
										assign node13213 = (inp[3]) ? node13249 : node13214;
											assign node13214 = (inp[13]) ? node13234 : node13215;
												assign node13215 = (inp[7]) ? node13227 : node13216;
													assign node13216 = (inp[9]) ? node13220 : node13217;
														assign node13217 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13220 = (inp[14]) ? 16'b0000000111111111 : node13221;
															assign node13221 = (inp[6]) ? 16'b0000001111111111 : node13222;
																assign node13222 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13227 = (inp[9]) ? node13231 : node13228;
														assign node13228 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node13231 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13234 = (inp[9]) ? node13244 : node13235;
													assign node13235 = (inp[14]) ? node13239 : node13236;
														assign node13236 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13239 = (inp[7]) ? node13241 : 16'b0000000111111111;
															assign node13241 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13244 = (inp[7]) ? 16'b0000000011111111 : node13245;
														assign node13245 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13249 = (inp[6]) ? node13263 : node13250;
												assign node13250 = (inp[14]) ? node13256 : node13251;
													assign node13251 = (inp[13]) ? 16'b0000000011111111 : node13252;
														assign node13252 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13256 = (inp[7]) ? node13260 : node13257;
														assign node13257 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13260 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13263 = (inp[9]) ? node13265 : 16'b0000000011111111;
													assign node13265 = (inp[14]) ? node13269 : node13266;
														assign node13266 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node13269 = (inp[5]) ? node13271 : 16'b0000000001111111;
															assign node13271 = (inp[13]) ? 16'b0000000000111111 : node13272;
																assign node13272 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13276 = (inp[7]) ? node13306 : node13277;
											assign node13277 = (inp[14]) ? node13293 : node13278;
												assign node13278 = (inp[13]) ? node13284 : node13279;
													assign node13279 = (inp[6]) ? 16'b0000000111111111 : node13280;
														assign node13280 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13284 = (inp[9]) ? node13288 : node13285;
														assign node13285 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node13288 = (inp[6]) ? node13290 : 16'b0000000011111111;
															assign node13290 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13293 = (inp[6]) ? node13301 : node13294;
													assign node13294 = (inp[5]) ? node13298 : node13295;
														assign node13295 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13298 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13301 = (inp[3]) ? node13303 : 16'b0000000001111111;
														assign node13303 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13306 = (inp[9]) ? node13330 : node13307;
												assign node13307 = (inp[13]) ? node13325 : node13308;
													assign node13308 = (inp[14]) ? node13314 : node13309;
														assign node13309 = (inp[5]) ? 16'b0000000011111111 : node13310;
															assign node13310 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13314 = (inp[3]) ? node13320 : node13315;
															assign node13315 = (inp[5]) ? node13317 : 16'b0000000011111111;
																assign node13317 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node13320 = (inp[6]) ? node13322 : 16'b0000000001111111;
																assign node13322 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13325 = (inp[14]) ? node13327 : 16'b0000000001111111;
														assign node13327 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13330 = (inp[14]) ? node13338 : node13331;
													assign node13331 = (inp[6]) ? node13335 : node13332;
														assign node13332 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13335 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13338 = (inp[5]) ? node13342 : node13339;
														assign node13339 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13342 = (inp[3]) ? node13344 : 16'b0000000000111111;
															assign node13344 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13347 = (inp[13]) ? node13415 : node13348;
										assign node13348 = (inp[5]) ? node13384 : node13349;
											assign node13349 = (inp[6]) ? node13367 : node13350;
												assign node13350 = (inp[7]) ? node13356 : node13351;
													assign node13351 = (inp[3]) ? node13353 : 16'b0000001111111111;
														assign node13353 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13356 = (inp[9]) ? node13362 : node13357;
														assign node13357 = (inp[14]) ? 16'b0000000011111111 : node13358;
															assign node13358 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13362 = (inp[3]) ? node13364 : 16'b0000000011111111;
															assign node13364 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13367 = (inp[14]) ? node13375 : node13368;
													assign node13368 = (inp[2]) ? node13372 : node13369;
														assign node13369 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13372 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13375 = (inp[7]) ? node13377 : 16'b0000000001111111;
														assign node13377 = (inp[2]) ? node13379 : 16'b0000000001111111;
															assign node13379 = (inp[3]) ? node13381 : 16'b0000000000111111;
																assign node13381 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node13384 = (inp[9]) ? node13400 : node13385;
												assign node13385 = (inp[14]) ? node13391 : node13386;
													assign node13386 = (inp[2]) ? node13388 : 16'b0000000011111111;
														assign node13388 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13391 = (inp[7]) ? node13395 : node13392;
														assign node13392 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13395 = (inp[3]) ? node13397 : 16'b0000000001111111;
															assign node13397 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13400 = (inp[7]) ? node13406 : node13401;
													assign node13401 = (inp[2]) ? node13403 : 16'b0000000001111111;
														assign node13403 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13406 = (inp[14]) ? 16'b0000000000011111 : node13407;
														assign node13407 = (inp[6]) ? node13409 : 16'b0000000001111111;
															assign node13409 = (inp[2]) ? node13411 : 16'b0000000000111111;
																assign node13411 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13415 = (inp[14]) ? node13457 : node13416;
											assign node13416 = (inp[3]) ? node13436 : node13417;
												assign node13417 = (inp[9]) ? node13425 : node13418;
													assign node13418 = (inp[7]) ? node13422 : node13419;
														assign node13419 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13422 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13425 = (inp[7]) ? node13429 : node13426;
														assign node13426 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13429 = (inp[6]) ? node13431 : 16'b0000000001111111;
															assign node13431 = (inp[5]) ? 16'b0000000000111111 : node13432;
																assign node13432 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13436 = (inp[5]) ? node13450 : node13437;
													assign node13437 = (inp[7]) ? node13443 : node13438;
														assign node13438 = (inp[2]) ? 16'b0000000001111111 : node13439;
															assign node13439 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13443 = (inp[9]) ? node13445 : 16'b0000000001111111;
															assign node13445 = (inp[6]) ? node13447 : 16'b0000000000111111;
																assign node13447 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13450 = (inp[6]) ? node13452 : 16'b0000000000111111;
														assign node13452 = (inp[7]) ? node13454 : 16'b0000000000011111;
															assign node13454 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node13457 = (inp[9]) ? node13477 : node13458;
												assign node13458 = (inp[7]) ? node13462 : node13459;
													assign node13459 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13462 = (inp[3]) ? node13472 : node13463;
														assign node13463 = (inp[2]) ? node13467 : node13464;
															assign node13464 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node13467 = (inp[5]) ? node13469 : 16'b0000000000111111;
																assign node13469 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node13472 = (inp[2]) ? 16'b0000000000011111 : node13473;
															assign node13473 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13477 = (inp[5]) ? 16'b0000000000011111 : node13478;
													assign node13478 = (inp[7]) ? node13480 : 16'b0000000000111111;
														assign node13480 = (inp[6]) ? 16'b0000000000011111 : node13481;
															assign node13481 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node13486 = (inp[5]) ? node13976 : node13487;
							assign node13487 = (inp[10]) ? node13717 : node13488;
								assign node13488 = (inp[7]) ? node13618 : node13489;
									assign node13489 = (inp[1]) ? node13565 : node13490;
										assign node13490 = (inp[14]) ? node13522 : node13491;
											assign node13491 = (inp[15]) ? node13507 : node13492;
												assign node13492 = (inp[13]) ? node13498 : node13493;
													assign node13493 = (inp[6]) ? 16'b0000011111111111 : node13494;
														assign node13494 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13498 = (inp[9]) ? node13504 : node13499;
														assign node13499 = (inp[3]) ? node13501 : 16'b0000011111111111;
															assign node13501 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13504 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node13507 = (inp[13]) ? node13513 : node13508;
													assign node13508 = (inp[9]) ? 16'b0000001111111111 : node13509;
														assign node13509 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13513 = (inp[3]) ? 16'b0000000111111111 : node13514;
														assign node13514 = (inp[9]) ? node13516 : 16'b0000001111111111;
															assign node13516 = (inp[2]) ? 16'b0000000111111111 : node13517;
																assign node13517 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node13522 = (inp[9]) ? node13542 : node13523;
												assign node13523 = (inp[13]) ? node13535 : node13524;
													assign node13524 = (inp[2]) ? node13532 : node13525;
														assign node13525 = (inp[6]) ? 16'b0000001111111111 : node13526;
															assign node13526 = (inp[15]) ? node13528 : 16'b0000011111111111;
																assign node13528 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13532 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node13535 = (inp[15]) ? node13539 : node13536;
														assign node13536 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node13539 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13542 = (inp[15]) ? node13554 : node13543;
													assign node13543 = (inp[2]) ? node13547 : node13544;
														assign node13544 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13547 = (inp[3]) ? 16'b0000000011111111 : node13548;
															assign node13548 = (inp[6]) ? node13550 : 16'b0000000111111111;
																assign node13550 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13554 = (inp[13]) ? node13562 : node13555;
														assign node13555 = (inp[2]) ? 16'b0000000011111111 : node13556;
															assign node13556 = (inp[6]) ? node13558 : 16'b0000000111111111;
																assign node13558 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13562 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13565 = (inp[15]) ? node13595 : node13566;
											assign node13566 = (inp[13]) ? node13582 : node13567;
												assign node13567 = (inp[14]) ? node13573 : node13568;
													assign node13568 = (inp[2]) ? node13570 : 16'b0000001111111111;
														assign node13570 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13573 = (inp[6]) ? node13579 : node13574;
														assign node13574 = (inp[3]) ? 16'b0000000111111111 : node13575;
															assign node13575 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13579 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node13582 = (inp[3]) ? node13586 : node13583;
													assign node13583 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13586 = (inp[2]) ? node13588 : 16'b0000000001111111;
														assign node13588 = (inp[14]) ? 16'b0000000011111111 : node13589;
															assign node13589 = (inp[6]) ? 16'b0000000011111111 : node13590;
																assign node13590 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13595 = (inp[14]) ? node13613 : node13596;
												assign node13596 = (inp[6]) ? node13606 : node13597;
													assign node13597 = (inp[3]) ? node13603 : node13598;
														assign node13598 = (inp[9]) ? 16'b0000000111111111 : node13599;
															assign node13599 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13603 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node13606 = (inp[13]) ? node13610 : node13607;
														assign node13607 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13610 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13613 = (inp[13]) ? 16'b0000000000011111 : node13614;
													assign node13614 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node13618 = (inp[9]) ? node13668 : node13619;
										assign node13619 = (inp[15]) ? node13643 : node13620;
											assign node13620 = (inp[13]) ? node13632 : node13621;
												assign node13621 = (inp[3]) ? node13627 : node13622;
													assign node13622 = (inp[2]) ? node13624 : 16'b0000001111111111;
														assign node13624 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13627 = (inp[14]) ? 16'b0000000111111111 : node13628;
														assign node13628 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13632 = (inp[14]) ? node13640 : node13633;
													assign node13633 = (inp[3]) ? 16'b0000000011111111 : node13634;
														assign node13634 = (inp[6]) ? node13636 : 16'b0000001111111111;
															assign node13636 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13640 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node13643 = (inp[3]) ? node13651 : node13644;
												assign node13644 = (inp[13]) ? node13646 : 16'b0000000111111111;
													assign node13646 = (inp[6]) ? node13648 : 16'b0000000111111111;
														assign node13648 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13651 = (inp[2]) ? node13657 : node13652;
													assign node13652 = (inp[1]) ? node13654 : 16'b0000000111111111;
														assign node13654 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13657 = (inp[1]) ? node13665 : node13658;
														assign node13658 = (inp[6]) ? node13660 : 16'b0000000011111111;
															assign node13660 = (inp[13]) ? 16'b0000000001111111 : node13661;
																assign node13661 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13665 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13668 = (inp[2]) ? node13694 : node13669;
											assign node13669 = (inp[6]) ? node13679 : node13670;
												assign node13670 = (inp[14]) ? node13674 : node13671;
													assign node13671 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node13674 = (inp[3]) ? 16'b0000000011111111 : node13675;
														assign node13675 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13679 = (inp[3]) ? node13689 : node13680;
													assign node13680 = (inp[15]) ? node13684 : node13681;
														assign node13681 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13684 = (inp[14]) ? node13686 : 16'b0000000011111111;
															assign node13686 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13689 = (inp[14]) ? 16'b0000000001111111 : node13690;
														assign node13690 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13694 = (inp[3]) ? node13704 : node13695;
												assign node13695 = (inp[15]) ? node13701 : node13696;
													assign node13696 = (inp[1]) ? node13698 : 16'b0000000011111111;
														assign node13698 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13701 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node13704 = (inp[1]) ? node13714 : node13705;
													assign node13705 = (inp[14]) ? node13707 : 16'b0000000001111111;
														assign node13707 = (inp[6]) ? node13709 : 16'b0000000001111111;
															assign node13709 = (inp[15]) ? 16'b0000000000111111 : node13710;
																assign node13710 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13714 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node13717 = (inp[14]) ? node13839 : node13718;
									assign node13718 = (inp[6]) ? node13788 : node13719;
										assign node13719 = (inp[9]) ? node13753 : node13720;
											assign node13720 = (inp[2]) ? node13742 : node13721;
												assign node13721 = (inp[3]) ? node13733 : node13722;
													assign node13722 = (inp[15]) ? node13730 : node13723;
														assign node13723 = (inp[1]) ? node13725 : 16'b0000111111111111;
															assign node13725 = (inp[7]) ? 16'b0000001111111111 : node13726;
																assign node13726 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13730 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13733 = (inp[7]) ? 16'b0000000111111111 : node13734;
														assign node13734 = (inp[13]) ? 16'b0000000111111111 : node13735;
															assign node13735 = (inp[15]) ? node13737 : 16'b0000001111111111;
																assign node13737 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13742 = (inp[7]) ? node13750 : node13743;
													assign node13743 = (inp[1]) ? node13745 : 16'b0000001111111111;
														assign node13745 = (inp[13]) ? node13747 : 16'b0000000111111111;
															assign node13747 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13750 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13753 = (inp[1]) ? node13767 : node13754;
												assign node13754 = (inp[13]) ? node13762 : node13755;
													assign node13755 = (inp[15]) ? node13757 : 16'b0000001111111111;
														assign node13757 = (inp[7]) ? 16'b0000000111111111 : node13758;
															assign node13758 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13762 = (inp[2]) ? 16'b0000000011111111 : node13763;
														assign node13763 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13767 = (inp[15]) ? node13781 : node13768;
													assign node13768 = (inp[3]) ? node13772 : node13769;
														assign node13769 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13772 = (inp[7]) ? node13778 : node13773;
															assign node13773 = (inp[13]) ? 16'b0000000011111111 : node13774;
																assign node13774 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node13778 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13781 = (inp[7]) ? node13785 : node13782;
														assign node13782 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13785 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13788 = (inp[15]) ? node13816 : node13789;
											assign node13789 = (inp[13]) ? node13799 : node13790;
												assign node13790 = (inp[9]) ? 16'b0000000011111111 : node13791;
													assign node13791 = (inp[1]) ? node13795 : node13792;
														assign node13792 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13795 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13799 = (inp[7]) ? node13809 : node13800;
													assign node13800 = (inp[1]) ? node13804 : node13801;
														assign node13801 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13804 = (inp[2]) ? 16'b0000000001111111 : node13805;
															assign node13805 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13809 = (inp[9]) ? node13813 : node13810;
														assign node13810 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13813 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13816 = (inp[3]) ? node13828 : node13817;
												assign node13817 = (inp[2]) ? node13823 : node13818;
													assign node13818 = (inp[1]) ? node13820 : 16'b0000000011111111;
														assign node13820 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13823 = (inp[1]) ? 16'b0000000000111111 : node13824;
														assign node13824 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node13828 = (inp[7]) ? node13834 : node13829;
													assign node13829 = (inp[1]) ? 16'b0000000001111111 : node13830;
														assign node13830 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13834 = (inp[1]) ? node13836 : 16'b0000000001111111;
														assign node13836 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13839 = (inp[7]) ? node13919 : node13840;
										assign node13840 = (inp[9]) ? node13886 : node13841;
											assign node13841 = (inp[3]) ? node13859 : node13842;
												assign node13842 = (inp[15]) ? node13852 : node13843;
													assign node13843 = (inp[6]) ? 16'b0000000111111111 : node13844;
														assign node13844 = (inp[1]) ? node13848 : node13845;
															assign node13845 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node13848 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13852 = (inp[13]) ? node13854 : 16'b0000000111111111;
														assign node13854 = (inp[1]) ? 16'b0000000001111111 : node13855;
															assign node13855 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13859 = (inp[13]) ? node13871 : node13860;
													assign node13860 = (inp[2]) ? node13866 : node13861;
														assign node13861 = (inp[1]) ? node13863 : 16'b0000000111111111;
															assign node13863 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13866 = (inp[1]) ? node13868 : 16'b0000000011111111;
															assign node13868 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13871 = (inp[2]) ? node13883 : node13872;
														assign node13872 = (inp[1]) ? node13878 : node13873;
															assign node13873 = (inp[15]) ? node13875 : 16'b0000000011111111;
																assign node13875 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node13878 = (inp[6]) ? 16'b0000000001111111 : node13879;
																assign node13879 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13883 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13886 = (inp[15]) ? node13900 : node13887;
												assign node13887 = (inp[13]) ? node13895 : node13888;
													assign node13888 = (inp[3]) ? 16'b0000000001111111 : node13889;
														assign node13889 = (inp[1]) ? node13891 : 16'b0000000111111111;
															assign node13891 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13895 = (inp[2]) ? node13897 : 16'b0000000001111111;
														assign node13897 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13900 = (inp[2]) ? node13910 : node13901;
													assign node13901 = (inp[1]) ? node13903 : 16'b0000000011111111;
														assign node13903 = (inp[13]) ? 16'b0000000000111111 : node13904;
															assign node13904 = (inp[3]) ? node13906 : 16'b0000000001111111;
																assign node13906 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13910 = (inp[1]) ? node13914 : node13911;
														assign node13911 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13914 = (inp[6]) ? node13916 : 16'b0000000000111111;
															assign node13916 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13919 = (inp[2]) ? node13947 : node13920;
											assign node13920 = (inp[6]) ? node13936 : node13921;
												assign node13921 = (inp[9]) ? node13933 : node13922;
													assign node13922 = (inp[3]) ? node13926 : node13923;
														assign node13923 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13926 = (inp[15]) ? 16'b0000000000111111 : node13927;
															assign node13927 = (inp[1]) ? node13929 : 16'b0000000011111111;
																assign node13929 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13933 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13936 = (inp[9]) ? node13942 : node13937;
													assign node13937 = (inp[13]) ? 16'b0000000000111111 : node13938;
														assign node13938 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13942 = (inp[13]) ? node13944 : 16'b0000000000111111;
														assign node13944 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node13947 = (inp[13]) ? node13957 : node13948;
												assign node13948 = (inp[6]) ? node13950 : 16'b0000000011111111;
													assign node13950 = (inp[15]) ? node13954 : node13951;
														assign node13951 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13954 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13957 = (inp[3]) ? node13963 : node13958;
													assign node13958 = (inp[1]) ? node13960 : 16'b0000000000111111;
														assign node13960 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node13963 = (inp[9]) ? node13969 : node13964;
														assign node13964 = (inp[6]) ? 16'b0000000000011111 : node13965;
															assign node13965 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node13969 = (inp[15]) ? node13971 : 16'b0000000000011111;
															assign node13971 = (inp[6]) ? 16'b0000000000001111 : node13972;
																assign node13972 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node13976 = (inp[2]) ? node14252 : node13977;
								assign node13977 = (inp[1]) ? node14119 : node13978;
									assign node13978 = (inp[14]) ? node14054 : node13979;
										assign node13979 = (inp[15]) ? node14017 : node13980;
											assign node13980 = (inp[3]) ? node13992 : node13981;
												assign node13981 = (inp[6]) ? node13989 : node13982;
													assign node13982 = (inp[9]) ? 16'b0000001111111111 : node13983;
														assign node13983 = (inp[7]) ? 16'b0000011111111111 : node13984;
															assign node13984 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node13989 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13992 = (inp[6]) ? node14006 : node13993;
													assign node13993 = (inp[7]) ? node13999 : node13994;
														assign node13994 = (inp[10]) ? node13996 : 16'b0000001111111111;
															assign node13996 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13999 = (inp[10]) ? 16'b0000000001111111 : node14000;
															assign node14000 = (inp[9]) ? 16'b0000000111111111 : node14001;
																assign node14001 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14006 = (inp[9]) ? node14014 : node14007;
														assign node14007 = (inp[13]) ? 16'b0000000011111111 : node14008;
															assign node14008 = (inp[10]) ? node14010 : 16'b0000000111111111;
																assign node14010 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14014 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node14017 = (inp[7]) ? node14039 : node14018;
												assign node14018 = (inp[6]) ? node14028 : node14019;
													assign node14019 = (inp[3]) ? node14025 : node14020;
														assign node14020 = (inp[10]) ? node14022 : 16'b0000011111111111;
															assign node14022 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14025 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14028 = (inp[9]) ? node14034 : node14029;
														assign node14029 = (inp[10]) ? 16'b0000000011111111 : node14030;
															assign node14030 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14034 = (inp[13]) ? node14036 : 16'b0000000011111111;
															assign node14036 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14039 = (inp[6]) ? node14047 : node14040;
													assign node14040 = (inp[10]) ? node14042 : 16'b0000000111111111;
														assign node14042 = (inp[13]) ? node14044 : 16'b0000000011111111;
															assign node14044 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14047 = (inp[9]) ? node14051 : node14048;
														assign node14048 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14051 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14054 = (inp[13]) ? node14084 : node14055;
											assign node14055 = (inp[15]) ? node14069 : node14056;
												assign node14056 = (inp[3]) ? 16'b0000000011111111 : node14057;
													assign node14057 = (inp[6]) ? node14063 : node14058;
														assign node14058 = (inp[7]) ? 16'b0000001111111111 : node14059;
															assign node14059 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node14063 = (inp[10]) ? 16'b0000000111111111 : node14064;
															assign node14064 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14069 = (inp[7]) ? node14075 : node14070;
													assign node14070 = (inp[9]) ? 16'b0000000011111111 : node14071;
														assign node14071 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14075 = (inp[9]) ? node14077 : 16'b0000000001111111;
														assign node14077 = (inp[3]) ? node14079 : 16'b0000000000111111;
															assign node14079 = (inp[6]) ? node14081 : 16'b0000000000111111;
																assign node14081 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14084 = (inp[15]) ? node14104 : node14085;
												assign node14085 = (inp[6]) ? node14097 : node14086;
													assign node14086 = (inp[10]) ? node14092 : node14087;
														assign node14087 = (inp[3]) ? node14089 : 16'b0000000111111111;
															assign node14089 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14092 = (inp[9]) ? 16'b0000000001111111 : node14093;
															assign node14093 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14097 = (inp[3]) ? node14099 : 16'b0000000001111111;
														assign node14099 = (inp[9]) ? 16'b0000000000111111 : node14100;
															assign node14100 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14104 = (inp[3]) ? node14114 : node14105;
													assign node14105 = (inp[10]) ? node14109 : node14106;
														assign node14106 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14109 = (inp[9]) ? node14111 : 16'b0000000001111111;
															assign node14111 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14114 = (inp[10]) ? node14116 : 16'b0000000000111111;
														assign node14116 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node14119 = (inp[6]) ? node14181 : node14120;
										assign node14120 = (inp[14]) ? node14162 : node14121;
											assign node14121 = (inp[9]) ? node14137 : node14122;
												assign node14122 = (inp[7]) ? node14132 : node14123;
													assign node14123 = (inp[3]) ? node14129 : node14124;
														assign node14124 = (inp[13]) ? 16'b0000000111111111 : node14125;
															assign node14125 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14129 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14132 = (inp[10]) ? node14134 : 16'b0000000111111111;
														assign node14134 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14137 = (inp[15]) ? node14151 : node14138;
													assign node14138 = (inp[10]) ? 16'b0000000001111111 : node14139;
														assign node14139 = (inp[3]) ? node14145 : node14140;
															assign node14140 = (inp[13]) ? node14142 : 16'b0000000111111111;
																assign node14142 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node14145 = (inp[7]) ? node14147 : 16'b0000000011111111;
																assign node14147 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14151 = (inp[7]) ? node14153 : 16'b0000000001111111;
														assign node14153 = (inp[13]) ? node14155 : 16'b0000000011111111;
															assign node14155 = (inp[10]) ? node14159 : node14156;
																assign node14156 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
																assign node14159 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14162 = (inp[9]) ? node14172 : node14163;
												assign node14163 = (inp[15]) ? 16'b0000000000111111 : node14164;
													assign node14164 = (inp[10]) ? 16'b0000000001111111 : node14165;
														assign node14165 = (inp[3]) ? node14167 : 16'b0000000011111111;
															assign node14167 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14172 = (inp[13]) ? node14176 : node14173;
													assign node14173 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node14176 = (inp[3]) ? node14178 : 16'b0000000000111111;
														assign node14178 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14181 = (inp[3]) ? node14217 : node14182;
											assign node14182 = (inp[13]) ? node14196 : node14183;
												assign node14183 = (inp[14]) ? node14189 : node14184;
													assign node14184 = (inp[10]) ? 16'b0000000011111111 : node14185;
														assign node14185 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14189 = (inp[9]) ? 16'b0000000001111111 : node14190;
														assign node14190 = (inp[10]) ? 16'b0000000001111111 : node14191;
															assign node14191 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14196 = (inp[9]) ? node14206 : node14197;
													assign node14197 = (inp[15]) ? node14203 : node14198;
														assign node14198 = (inp[14]) ? 16'b0000000001111111 : node14199;
															assign node14199 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14203 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node14206 = (inp[10]) ? node14212 : node14207;
														assign node14207 = (inp[7]) ? 16'b0000000000111111 : node14208;
															assign node14208 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14212 = (inp[14]) ? 16'b0000000000011111 : node14213;
															assign node14213 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14217 = (inp[13]) ? node14237 : node14218;
												assign node14218 = (inp[14]) ? node14230 : node14219;
													assign node14219 = (inp[15]) ? node14223 : node14220;
														assign node14220 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14223 = (inp[10]) ? 16'b0000000000111111 : node14224;
															assign node14224 = (inp[9]) ? node14226 : 16'b0000000001111111;
																assign node14226 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14230 = (inp[15]) ? node14234 : node14231;
														assign node14231 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14234 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14237 = (inp[10]) ? node14245 : node14238;
													assign node14238 = (inp[7]) ? node14240 : 16'b0000000001111111;
														assign node14240 = (inp[15]) ? node14242 : 16'b0000000000111111;
															assign node14242 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node14245 = (inp[15]) ? node14247 : 16'b0000000000011111;
														assign node14247 = (inp[14]) ? node14249 : 16'b0000000000001111;
															assign node14249 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node14252 = (inp[9]) ? node14376 : node14253;
									assign node14253 = (inp[14]) ? node14303 : node14254;
										assign node14254 = (inp[10]) ? node14282 : node14255;
											assign node14255 = (inp[6]) ? node14263 : node14256;
												assign node14256 = (inp[3]) ? node14258 : 16'b0000000111111111;
													assign node14258 = (inp[7]) ? 16'b0000000011111111 : node14259;
														assign node14259 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14263 = (inp[3]) ? node14275 : node14264;
													assign node14264 = (inp[15]) ? node14272 : node14265;
														assign node14265 = (inp[13]) ? 16'b0000000011111111 : node14266;
															assign node14266 = (inp[7]) ? node14268 : 16'b0000000111111111;
																assign node14268 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14272 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14275 = (inp[7]) ? node14279 : node14276;
														assign node14276 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14279 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14282 = (inp[6]) ? node14294 : node14283;
												assign node14283 = (inp[15]) ? node14285 : 16'b0000000111111111;
													assign node14285 = (inp[1]) ? node14291 : node14286;
														assign node14286 = (inp[7]) ? node14288 : 16'b0000000011111111;
															assign node14288 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14291 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14294 = (inp[13]) ? node14298 : node14295;
													assign node14295 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node14298 = (inp[1]) ? 16'b0000000000111111 : node14299;
														assign node14299 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14303 = (inp[7]) ? node14349 : node14304;
											assign node14304 = (inp[3]) ? node14320 : node14305;
												assign node14305 = (inp[10]) ? node14311 : node14306;
													assign node14306 = (inp[13]) ? 16'b0000000011111111 : node14307;
														assign node14307 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14311 = (inp[15]) ? node14317 : node14312;
														assign node14312 = (inp[6]) ? 16'b0000000001111111 : node14313;
															assign node14313 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node14317 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14320 = (inp[13]) ? node14334 : node14321;
													assign node14321 = (inp[6]) ? node14329 : node14322;
														assign node14322 = (inp[10]) ? node14324 : 16'b0000000011111111;
															assign node14324 = (inp[15]) ? node14326 : 16'b0000000001111111;
																assign node14326 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14329 = (inp[15]) ? 16'b0000000000111111 : node14330;
															assign node14330 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14334 = (inp[1]) ? node14340 : node14335;
														assign node14335 = (inp[15]) ? node14337 : 16'b0000000001111111;
															assign node14337 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14340 = (inp[6]) ? node14344 : node14341;
															assign node14341 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node14344 = (inp[15]) ? node14346 : 16'b0000000000011111;
																assign node14346 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node14349 = (inp[10]) ? node14365 : node14350;
												assign node14350 = (inp[1]) ? node14360 : node14351;
													assign node14351 = (inp[15]) ? 16'b0000000000111111 : node14352;
														assign node14352 = (inp[6]) ? node14354 : 16'b0000000001111111;
															assign node14354 = (inp[13]) ? node14356 : 16'b0000000001111111;
																assign node14356 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14360 = (inp[3]) ? 16'b0000000000111111 : node14361;
														assign node14361 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14365 = (inp[15]) ? node14373 : node14366;
													assign node14366 = (inp[6]) ? node14368 : 16'b0000000000111111;
														assign node14368 = (inp[3]) ? 16'b0000000000011111 : node14369;
															assign node14369 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14373 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node14376 = (inp[7]) ? node14444 : node14377;
										assign node14377 = (inp[6]) ? node14407 : node14378;
											assign node14378 = (inp[1]) ? node14386 : node14379;
												assign node14379 = (inp[13]) ? node14383 : node14380;
													assign node14380 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node14383 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14386 = (inp[13]) ? node14394 : node14387;
													assign node14387 = (inp[15]) ? 16'b0000000000111111 : node14388;
														assign node14388 = (inp[3]) ? 16'b0000000001111111 : node14389;
															assign node14389 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14394 = (inp[3]) ? node14402 : node14395;
														assign node14395 = (inp[10]) ? 16'b0000000000111111 : node14396;
															assign node14396 = (inp[15]) ? node14398 : 16'b0000000001111111;
																assign node14398 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14402 = (inp[10]) ? 16'b0000000000011111 : node14403;
															assign node14403 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14407 = (inp[15]) ? node14425 : node14408;
												assign node14408 = (inp[14]) ? node14420 : node14409;
													assign node14409 = (inp[13]) ? node14417 : node14410;
														assign node14410 = (inp[10]) ? node14412 : 16'b0000000001111111;
															assign node14412 = (inp[1]) ? node14414 : 16'b0000000001111111;
																assign node14414 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14417 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14420 = (inp[10]) ? node14422 : 16'b0000000000111111;
														assign node14422 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14425 = (inp[1]) ? node14433 : node14426;
													assign node14426 = (inp[3]) ? node14430 : node14427;
														assign node14427 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14430 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14433 = (inp[13]) ? node14439 : node14434;
														assign node14434 = (inp[3]) ? 16'b0000000000011111 : node14435;
															assign node14435 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14439 = (inp[10]) ? 16'b0000000000001111 : node14440;
															assign node14440 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14444 = (inp[3]) ? node14484 : node14445;
											assign node14445 = (inp[13]) ? node14463 : node14446;
												assign node14446 = (inp[6]) ? node14454 : node14447;
													assign node14447 = (inp[15]) ? node14449 : 16'b0000000011111111;
														assign node14449 = (inp[1]) ? node14451 : 16'b0000000001111111;
															assign node14451 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14454 = (inp[15]) ? node14458 : node14455;
														assign node14455 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14458 = (inp[10]) ? node14460 : 16'b0000000000111111;
															assign node14460 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14463 = (inp[14]) ? node14471 : node14464;
													assign node14464 = (inp[1]) ? node14466 : 16'b0000000000111111;
														assign node14466 = (inp[15]) ? node14468 : 16'b0000000000111111;
															assign node14468 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14471 = (inp[1]) ? node14479 : node14472;
														assign node14472 = (inp[15]) ? 16'b0000000000011111 : node14473;
															assign node14473 = (inp[10]) ? node14475 : 16'b0000000000111111;
																assign node14475 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14479 = (inp[6]) ? 16'b0000000000000111 : node14480;
															assign node14480 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node14484 = (inp[10]) ? node14498 : node14485;
												assign node14485 = (inp[14]) ? node14491 : node14486;
													assign node14486 = (inp[6]) ? node14488 : 16'b0000000001111111;
														assign node14488 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node14491 = (inp[1]) ? node14493 : 16'b0000000000111111;
														assign node14493 = (inp[15]) ? 16'b0000000000001111 : node14494;
															assign node14494 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node14498 = (inp[13]) ? node14506 : node14499;
													assign node14499 = (inp[14]) ? node14501 : 16'b0000000000011111;
														assign node14501 = (inp[1]) ? 16'b0000000000000111 : node14502;
															assign node14502 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node14506 = (inp[14]) ? node14508 : 16'b0000000000001111;
														assign node14508 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000001111;
					assign node14511 = (inp[15]) ? node15601 : node14512;
						assign node14512 = (inp[6]) ? node15032 : node14513;
							assign node14513 = (inp[3]) ? node14755 : node14514;
								assign node14514 = (inp[10]) ? node14634 : node14515;
									assign node14515 = (inp[14]) ? node14581 : node14516;
										assign node14516 = (inp[11]) ? node14544 : node14517;
											assign node14517 = (inp[9]) ? node14533 : node14518;
												assign node14518 = (inp[13]) ? node14528 : node14519;
													assign node14519 = (inp[7]) ? node14525 : node14520;
														assign node14520 = (inp[5]) ? 16'b0000011111111111 : node14521;
															assign node14521 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node14525 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14528 = (inp[5]) ? 16'b0000001111111111 : node14529;
														assign node14529 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node14533 = (inp[1]) ? node14535 : 16'b0000001111111111;
													assign node14535 = (inp[13]) ? node14537 : 16'b0000001111111111;
														assign node14537 = (inp[7]) ? node14539 : 16'b0000000111111111;
															assign node14539 = (inp[5]) ? 16'b0000000011111111 : node14540;
																assign node14540 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14544 = (inp[13]) ? node14562 : node14545;
												assign node14545 = (inp[7]) ? node14555 : node14546;
													assign node14546 = (inp[9]) ? node14552 : node14547;
														assign node14547 = (inp[2]) ? 16'b0000001111111111 : node14548;
															assign node14548 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node14552 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14555 = (inp[5]) ? 16'b0000000111111111 : node14556;
														assign node14556 = (inp[1]) ? 16'b0000000111111111 : node14557;
															assign node14557 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node14562 = (inp[1]) ? node14570 : node14563;
													assign node14563 = (inp[9]) ? 16'b0000000111111111 : node14564;
														assign node14564 = (inp[7]) ? 16'b0000000111111111 : node14565;
															assign node14565 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14570 = (inp[2]) ? node14578 : node14571;
														assign node14571 = (inp[9]) ? node14573 : 16'b0000000111111111;
															assign node14573 = (inp[5]) ? 16'b0000000011111111 : node14574;
																assign node14574 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14578 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node14581 = (inp[9]) ? node14607 : node14582;
											assign node14582 = (inp[1]) ? node14594 : node14583;
												assign node14583 = (inp[7]) ? node14589 : node14584;
													assign node14584 = (inp[11]) ? node14586 : 16'b0000001111111111;
														assign node14586 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14589 = (inp[2]) ? node14591 : 16'b0000000111111111;
														assign node14591 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node14594 = (inp[5]) ? node14596 : 16'b0000000111111111;
													assign node14596 = (inp[13]) ? node14604 : node14597;
														assign node14597 = (inp[11]) ? 16'b0000000011111111 : node14598;
															assign node14598 = (inp[7]) ? 16'b0000000111111111 : node14599;
																assign node14599 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14604 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14607 = (inp[7]) ? node14615 : node14608;
												assign node14608 = (inp[5]) ? node14610 : 16'b0000000111111111;
													assign node14610 = (inp[1]) ? 16'b0000000001111111 : node14611;
														assign node14611 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14615 = (inp[13]) ? node14625 : node14616;
													assign node14616 = (inp[1]) ? node14618 : 16'b0000000111111111;
														assign node14618 = (inp[2]) ? 16'b0000000001111111 : node14619;
															assign node14619 = (inp[11]) ? node14621 : 16'b0000000011111111;
																assign node14621 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14625 = (inp[2]) ? node14629 : node14626;
														assign node14626 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14629 = (inp[1]) ? node14631 : 16'b0000000001111111;
															assign node14631 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node14634 = (inp[5]) ? node14696 : node14635;
										assign node14635 = (inp[1]) ? node14665 : node14636;
											assign node14636 = (inp[13]) ? node14654 : node14637;
												assign node14637 = (inp[11]) ? node14645 : node14638;
													assign node14638 = (inp[9]) ? node14642 : node14639;
														assign node14639 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node14642 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14645 = (inp[7]) ? node14647 : 16'b0000001111111111;
														assign node14647 = (inp[9]) ? 16'b0000000001111111 : node14648;
															assign node14648 = (inp[14]) ? node14650 : 16'b0000000111111111;
																assign node14650 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14654 = (inp[2]) ? node14656 : 16'b0000000111111111;
													assign node14656 = (inp[11]) ? 16'b0000000011111111 : node14657;
														assign node14657 = (inp[14]) ? node14659 : 16'b0000000111111111;
															assign node14659 = (inp[7]) ? 16'b0000000011111111 : node14660;
																assign node14660 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14665 = (inp[9]) ? node14685 : node14666;
												assign node14666 = (inp[11]) ? node14676 : node14667;
													assign node14667 = (inp[13]) ? node14671 : node14668;
														assign node14668 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14671 = (inp[14]) ? node14673 : 16'b0000000111111111;
															assign node14673 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node14676 = (inp[13]) ? node14680 : node14677;
														assign node14677 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14680 = (inp[7]) ? 16'b0000000001111111 : node14681;
															assign node14681 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14685 = (inp[7]) ? node14687 : 16'b0000000011111111;
													assign node14687 = (inp[11]) ? node14691 : node14688;
														assign node14688 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14691 = (inp[14]) ? 16'b0000000000111111 : node14692;
															assign node14692 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14696 = (inp[7]) ? node14718 : node14697;
											assign node14697 = (inp[14]) ? node14707 : node14698;
												assign node14698 = (inp[9]) ? 16'b0000000011111111 : node14699;
													assign node14699 = (inp[11]) ? node14701 : 16'b0000000111111111;
														assign node14701 = (inp[13]) ? 16'b0000000011111111 : node14702;
															assign node14702 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14707 = (inp[11]) ? 16'b0000000001111111 : node14708;
													assign node14708 = (inp[1]) ? node14712 : node14709;
														assign node14709 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14712 = (inp[13]) ? 16'b0000000001111111 : node14713;
															assign node14713 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14718 = (inp[2]) ? node14732 : node14719;
												assign node14719 = (inp[1]) ? node14729 : node14720;
													assign node14720 = (inp[14]) ? node14726 : node14721;
														assign node14721 = (inp[11]) ? 16'b0000000011111111 : node14722;
															assign node14722 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14726 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14729 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node14732 = (inp[13]) ? node14746 : node14733;
													assign node14733 = (inp[9]) ? node14741 : node14734;
														assign node14734 = (inp[14]) ? node14736 : 16'b0000000011111111;
															assign node14736 = (inp[1]) ? 16'b0000000001111111 : node14737;
																assign node14737 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14741 = (inp[14]) ? 16'b0000000000111111 : node14742;
															assign node14742 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14746 = (inp[1]) ? node14750 : node14747;
														assign node14747 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node14750 = (inp[11]) ? node14752 : 16'b0000000000011111;
															assign node14752 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node14755 = (inp[13]) ? node14907 : node14756;
									assign node14756 = (inp[14]) ? node14838 : node14757;
										assign node14757 = (inp[7]) ? node14803 : node14758;
											assign node14758 = (inp[2]) ? node14780 : node14759;
												assign node14759 = (inp[1]) ? node14775 : node14760;
													assign node14760 = (inp[5]) ? node14768 : node14761;
														assign node14761 = (inp[10]) ? 16'b0000001111111111 : node14762;
															assign node14762 = (inp[11]) ? node14764 : 16'b0000011111111111;
																assign node14764 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node14768 = (inp[10]) ? 16'b0000000111111111 : node14769;
															assign node14769 = (inp[9]) ? node14771 : 16'b0000001111111111;
																assign node14771 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14775 = (inp[5]) ? 16'b0000000011111111 : node14776;
														assign node14776 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node14780 = (inp[5]) ? node14790 : node14781;
													assign node14781 = (inp[9]) ? node14785 : node14782;
														assign node14782 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node14785 = (inp[10]) ? node14787 : 16'b0000000111111111;
															assign node14787 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14790 = (inp[11]) ? node14798 : node14791;
														assign node14791 = (inp[9]) ? 16'b0000000011111111 : node14792;
															assign node14792 = (inp[10]) ? node14794 : 16'b0000000111111111;
																assign node14794 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14798 = (inp[9]) ? 16'b0000000001111111 : node14799;
															assign node14799 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14803 = (inp[11]) ? node14825 : node14804;
												assign node14804 = (inp[9]) ? node14814 : node14805;
													assign node14805 = (inp[5]) ? 16'b0000000011111111 : node14806;
														assign node14806 = (inp[1]) ? 16'b0000000111111111 : node14807;
															assign node14807 = (inp[10]) ? node14809 : 16'b0000001111111111;
																assign node14809 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14814 = (inp[10]) ? node14818 : node14815;
														assign node14815 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14818 = (inp[2]) ? node14820 : 16'b0000000011111111;
															assign node14820 = (inp[1]) ? 16'b0000000001111111 : node14821;
																assign node14821 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14825 = (inp[2]) ? node14833 : node14826;
													assign node14826 = (inp[5]) ? node14830 : node14827;
														assign node14827 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14830 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14833 = (inp[9]) ? node14835 : 16'b0000000001111111;
														assign node14835 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14838 = (inp[5]) ? node14874 : node14839;
											assign node14839 = (inp[10]) ? node14859 : node14840;
												assign node14840 = (inp[9]) ? node14850 : node14841;
													assign node14841 = (inp[7]) ? node14845 : node14842;
														assign node14842 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node14845 = (inp[2]) ? node14847 : 16'b0000000111111111;
															assign node14847 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14850 = (inp[1]) ? node14856 : node14851;
														assign node14851 = (inp[2]) ? 16'b0000000011111111 : node14852;
															assign node14852 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14856 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14859 = (inp[1]) ? node14865 : node14860;
													assign node14860 = (inp[2]) ? node14862 : 16'b0000000011111111;
														assign node14862 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14865 = (inp[11]) ? node14867 : 16'b0000000011111111;
														assign node14867 = (inp[7]) ? node14871 : node14868;
															assign node14868 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node14871 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14874 = (inp[10]) ? node14894 : node14875;
												assign node14875 = (inp[1]) ? node14883 : node14876;
													assign node14876 = (inp[2]) ? node14880 : node14877;
														assign node14877 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14880 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14883 = (inp[7]) ? node14887 : node14884;
														assign node14884 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14887 = (inp[11]) ? node14889 : 16'b0000000001111111;
															assign node14889 = (inp[2]) ? 16'b0000000000111111 : node14890;
																assign node14890 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14894 = (inp[1]) ? node14902 : node14895;
													assign node14895 = (inp[7]) ? node14897 : 16'b0000000001111111;
														assign node14897 = (inp[9]) ? node14899 : 16'b0000000001111111;
															assign node14899 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14902 = (inp[2]) ? node14904 : 16'b0000000000111111;
														assign node14904 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node14907 = (inp[11]) ? node14953 : node14908;
										assign node14908 = (inp[1]) ? node14928 : node14909;
											assign node14909 = (inp[7]) ? node14919 : node14910;
												assign node14910 = (inp[14]) ? node14914 : node14911;
													assign node14911 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14914 = (inp[5]) ? 16'b0000000011111111 : node14915;
														assign node14915 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node14919 = (inp[10]) ? node14925 : node14920;
													assign node14920 = (inp[14]) ? 16'b0000000011111111 : node14921;
														assign node14921 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14925 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14928 = (inp[7]) ? node14938 : node14929;
												assign node14929 = (inp[9]) ? node14933 : node14930;
													assign node14930 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14933 = (inp[5]) ? 16'b0000000000111111 : node14934;
														assign node14934 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14938 = (inp[10]) ? node14946 : node14939;
													assign node14939 = (inp[14]) ? node14941 : 16'b0000000001111111;
														assign node14941 = (inp[5]) ? 16'b0000000000111111 : node14942;
															assign node14942 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14946 = (inp[5]) ? node14948 : 16'b0000000000111111;
														assign node14948 = (inp[14]) ? node14950 : 16'b0000000000111111;
															assign node14950 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14953 = (inp[7]) ? node14991 : node14954;
											assign node14954 = (inp[14]) ? node14972 : node14955;
												assign node14955 = (inp[9]) ? node14965 : node14956;
													assign node14956 = (inp[2]) ? node14962 : node14957;
														assign node14957 = (inp[1]) ? 16'b0000000011111111 : node14958;
															assign node14958 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14962 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14965 = (inp[5]) ? node14969 : node14966;
														assign node14966 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14969 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node14972 = (inp[9]) ? node14978 : node14973;
													assign node14973 = (inp[5]) ? node14975 : 16'b0000000001111111;
														assign node14975 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14978 = (inp[5]) ? node14986 : node14979;
														assign node14979 = (inp[1]) ? 16'b0000000000111111 : node14980;
															assign node14980 = (inp[2]) ? node14982 : 16'b0000000001111111;
																assign node14982 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14986 = (inp[2]) ? node14988 : 16'b0000000000111111;
															assign node14988 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14991 = (inp[2]) ? node15011 : node14992;
												assign node14992 = (inp[10]) ? node15004 : node14993;
													assign node14993 = (inp[5]) ? node15001 : node14994;
														assign node14994 = (inp[14]) ? 16'b0000000001111111 : node14995;
															assign node14995 = (inp[1]) ? node14997 : 16'b0000000011111111;
																assign node14997 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15001 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15004 = (inp[5]) ? node15006 : 16'b0000000000111111;
														assign node15006 = (inp[14]) ? 16'b0000000000011111 : node15007;
															assign node15007 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15011 = (inp[1]) ? node15023 : node15012;
													assign node15012 = (inp[14]) ? node15016 : node15013;
														assign node15013 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15016 = (inp[5]) ? 16'b0000000000011111 : node15017;
															assign node15017 = (inp[10]) ? node15019 : 16'b0000000000111111;
																assign node15019 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15023 = (inp[9]) ? node15029 : node15024;
														assign node15024 = (inp[10]) ? 16'b0000000000011111 : node15025;
															assign node15025 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15029 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node15032 = (inp[2]) ? node15302 : node15033;
								assign node15033 = (inp[11]) ? node15163 : node15034;
									assign node15034 = (inp[14]) ? node15084 : node15035;
										assign node15035 = (inp[3]) ? node15061 : node15036;
											assign node15036 = (inp[7]) ? node15052 : node15037;
												assign node15037 = (inp[10]) ? node15045 : node15038;
													assign node15038 = (inp[1]) ? 16'b0000001111111111 : node15039;
														assign node15039 = (inp[13]) ? 16'b0000001111111111 : node15040;
															assign node15040 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node15045 = (inp[5]) ? 16'b0000000111111111 : node15046;
														assign node15046 = (inp[1]) ? node15048 : 16'b0000001111111111;
															assign node15048 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15052 = (inp[10]) ? node15058 : node15053;
													assign node15053 = (inp[13]) ? 16'b0000000111111111 : node15054;
														assign node15054 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node15058 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15061 = (inp[13]) ? node15071 : node15062;
												assign node15062 = (inp[9]) ? node15064 : 16'b0000000111111111;
													assign node15064 = (inp[7]) ? 16'b0000000011111111 : node15065;
														assign node15065 = (inp[10]) ? node15067 : 16'b0000000111111111;
															assign node15067 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15071 = (inp[9]) ? node15077 : node15072;
													assign node15072 = (inp[10]) ? 16'b0000000011111111 : node15073;
														assign node15073 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15077 = (inp[7]) ? node15081 : node15078;
														assign node15078 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15081 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15084 = (inp[5]) ? node15122 : node15085;
											assign node15085 = (inp[3]) ? node15109 : node15086;
												assign node15086 = (inp[7]) ? node15096 : node15087;
													assign node15087 = (inp[1]) ? node15093 : node15088;
														assign node15088 = (inp[10]) ? 16'b0000000111111111 : node15089;
															assign node15089 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15093 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15096 = (inp[9]) ? node15104 : node15097;
														assign node15097 = (inp[10]) ? 16'b0000000011111111 : node15098;
															assign node15098 = (inp[13]) ? node15100 : 16'b0000000111111111;
																assign node15100 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15104 = (inp[10]) ? node15106 : 16'b0000000011111111;
															assign node15106 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15109 = (inp[1]) ? node15115 : node15110;
													assign node15110 = (inp[7]) ? node15112 : 16'b0000000011111111;
														assign node15112 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15115 = (inp[7]) ? node15119 : node15116;
														assign node15116 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15119 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15122 = (inp[7]) ? node15146 : node15123;
												assign node15123 = (inp[1]) ? node15135 : node15124;
													assign node15124 = (inp[9]) ? node15132 : node15125;
														assign node15125 = (inp[10]) ? node15127 : 16'b0000000111111111;
															assign node15127 = (inp[3]) ? 16'b0000000011111111 : node15128;
																assign node15128 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15132 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node15135 = (inp[3]) ? node15139 : node15136;
														assign node15136 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15139 = (inp[13]) ? 16'b0000000000111111 : node15140;
															assign node15140 = (inp[9]) ? node15142 : 16'b0000000001111111;
																assign node15142 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15146 = (inp[9]) ? node15152 : node15147;
													assign node15147 = (inp[3]) ? node15149 : 16'b0000000001111111;
														assign node15149 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15152 = (inp[1]) ? node15160 : node15153;
														assign node15153 = (inp[13]) ? node15155 : 16'b0000000011111111;
															assign node15155 = (inp[3]) ? 16'b0000000000111111 : node15156;
																assign node15156 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15160 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node15163 = (inp[3]) ? node15243 : node15164;
										assign node15164 = (inp[14]) ? node15202 : node15165;
											assign node15165 = (inp[9]) ? node15181 : node15166;
												assign node15166 = (inp[5]) ? node15174 : node15167;
													assign node15167 = (inp[1]) ? node15171 : node15168;
														assign node15168 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15171 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15174 = (inp[13]) ? 16'b0000000001111111 : node15175;
														assign node15175 = (inp[7]) ? 16'b0000000011111111 : node15176;
															assign node15176 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15181 = (inp[7]) ? node15191 : node15182;
													assign node15182 = (inp[5]) ? 16'b0000000001111111 : node15183;
														assign node15183 = (inp[13]) ? 16'b0000000011111111 : node15184;
															assign node15184 = (inp[10]) ? node15186 : 16'b0000000111111111;
																assign node15186 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15191 = (inp[10]) ? node15193 : 16'b0000000001111111;
														assign node15193 = (inp[5]) ? node15199 : node15194;
															assign node15194 = (inp[1]) ? node15196 : 16'b0000000001111111;
																assign node15196 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node15199 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node15202 = (inp[1]) ? node15222 : node15203;
												assign node15203 = (inp[10]) ? node15209 : node15204;
													assign node15204 = (inp[9]) ? 16'b0000000011111111 : node15205;
														assign node15205 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15209 = (inp[7]) ? node15217 : node15210;
														assign node15210 = (inp[5]) ? node15212 : 16'b0000000011111111;
															assign node15212 = (inp[13]) ? 16'b0000000001111111 : node15213;
																assign node15213 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15217 = (inp[5]) ? 16'b0000000000111111 : node15218;
															assign node15218 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15222 = (inp[13]) ? node15230 : node15223;
													assign node15223 = (inp[7]) ? 16'b0000000001111111 : node15224;
														assign node15224 = (inp[10]) ? 16'b0000000001111111 : node15225;
															assign node15225 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15230 = (inp[10]) ? node15236 : node15231;
														assign node15231 = (inp[7]) ? node15233 : 16'b0000000001111111;
															assign node15233 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15236 = (inp[9]) ? 16'b0000000000011111 : node15237;
															assign node15237 = (inp[7]) ? 16'b0000000000111111 : node15238;
																assign node15238 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15243 = (inp[14]) ? node15277 : node15244;
											assign node15244 = (inp[7]) ? node15262 : node15245;
												assign node15245 = (inp[10]) ? node15251 : node15246;
													assign node15246 = (inp[13]) ? 16'b0000000011111111 : node15247;
														assign node15247 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15251 = (inp[9]) ? node15259 : node15252;
														assign node15252 = (inp[1]) ? node15254 : 16'b0000000011111111;
															assign node15254 = (inp[5]) ? 16'b0000000001111111 : node15255;
																assign node15255 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15259 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15262 = (inp[10]) ? node15264 : 16'b0000000001111111;
													assign node15264 = (inp[1]) ? node15270 : node15265;
														assign node15265 = (inp[13]) ? 16'b0000000000111111 : node15266;
															assign node15266 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15270 = (inp[9]) ? node15272 : 16'b0000000000111111;
															assign node15272 = (inp[13]) ? 16'b0000000000011111 : node15273;
																assign node15273 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node15277 = (inp[13]) ? node15287 : node15278;
												assign node15278 = (inp[1]) ? node15280 : 16'b0000000001111111;
													assign node15280 = (inp[10]) ? 16'b0000000000111111 : node15281;
														assign node15281 = (inp[9]) ? node15283 : 16'b0000000001111111;
															assign node15283 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15287 = (inp[5]) ? node15293 : node15288;
													assign node15288 = (inp[1]) ? 16'b0000000000111111 : node15289;
														assign node15289 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15293 = (inp[1]) ? 16'b0000000000011111 : node15294;
														assign node15294 = (inp[10]) ? 16'b0000000000011111 : node15295;
															assign node15295 = (inp[7]) ? 16'b0000000000111111 : node15296;
																assign node15296 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node15302 = (inp[14]) ? node15430 : node15303;
									assign node15303 = (inp[5]) ? node15359 : node15304;
										assign node15304 = (inp[11]) ? node15328 : node15305;
											assign node15305 = (inp[3]) ? node15315 : node15306;
												assign node15306 = (inp[10]) ? node15308 : 16'b0000000111111111;
													assign node15308 = (inp[13]) ? 16'b0000000001111111 : node15309;
														assign node15309 = (inp[1]) ? node15311 : 16'b0000000111111111;
															assign node15311 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15315 = (inp[10]) ? node15323 : node15316;
													assign node15316 = (inp[7]) ? node15320 : node15317;
														assign node15317 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15320 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15323 = (inp[13]) ? 16'b0000000001111111 : node15324;
														assign node15324 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15328 = (inp[1]) ? node15346 : node15329;
												assign node15329 = (inp[7]) ? node15337 : node15330;
													assign node15330 = (inp[3]) ? node15332 : 16'b0000000011111111;
														assign node15332 = (inp[9]) ? node15334 : 16'b0000000011111111;
															assign node15334 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15337 = (inp[3]) ? node15341 : node15338;
														assign node15338 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15341 = (inp[9]) ? node15343 : 16'b0000000001111111;
															assign node15343 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15346 = (inp[10]) ? node15352 : node15347;
													assign node15347 = (inp[9]) ? 16'b0000000001111111 : node15348;
														assign node15348 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15352 = (inp[9]) ? 16'b0000000000111111 : node15353;
														assign node15353 = (inp[13]) ? node15355 : 16'b0000000001111111;
															assign node15355 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15359 = (inp[3]) ? node15399 : node15360;
											assign node15360 = (inp[13]) ? node15380 : node15361;
												assign node15361 = (inp[11]) ? node15371 : node15362;
													assign node15362 = (inp[7]) ? 16'b0000000001111111 : node15363;
														assign node15363 = (inp[10]) ? node15365 : 16'b0000000111111111;
															assign node15365 = (inp[1]) ? 16'b0000000011111111 : node15366;
																assign node15366 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15371 = (inp[1]) ? node15377 : node15372;
														assign node15372 = (inp[9]) ? node15374 : 16'b0000000011111111;
															assign node15374 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15377 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15380 = (inp[1]) ? node15394 : node15381;
													assign node15381 = (inp[9]) ? node15383 : 16'b0000000001111111;
														assign node15383 = (inp[10]) ? node15389 : node15384;
															assign node15384 = (inp[7]) ? node15386 : 16'b0000000001111111;
																assign node15386 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node15389 = (inp[7]) ? 16'b0000000000111111 : node15390;
																assign node15390 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15394 = (inp[10]) ? 16'b0000000000111111 : node15395;
														assign node15395 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15399 = (inp[10]) ? node15415 : node15400;
												assign node15400 = (inp[11]) ? node15406 : node15401;
													assign node15401 = (inp[13]) ? node15403 : 16'b0000000011111111;
														assign node15403 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15406 = (inp[7]) ? 16'b0000000000111111 : node15407;
														assign node15407 = (inp[9]) ? 16'b0000000000111111 : node15408;
															assign node15408 = (inp[13]) ? node15410 : 16'b0000000001111111;
																assign node15410 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15415 = (inp[9]) ? node15421 : node15416;
													assign node15416 = (inp[7]) ? node15418 : 16'b0000000000111111;
														assign node15418 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node15421 = (inp[1]) ? node15423 : 16'b0000000000011111;
														assign node15423 = (inp[13]) ? 16'b0000000000001111 : node15424;
															assign node15424 = (inp[11]) ? 16'b0000000000001111 : node15425;
																assign node15425 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node15430 = (inp[5]) ? node15526 : node15431;
										assign node15431 = (inp[11]) ? node15465 : node15432;
											assign node15432 = (inp[10]) ? node15448 : node15433;
												assign node15433 = (inp[7]) ? node15443 : node15434;
													assign node15434 = (inp[13]) ? node15440 : node15435;
														assign node15435 = (inp[9]) ? 16'b0000000011111111 : node15436;
															assign node15436 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15440 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15443 = (inp[13]) ? 16'b0000000000111111 : node15444;
														assign node15444 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node15448 = (inp[13]) ? node15460 : node15449;
													assign node15449 = (inp[7]) ? node15453 : node15450;
														assign node15450 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15453 = (inp[1]) ? 16'b0000000000111111 : node15454;
															assign node15454 = (inp[9]) ? node15456 : 16'b0000000001111111;
																assign node15456 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15460 = (inp[3]) ? 16'b0000000000011111 : node15461;
														assign node15461 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15465 = (inp[7]) ? node15501 : node15466;
												assign node15466 = (inp[3]) ? node15478 : node15467;
													assign node15467 = (inp[1]) ? node15471 : node15468;
														assign node15468 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15471 = (inp[10]) ? node15473 : 16'b0000000001111111;
															assign node15473 = (inp[13]) ? 16'b0000000000111111 : node15474;
																assign node15474 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15478 = (inp[10]) ? node15488 : node15479;
														assign node15479 = (inp[13]) ? node15483 : node15480;
															assign node15480 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node15483 = (inp[1]) ? 16'b0000000000111111 : node15484;
																assign node15484 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15488 = (inp[1]) ? node15496 : node15489;
															assign node15489 = (inp[9]) ? node15493 : node15490;
																assign node15490 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
																assign node15493 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node15496 = (inp[13]) ? 16'b0000000000011111 : node15497;
																assign node15497 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15501 = (inp[9]) ? node15517 : node15502;
													assign node15502 = (inp[3]) ? node15506 : node15503;
														assign node15503 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node15506 = (inp[10]) ? node15512 : node15507;
															assign node15507 = (inp[1]) ? node15509 : 16'b0000000000111111;
																assign node15509 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node15512 = (inp[1]) ? 16'b0000000000011111 : node15513;
																assign node15513 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15517 = (inp[3]) ? 16'b0000000000001111 : node15518;
														assign node15518 = (inp[1]) ? node15520 : 16'b0000000000111111;
															assign node15520 = (inp[13]) ? node15522 : 16'b0000000000011111;
																assign node15522 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node15526 = (inp[1]) ? node15568 : node15527;
											assign node15527 = (inp[13]) ? node15547 : node15528;
												assign node15528 = (inp[9]) ? node15536 : node15529;
													assign node15529 = (inp[10]) ? node15533 : node15530;
														assign node15530 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15533 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15536 = (inp[7]) ? node15540 : node15537;
														assign node15537 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15540 = (inp[3]) ? 16'b0000000000001111 : node15541;
															assign node15541 = (inp[11]) ? node15543 : 16'b0000000000111111;
																assign node15543 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15547 = (inp[11]) ? node15557 : node15548;
													assign node15548 = (inp[9]) ? node15550 : 16'b0000000000111111;
														assign node15550 = (inp[10]) ? 16'b0000000000011111 : node15551;
															assign node15551 = (inp[3]) ? node15553 : 16'b0000000000111111;
																assign node15553 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15557 = (inp[9]) ? node15565 : node15558;
														assign node15558 = (inp[10]) ? node15560 : 16'b0000000000111111;
															assign node15560 = (inp[7]) ? 16'b0000000000011111 : node15561;
																assign node15561 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15565 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node15568 = (inp[7]) ? node15586 : node15569;
												assign node15569 = (inp[13]) ? node15581 : node15570;
													assign node15570 = (inp[11]) ? node15576 : node15571;
														assign node15571 = (inp[10]) ? node15573 : 16'b0000000001111111;
															assign node15573 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15576 = (inp[10]) ? 16'b0000000000011111 : node15577;
															assign node15577 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15581 = (inp[10]) ? node15583 : 16'b0000000000011111;
														assign node15583 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node15586 = (inp[13]) ? node15594 : node15587;
													assign node15587 = (inp[10]) ? node15589 : 16'b0000000000011111;
														assign node15589 = (inp[9]) ? 16'b0000000000001111 : node15590;
															assign node15590 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15594 = (inp[10]) ? node15596 : 16'b0000000000001111;
														assign node15596 = (inp[11]) ? 16'b0000000000000111 : node15597;
															assign node15597 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node15601 = (inp[10]) ? node16131 : node15602;
							assign node15602 = (inp[7]) ? node15870 : node15603;
								assign node15603 = (inp[5]) ? node15747 : node15604;
									assign node15604 = (inp[13]) ? node15686 : node15605;
										assign node15605 = (inp[2]) ? node15647 : node15606;
											assign node15606 = (inp[6]) ? node15630 : node15607;
												assign node15607 = (inp[14]) ? node15619 : node15608;
													assign node15608 = (inp[1]) ? node15612 : node15609;
														assign node15609 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15612 = (inp[9]) ? node15614 : 16'b0000001111111111;
															assign node15614 = (inp[3]) ? 16'b0000000111111111 : node15615;
																assign node15615 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15619 = (inp[3]) ? node15625 : node15620;
														assign node15620 = (inp[9]) ? node15622 : 16'b0000001111111111;
															assign node15622 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15625 = (inp[9]) ? node15627 : 16'b0000000111111111;
															assign node15627 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15630 = (inp[1]) ? node15640 : node15631;
													assign node15631 = (inp[14]) ? node15637 : node15632;
														assign node15632 = (inp[11]) ? node15634 : 16'b0000001111111111;
															assign node15634 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15637 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15640 = (inp[11]) ? node15644 : node15641;
														assign node15641 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15644 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node15647 = (inp[1]) ? node15667 : node15648;
												assign node15648 = (inp[11]) ? node15658 : node15649;
													assign node15649 = (inp[14]) ? node15651 : 16'b0000011111111111;
														assign node15651 = (inp[3]) ? node15655 : node15652;
															assign node15652 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node15655 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15658 = (inp[3]) ? 16'b0000000011111111 : node15659;
														assign node15659 = (inp[14]) ? node15661 : 16'b0000000111111111;
															assign node15661 = (inp[9]) ? 16'b0000000011111111 : node15662;
																assign node15662 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15667 = (inp[11]) ? node15679 : node15668;
													assign node15668 = (inp[3]) ? node15672 : node15669;
														assign node15669 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15672 = (inp[9]) ? 16'b0000000000111111 : node15673;
															assign node15673 = (inp[14]) ? node15675 : 16'b0000000011111111;
																assign node15675 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15679 = (inp[14]) ? node15681 : 16'b0000000001111111;
														assign node15681 = (inp[3]) ? node15683 : 16'b0000000001111111;
															assign node15683 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15686 = (inp[9]) ? node15720 : node15687;
											assign node15687 = (inp[6]) ? node15703 : node15688;
												assign node15688 = (inp[2]) ? node15694 : node15689;
													assign node15689 = (inp[11]) ? 16'b0000000111111111 : node15690;
														assign node15690 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15694 = (inp[14]) ? 16'b0000000011111111 : node15695;
														assign node15695 = (inp[3]) ? 16'b0000000011111111 : node15696;
															assign node15696 = (inp[11]) ? node15698 : 16'b0000000111111111;
																assign node15698 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15703 = (inp[11]) ? node15709 : node15704;
													assign node15704 = (inp[2]) ? node15706 : 16'b0000000111111111;
														assign node15706 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15709 = (inp[2]) ? node15715 : node15710;
														assign node15710 = (inp[14]) ? 16'b0000000001111111 : node15711;
															assign node15711 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15715 = (inp[14]) ? node15717 : 16'b0000000001111111;
															assign node15717 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15720 = (inp[14]) ? node15722 : 16'b0000000011111111;
												assign node15722 = (inp[2]) ? node15736 : node15723;
													assign node15723 = (inp[6]) ? 16'b0000000000111111 : node15724;
														assign node15724 = (inp[3]) ? node15730 : node15725;
															assign node15725 = (inp[1]) ? node15727 : 16'b0000000011111111;
																assign node15727 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node15730 = (inp[11]) ? node15732 : 16'b0000000001111111;
																assign node15732 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15736 = (inp[1]) ? node15740 : node15737;
														assign node15737 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15740 = (inp[3]) ? 16'b0000000000011111 : node15741;
															assign node15741 = (inp[6]) ? node15743 : 16'b0000000000111111;
																assign node15743 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node15747 = (inp[13]) ? node15817 : node15748;
										assign node15748 = (inp[14]) ? node15784 : node15749;
											assign node15749 = (inp[9]) ? node15765 : node15750;
												assign node15750 = (inp[3]) ? node15758 : node15751;
													assign node15751 = (inp[6]) ? node15753 : 16'b0000001111111111;
														assign node15753 = (inp[1]) ? node15755 : 16'b0000000111111111;
															assign node15755 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15758 = (inp[11]) ? 16'b0000000011111111 : node15759;
														assign node15759 = (inp[2]) ? node15761 : 16'b0000000011111111;
															assign node15761 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15765 = (inp[11]) ? node15771 : node15766;
													assign node15766 = (inp[6]) ? node15768 : 16'b0000000011111111;
														assign node15768 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node15771 = (inp[2]) ? node15779 : node15772;
														assign node15772 = (inp[1]) ? 16'b0000000001111111 : node15773;
															assign node15773 = (inp[3]) ? node15775 : 16'b0000000011111111;
																assign node15775 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15779 = (inp[6]) ? node15781 : 16'b0000000001111111;
															assign node15781 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15784 = (inp[3]) ? node15800 : node15785;
												assign node15785 = (inp[11]) ? node15793 : node15786;
													assign node15786 = (inp[2]) ? node15788 : 16'b0000000011111111;
														assign node15788 = (inp[9]) ? node15790 : 16'b0000000011111111;
															assign node15790 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15793 = (inp[1]) ? node15797 : node15794;
														assign node15794 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15797 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15800 = (inp[11]) ? node15812 : node15801;
													assign node15801 = (inp[9]) ? node15805 : node15802;
														assign node15802 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15805 = (inp[6]) ? node15807 : 16'b0000000001111111;
															assign node15807 = (inp[1]) ? 16'b0000000000111111 : node15808;
																assign node15808 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15812 = (inp[1]) ? node15814 : 16'b0000000001111111;
														assign node15814 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node15817 = (inp[2]) ? node15847 : node15818;
											assign node15818 = (inp[6]) ? node15832 : node15819;
												assign node15819 = (inp[3]) ? node15825 : node15820;
													assign node15820 = (inp[1]) ? node15822 : 16'b0000000111111111;
														assign node15822 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15825 = (inp[1]) ? node15827 : 16'b0000000001111111;
														assign node15827 = (inp[11]) ? node15829 : 16'b0000000001111111;
															assign node15829 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15832 = (inp[1]) ? node15838 : node15833;
													assign node15833 = (inp[14]) ? 16'b0000000001111111 : node15834;
														assign node15834 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15838 = (inp[11]) ? 16'b0000000000111111 : node15839;
														assign node15839 = (inp[9]) ? node15841 : 16'b0000000001111111;
															assign node15841 = (inp[3]) ? 16'b0000000000111111 : node15842;
																assign node15842 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15847 = (inp[9]) ? node15859 : node15848;
												assign node15848 = (inp[14]) ? node15854 : node15849;
													assign node15849 = (inp[3]) ? node15851 : 16'b0000000001111111;
														assign node15851 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15854 = (inp[6]) ? node15856 : 16'b0000000000111111;
														assign node15856 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15859 = (inp[6]) ? node15861 : 16'b0000000001111111;
													assign node15861 = (inp[11]) ? node15863 : 16'b0000000000011111;
														assign node15863 = (inp[3]) ? node15865 : 16'b0000000000011111;
															assign node15865 = (inp[14]) ? node15867 : 16'b0000000000001111;
																assign node15867 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node15870 = (inp[1]) ? node15978 : node15871;
									assign node15871 = (inp[2]) ? node15913 : node15872;
										assign node15872 = (inp[14]) ? node15890 : node15873;
											assign node15873 = (inp[5]) ? node15885 : node15874;
												assign node15874 = (inp[6]) ? node15880 : node15875;
													assign node15875 = (inp[11]) ? 16'b0000000111111111 : node15876;
														assign node15876 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15880 = (inp[9]) ? 16'b0000000011111111 : node15881;
														assign node15881 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15885 = (inp[6]) ? 16'b0000000001111111 : node15886;
													assign node15886 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15890 = (inp[11]) ? node15902 : node15891;
												assign node15891 = (inp[9]) ? node15893 : 16'b0000000011111111;
													assign node15893 = (inp[3]) ? node15899 : node15894;
														assign node15894 = (inp[13]) ? node15896 : 16'b0000000011111111;
															assign node15896 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15899 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15902 = (inp[6]) ? node15906 : node15903;
													assign node15903 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15906 = (inp[5]) ? 16'b0000000000111111 : node15907;
														assign node15907 = (inp[13]) ? node15909 : 16'b0000000001111111;
															assign node15909 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node15913 = (inp[14]) ? node15947 : node15914;
											assign node15914 = (inp[6]) ? node15928 : node15915;
												assign node15915 = (inp[9]) ? node15923 : node15916;
													assign node15916 = (inp[5]) ? 16'b0000000011111111 : node15917;
														assign node15917 = (inp[13]) ? node15919 : 16'b0000000111111111;
															assign node15919 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15923 = (inp[13]) ? node15925 : 16'b0000000011111111;
														assign node15925 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15928 = (inp[3]) ? node15940 : node15929;
													assign node15929 = (inp[5]) ? node15935 : node15930;
														assign node15930 = (inp[11]) ? node15932 : 16'b0000000011111111;
															assign node15932 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15935 = (inp[9]) ? node15937 : 16'b0000000001111111;
															assign node15937 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15940 = (inp[5]) ? node15944 : node15941;
														assign node15941 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15944 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node15947 = (inp[9]) ? node15959 : node15948;
												assign node15948 = (inp[3]) ? 16'b0000000000111111 : node15949;
													assign node15949 = (inp[5]) ? node15951 : 16'b0000000011111111;
														assign node15951 = (inp[13]) ? 16'b0000000000111111 : node15952;
															assign node15952 = (inp[11]) ? 16'b0000000000111111 : node15953;
																assign node15953 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node15959 = (inp[6]) ? node15969 : node15960;
													assign node15960 = (inp[11]) ? node15966 : node15961;
														assign node15961 = (inp[3]) ? 16'b0000000000111111 : node15962;
															assign node15962 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15966 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15969 = (inp[5]) ? node15973 : node15970;
														assign node15970 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15973 = (inp[11]) ? node15975 : 16'b0000000000011111;
															assign node15975 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node15978 = (inp[6]) ? node16046 : node15979;
										assign node15979 = (inp[14]) ? node16005 : node15980;
											assign node15980 = (inp[9]) ? node15992 : node15981;
												assign node15981 = (inp[2]) ? node15987 : node15982;
													assign node15982 = (inp[5]) ? node15984 : 16'b0000000011111111;
														assign node15984 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node15987 = (inp[11]) ? node15989 : 16'b0000000011111111;
														assign node15989 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15992 = (inp[3]) ? node16000 : node15993;
													assign node15993 = (inp[11]) ? node15997 : node15994;
														assign node15994 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15997 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16000 = (inp[2]) ? 16'b0000000000111111 : node16001;
														assign node16001 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16005 = (inp[5]) ? node16025 : node16006;
												assign node16006 = (inp[13]) ? node16016 : node16007;
													assign node16007 = (inp[11]) ? node16011 : node16008;
														assign node16008 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16011 = (inp[9]) ? node16013 : 16'b0000000001111111;
															assign node16013 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16016 = (inp[11]) ? node16018 : 16'b0000000001111111;
														assign node16018 = (inp[9]) ? node16020 : 16'b0000000000111111;
															assign node16020 = (inp[2]) ? 16'b0000000000001111 : node16021;
																assign node16021 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16025 = (inp[2]) ? node16033 : node16026;
													assign node16026 = (inp[11]) ? node16030 : node16027;
														assign node16027 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16030 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16033 = (inp[11]) ? node16041 : node16034;
														assign node16034 = (inp[9]) ? node16036 : 16'b0000000000111111;
															assign node16036 = (inp[13]) ? 16'b0000000000011111 : node16037;
																assign node16037 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16041 = (inp[3]) ? node16043 : 16'b0000000000011111;
															assign node16043 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node16046 = (inp[5]) ? node16092 : node16047;
											assign node16047 = (inp[13]) ? node16069 : node16048;
												assign node16048 = (inp[14]) ? node16060 : node16049;
													assign node16049 = (inp[11]) ? node16057 : node16050;
														assign node16050 = (inp[3]) ? 16'b0000000001111111 : node16051;
															assign node16051 = (inp[9]) ? node16053 : 16'b0000000011111111;
																assign node16053 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16057 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16060 = (inp[9]) ? node16064 : node16061;
														assign node16061 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16064 = (inp[3]) ? node16066 : 16'b0000000000111111;
															assign node16066 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16069 = (inp[14]) ? node16079 : node16070;
													assign node16070 = (inp[11]) ? node16074 : node16071;
														assign node16071 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node16074 = (inp[3]) ? 16'b0000000000011111 : node16075;
															assign node16075 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16079 = (inp[9]) ? node16085 : node16080;
														assign node16080 = (inp[3]) ? node16082 : 16'b0000000001111111;
															assign node16082 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16085 = (inp[3]) ? node16087 : 16'b0000000000001111;
															assign node16087 = (inp[2]) ? node16089 : 16'b0000000000001111;
																assign node16089 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node16092 = (inp[11]) ? node16106 : node16093;
												assign node16093 = (inp[14]) ? node16095 : 16'b0000000000111111;
													assign node16095 = (inp[2]) ? node16099 : node16096;
														assign node16096 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16099 = (inp[9]) ? node16101 : 16'b0000000000011111;
															assign node16101 = (inp[3]) ? node16103 : 16'b0000000000001111;
																assign node16103 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node16106 = (inp[13]) ? node16118 : node16107;
													assign node16107 = (inp[3]) ? node16109 : 16'b0000000000011111;
														assign node16109 = (inp[9]) ? node16115 : node16110;
															assign node16110 = (inp[14]) ? node16112 : 16'b0000000000011111;
																assign node16112 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node16115 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node16118 = (inp[2]) ? node16124 : node16119;
														assign node16119 = (inp[9]) ? 16'b0000000000001111 : node16120;
															assign node16120 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16124 = (inp[9]) ? 16'b0000000000000011 : node16125;
															assign node16125 = (inp[3]) ? node16127 : 16'b0000000000001111;
																assign node16127 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node16131 = (inp[3]) ? node16399 : node16132;
								assign node16132 = (inp[13]) ? node16250 : node16133;
									assign node16133 = (inp[11]) ? node16179 : node16134;
										assign node16134 = (inp[7]) ? node16154 : node16135;
											assign node16135 = (inp[1]) ? node16151 : node16136;
												assign node16136 = (inp[14]) ? node16146 : node16137;
													assign node16137 = (inp[5]) ? node16143 : node16138;
														assign node16138 = (inp[6]) ? 16'b0000000111111111 : node16139;
															assign node16139 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16143 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16146 = (inp[2]) ? 16'b0000000001111111 : node16147;
														assign node16147 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16151 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16154 = (inp[6]) ? node16164 : node16155;
												assign node16155 = (inp[1]) ? node16161 : node16156;
													assign node16156 = (inp[2]) ? node16158 : 16'b0000000111111111;
														assign node16158 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16161 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node16164 = (inp[2]) ? node16174 : node16165;
													assign node16165 = (inp[14]) ? node16171 : node16166;
														assign node16166 = (inp[9]) ? node16168 : 16'b0000000011111111;
															assign node16168 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16171 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16174 = (inp[9]) ? 16'b0000000000011111 : node16175;
														assign node16175 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node16179 = (inp[14]) ? node16201 : node16180;
											assign node16180 = (inp[6]) ? node16196 : node16181;
												assign node16181 = (inp[1]) ? node16189 : node16182;
													assign node16182 = (inp[9]) ? node16186 : node16183;
														assign node16183 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16186 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16189 = (inp[9]) ? node16191 : 16'b0000000001111111;
														assign node16191 = (inp[7]) ? 16'b0000000001111111 : node16192;
															assign node16192 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16196 = (inp[2]) ? node16198 : 16'b0000000001111111;
													assign node16198 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node16201 = (inp[5]) ? node16225 : node16202;
												assign node16202 = (inp[1]) ? node16214 : node16203;
													assign node16203 = (inp[2]) ? node16211 : node16204;
														assign node16204 = (inp[6]) ? node16206 : 16'b0000000011111111;
															assign node16206 = (inp[9]) ? 16'b0000000001111111 : node16207;
																assign node16207 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16211 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16214 = (inp[9]) ? node16222 : node16215;
														assign node16215 = (inp[7]) ? node16219 : node16216;
															assign node16216 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node16219 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16222 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16225 = (inp[2]) ? node16237 : node16226;
													assign node16226 = (inp[1]) ? node16232 : node16227;
														assign node16227 = (inp[9]) ? 16'b0000000000111111 : node16228;
															assign node16228 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16232 = (inp[6]) ? 16'b0000000000011111 : node16233;
															assign node16233 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16237 = (inp[9]) ? node16245 : node16238;
														assign node16238 = (inp[7]) ? 16'b0000000000011111 : node16239;
															assign node16239 = (inp[1]) ? node16241 : 16'b0000000000111111;
																assign node16241 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16245 = (inp[7]) ? 16'b0000000000001111 : node16246;
															assign node16246 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node16250 = (inp[7]) ? node16308 : node16251;
										assign node16251 = (inp[11]) ? node16277 : node16252;
											assign node16252 = (inp[2]) ? node16270 : node16253;
												assign node16253 = (inp[6]) ? node16259 : node16254;
													assign node16254 = (inp[14]) ? node16256 : 16'b0000000111111111;
														assign node16256 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16259 = (inp[9]) ? node16263 : node16260;
														assign node16260 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16263 = (inp[14]) ? node16265 : 16'b0000000001111111;
															assign node16265 = (inp[1]) ? 16'b0000000000111111 : node16266;
																assign node16266 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16270 = (inp[14]) ? node16272 : 16'b0000000001111111;
													assign node16272 = (inp[9]) ? node16274 : 16'b0000000001111111;
														assign node16274 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node16277 = (inp[9]) ? node16299 : node16278;
												assign node16278 = (inp[1]) ? node16290 : node16279;
													assign node16279 = (inp[2]) ? node16285 : node16280;
														assign node16280 = (inp[14]) ? 16'b0000000001111111 : node16281;
															assign node16281 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16285 = (inp[14]) ? node16287 : 16'b0000000001111111;
															assign node16287 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16290 = (inp[14]) ? node16296 : node16291;
														assign node16291 = (inp[6]) ? 16'b0000000000111111 : node16292;
															assign node16292 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16296 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16299 = (inp[1]) ? node16303 : node16300;
													assign node16300 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node16303 = (inp[5]) ? node16305 : 16'b0000000000011111;
														assign node16305 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node16308 = (inp[9]) ? node16348 : node16309;
											assign node16309 = (inp[6]) ? node16327 : node16310;
												assign node16310 = (inp[11]) ? node16314 : node16311;
													assign node16311 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16314 = (inp[5]) ? node16322 : node16315;
														assign node16315 = (inp[1]) ? node16317 : 16'b0000000001111111;
															assign node16317 = (inp[2]) ? 16'b0000000000111111 : node16318;
																assign node16318 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16322 = (inp[14]) ? 16'b0000000000111111 : node16323;
															assign node16323 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node16327 = (inp[14]) ? node16337 : node16328;
													assign node16328 = (inp[2]) ? node16332 : node16329;
														assign node16329 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16332 = (inp[11]) ? node16334 : 16'b0000000000111111;
															assign node16334 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16337 = (inp[1]) ? node16341 : node16338;
														assign node16338 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16341 = (inp[5]) ? 16'b0000000000001111 : node16342;
															assign node16342 = (inp[11]) ? node16344 : 16'b0000000000011111;
																assign node16344 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node16348 = (inp[5]) ? node16366 : node16349;
												assign node16349 = (inp[14]) ? 16'b0000000000011111 : node16350;
													assign node16350 = (inp[2]) ? node16352 : 16'b0000000001111111;
														assign node16352 = (inp[6]) ? node16358 : node16353;
															assign node16353 = (inp[11]) ? 16'b0000000000111111 : node16354;
																assign node16354 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node16358 = (inp[11]) ? node16362 : node16359;
																assign node16359 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
																assign node16362 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16366 = (inp[1]) ? node16388 : node16367;
													assign node16367 = (inp[11]) ? node16381 : node16368;
														assign node16368 = (inp[14]) ? node16374 : node16369;
															assign node16369 = (inp[2]) ? node16371 : 16'b0000000000111111;
																assign node16371 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node16374 = (inp[2]) ? node16378 : node16375;
																assign node16375 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
																assign node16378 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16381 = (inp[14]) ? node16383 : 16'b0000000000011111;
															assign node16383 = (inp[6]) ? 16'b0000000000001111 : node16384;
																assign node16384 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node16388 = (inp[14]) ? node16396 : node16389;
														assign node16389 = (inp[2]) ? 16'b0000000000001111 : node16390;
															assign node16390 = (inp[11]) ? node16392 : 16'b0000000000011111;
																assign node16392 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16396 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000000111;
								assign node16399 = (inp[7]) ? node16527 : node16400;
									assign node16400 = (inp[6]) ? node16468 : node16401;
										assign node16401 = (inp[11]) ? node16433 : node16402;
											assign node16402 = (inp[14]) ? node16416 : node16403;
												assign node16403 = (inp[13]) ? node16411 : node16404;
													assign node16404 = (inp[9]) ? node16408 : node16405;
														assign node16405 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node16408 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16411 = (inp[1]) ? 16'b0000000001111111 : node16412;
														assign node16412 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16416 = (inp[1]) ? node16428 : node16417;
													assign node16417 = (inp[9]) ? node16419 : 16'b0000000001111111;
														assign node16419 = (inp[13]) ? node16425 : node16420;
															assign node16420 = (inp[5]) ? node16422 : 16'b0000000001111111;
																assign node16422 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node16425 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16428 = (inp[9]) ? node16430 : 16'b0000000000111111;
														assign node16430 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node16433 = (inp[13]) ? node16451 : node16434;
												assign node16434 = (inp[1]) ? node16440 : node16435;
													assign node16435 = (inp[14]) ? node16437 : 16'b0000000011111111;
														assign node16437 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16440 = (inp[14]) ? node16444 : node16441;
														assign node16441 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16444 = (inp[5]) ? node16446 : 16'b0000000000111111;
															assign node16446 = (inp[9]) ? 16'b0000000000011111 : node16447;
																assign node16447 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16451 = (inp[9]) ? node16461 : node16452;
													assign node16452 = (inp[1]) ? node16456 : node16453;
														assign node16453 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16456 = (inp[5]) ? 16'b0000000000011111 : node16457;
															assign node16457 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16461 = (inp[1]) ? node16463 : 16'b0000000000011111;
														assign node16463 = (inp[5]) ? 16'b0000000000001111 : node16464;
															assign node16464 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node16468 = (inp[2]) ? node16488 : node16469;
											assign node16469 = (inp[14]) ? node16477 : node16470;
												assign node16470 = (inp[1]) ? 16'b0000000000111111 : node16471;
													assign node16471 = (inp[9]) ? node16473 : 16'b0000000001111111;
														assign node16473 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16477 = (inp[1]) ? node16483 : node16478;
													assign node16478 = (inp[9]) ? node16480 : 16'b0000000000111111;
														assign node16480 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16483 = (inp[13]) ? node16485 : 16'b0000000000111111;
														assign node16485 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node16488 = (inp[5]) ? node16506 : node16489;
												assign node16489 = (inp[1]) ? node16495 : node16490;
													assign node16490 = (inp[9]) ? node16492 : 16'b0000000001111111;
														assign node16492 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16495 = (inp[13]) ? node16501 : node16496;
														assign node16496 = (inp[9]) ? node16498 : 16'b0000000000111111;
															assign node16498 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16501 = (inp[11]) ? node16503 : 16'b0000000000011111;
															assign node16503 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16506 = (inp[14]) ? node16518 : node16507;
													assign node16507 = (inp[11]) ? node16513 : node16508;
														assign node16508 = (inp[1]) ? 16'b0000000000011111 : node16509;
															assign node16509 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16513 = (inp[9]) ? node16515 : 16'b0000000000011111;
															assign node16515 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node16518 = (inp[13]) ? node16522 : node16519;
														assign node16519 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16522 = (inp[1]) ? node16524 : 16'b0000000000001111;
															assign node16524 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node16527 = (inp[14]) ? node16589 : node16528;
										assign node16528 = (inp[11]) ? node16558 : node16529;
											assign node16529 = (inp[9]) ? node16541 : node16530;
												assign node16530 = (inp[6]) ? node16532 : 16'b0000000001111111;
													assign node16532 = (inp[1]) ? node16538 : node16533;
														assign node16533 = (inp[5]) ? 16'b0000000000111111 : node16534;
															assign node16534 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16538 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node16541 = (inp[5]) ? node16553 : node16542;
													assign node16542 = (inp[1]) ? node16546 : node16543;
														assign node16543 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16546 = (inp[2]) ? 16'b0000000000011111 : node16547;
															assign node16547 = (inp[6]) ? node16549 : 16'b0000000000111111;
																assign node16549 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16553 = (inp[2]) ? node16555 : 16'b0000000000011111;
														assign node16555 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node16558 = (inp[1]) ? node16574 : node16559;
												assign node16559 = (inp[6]) ? node16567 : node16560;
													assign node16560 = (inp[5]) ? node16562 : 16'b0000000001111111;
														assign node16562 = (inp[9]) ? 16'b0000000000011111 : node16563;
															assign node16563 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16567 = (inp[9]) ? node16571 : node16568;
														assign node16568 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16571 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16574 = (inp[13]) ? node16580 : node16575;
													assign node16575 = (inp[5]) ? node16577 : 16'b0000000000011111;
														assign node16577 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node16580 = (inp[9]) ? node16584 : node16581;
														assign node16581 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16584 = (inp[6]) ? 16'b0000000000000111 : node16585;
															assign node16585 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node16589 = (inp[11]) ? node16621 : node16590;
											assign node16590 = (inp[5]) ? node16606 : node16591;
												assign node16591 = (inp[2]) ? node16597 : node16592;
													assign node16592 = (inp[13]) ? node16594 : 16'b0000000001111111;
														assign node16594 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node16597 = (inp[9]) ? node16601 : node16598;
														assign node16598 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node16601 = (inp[13]) ? node16603 : 16'b0000000000011111;
															assign node16603 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node16606 = (inp[9]) ? node16614 : node16607;
													assign node16607 = (inp[2]) ? node16609 : 16'b0000000000111111;
														assign node16609 = (inp[1]) ? node16611 : 16'b0000000000011111;
															assign node16611 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node16614 = (inp[1]) ? node16618 : node16615;
														assign node16615 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node16618 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node16621 = (inp[2]) ? node16631 : node16622;
												assign node16622 = (inp[6]) ? node16628 : node16623;
													assign node16623 = (inp[9]) ? node16625 : 16'b0000000000011111;
														assign node16625 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node16628 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000000111;
												assign node16631 = (inp[1]) ? node16639 : node16632;
													assign node16632 = (inp[6]) ? 16'b0000000000000111 : node16633;
														assign node16633 = (inp[9]) ? node16635 : 16'b0000000000001111;
															assign node16635 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node16639 = (inp[6]) ? 16'b0000000000000001 : 16'b0000000000000011;
		assign node16642 = (inp[3]) ? node24980 : node16643;
			assign node16643 = (inp[6]) ? node20771 : node16644;
				assign node16644 = (inp[1]) ? node18706 : node16645;
					assign node16645 = (inp[15]) ? node17773 : node16646;
						assign node16646 = (inp[12]) ? node17220 : node16647;
							assign node16647 = (inp[5]) ? node16933 : node16648;
								assign node16648 = (inp[8]) ? node16802 : node16649;
									assign node16649 = (inp[4]) ? node16727 : node16650;
										assign node16650 = (inp[11]) ? node16686 : node16651;
											assign node16651 = (inp[9]) ? node16671 : node16652;
												assign node16652 = (inp[13]) ? node16658 : node16653;
													assign node16653 = (inp[10]) ? 16'b0011111111111111 : node16654;
														assign node16654 = (inp[14]) ? 16'b0011111111111111 : 16'b0111111111111111;
													assign node16658 = (inp[2]) ? 16'b0000111111111111 : node16659;
														assign node16659 = (inp[7]) ? node16665 : node16660;
															assign node16660 = (inp[14]) ? 16'b0001111111111111 : node16661;
																assign node16661 = (inp[10]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node16665 = (inp[14]) ? 16'b0000111111111111 : node16666;
																assign node16666 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node16671 = (inp[13]) ? node16681 : node16672;
													assign node16672 = (inp[14]) ? 16'b0000111111111111 : node16673;
														assign node16673 = (inp[2]) ? node16675 : 16'b0011111111111111;
															assign node16675 = (inp[7]) ? 16'b0000111111111111 : node16676;
																assign node16676 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node16681 = (inp[14]) ? 16'b0000011111111111 : node16682;
														assign node16682 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node16686 = (inp[14]) ? node16708 : node16687;
												assign node16687 = (inp[2]) ? node16697 : node16688;
													assign node16688 = (inp[9]) ? node16694 : node16689;
														assign node16689 = (inp[7]) ? 16'b0000111111111111 : node16690;
															assign node16690 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node16694 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16697 = (inp[10]) ? node16705 : node16698;
														assign node16698 = (inp[9]) ? node16702 : node16699;
															assign node16699 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node16702 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16705 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16708 = (inp[10]) ? node16720 : node16709;
													assign node16709 = (inp[7]) ? node16715 : node16710;
														assign node16710 = (inp[13]) ? node16712 : 16'b0000111111111111;
															assign node16712 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16715 = (inp[13]) ? node16717 : 16'b0000011111111111;
															assign node16717 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16720 = (inp[2]) ? 16'b0000001111111111 : node16721;
														assign node16721 = (inp[9]) ? 16'b0000001111111111 : node16722;
															assign node16722 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node16727 = (inp[10]) ? node16765 : node16728;
											assign node16728 = (inp[7]) ? node16746 : node16729;
												assign node16729 = (inp[2]) ? node16741 : node16730;
													assign node16730 = (inp[9]) ? node16738 : node16731;
														assign node16731 = (inp[13]) ? 16'b0000111111111111 : node16732;
															assign node16732 = (inp[11]) ? 16'b0001111111111111 : node16733;
																assign node16733 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node16738 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16741 = (inp[13]) ? 16'b0000011111111111 : node16742;
														assign node16742 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node16746 = (inp[11]) ? node16758 : node16747;
													assign node16747 = (inp[2]) ? node16755 : node16748;
														assign node16748 = (inp[13]) ? node16750 : 16'b0000111111111111;
															assign node16750 = (inp[9]) ? 16'b0000011111111111 : node16751;
																assign node16751 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16755 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16758 = (inp[9]) ? node16762 : node16759;
														assign node16759 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16762 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node16765 = (inp[14]) ? node16787 : node16766;
												assign node16766 = (inp[11]) ? node16780 : node16767;
													assign node16767 = (inp[13]) ? node16775 : node16768;
														assign node16768 = (inp[9]) ? node16770 : 16'b0001111111111111;
															assign node16770 = (inp[2]) ? 16'b0000011111111111 : node16771;
																assign node16771 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16775 = (inp[7]) ? node16777 : 16'b0000011111111111;
															assign node16777 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16780 = (inp[7]) ? node16784 : node16781;
														assign node16781 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16784 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16787 = (inp[13]) ? node16793 : node16788;
													assign node16788 = (inp[2]) ? node16790 : 16'b0000011111111111;
														assign node16790 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16793 = (inp[7]) ? node16797 : node16794;
														assign node16794 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node16797 = (inp[2]) ? node16799 : 16'b0000000111111111;
															assign node16799 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node16802 = (inp[13]) ? node16872 : node16803;
										assign node16803 = (inp[2]) ? node16833 : node16804;
											assign node16804 = (inp[7]) ? node16824 : node16805;
												assign node16805 = (inp[11]) ? node16813 : node16806;
													assign node16806 = (inp[4]) ? node16810 : node16807;
														assign node16807 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node16810 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16813 = (inp[14]) ? node16821 : node16814;
														assign node16814 = (inp[9]) ? 16'b0000011111111111 : node16815;
															assign node16815 = (inp[10]) ? node16817 : 16'b0000111111111111;
																assign node16817 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16821 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16824 = (inp[14]) ? node16828 : node16825;
													assign node16825 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16828 = (inp[10]) ? node16830 : 16'b0000011111111111;
														assign node16830 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node16833 = (inp[10]) ? node16857 : node16834;
												assign node16834 = (inp[11]) ? node16848 : node16835;
													assign node16835 = (inp[14]) ? node16843 : node16836;
														assign node16836 = (inp[9]) ? node16840 : node16837;
															assign node16837 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node16840 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16843 = (inp[9]) ? node16845 : 16'b0000011111111111;
															assign node16845 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16848 = (inp[4]) ? node16854 : node16849;
														assign node16849 = (inp[9]) ? 16'b0000001111111111 : node16850;
															assign node16850 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16854 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16857 = (inp[4]) ? node16863 : node16858;
													assign node16858 = (inp[7]) ? node16860 : 16'b0000001111111111;
														assign node16860 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16863 = (inp[11]) ? node16869 : node16864;
														assign node16864 = (inp[14]) ? 16'b0000000111111111 : node16865;
															assign node16865 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16869 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node16872 = (inp[9]) ? node16910 : node16873;
											assign node16873 = (inp[10]) ? node16889 : node16874;
												assign node16874 = (inp[2]) ? 16'b0000001111111111 : node16875;
													assign node16875 = (inp[14]) ? node16881 : node16876;
														assign node16876 = (inp[7]) ? node16878 : 16'b0001111111111111;
															assign node16878 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16881 = (inp[7]) ? 16'b0000001111111111 : node16882;
															assign node16882 = (inp[4]) ? 16'b0000011111111111 : node16883;
																assign node16883 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node16889 = (inp[4]) ? node16895 : node16890;
													assign node16890 = (inp[11]) ? 16'b0000001111111111 : node16891;
														assign node16891 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16895 = (inp[2]) ? node16903 : node16896;
														assign node16896 = (inp[14]) ? 16'b0000000111111111 : node16897;
															assign node16897 = (inp[11]) ? 16'b0000001111111111 : node16898;
																assign node16898 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16903 = (inp[7]) ? 16'b0000000011111111 : node16904;
															assign node16904 = (inp[11]) ? node16906 : 16'b0000000111111111;
																assign node16906 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16910 = (inp[7]) ? node16922 : node16911;
												assign node16911 = (inp[10]) ? node16919 : node16912;
													assign node16912 = (inp[14]) ? node16914 : 16'b0000011111111111;
														assign node16914 = (inp[2]) ? node16916 : 16'b0000001111111111;
															assign node16916 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16919 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node16922 = (inp[11]) ? node16926 : node16923;
													assign node16923 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16926 = (inp[4]) ? node16928 : 16'b0000000011111111;
														assign node16928 = (inp[10]) ? node16930 : 16'b0000000001111111;
															assign node16930 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node16933 = (inp[7]) ? node17087 : node16934;
									assign node16934 = (inp[9]) ? node17008 : node16935;
										assign node16935 = (inp[14]) ? node16977 : node16936;
											assign node16936 = (inp[8]) ? node16960 : node16937;
												assign node16937 = (inp[4]) ? node16945 : node16938;
													assign node16938 = (inp[11]) ? node16940 : 16'b0001111111111111;
														assign node16940 = (inp[2]) ? 16'b0000011111111111 : node16941;
															assign node16941 = (inp[13]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node16945 = (inp[13]) ? node16955 : node16946;
														assign node16946 = (inp[10]) ? node16952 : node16947;
															assign node16947 = (inp[11]) ? 16'b0000111111111111 : node16948;
																assign node16948 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node16952 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16955 = (inp[2]) ? node16957 : 16'b0000011111111111;
															assign node16957 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16960 = (inp[11]) ? node16972 : node16961;
													assign node16961 = (inp[10]) ? node16969 : node16962;
														assign node16962 = (inp[4]) ? node16964 : 16'b0000111111111111;
															assign node16964 = (inp[2]) ? 16'b0000001111111111 : node16965;
																assign node16965 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16969 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16972 = (inp[13]) ? node16974 : 16'b0000001111111111;
														assign node16974 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node16977 = (inp[10]) ? node16995 : node16978;
												assign node16978 = (inp[11]) ? node16986 : node16979;
													assign node16979 = (inp[8]) ? node16983 : node16980;
														assign node16980 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node16983 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16986 = (inp[4]) ? node16990 : node16987;
														assign node16987 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16990 = (inp[2]) ? 16'b0000001111111111 : node16991;
															assign node16991 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16995 = (inp[13]) ? node17003 : node16996;
													assign node16996 = (inp[11]) ? 16'b0000000111111111 : node16997;
														assign node16997 = (inp[2]) ? node16999 : 16'b0000011111111111;
															assign node16999 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node17003 = (inp[11]) ? node17005 : 16'b0000000111111111;
														assign node17005 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17008 = (inp[13]) ? node17048 : node17009;
											assign node17009 = (inp[11]) ? node17033 : node17010;
												assign node17010 = (inp[2]) ? node17020 : node17011;
													assign node17011 = (inp[14]) ? 16'b0000011111111111 : node17012;
														assign node17012 = (inp[8]) ? node17014 : 16'b0000111111111111;
															assign node17014 = (inp[10]) ? 16'b0000011111111111 : node17015;
																assign node17015 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node17020 = (inp[4]) ? node17028 : node17021;
														assign node17021 = (inp[8]) ? node17023 : 16'b0000011111111111;
															assign node17023 = (inp[10]) ? 16'b0000001111111111 : node17024;
																assign node17024 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17028 = (inp[10]) ? node17030 : 16'b0000001111111111;
															assign node17030 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17033 = (inp[8]) ? node17043 : node17034;
													assign node17034 = (inp[14]) ? node17038 : node17035;
														assign node17035 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node17038 = (inp[4]) ? node17040 : 16'b0000001111111111;
															assign node17040 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17043 = (inp[10]) ? 16'b0000000111111111 : node17044;
														assign node17044 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17048 = (inp[8]) ? node17072 : node17049;
												assign node17049 = (inp[10]) ? node17057 : node17050;
													assign node17050 = (inp[11]) ? node17054 : node17051;
														assign node17051 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17054 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17057 = (inp[4]) ? node17065 : node17058;
														assign node17058 = (inp[11]) ? node17062 : node17059;
															assign node17059 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node17062 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17065 = (inp[2]) ? node17067 : 16'b0000000111111111;
															assign node17067 = (inp[11]) ? 16'b0000000011111111 : node17068;
																assign node17068 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17072 = (inp[10]) ? node17080 : node17073;
													assign node17073 = (inp[11]) ? node17075 : 16'b0000001111111111;
														assign node17075 = (inp[4]) ? 16'b0000000011111111 : node17076;
															assign node17076 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17080 = (inp[11]) ? 16'b0000000001111111 : node17081;
														assign node17081 = (inp[4]) ? node17083 : 16'b0000000111111111;
															assign node17083 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node17087 = (inp[13]) ? node17157 : node17088;
										assign node17088 = (inp[2]) ? node17118 : node17089;
											assign node17089 = (inp[11]) ? node17103 : node17090;
												assign node17090 = (inp[4]) ? node17100 : node17091;
													assign node17091 = (inp[10]) ? node17097 : node17092;
														assign node17092 = (inp[8]) ? node17094 : 16'b0000111111111111;
															assign node17094 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17097 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17100 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17103 = (inp[10]) ? node17111 : node17104;
													assign node17104 = (inp[8]) ? 16'b0000001111111111 : node17105;
														assign node17105 = (inp[14]) ? 16'b0000001111111111 : node17106;
															assign node17106 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node17111 = (inp[9]) ? 16'b0000000111111111 : node17112;
														assign node17112 = (inp[8]) ? node17114 : 16'b0000001111111111;
															assign node17114 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17118 = (inp[11]) ? node17134 : node17119;
												assign node17119 = (inp[4]) ? node17127 : node17120;
													assign node17120 = (inp[8]) ? node17122 : 16'b0000001111111111;
														assign node17122 = (inp[9]) ? node17124 : 16'b0000001111111111;
															assign node17124 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17127 = (inp[9]) ? node17131 : node17128;
														assign node17128 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17131 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17134 = (inp[9]) ? node17146 : node17135;
													assign node17135 = (inp[10]) ? node17141 : node17136;
														assign node17136 = (inp[14]) ? node17138 : 16'b0000001111111111;
															assign node17138 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17141 = (inp[14]) ? node17143 : 16'b0000000111111111;
															assign node17143 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17146 = (inp[4]) ? node17154 : node17147;
														assign node17147 = (inp[14]) ? node17149 : 16'b0000000111111111;
															assign node17149 = (inp[8]) ? 16'b0000000011111111 : node17150;
																assign node17150 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17154 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17157 = (inp[14]) ? node17187 : node17158;
											assign node17158 = (inp[8]) ? node17178 : node17159;
												assign node17159 = (inp[9]) ? node17173 : node17160;
													assign node17160 = (inp[4]) ? node17166 : node17161;
														assign node17161 = (inp[2]) ? node17163 : 16'b0000011111111111;
															assign node17163 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17166 = (inp[2]) ? node17168 : 16'b0000001111111111;
															assign node17168 = (inp[10]) ? 16'b0000000111111111 : node17169;
																assign node17169 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17173 = (inp[11]) ? 16'b0000000011111111 : node17174;
														assign node17174 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17178 = (inp[11]) ? node17180 : 16'b0000000111111111;
													assign node17180 = (inp[2]) ? node17184 : node17181;
														assign node17181 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17184 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node17187 = (inp[10]) ? node17203 : node17188;
												assign node17188 = (inp[8]) ? node17198 : node17189;
													assign node17189 = (inp[11]) ? node17195 : node17190;
														assign node17190 = (inp[2]) ? node17192 : 16'b0000001111111111;
															assign node17192 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17195 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17198 = (inp[4]) ? node17200 : 16'b0000000011111111;
														assign node17200 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node17203 = (inp[4]) ? node17211 : node17204;
													assign node17204 = (inp[11]) ? node17208 : node17205;
														assign node17205 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17208 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17211 = (inp[2]) ? node17215 : node17212;
														assign node17212 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17215 = (inp[8]) ? 16'b0000000000111111 : node17216;
															assign node17216 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node17220 = (inp[2]) ? node17536 : node17221;
								assign node17221 = (inp[8]) ? node17381 : node17222;
									assign node17222 = (inp[11]) ? node17308 : node17223;
										assign node17223 = (inp[5]) ? node17263 : node17224;
											assign node17224 = (inp[10]) ? node17240 : node17225;
												assign node17225 = (inp[7]) ? node17233 : node17226;
													assign node17226 = (inp[14]) ? node17228 : 16'b0001111111111111;
														assign node17228 = (inp[9]) ? node17230 : 16'b0000111111111111;
															assign node17230 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node17233 = (inp[9]) ? node17237 : node17234;
														assign node17234 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17237 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node17240 = (inp[7]) ? node17256 : node17241;
													assign node17241 = (inp[13]) ? node17249 : node17242;
														assign node17242 = (inp[4]) ? node17244 : 16'b0000111111111111;
															assign node17244 = (inp[9]) ? 16'b0000011111111111 : node17245;
																assign node17245 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17249 = (inp[9]) ? node17251 : 16'b0000011111111111;
															assign node17251 = (inp[4]) ? 16'b0000001111111111 : node17252;
																assign node17252 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17256 = (inp[4]) ? node17260 : node17257;
														assign node17257 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17260 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17263 = (inp[14]) ? node17289 : node17264;
												assign node17264 = (inp[7]) ? node17274 : node17265;
													assign node17265 = (inp[13]) ? node17271 : node17266;
														assign node17266 = (inp[9]) ? 16'b0000111111111111 : node17267;
															assign node17267 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node17271 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17274 = (inp[9]) ? node17282 : node17275;
														assign node17275 = (inp[10]) ? 16'b0000001111111111 : node17276;
															assign node17276 = (inp[4]) ? node17278 : 16'b0000011111111111;
																assign node17278 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17282 = (inp[13]) ? node17284 : 16'b0000001111111111;
															assign node17284 = (inp[10]) ? node17286 : 16'b0000000111111111;
																assign node17286 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17289 = (inp[13]) ? node17299 : node17290;
													assign node17290 = (inp[4]) ? node17294 : node17291;
														assign node17291 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17294 = (inp[10]) ? 16'b0000000111111111 : node17295;
															assign node17295 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17299 = (inp[9]) ? node17303 : node17300;
														assign node17300 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17303 = (inp[4]) ? 16'b0000000011111111 : node17304;
															assign node17304 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17308 = (inp[7]) ? node17346 : node17309;
											assign node17309 = (inp[5]) ? node17331 : node17310;
												assign node17310 = (inp[4]) ? node17318 : node17311;
													assign node17311 = (inp[9]) ? node17315 : node17312;
														assign node17312 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17315 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17318 = (inp[9]) ? node17324 : node17319;
														assign node17319 = (inp[14]) ? 16'b0000001111111111 : node17320;
															assign node17320 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17324 = (inp[14]) ? 16'b0000000111111111 : node17325;
															assign node17325 = (inp[10]) ? node17327 : 16'b0000001111111111;
																assign node17327 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17331 = (inp[4]) ? node17339 : node17332;
													assign node17332 = (inp[14]) ? node17334 : 16'b0000001111111111;
														assign node17334 = (inp[13]) ? node17336 : 16'b0000001111111111;
															assign node17336 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17339 = (inp[13]) ? 16'b0000000011111111 : node17340;
														assign node17340 = (inp[10]) ? 16'b0000000111111111 : node17341;
															assign node17341 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node17346 = (inp[9]) ? node17366 : node17347;
												assign node17347 = (inp[5]) ? node17357 : node17348;
													assign node17348 = (inp[14]) ? node17354 : node17349;
														assign node17349 = (inp[13]) ? 16'b0000001111111111 : node17350;
															assign node17350 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17354 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17357 = (inp[14]) ? 16'b0000000111111111 : node17358;
														assign node17358 = (inp[13]) ? node17360 : 16'b0000001111111111;
															assign node17360 = (inp[4]) ? 16'b0000000111111111 : node17361;
																assign node17361 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17366 = (inp[5]) ? node17376 : node17367;
													assign node17367 = (inp[14]) ? node17373 : node17368;
														assign node17368 = (inp[10]) ? 16'b0000000111111111 : node17369;
															assign node17369 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17373 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node17376 = (inp[13]) ? 16'b0000000001111111 : node17377;
														assign node17377 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node17381 = (inp[13]) ? node17463 : node17382;
										assign node17382 = (inp[7]) ? node17430 : node17383;
											assign node17383 = (inp[11]) ? node17405 : node17384;
												assign node17384 = (inp[9]) ? node17400 : node17385;
													assign node17385 = (inp[4]) ? node17395 : node17386;
														assign node17386 = (inp[14]) ? node17392 : node17387;
															assign node17387 = (inp[10]) ? 16'b0000111111111111 : node17388;
																assign node17388 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
															assign node17392 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17395 = (inp[5]) ? node17397 : 16'b0000011111111111;
															assign node17397 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17400 = (inp[5]) ? 16'b0000001111111111 : node17401;
														assign node17401 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node17405 = (inp[14]) ? node17415 : node17406;
													assign node17406 = (inp[5]) ? 16'b0000000111111111 : node17407;
														assign node17407 = (inp[4]) ? node17411 : node17408;
															assign node17408 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node17411 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17415 = (inp[4]) ? node17423 : node17416;
														assign node17416 = (inp[5]) ? 16'b0000000111111111 : node17417;
															assign node17417 = (inp[9]) ? node17419 : 16'b0000001111111111;
																assign node17419 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17423 = (inp[9]) ? 16'b0000000011111111 : node17424;
															assign node17424 = (inp[5]) ? node17426 : 16'b0000000111111111;
																assign node17426 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17430 = (inp[5]) ? node17446 : node17431;
												assign node17431 = (inp[9]) ? node17437 : node17432;
													assign node17432 = (inp[4]) ? 16'b0000001111111111 : node17433;
														assign node17433 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17437 = (inp[14]) ? node17441 : node17438;
														assign node17438 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17441 = (inp[11]) ? node17443 : 16'b0000000111111111;
															assign node17443 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17446 = (inp[10]) ? node17458 : node17447;
													assign node17447 = (inp[14]) ? node17451 : node17448;
														assign node17448 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17451 = (inp[11]) ? 16'b0000000111111111 : node17452;
															assign node17452 = (inp[9]) ? 16'b0000000111111111 : node17453;
																assign node17453 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17458 = (inp[14]) ? 16'b0000000011111111 : node17459;
														assign node17459 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17463 = (inp[14]) ? node17497 : node17464;
											assign node17464 = (inp[9]) ? node17478 : node17465;
												assign node17465 = (inp[7]) ? node17473 : node17466;
													assign node17466 = (inp[4]) ? node17468 : 16'b0000011111111111;
														assign node17468 = (inp[11]) ? node17470 : 16'b0000001111111111;
															assign node17470 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17473 = (inp[11]) ? 16'b0000000111111111 : node17474;
														assign node17474 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17478 = (inp[4]) ? node17486 : node17479;
													assign node17479 = (inp[7]) ? node17481 : 16'b0000000111111111;
														assign node17481 = (inp[11]) ? node17483 : 16'b0000000111111111;
															assign node17483 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17486 = (inp[11]) ? node17492 : node17487;
														assign node17487 = (inp[10]) ? node17489 : 16'b0000000111111111;
															assign node17489 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17492 = (inp[10]) ? 16'b0000000011111111 : node17493;
															assign node17493 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17497 = (inp[9]) ? node17519 : node17498;
												assign node17498 = (inp[4]) ? node17508 : node17499;
													assign node17499 = (inp[5]) ? node17505 : node17500;
														assign node17500 = (inp[7]) ? node17502 : 16'b0000001111111111;
															assign node17502 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17505 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node17508 = (inp[7]) ? node17516 : node17509;
														assign node17509 = (inp[11]) ? node17511 : 16'b0000000111111111;
															assign node17511 = (inp[10]) ? 16'b0000000011111111 : node17512;
																assign node17512 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17516 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17519 = (inp[4]) ? node17529 : node17520;
													assign node17520 = (inp[5]) ? node17526 : node17521;
														assign node17521 = (inp[10]) ? 16'b0000000011111111 : node17522;
															assign node17522 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17526 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17529 = (inp[11]) ? node17533 : node17530;
														assign node17530 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17533 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node17536 = (inp[10]) ? node17650 : node17537;
									assign node17537 = (inp[5]) ? node17591 : node17538;
										assign node17538 = (inp[8]) ? node17568 : node17539;
											assign node17539 = (inp[14]) ? node17555 : node17540;
												assign node17540 = (inp[11]) ? node17548 : node17541;
													assign node17541 = (inp[4]) ? node17545 : node17542;
														assign node17542 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17545 = (inp[13]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node17548 = (inp[7]) ? 16'b0000001111111111 : node17549;
														assign node17549 = (inp[13]) ? node17551 : 16'b0000011111111111;
															assign node17551 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17555 = (inp[9]) ? node17563 : node17556;
													assign node17556 = (inp[11]) ? node17560 : node17557;
														assign node17557 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17560 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17563 = (inp[7]) ? 16'b0000000111111111 : node17564;
														assign node17564 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17568 = (inp[4]) ? node17578 : node17569;
												assign node17569 = (inp[7]) ? node17575 : node17570;
													assign node17570 = (inp[14]) ? 16'b0000000111111111 : node17571;
														assign node17571 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17575 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node17578 = (inp[11]) ? node17584 : node17579;
													assign node17579 = (inp[14]) ? node17581 : 16'b0000001111111111;
														assign node17581 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17584 = (inp[14]) ? 16'b0000000011111111 : node17585;
														assign node17585 = (inp[13]) ? 16'b0000000011111111 : node17586;
															assign node17586 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17591 = (inp[9]) ? node17619 : node17592;
											assign node17592 = (inp[8]) ? node17610 : node17593;
												assign node17593 = (inp[13]) ? node17605 : node17594;
													assign node17594 = (inp[11]) ? node17598 : node17595;
														assign node17595 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17598 = (inp[7]) ? node17600 : 16'b0000001111111111;
															assign node17600 = (inp[4]) ? 16'b0000000111111111 : node17601;
																assign node17601 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17605 = (inp[7]) ? 16'b0000000111111111 : node17606;
														assign node17606 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17610 = (inp[13]) ? node17612 : 16'b0000000111111111;
													assign node17612 = (inp[11]) ? node17616 : node17613;
														assign node17613 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node17616 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17619 = (inp[11]) ? node17641 : node17620;
												assign node17620 = (inp[14]) ? node17634 : node17621;
													assign node17621 = (inp[7]) ? node17627 : node17622;
														assign node17622 = (inp[13]) ? 16'b0000000111111111 : node17623;
															assign node17623 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17627 = (inp[13]) ? 16'b0000000011111111 : node17628;
															assign node17628 = (inp[8]) ? node17630 : 16'b0000000111111111;
																assign node17630 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17634 = (inp[13]) ? node17638 : node17635;
														assign node17635 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17638 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17641 = (inp[8]) ? 16'b0000000001111111 : node17642;
													assign node17642 = (inp[7]) ? node17644 : 16'b0000000011111111;
														assign node17644 = (inp[13]) ? 16'b0000000001111111 : node17645;
															assign node17645 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node17650 = (inp[9]) ? node17708 : node17651;
										assign node17651 = (inp[8]) ? node17681 : node17652;
											assign node17652 = (inp[4]) ? node17666 : node17653;
												assign node17653 = (inp[14]) ? node17659 : node17654;
													assign node17654 = (inp[11]) ? 16'b0000001111111111 : node17655;
														assign node17655 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node17659 = (inp[7]) ? 16'b0000000111111111 : node17660;
														assign node17660 = (inp[11]) ? node17662 : 16'b0000001111111111;
															assign node17662 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17666 = (inp[14]) ? node17676 : node17667;
													assign node17667 = (inp[13]) ? 16'b0000000111111111 : node17668;
														assign node17668 = (inp[7]) ? node17670 : 16'b0000001111111111;
															assign node17670 = (inp[5]) ? 16'b0000000111111111 : node17671;
																assign node17671 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17676 = (inp[13]) ? 16'b0000000011111111 : node17677;
														assign node17677 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17681 = (inp[14]) ? node17697 : node17682;
												assign node17682 = (inp[13]) ? node17690 : node17683;
													assign node17683 = (inp[11]) ? node17687 : node17684;
														assign node17684 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17687 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node17690 = (inp[7]) ? 16'b0000000000111111 : node17691;
														assign node17691 = (inp[5]) ? node17693 : 16'b0000000011111111;
															assign node17693 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17697 = (inp[11]) ? 16'b0000000001111111 : node17698;
													assign node17698 = (inp[4]) ? node17700 : 16'b0000000011111111;
														assign node17700 = (inp[5]) ? 16'b0000000001111111 : node17701;
															assign node17701 = (inp[7]) ? node17703 : 16'b0000000011111111;
																assign node17703 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17708 = (inp[7]) ? node17740 : node17709;
											assign node17709 = (inp[14]) ? node17725 : node17710;
												assign node17710 = (inp[13]) ? node17720 : node17711;
													assign node17711 = (inp[8]) ? node17715 : node17712;
														assign node17712 = (inp[11]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node17715 = (inp[4]) ? node17717 : 16'b0000000111111111;
															assign node17717 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17720 = (inp[8]) ? 16'b0000000011111111 : node17721;
														assign node17721 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17725 = (inp[13]) ? node17731 : node17726;
													assign node17726 = (inp[5]) ? 16'b0000000001111111 : node17727;
														assign node17727 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17731 = (inp[5]) ? node17737 : node17732;
														assign node17732 = (inp[11]) ? 16'b0000000001111111 : node17733;
															assign node17733 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17737 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node17740 = (inp[4]) ? node17758 : node17741;
												assign node17741 = (inp[8]) ? node17751 : node17742;
													assign node17742 = (inp[5]) ? node17746 : node17743;
														assign node17743 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17746 = (inp[14]) ? 16'b0000000001111111 : node17747;
															assign node17747 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17751 = (inp[13]) ? 16'b0000000000111111 : node17752;
														assign node17752 = (inp[5]) ? 16'b0000000001111111 : node17753;
															assign node17753 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17758 = (inp[13]) ? node17764 : node17759;
													assign node17759 = (inp[14]) ? node17761 : 16'b0000000001111111;
														assign node17761 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node17764 = (inp[11]) ? node17766 : 16'b0000000001111111;
														assign node17766 = (inp[5]) ? 16'b0000000000011111 : node17767;
															assign node17767 = (inp[14]) ? node17769 : 16'b0000000000111111;
																assign node17769 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node17773 = (inp[13]) ? node18273 : node17774;
							assign node17774 = (inp[10]) ? node18036 : node17775;
								assign node17775 = (inp[4]) ? node17907 : node17776;
									assign node17776 = (inp[9]) ? node17834 : node17777;
										assign node17777 = (inp[2]) ? node17817 : node17778;
											assign node17778 = (inp[11]) ? node17802 : node17779;
												assign node17779 = (inp[14]) ? node17797 : node17780;
													assign node17780 = (inp[8]) ? node17790 : node17781;
														assign node17781 = (inp[5]) ? node17785 : node17782;
															assign node17782 = (inp[7]) ? 16'b0001111111111111 : 16'b0011111111111111;
															assign node17785 = (inp[7]) ? 16'b0000111111111111 : node17786;
																assign node17786 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node17790 = (inp[7]) ? 16'b0000011111111111 : node17791;
															assign node17791 = (inp[12]) ? 16'b0000111111111111 : node17792;
																assign node17792 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node17797 = (inp[7]) ? 16'b0000011111111111 : node17798;
														assign node17798 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node17802 = (inp[12]) ? node17810 : node17803;
													assign node17803 = (inp[5]) ? node17805 : 16'b0000111111111111;
														assign node17805 = (inp[7]) ? node17807 : 16'b0000011111111111;
															assign node17807 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17810 = (inp[8]) ? node17812 : 16'b0000001111111111;
														assign node17812 = (inp[14]) ? node17814 : 16'b0000001111111111;
															assign node17814 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17817 = (inp[5]) ? node17825 : node17818;
												assign node17818 = (inp[8]) ? node17820 : 16'b0000011111111111;
													assign node17820 = (inp[14]) ? 16'b0000001111111111 : node17821;
														assign node17821 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node17825 = (inp[12]) ? node17831 : node17826;
													assign node17826 = (inp[14]) ? node17828 : 16'b0000011111111111;
														assign node17828 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17831 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17834 = (inp[12]) ? node17868 : node17835;
											assign node17835 = (inp[5]) ? node17853 : node17836;
												assign node17836 = (inp[8]) ? node17846 : node17837;
													assign node17837 = (inp[11]) ? node17843 : node17838;
														assign node17838 = (inp[7]) ? node17840 : 16'b0000111111111111;
															assign node17840 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17843 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17846 = (inp[7]) ? node17848 : 16'b0000011111111111;
														assign node17848 = (inp[14]) ? 16'b0000000111111111 : node17849;
															assign node17849 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17853 = (inp[7]) ? node17863 : node17854;
													assign node17854 = (inp[14]) ? node17858 : node17855;
														assign node17855 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17858 = (inp[8]) ? 16'b0000000111111111 : node17859;
															assign node17859 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17863 = (inp[2]) ? node17865 : 16'b0000000111111111;
														assign node17865 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17868 = (inp[7]) ? node17886 : node17869;
												assign node17869 = (inp[14]) ? node17875 : node17870;
													assign node17870 = (inp[5]) ? node17872 : 16'b0000001111111111;
														assign node17872 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17875 = (inp[5]) ? node17879 : node17876;
														assign node17876 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17879 = (inp[8]) ? 16'b0000000111111111 : node17880;
															assign node17880 = (inp[11]) ? 16'b0000000111111111 : node17881;
																assign node17881 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17886 = (inp[5]) ? node17898 : node17887;
													assign node17887 = (inp[2]) ? node17895 : node17888;
														assign node17888 = (inp[11]) ? node17890 : 16'b0000000111111111;
															assign node17890 = (inp[14]) ? node17892 : 16'b0000000111111111;
																assign node17892 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17895 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17898 = (inp[2]) ? node17902 : node17899;
														assign node17899 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17902 = (inp[14]) ? node17904 : 16'b0000000011111111;
															assign node17904 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node17907 = (inp[11]) ? node17963 : node17908;
										assign node17908 = (inp[14]) ? node17934 : node17909;
											assign node17909 = (inp[5]) ? node17925 : node17910;
												assign node17910 = (inp[8]) ? node17920 : node17911;
													assign node17911 = (inp[12]) ? node17913 : 16'b0000111111111111;
														assign node17913 = (inp[9]) ? node17915 : 16'b0000011111111111;
															assign node17915 = (inp[2]) ? 16'b0000001111111111 : node17916;
																assign node17916 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17920 = (inp[12]) ? 16'b0000000111111111 : node17921;
														assign node17921 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node17925 = (inp[9]) ? node17927 : 16'b0000001111111111;
													assign node17927 = (inp[12]) ? node17931 : node17928;
														assign node17928 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17931 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17934 = (inp[2]) ? node17956 : node17935;
												assign node17935 = (inp[7]) ? node17949 : node17936;
													assign node17936 = (inp[5]) ? node17942 : node17937;
														assign node17937 = (inp[9]) ? node17939 : 16'b0000011111111111;
															assign node17939 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17942 = (inp[8]) ? 16'b0000000111111111 : node17943;
															assign node17943 = (inp[12]) ? node17945 : 16'b0000001111111111;
																assign node17945 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17949 = (inp[9]) ? node17953 : node17950;
														assign node17950 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17953 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17956 = (inp[7]) ? node17958 : 16'b0000000111111111;
													assign node17958 = (inp[12]) ? node17960 : 16'b0000000111111111;
														assign node17960 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node17963 = (inp[7]) ? node17997 : node17964;
											assign node17964 = (inp[12]) ? node17980 : node17965;
												assign node17965 = (inp[5]) ? node17975 : node17966;
													assign node17966 = (inp[8]) ? node17972 : node17967;
														assign node17967 = (inp[2]) ? 16'b0000001111111111 : node17968;
															assign node17968 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17972 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node17975 = (inp[2]) ? 16'b0000000111111111 : node17976;
														assign node17976 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17980 = (inp[2]) ? node17994 : node17981;
													assign node17981 = (inp[9]) ? node17989 : node17982;
														assign node17982 = (inp[14]) ? 16'b0000000111111111 : node17983;
															assign node17983 = (inp[8]) ? node17985 : 16'b0000001111111111;
																assign node17985 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17989 = (inp[5]) ? node17991 : 16'b0000000111111111;
															assign node17991 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17994 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17997 = (inp[14]) ? node18021 : node17998;
												assign node17998 = (inp[9]) ? node18014 : node17999;
													assign node17999 = (inp[12]) ? node18009 : node18000;
														assign node18000 = (inp[5]) ? node18006 : node18001;
															assign node18001 = (inp[2]) ? node18003 : 16'b0000001111111111;
																assign node18003 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node18006 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18009 = (inp[8]) ? node18011 : 16'b0000000111111111;
															assign node18011 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18014 = (inp[8]) ? node18018 : node18015;
														assign node18015 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18018 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18021 = (inp[12]) ? node18029 : node18022;
													assign node18022 = (inp[8]) ? node18026 : node18023;
														assign node18023 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18026 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18029 = (inp[5]) ? node18033 : node18030;
														assign node18030 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18033 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node18036 = (inp[11]) ? node18148 : node18037;
									assign node18037 = (inp[7]) ? node18087 : node18038;
										assign node18038 = (inp[5]) ? node18062 : node18039;
											assign node18039 = (inp[12]) ? node18055 : node18040;
												assign node18040 = (inp[9]) ? node18050 : node18041;
													assign node18041 = (inp[14]) ? node18045 : node18042;
														assign node18042 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node18045 = (inp[2]) ? node18047 : 16'b0000011111111111;
															assign node18047 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18050 = (inp[2]) ? 16'b0000001111111111 : node18051;
														assign node18051 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18055 = (inp[9]) ? node18057 : 16'b0000001111111111;
													assign node18057 = (inp[2]) ? 16'b0000000111111111 : node18058;
														assign node18058 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node18062 = (inp[12]) ? node18078 : node18063;
												assign node18063 = (inp[14]) ? node18073 : node18064;
													assign node18064 = (inp[4]) ? node18070 : node18065;
														assign node18065 = (inp[2]) ? 16'b0000001111111111 : node18066;
															assign node18066 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18070 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18073 = (inp[8]) ? 16'b0000000011111111 : node18074;
														assign node18074 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18078 = (inp[8]) ? 16'b0000000011111111 : node18079;
													assign node18079 = (inp[9]) ? node18081 : 16'b0000000111111111;
														assign node18081 = (inp[4]) ? node18083 : 16'b0000000111111111;
															assign node18083 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18087 = (inp[9]) ? node18117 : node18088;
											assign node18088 = (inp[14]) ? node18104 : node18089;
												assign node18089 = (inp[2]) ? node18099 : node18090;
													assign node18090 = (inp[5]) ? node18094 : node18091;
														assign node18091 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18094 = (inp[4]) ? node18096 : 16'b0000001111111111;
															assign node18096 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18099 = (inp[12]) ? node18101 : 16'b0000001111111111;
														assign node18101 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18104 = (inp[4]) ? node18106 : 16'b0000000111111111;
													assign node18106 = (inp[12]) ? node18114 : node18107;
														assign node18107 = (inp[5]) ? 16'b0000000011111111 : node18108;
															assign node18108 = (inp[2]) ? 16'b0000000111111111 : node18109;
																assign node18109 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18114 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18117 = (inp[8]) ? node18129 : node18118;
												assign node18118 = (inp[2]) ? node18120 : 16'b0000000111111111;
													assign node18120 = (inp[14]) ? 16'b0000000011111111 : node18121;
														assign node18121 = (inp[4]) ? 16'b0000000011111111 : node18122;
															assign node18122 = (inp[12]) ? node18124 : 16'b0000000111111111;
																assign node18124 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18129 = (inp[4]) ? node18137 : node18130;
													assign node18130 = (inp[12]) ? node18134 : node18131;
														assign node18131 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18134 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18137 = (inp[2]) ? node18141 : node18138;
														assign node18138 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node18141 = (inp[14]) ? node18143 : 16'b0000000001111111;
															assign node18143 = (inp[12]) ? node18145 : 16'b0000000000111111;
																assign node18145 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node18148 = (inp[14]) ? node18220 : node18149;
										assign node18149 = (inp[9]) ? node18191 : node18150;
											assign node18150 = (inp[2]) ? node18170 : node18151;
												assign node18151 = (inp[8]) ? node18159 : node18152;
													assign node18152 = (inp[4]) ? 16'b0000001111111111 : node18153;
														assign node18153 = (inp[5]) ? node18155 : 16'b0000011111111111;
															assign node18155 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18159 = (inp[12]) ? node18167 : node18160;
														assign node18160 = (inp[5]) ? node18162 : 16'b0000001111111111;
															assign node18162 = (inp[7]) ? 16'b0000000111111111 : node18163;
																assign node18163 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18167 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node18170 = (inp[8]) ? node18178 : node18171;
													assign node18171 = (inp[12]) ? node18175 : node18172;
														assign node18172 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18175 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18178 = (inp[7]) ? node18186 : node18179;
														assign node18179 = (inp[5]) ? node18181 : 16'b0000001111111111;
															assign node18181 = (inp[4]) ? 16'b0000000011111111 : node18182;
																assign node18182 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18186 = (inp[5]) ? node18188 : 16'b0000000011111111;
															assign node18188 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18191 = (inp[7]) ? node18201 : node18192;
												assign node18192 = (inp[5]) ? 16'b0000000011111111 : node18193;
													assign node18193 = (inp[8]) ? 16'b0000000011111111 : node18194;
														assign node18194 = (inp[2]) ? node18196 : 16'b0000000111111111;
															assign node18196 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18201 = (inp[4]) ? node18215 : node18202;
													assign node18202 = (inp[12]) ? node18208 : node18203;
														assign node18203 = (inp[5]) ? node18205 : 16'b0000000111111111;
															assign node18205 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node18208 = (inp[8]) ? 16'b0000000001111111 : node18209;
															assign node18209 = (inp[5]) ? node18211 : 16'b0000000011111111;
																assign node18211 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18215 = (inp[2]) ? node18217 : 16'b0000000001111111;
														assign node18217 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node18220 = (inp[4]) ? node18246 : node18221;
											assign node18221 = (inp[2]) ? node18231 : node18222;
												assign node18222 = (inp[7]) ? 16'b0000000011111111 : node18223;
													assign node18223 = (inp[9]) ? node18227 : node18224;
														assign node18224 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18227 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18231 = (inp[7]) ? node18243 : node18232;
													assign node18232 = (inp[9]) ? node18236 : node18233;
														assign node18233 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node18236 = (inp[5]) ? node18238 : 16'b0000000011111111;
															assign node18238 = (inp[12]) ? 16'b0000000001111111 : node18239;
																assign node18239 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18243 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18246 = (inp[12]) ? node18260 : node18247;
												assign node18247 = (inp[5]) ? node18255 : node18248;
													assign node18248 = (inp[8]) ? node18252 : node18249;
														assign node18249 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18252 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node18255 = (inp[9]) ? 16'b0000000000111111 : node18256;
														assign node18256 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18260 = (inp[2]) ? 16'b0000000000111111 : node18261;
													assign node18261 = (inp[7]) ? node18267 : node18262;
														assign node18262 = (inp[8]) ? 16'b0000000001111111 : node18263;
															assign node18263 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18267 = (inp[9]) ? node18269 : 16'b0000000001111111;
															assign node18269 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node18273 = (inp[5]) ? node18503 : node18274;
								assign node18274 = (inp[8]) ? node18392 : node18275;
									assign node18275 = (inp[7]) ? node18343 : node18276;
										assign node18276 = (inp[12]) ? node18310 : node18277;
											assign node18277 = (inp[14]) ? node18293 : node18278;
												assign node18278 = (inp[10]) ? node18286 : node18279;
													assign node18279 = (inp[9]) ? node18283 : node18280;
														assign node18280 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node18283 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18286 = (inp[9]) ? node18290 : node18287;
														assign node18287 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18290 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18293 = (inp[2]) ? node18301 : node18294;
													assign node18294 = (inp[4]) ? node18298 : node18295;
														assign node18295 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node18298 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18301 = (inp[11]) ? node18307 : node18302;
														assign node18302 = (inp[4]) ? 16'b0000000111111111 : node18303;
															assign node18303 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18307 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18310 = (inp[10]) ? node18332 : node18311;
												assign node18311 = (inp[4]) ? node18321 : node18312;
													assign node18312 = (inp[14]) ? node18316 : node18313;
														assign node18313 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18316 = (inp[2]) ? node18318 : 16'b0000001111111111;
															assign node18318 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18321 = (inp[2]) ? node18327 : node18322;
														assign node18322 = (inp[9]) ? 16'b0000000111111111 : node18323;
															assign node18323 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18327 = (inp[11]) ? 16'b0000000011111111 : node18328;
															assign node18328 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18332 = (inp[2]) ? node18338 : node18333;
													assign node18333 = (inp[9]) ? node18335 : 16'b0000000111111111;
														assign node18335 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18338 = (inp[14]) ? 16'b0000000011111111 : node18339;
														assign node18339 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18343 = (inp[10]) ? node18365 : node18344;
											assign node18344 = (inp[11]) ? node18352 : node18345;
												assign node18345 = (inp[4]) ? node18347 : 16'b0000001111111111;
													assign node18347 = (inp[2]) ? 16'b0000000111111111 : node18348;
														assign node18348 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node18352 = (inp[14]) ? node18360 : node18353;
													assign node18353 = (inp[4]) ? 16'b0000000111111111 : node18354;
														assign node18354 = (inp[9]) ? 16'b0000000111111111 : node18355;
															assign node18355 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18360 = (inp[12]) ? node18362 : 16'b0000000111111111;
														assign node18362 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18365 = (inp[14]) ? node18379 : node18366;
												assign node18366 = (inp[2]) ? node18372 : node18367;
													assign node18367 = (inp[12]) ? 16'b0000000011111111 : node18368;
														assign node18368 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18372 = (inp[11]) ? node18376 : node18373;
														assign node18373 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18376 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18379 = (inp[4]) ? node18385 : node18380;
													assign node18380 = (inp[11]) ? 16'b0000000011111111 : node18381;
														assign node18381 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18385 = (inp[11]) ? 16'b0000000001111111 : node18386;
														assign node18386 = (inp[9]) ? 16'b0000000001111111 : node18387;
															assign node18387 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node18392 = (inp[14]) ? node18450 : node18393;
										assign node18393 = (inp[12]) ? node18411 : node18394;
											assign node18394 = (inp[10]) ? node18402 : node18395;
												assign node18395 = (inp[2]) ? 16'b0000000111111111 : node18396;
													assign node18396 = (inp[11]) ? node18398 : 16'b0000001111111111;
														assign node18398 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18402 = (inp[4]) ? 16'b0000000011111111 : node18403;
													assign node18403 = (inp[7]) ? node18405 : 16'b0000000111111111;
														assign node18405 = (inp[9]) ? 16'b0000000011111111 : node18406;
															assign node18406 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18411 = (inp[9]) ? node18429 : node18412;
												assign node18412 = (inp[4]) ? node18422 : node18413;
													assign node18413 = (inp[7]) ? node18417 : node18414;
														assign node18414 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node18417 = (inp[11]) ? node18419 : 16'b0000000111111111;
															assign node18419 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18422 = (inp[7]) ? node18426 : node18423;
														assign node18423 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18426 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18429 = (inp[2]) ? node18441 : node18430;
													assign node18430 = (inp[11]) ? node18438 : node18431;
														assign node18431 = (inp[10]) ? node18433 : 16'b0000000111111111;
															assign node18433 = (inp[4]) ? 16'b0000000011111111 : node18434;
																assign node18434 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18438 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18441 = (inp[7]) ? node18445 : node18442;
														assign node18442 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18445 = (inp[11]) ? 16'b0000000000011111 : node18446;
															assign node18446 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node18450 = (inp[9]) ? node18480 : node18451;
											assign node18451 = (inp[12]) ? node18463 : node18452;
												assign node18452 = (inp[7]) ? node18456 : node18453;
													assign node18453 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18456 = (inp[11]) ? node18460 : node18457;
														assign node18457 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18460 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18463 = (inp[11]) ? node18471 : node18464;
													assign node18464 = (inp[4]) ? node18468 : node18465;
														assign node18465 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18468 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node18471 = (inp[10]) ? node18475 : node18472;
														assign node18472 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18475 = (inp[4]) ? node18477 : 16'b0000000001111111;
															assign node18477 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18480 = (inp[7]) ? node18490 : node18481;
												assign node18481 = (inp[12]) ? 16'b0000000001111111 : node18482;
													assign node18482 = (inp[4]) ? node18486 : node18483;
														assign node18483 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18486 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18490 = (inp[4]) ? node18494 : node18491;
													assign node18491 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18494 = (inp[11]) ? node18500 : node18495;
														assign node18495 = (inp[10]) ? 16'b0000000000111111 : node18496;
															assign node18496 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18500 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node18503 = (inp[4]) ? node18583 : node18504;
									assign node18504 = (inp[11]) ? node18560 : node18505;
										assign node18505 = (inp[12]) ? node18527 : node18506;
											assign node18506 = (inp[7]) ? node18514 : node18507;
												assign node18507 = (inp[9]) ? 16'b0000000111111111 : node18508;
													assign node18508 = (inp[14]) ? node18510 : 16'b0000001111111111;
														assign node18510 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18514 = (inp[14]) ? 16'b0000000011111111 : node18515;
													assign node18515 = (inp[9]) ? node18523 : node18516;
														assign node18516 = (inp[8]) ? node18518 : 16'b0000001111111111;
															assign node18518 = (inp[2]) ? node18520 : 16'b0000001111111111;
																assign node18520 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18523 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18527 = (inp[8]) ? node18539 : node18528;
												assign node18528 = (inp[14]) ? node18532 : node18529;
													assign node18529 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node18532 = (inp[10]) ? node18536 : node18533;
														assign node18533 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18536 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18539 = (inp[10]) ? node18553 : node18540;
													assign node18540 = (inp[9]) ? node18546 : node18541;
														assign node18541 = (inp[2]) ? 16'b0000000011111111 : node18542;
															assign node18542 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18546 = (inp[7]) ? 16'b0000000001111111 : node18547;
															assign node18547 = (inp[14]) ? 16'b0000000001111111 : node18548;
																assign node18548 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18553 = (inp[9]) ? node18557 : node18554;
														assign node18554 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18557 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node18560 = (inp[7]) ? node18572 : node18561;
											assign node18561 = (inp[9]) ? node18565 : node18562;
												assign node18562 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18565 = (inp[10]) ? node18567 : 16'b0000000011111111;
													assign node18567 = (inp[14]) ? 16'b0000000000111111 : node18568;
														assign node18568 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18572 = (inp[12]) ? node18576 : node18573;
												assign node18573 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18576 = (inp[8]) ? 16'b0000000000011111 : node18577;
													assign node18577 = (inp[9]) ? 16'b0000000001111111 : node18578;
														assign node18578 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node18583 = (inp[7]) ? node18635 : node18584;
										assign node18584 = (inp[8]) ? node18612 : node18585;
											assign node18585 = (inp[9]) ? node18597 : node18586;
												assign node18586 = (inp[14]) ? 16'b0000000011111111 : node18587;
													assign node18587 = (inp[10]) ? node18593 : node18588;
														assign node18588 = (inp[11]) ? 16'b0000000111111111 : node18589;
															assign node18589 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18593 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18597 = (inp[12]) ? node18605 : node18598;
													assign node18598 = (inp[14]) ? node18602 : node18599;
														assign node18599 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node18602 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18605 = (inp[11]) ? 16'b0000000001111111 : node18606;
														assign node18606 = (inp[2]) ? 16'b0000000001111111 : node18607;
															assign node18607 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18612 = (inp[10]) ? node18624 : node18613;
												assign node18613 = (inp[9]) ? node18615 : 16'b0000000000111111;
													assign node18615 = (inp[11]) ? node18617 : 16'b0000000011111111;
														assign node18617 = (inp[12]) ? 16'b0000000001111111 : node18618;
															assign node18618 = (inp[2]) ? 16'b0000000001111111 : node18619;
																assign node18619 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18624 = (inp[12]) ? node18628 : node18625;
													assign node18625 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18628 = (inp[11]) ? node18632 : node18629;
														assign node18629 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18632 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node18635 = (inp[14]) ? node18673 : node18636;
											assign node18636 = (inp[2]) ? node18658 : node18637;
												assign node18637 = (inp[12]) ? node18643 : node18638;
													assign node18638 = (inp[9]) ? 16'b0000000011111111 : node18639;
														assign node18639 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18643 = (inp[11]) ? node18651 : node18644;
														assign node18644 = (inp[10]) ? node18646 : 16'b0000000011111111;
															assign node18646 = (inp[9]) ? 16'b0000000001111111 : node18647;
																assign node18647 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18651 = (inp[10]) ? node18655 : node18652;
															assign node18652 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node18655 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node18658 = (inp[10]) ? node18664 : node18659;
													assign node18659 = (inp[9]) ? node18661 : 16'b0000000001111111;
														assign node18661 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node18664 = (inp[8]) ? node18670 : node18665;
														assign node18665 = (inp[12]) ? 16'b0000000000111111 : node18666;
															assign node18666 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18670 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node18673 = (inp[12]) ? node18685 : node18674;
												assign node18674 = (inp[10]) ? node18680 : node18675;
													assign node18675 = (inp[9]) ? node18677 : 16'b0000000001111111;
														assign node18677 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18680 = (inp[2]) ? node18682 : 16'b0000000000111111;
														assign node18682 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node18685 = (inp[11]) ? node18693 : node18686;
													assign node18686 = (inp[10]) ? node18688 : 16'b0000000000111111;
														assign node18688 = (inp[2]) ? 16'b0000000000011111 : node18689;
															assign node18689 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node18693 = (inp[2]) ? node18701 : node18694;
														assign node18694 = (inp[8]) ? node18696 : 16'b0000000000111111;
															assign node18696 = (inp[9]) ? node18698 : 16'b0000000000011111;
																assign node18698 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node18701 = (inp[8]) ? node18703 : 16'b0000000000001111;
															assign node18703 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node18706 = (inp[13]) ? node19716 : node18707;
						assign node18707 = (inp[12]) ? node19225 : node18708;
							assign node18708 = (inp[7]) ? node18992 : node18709;
								assign node18709 = (inp[8]) ? node18853 : node18710;
									assign node18710 = (inp[14]) ? node18778 : node18711;
										assign node18711 = (inp[5]) ? node18745 : node18712;
											assign node18712 = (inp[11]) ? node18734 : node18713;
												assign node18713 = (inp[4]) ? node18727 : node18714;
													assign node18714 = (inp[10]) ? node18722 : node18715;
														assign node18715 = (inp[15]) ? node18717 : 16'b0001111111111111;
															assign node18717 = (inp[9]) ? 16'b0000111111111111 : node18718;
																assign node18718 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node18722 = (inp[9]) ? 16'b0000011111111111 : node18723;
															assign node18723 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node18727 = (inp[2]) ? 16'b0000011111111111 : node18728;
														assign node18728 = (inp[9]) ? 16'b0000001111111111 : node18729;
															assign node18729 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node18734 = (inp[2]) ? node18740 : node18735;
													assign node18735 = (inp[15]) ? node18737 : 16'b0000011111111111;
														assign node18737 = (inp[4]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node18740 = (inp[10]) ? 16'b0000001111111111 : node18741;
														assign node18741 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node18745 = (inp[4]) ? node18759 : node18746;
												assign node18746 = (inp[11]) ? node18752 : node18747;
													assign node18747 = (inp[10]) ? node18749 : 16'b0000111111111111;
														assign node18749 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node18752 = (inp[2]) ? 16'b0000001111111111 : node18753;
														assign node18753 = (inp[15]) ? node18755 : 16'b0000011111111111;
															assign node18755 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18759 = (inp[11]) ? node18769 : node18760;
													assign node18760 = (inp[2]) ? node18766 : node18761;
														assign node18761 = (inp[9]) ? node18763 : 16'b0000011111111111;
															assign node18763 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18766 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18769 = (inp[15]) ? node18773 : node18770;
														assign node18770 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18773 = (inp[2]) ? node18775 : 16'b0000000111111111;
															assign node18775 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18778 = (inp[5]) ? node18810 : node18779;
											assign node18779 = (inp[2]) ? node18793 : node18780;
												assign node18780 = (inp[9]) ? node18788 : node18781;
													assign node18781 = (inp[4]) ? 16'b0000011111111111 : node18782;
														assign node18782 = (inp[15]) ? 16'b0000011111111111 : node18783;
															assign node18783 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node18788 = (inp[10]) ? node18790 : 16'b0000011111111111;
														assign node18790 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node18793 = (inp[9]) ? node18801 : node18794;
													assign node18794 = (inp[15]) ? node18798 : node18795;
														assign node18795 = (inp[4]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node18798 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18801 = (inp[11]) ? node18805 : node18802;
														assign node18802 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18805 = (inp[10]) ? node18807 : 16'b0000000111111111;
															assign node18807 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18810 = (inp[15]) ? node18836 : node18811;
												assign node18811 = (inp[10]) ? node18823 : node18812;
													assign node18812 = (inp[4]) ? node18816 : node18813;
														assign node18813 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18816 = (inp[11]) ? 16'b0000001111111111 : node18817;
															assign node18817 = (inp[2]) ? 16'b0000001111111111 : node18818;
																assign node18818 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18823 = (inp[4]) ? node18829 : node18824;
														assign node18824 = (inp[11]) ? node18826 : 16'b0000001111111111;
															assign node18826 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18829 = (inp[2]) ? node18831 : 16'b0000000111111111;
															assign node18831 = (inp[11]) ? 16'b0000000011111111 : node18832;
																assign node18832 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18836 = (inp[9]) ? 16'b0000000011111111 : node18837;
													assign node18837 = (inp[2]) ? node18849 : node18838;
														assign node18838 = (inp[4]) ? node18844 : node18839;
															assign node18839 = (inp[10]) ? node18841 : 16'b0000001111111111;
																assign node18841 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node18844 = (inp[10]) ? node18846 : 16'b0000000111111111;
																assign node18846 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18849 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node18853 = (inp[4]) ? node18923 : node18854;
										assign node18854 = (inp[2]) ? node18888 : node18855;
											assign node18855 = (inp[11]) ? node18871 : node18856;
												assign node18856 = (inp[9]) ? node18864 : node18857;
													assign node18857 = (inp[10]) ? node18859 : 16'b0000111111111111;
														assign node18859 = (inp[5]) ? node18861 : 16'b0000011111111111;
															assign node18861 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18864 = (inp[10]) ? 16'b0000001111111111 : node18865;
														assign node18865 = (inp[14]) ? node18867 : 16'b0000011111111111;
															assign node18867 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node18871 = (inp[10]) ? node18879 : node18872;
													assign node18872 = (inp[5]) ? 16'b0000001111111111 : node18873;
														assign node18873 = (inp[15]) ? node18875 : 16'b0000011111111111;
															assign node18875 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18879 = (inp[14]) ? node18885 : node18880;
														assign node18880 = (inp[5]) ? 16'b0000000111111111 : node18881;
															assign node18881 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18885 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18888 = (inp[5]) ? node18902 : node18889;
												assign node18889 = (inp[15]) ? node18893 : node18890;
													assign node18890 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18893 = (inp[10]) ? node18897 : node18894;
														assign node18894 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18897 = (inp[9]) ? node18899 : 16'b0000000111111111;
															assign node18899 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18902 = (inp[10]) ? node18912 : node18903;
													assign node18903 = (inp[14]) ? node18909 : node18904;
														assign node18904 = (inp[9]) ? node18906 : 16'b0000001111111111;
															assign node18906 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18909 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18912 = (inp[9]) ? node18920 : node18913;
														assign node18913 = (inp[14]) ? 16'b0000000011111111 : node18914;
															assign node18914 = (inp[11]) ? node18916 : 16'b0000000111111111;
																assign node18916 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18920 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node18923 = (inp[11]) ? node18957 : node18924;
											assign node18924 = (inp[14]) ? node18942 : node18925;
												assign node18925 = (inp[2]) ? node18933 : node18926;
													assign node18926 = (inp[5]) ? node18928 : 16'b0000001111111111;
														assign node18928 = (inp[10]) ? 16'b0000000111111111 : node18929;
															assign node18929 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18933 = (inp[9]) ? node18937 : node18934;
														assign node18934 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node18937 = (inp[10]) ? node18939 : 16'b0000000111111111;
															assign node18939 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18942 = (inp[15]) ? node18944 : 16'b0000000111111111;
													assign node18944 = (inp[2]) ? node18952 : node18945;
														assign node18945 = (inp[9]) ? node18947 : 16'b0000001111111111;
															assign node18947 = (inp[10]) ? 16'b0000000011111111 : node18948;
																assign node18948 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18952 = (inp[10]) ? node18954 : 16'b0000000011111111;
															assign node18954 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18957 = (inp[15]) ? node18973 : node18958;
												assign node18958 = (inp[10]) ? node18964 : node18959;
													assign node18959 = (inp[9]) ? 16'b0000000111111111 : node18960;
														assign node18960 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18964 = (inp[9]) ? node18968 : node18965;
														assign node18965 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18968 = (inp[5]) ? node18970 : 16'b0000000011111111;
															assign node18970 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18973 = (inp[2]) ? node18981 : node18974;
													assign node18974 = (inp[10]) ? node18978 : node18975;
														assign node18975 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18978 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18981 = (inp[5]) ? node18987 : node18982;
														assign node18982 = (inp[9]) ? node18984 : 16'b0000000001111111;
															assign node18984 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18987 = (inp[14]) ? node18989 : 16'b0000000000111111;
															assign node18989 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node18992 = (inp[9]) ? node19124 : node18993;
									assign node18993 = (inp[14]) ? node19059 : node18994;
										assign node18994 = (inp[11]) ? node19026 : node18995;
											assign node18995 = (inp[5]) ? node19011 : node18996;
												assign node18996 = (inp[15]) ? 16'b0000001111111111 : node18997;
													assign node18997 = (inp[10]) ? node19003 : node18998;
														assign node18998 = (inp[8]) ? 16'b0000011111111111 : node18999;
															assign node18999 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19003 = (inp[4]) ? 16'b0000001111111111 : node19004;
															assign node19004 = (inp[2]) ? node19006 : 16'b0000111111111111;
																assign node19006 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19011 = (inp[15]) ? node19021 : node19012;
													assign node19012 = (inp[2]) ? node19018 : node19013;
														assign node19013 = (inp[8]) ? 16'b0000001111111111 : node19014;
															assign node19014 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19018 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19021 = (inp[10]) ? 16'b0000000111111111 : node19022;
														assign node19022 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node19026 = (inp[4]) ? node19040 : node19027;
												assign node19027 = (inp[5]) ? node19035 : node19028;
													assign node19028 = (inp[2]) ? 16'b0000001111111111 : node19029;
														assign node19029 = (inp[8]) ? node19031 : 16'b0000111111111111;
															assign node19031 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19035 = (inp[15]) ? 16'b0000000011111111 : node19036;
														assign node19036 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19040 = (inp[8]) ? node19048 : node19041;
													assign node19041 = (inp[10]) ? node19045 : node19042;
														assign node19042 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19045 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19048 = (inp[15]) ? node19052 : node19049;
														assign node19049 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19052 = (inp[5]) ? node19054 : 16'b0000000011111111;
															assign node19054 = (inp[2]) ? 16'b0000000001111111 : node19055;
																assign node19055 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19059 = (inp[4]) ? node19081 : node19060;
											assign node19060 = (inp[10]) ? node19076 : node19061;
												assign node19061 = (inp[15]) ? node19069 : node19062;
													assign node19062 = (inp[5]) ? node19064 : 16'b0000001111111111;
														assign node19064 = (inp[11]) ? node19066 : 16'b0000001111111111;
															assign node19066 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19069 = (inp[5]) ? 16'b0000000111111111 : node19070;
														assign node19070 = (inp[8]) ? 16'b0000000111111111 : node19071;
															assign node19071 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19076 = (inp[8]) ? node19078 : 16'b0000000111111111;
													assign node19078 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19081 = (inp[5]) ? node19105 : node19082;
												assign node19082 = (inp[8]) ? node19092 : node19083;
													assign node19083 = (inp[10]) ? node19087 : node19084;
														assign node19084 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19087 = (inp[2]) ? 16'b0000000011111111 : node19088;
															assign node19088 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19092 = (inp[10]) ? node19098 : node19093;
														assign node19093 = (inp[2]) ? 16'b0000000011111111 : node19094;
															assign node19094 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19098 = (inp[15]) ? 16'b0000000001111111 : node19099;
															assign node19099 = (inp[11]) ? 16'b0000000001111111 : node19100;
																assign node19100 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19105 = (inp[11]) ? node19117 : node19106;
													assign node19106 = (inp[8]) ? node19110 : node19107;
														assign node19107 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19110 = (inp[15]) ? node19112 : 16'b0000000011111111;
															assign node19112 = (inp[2]) ? 16'b0000000001111111 : node19113;
																assign node19113 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19117 = (inp[8]) ? 16'b0000000000111111 : node19118;
														assign node19118 = (inp[2]) ? 16'b0000000001111111 : node19119;
															assign node19119 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node19124 = (inp[11]) ? node19172 : node19125;
										assign node19125 = (inp[10]) ? node19149 : node19126;
											assign node19126 = (inp[8]) ? node19136 : node19127;
												assign node19127 = (inp[4]) ? node19131 : node19128;
													assign node19128 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19131 = (inp[15]) ? node19133 : 16'b0000000111111111;
														assign node19133 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19136 = (inp[15]) ? node19144 : node19137;
													assign node19137 = (inp[2]) ? node19139 : 16'b0000001111111111;
														assign node19139 = (inp[5]) ? 16'b0000000011111111 : node19140;
															assign node19140 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19144 = (inp[2]) ? node19146 : 16'b0000000011111111;
														assign node19146 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19149 = (inp[4]) ? node19163 : node19150;
												assign node19150 = (inp[2]) ? node19156 : node19151;
													assign node19151 = (inp[15]) ? node19153 : 16'b0000000111111111;
														assign node19153 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19156 = (inp[8]) ? node19158 : 16'b0000000011111111;
														assign node19158 = (inp[15]) ? 16'b0000000011111111 : node19159;
															assign node19159 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19163 = (inp[8]) ? 16'b0000000001111111 : node19164;
													assign node19164 = (inp[14]) ? node19168 : node19165;
														assign node19165 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19168 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19172 = (inp[5]) ? node19198 : node19173;
											assign node19173 = (inp[4]) ? node19181 : node19174;
												assign node19174 = (inp[15]) ? 16'b0000000011111111 : node19175;
													assign node19175 = (inp[2]) ? node19177 : 16'b0000000111111111;
														assign node19177 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19181 = (inp[10]) ? node19191 : node19182;
													assign node19182 = (inp[15]) ? node19186 : node19183;
														assign node19183 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19186 = (inp[14]) ? 16'b0000000001111111 : node19187;
															assign node19187 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19191 = (inp[2]) ? node19195 : node19192;
														assign node19192 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19195 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node19198 = (inp[14]) ? node19212 : node19199;
												assign node19199 = (inp[10]) ? node19205 : node19200;
													assign node19200 = (inp[15]) ? node19202 : 16'b0000001111111111;
														assign node19202 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19205 = (inp[15]) ? 16'b0000000001111111 : node19206;
														assign node19206 = (inp[8]) ? 16'b0000000001111111 : node19207;
															assign node19207 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19212 = (inp[8]) ? node19218 : node19213;
													assign node19213 = (inp[4]) ? node19215 : 16'b0000000001111111;
														assign node19215 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19218 = (inp[10]) ? 16'b0000000000111111 : node19219;
														assign node19219 = (inp[15]) ? 16'b0000000000111111 : node19220;
															assign node19220 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node19225 = (inp[15]) ? node19495 : node19226;
								assign node19226 = (inp[2]) ? node19358 : node19227;
									assign node19227 = (inp[5]) ? node19293 : node19228;
										assign node19228 = (inp[10]) ? node19266 : node19229;
											assign node19229 = (inp[8]) ? node19243 : node19230;
												assign node19230 = (inp[7]) ? node19236 : node19231;
													assign node19231 = (inp[4]) ? 16'b0000011111111111 : node19232;
														assign node19232 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node19236 = (inp[9]) ? node19240 : node19237;
														assign node19237 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19240 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19243 = (inp[9]) ? node19255 : node19244;
													assign node19244 = (inp[4]) ? node19248 : node19245;
														assign node19245 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19248 = (inp[7]) ? node19250 : 16'b0000001111111111;
															assign node19250 = (inp[11]) ? 16'b0000000111111111 : node19251;
																assign node19251 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19255 = (inp[11]) ? node19263 : node19256;
														assign node19256 = (inp[14]) ? node19258 : 16'b0000001111111111;
															assign node19258 = (inp[4]) ? 16'b0000000111111111 : node19259;
																assign node19259 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19263 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node19266 = (inp[8]) ? node19276 : node19267;
												assign node19267 = (inp[11]) ? node19269 : 16'b0000001111111111;
													assign node19269 = (inp[14]) ? node19273 : node19270;
														assign node19270 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19273 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19276 = (inp[4]) ? node19278 : 16'b0000000111111111;
													assign node19278 = (inp[14]) ? node19290 : node19279;
														assign node19279 = (inp[11]) ? node19285 : node19280;
															assign node19280 = (inp[9]) ? 16'b0000000111111111 : node19281;
																assign node19281 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node19285 = (inp[7]) ? 16'b0000000011111111 : node19286;
																assign node19286 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19290 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19293 = (inp[14]) ? node19331 : node19294;
											assign node19294 = (inp[11]) ? node19314 : node19295;
												assign node19295 = (inp[8]) ? node19303 : node19296;
													assign node19296 = (inp[4]) ? node19300 : node19297;
														assign node19297 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19300 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19303 = (inp[9]) ? 16'b0000000001111111 : node19304;
														assign node19304 = (inp[10]) ? node19310 : node19305;
															assign node19305 = (inp[7]) ? node19307 : 16'b0000001111111111;
																assign node19307 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node19310 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19314 = (inp[7]) ? node19324 : node19315;
													assign node19315 = (inp[10]) ? node19319 : node19316;
														assign node19316 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19319 = (inp[9]) ? node19321 : 16'b0000000111111111;
															assign node19321 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19324 = (inp[8]) ? 16'b0000000011111111 : node19325;
														assign node19325 = (inp[4]) ? node19327 : 16'b0000000111111111;
															assign node19327 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19331 = (inp[7]) ? node19341 : node19332;
												assign node19332 = (inp[8]) ? 16'b0000000011111111 : node19333;
													assign node19333 = (inp[9]) ? node19337 : node19334;
														assign node19334 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node19337 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19341 = (inp[9]) ? node19353 : node19342;
													assign node19342 = (inp[10]) ? node19350 : node19343;
														assign node19343 = (inp[4]) ? node19345 : 16'b0000000111111111;
															assign node19345 = (inp[8]) ? 16'b0000000011111111 : node19346;
																assign node19346 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19350 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19353 = (inp[10]) ? node19355 : 16'b0000000001111111;
														assign node19355 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node19358 = (inp[5]) ? node19444 : node19359;
										assign node19359 = (inp[4]) ? node19407 : node19360;
											assign node19360 = (inp[10]) ? node19388 : node19361;
												assign node19361 = (inp[8]) ? node19373 : node19362;
													assign node19362 = (inp[9]) ? node19370 : node19363;
														assign node19363 = (inp[7]) ? node19365 : 16'b0000011111111111;
															assign node19365 = (inp[14]) ? 16'b0000001111111111 : node19366;
																assign node19366 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19370 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19373 = (inp[7]) ? node19381 : node19374;
														assign node19374 = (inp[11]) ? node19378 : node19375;
															assign node19375 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node19378 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19381 = (inp[9]) ? node19383 : 16'b0000000111111111;
															assign node19383 = (inp[14]) ? 16'b0000000001111111 : node19384;
																assign node19384 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19388 = (inp[7]) ? node19404 : node19389;
													assign node19389 = (inp[14]) ? node19393 : node19390;
														assign node19390 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node19393 = (inp[8]) ? node19399 : node19394;
															assign node19394 = (inp[11]) ? node19396 : 16'b0000000111111111;
																assign node19396 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node19399 = (inp[9]) ? 16'b0000000011111111 : node19400;
																assign node19400 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19404 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19407 = (inp[8]) ? node19425 : node19408;
												assign node19408 = (inp[7]) ? node19416 : node19409;
													assign node19409 = (inp[11]) ? node19413 : node19410;
														assign node19410 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19413 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19416 = (inp[9]) ? node19420 : node19417;
														assign node19417 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node19420 = (inp[11]) ? node19422 : 16'b0000000011111111;
															assign node19422 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19425 = (inp[10]) ? node19433 : node19426;
													assign node19426 = (inp[7]) ? node19428 : 16'b0000000011111111;
														assign node19428 = (inp[14]) ? node19430 : 16'b0000000011111111;
															assign node19430 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19433 = (inp[14]) ? node19439 : node19434;
														assign node19434 = (inp[11]) ? node19436 : 16'b0000000011111111;
															assign node19436 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19439 = (inp[9]) ? node19441 : 16'b0000000001111111;
															assign node19441 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19444 = (inp[11]) ? node19464 : node19445;
											assign node19445 = (inp[9]) ? node19455 : node19446;
												assign node19446 = (inp[4]) ? 16'b0000000011111111 : node19447;
													assign node19447 = (inp[7]) ? node19449 : 16'b0000000111111111;
														assign node19449 = (inp[10]) ? node19451 : 16'b0000000111111111;
															assign node19451 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19455 = (inp[14]) ? node19459 : node19456;
													assign node19456 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node19459 = (inp[7]) ? 16'b0000000001111111 : node19460;
														assign node19460 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19464 = (inp[9]) ? node19482 : node19465;
												assign node19465 = (inp[14]) ? node19471 : node19466;
													assign node19466 = (inp[4]) ? 16'b0000000001111111 : node19467;
														assign node19467 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19471 = (inp[10]) ? node19475 : node19472;
														assign node19472 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19475 = (inp[7]) ? node19477 : 16'b0000000001111111;
															assign node19477 = (inp[8]) ? 16'b0000000000111111 : node19478;
																assign node19478 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19482 = (inp[10]) ? node19492 : node19483;
													assign node19483 = (inp[7]) ? node19485 : 16'b0000000001111111;
														assign node19485 = (inp[14]) ? node19487 : 16'b0000000001111111;
															assign node19487 = (inp[4]) ? node19489 : 16'b0000000000111111;
																assign node19489 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19492 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node19495 = (inp[11]) ? node19603 : node19496;
									assign node19496 = (inp[5]) ? node19550 : node19497;
										assign node19497 = (inp[2]) ? node19521 : node19498;
											assign node19498 = (inp[7]) ? node19510 : node19499;
												assign node19499 = (inp[8]) ? node19503 : node19500;
													assign node19500 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node19503 = (inp[10]) ? node19505 : 16'b0000001111111111;
														assign node19505 = (inp[14]) ? 16'b0000000111111111 : node19506;
															assign node19506 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19510 = (inp[10]) ? node19516 : node19511;
													assign node19511 = (inp[8]) ? 16'b0000000111111111 : node19512;
														assign node19512 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19516 = (inp[14]) ? node19518 : 16'b0000000011111111;
														assign node19518 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node19521 = (inp[14]) ? node19533 : node19522;
												assign node19522 = (inp[10]) ? node19524 : 16'b0000000111111111;
													assign node19524 = (inp[4]) ? 16'b0000000001111111 : node19525;
														assign node19525 = (inp[8]) ? 16'b0000000011111111 : node19526;
															assign node19526 = (inp[9]) ? node19528 : 16'b0000000111111111;
																assign node19528 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19533 = (inp[4]) ? node19541 : node19534;
													assign node19534 = (inp[9]) ? node19538 : node19535;
														assign node19535 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19538 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19541 = (inp[8]) ? 16'b0000000001111111 : node19542;
														assign node19542 = (inp[10]) ? node19544 : 16'b0000000011111111;
															assign node19544 = (inp[7]) ? 16'b0000000001111111 : node19545;
																assign node19545 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19550 = (inp[7]) ? node19580 : node19551;
											assign node19551 = (inp[8]) ? node19565 : node19552;
												assign node19552 = (inp[10]) ? node19558 : node19553;
													assign node19553 = (inp[14]) ? 16'b0000000111111111 : node19554;
														assign node19554 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19558 = (inp[9]) ? node19560 : 16'b0000000111111111;
														assign node19560 = (inp[2]) ? node19562 : 16'b0000000011111111;
															assign node19562 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19565 = (inp[2]) ? node19575 : node19566;
													assign node19566 = (inp[4]) ? node19568 : 16'b0000000011111111;
														assign node19568 = (inp[9]) ? 16'b0000000001111111 : node19569;
															assign node19569 = (inp[10]) ? node19571 : 16'b0000000011111111;
																assign node19571 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19575 = (inp[10]) ? node19577 : 16'b0000000011111111;
														assign node19577 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19580 = (inp[10]) ? node19594 : node19581;
												assign node19581 = (inp[14]) ? node19583 : 16'b0000000011111111;
													assign node19583 = (inp[8]) ? node19591 : node19584;
														assign node19584 = (inp[9]) ? 16'b0000000001111111 : node19585;
															assign node19585 = (inp[4]) ? node19587 : 16'b0000000011111111;
																assign node19587 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19591 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node19594 = (inp[14]) ? 16'b0000000000111111 : node19595;
													assign node19595 = (inp[2]) ? node19597 : 16'b0000000001111111;
														assign node19597 = (inp[9]) ? 16'b0000000000111111 : node19598;
															assign node19598 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node19603 = (inp[7]) ? node19667 : node19604;
										assign node19604 = (inp[9]) ? node19626 : node19605;
											assign node19605 = (inp[10]) ? node19617 : node19606;
												assign node19606 = (inp[2]) ? node19612 : node19607;
													assign node19607 = (inp[5]) ? 16'b0000000111111111 : node19608;
														assign node19608 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19612 = (inp[14]) ? 16'b0000000011111111 : node19613;
														assign node19613 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19617 = (inp[5]) ? node19619 : 16'b0000000011111111;
													assign node19619 = (inp[2]) ? node19623 : node19620;
														assign node19620 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19623 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19626 = (inp[5]) ? node19650 : node19627;
												assign node19627 = (inp[4]) ? node19641 : node19628;
													assign node19628 = (inp[8]) ? node19636 : node19629;
														assign node19629 = (inp[10]) ? node19631 : 16'b0000000111111111;
															assign node19631 = (inp[2]) ? node19633 : 16'b0000000011111111;
																assign node19633 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19636 = (inp[10]) ? 16'b0000000001111111 : node19637;
															assign node19637 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19641 = (inp[10]) ? 16'b0000000000111111 : node19642;
														assign node19642 = (inp[14]) ? node19644 : 16'b0000000011111111;
															assign node19644 = (inp[8]) ? node19646 : 16'b0000000001111111;
																assign node19646 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19650 = (inp[14]) ? node19658 : node19651;
													assign node19651 = (inp[8]) ? node19655 : node19652;
														assign node19652 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19655 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19658 = (inp[4]) ? 16'b0000000000111111 : node19659;
														assign node19659 = (inp[10]) ? node19661 : 16'b0000000000111111;
															assign node19661 = (inp[8]) ? node19663 : 16'b0000000000111111;
																assign node19663 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19667 = (inp[10]) ? node19699 : node19668;
											assign node19668 = (inp[9]) ? node19684 : node19669;
												assign node19669 = (inp[8]) ? node19679 : node19670;
													assign node19670 = (inp[2]) ? node19672 : 16'b0000000011111111;
														assign node19672 = (inp[4]) ? node19674 : 16'b0000000011111111;
															assign node19674 = (inp[5]) ? 16'b0000000001111111 : node19675;
																assign node19675 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19679 = (inp[2]) ? 16'b0000000000111111 : node19680;
														assign node19680 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19684 = (inp[4]) ? node19686 : 16'b0000000001111111;
													assign node19686 = (inp[2]) ? node19694 : node19687;
														assign node19687 = (inp[5]) ? 16'b0000000000111111 : node19688;
															assign node19688 = (inp[14]) ? node19690 : 16'b0000000001111111;
																assign node19690 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19694 = (inp[8]) ? node19696 : 16'b0000000000111111;
															assign node19696 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node19699 = (inp[8]) ? node19707 : node19700;
												assign node19700 = (inp[4]) ? node19704 : node19701;
													assign node19701 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19704 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node19707 = (inp[9]) ? node19713 : node19708;
													assign node19708 = (inp[14]) ? node19710 : 16'b0000000000111111;
														assign node19710 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node19713 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node19716 = (inp[7]) ? node20232 : node19717;
							assign node19717 = (inp[2]) ? node19983 : node19718;
								assign node19718 = (inp[12]) ? node19860 : node19719;
									assign node19719 = (inp[4]) ? node19787 : node19720;
										assign node19720 = (inp[8]) ? node19752 : node19721;
											assign node19721 = (inp[9]) ? node19737 : node19722;
												assign node19722 = (inp[5]) ? node19732 : node19723;
													assign node19723 = (inp[10]) ? 16'b0000011111111111 : node19724;
														assign node19724 = (inp[11]) ? node19726 : 16'b0000111111111111;
															assign node19726 = (inp[14]) ? 16'b0000001111111111 : node19727;
																assign node19727 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node19732 = (inp[10]) ? 16'b0000001111111111 : node19733;
														assign node19733 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19737 = (inp[5]) ? node19749 : node19738;
													assign node19738 = (inp[11]) ? node19746 : node19739;
														assign node19739 = (inp[10]) ? 16'b0000001111111111 : node19740;
															assign node19740 = (inp[15]) ? node19742 : 16'b0000011111111111;
																assign node19742 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19746 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19749 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node19752 = (inp[11]) ? node19766 : node19753;
												assign node19753 = (inp[14]) ? node19757 : node19754;
													assign node19754 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19757 = (inp[15]) ? node19763 : node19758;
														assign node19758 = (inp[10]) ? 16'b0000000111111111 : node19759;
															assign node19759 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19763 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19766 = (inp[9]) ? node19778 : node19767;
													assign node19767 = (inp[15]) ? node19773 : node19768;
														assign node19768 = (inp[14]) ? 16'b0000000111111111 : node19769;
															assign node19769 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19773 = (inp[10]) ? node19775 : 16'b0000000111111111;
															assign node19775 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19778 = (inp[5]) ? node19784 : node19779;
														assign node19779 = (inp[10]) ? 16'b0000000011111111 : node19780;
															assign node19780 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19784 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19787 = (inp[9]) ? node19829 : node19788;
											assign node19788 = (inp[10]) ? node19806 : node19789;
												assign node19789 = (inp[15]) ? node19799 : node19790;
													assign node19790 = (inp[14]) ? node19794 : node19791;
														assign node19791 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19794 = (inp[5]) ? 16'b0000000011111111 : node19795;
															assign node19795 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19799 = (inp[5]) ? 16'b0000000111111111 : node19800;
														assign node19800 = (inp[14]) ? 16'b0000000111111111 : node19801;
															assign node19801 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19806 = (inp[15]) ? node19820 : node19807;
													assign node19807 = (inp[8]) ? node19813 : node19808;
														assign node19808 = (inp[14]) ? 16'b0000000111111111 : node19809;
															assign node19809 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19813 = (inp[5]) ? 16'b0000000011111111 : node19814;
															assign node19814 = (inp[11]) ? node19816 : 16'b0000001111111111;
																assign node19816 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19820 = (inp[5]) ? node19826 : node19821;
														assign node19821 = (inp[11]) ? 16'b0000000011111111 : node19822;
															assign node19822 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19826 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node19829 = (inp[11]) ? node19845 : node19830;
												assign node19830 = (inp[5]) ? node19838 : node19831;
													assign node19831 = (inp[15]) ? 16'b0000000111111111 : node19832;
														assign node19832 = (inp[10]) ? node19834 : 16'b0000011111111111;
															assign node19834 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19838 = (inp[8]) ? node19842 : node19839;
														assign node19839 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19842 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19845 = (inp[15]) ? node19853 : node19846;
													assign node19846 = (inp[14]) ? node19848 : 16'b0000000111111111;
														assign node19848 = (inp[5]) ? 16'b0000000001111111 : node19849;
															assign node19849 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19853 = (inp[10]) ? node19855 : 16'b0000000011111111;
														assign node19855 = (inp[14]) ? 16'b0000000000111111 : node19856;
															assign node19856 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node19860 = (inp[9]) ? node19920 : node19861;
										assign node19861 = (inp[5]) ? node19897 : node19862;
											assign node19862 = (inp[10]) ? node19880 : node19863;
												assign node19863 = (inp[15]) ? node19871 : node19864;
													assign node19864 = (inp[8]) ? node19868 : node19865;
														assign node19865 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19868 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19871 = (inp[4]) ? node19877 : node19872;
														assign node19872 = (inp[14]) ? 16'b0000000111111111 : node19873;
															assign node19873 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19877 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19880 = (inp[4]) ? node19894 : node19881;
													assign node19881 = (inp[14]) ? node19887 : node19882;
														assign node19882 = (inp[8]) ? 16'b0000000111111111 : node19883;
															assign node19883 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19887 = (inp[15]) ? 16'b0000000011111111 : node19888;
															assign node19888 = (inp[8]) ? node19890 : 16'b0000000111111111;
																assign node19890 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19894 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19897 = (inp[14]) ? node19909 : node19898;
												assign node19898 = (inp[15]) ? node19900 : 16'b0000000111111111;
													assign node19900 = (inp[4]) ? node19904 : node19901;
														assign node19901 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19904 = (inp[10]) ? node19906 : 16'b0000000011111111;
															assign node19906 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19909 = (inp[8]) ? node19911 : 16'b0000000111111111;
													assign node19911 = (inp[15]) ? 16'b0000000001111111 : node19912;
														assign node19912 = (inp[4]) ? node19914 : 16'b0000000111111111;
															assign node19914 = (inp[11]) ? 16'b0000000001111111 : node19915;
																assign node19915 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19920 = (inp[8]) ? node19956 : node19921;
											assign node19921 = (inp[5]) ? node19937 : node19922;
												assign node19922 = (inp[14]) ? node19928 : node19923;
													assign node19923 = (inp[11]) ? node19925 : 16'b0000000111111111;
														assign node19925 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19928 = (inp[10]) ? node19934 : node19929;
														assign node19929 = (inp[4]) ? 16'b0000000011111111 : node19930;
															assign node19930 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19934 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19937 = (inp[4]) ? node19951 : node19938;
													assign node19938 = (inp[15]) ? node19944 : node19939;
														assign node19939 = (inp[10]) ? 16'b0000000011111111 : node19940;
															assign node19940 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19944 = (inp[10]) ? node19946 : 16'b0000000011111111;
															assign node19946 = (inp[11]) ? 16'b0000000001111111 : node19947;
																assign node19947 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19951 = (inp[11]) ? node19953 : 16'b0000000001111111;
														assign node19953 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node19956 = (inp[10]) ? node19970 : node19957;
												assign node19957 = (inp[15]) ? node19961 : node19958;
													assign node19958 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19961 = (inp[14]) ? node19967 : node19962;
														assign node19962 = (inp[11]) ? node19964 : 16'b0000000011111111;
															assign node19964 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19967 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19970 = (inp[15]) ? node19974 : node19971;
													assign node19971 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19974 = (inp[4]) ? node19976 : 16'b0000000000111111;
														assign node19976 = (inp[11]) ? node19978 : 16'b0000000000111111;
															assign node19978 = (inp[14]) ? node19980 : 16'b0000000000011111;
																assign node19980 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node19983 = (inp[11]) ? node20093 : node19984;
									assign node19984 = (inp[9]) ? node20042 : node19985;
										assign node19985 = (inp[12]) ? node20017 : node19986;
											assign node19986 = (inp[15]) ? node20002 : node19987;
												assign node19987 = (inp[4]) ? node19993 : node19988;
													assign node19988 = (inp[8]) ? node19990 : 16'b0000001111111111;
														assign node19990 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19993 = (inp[8]) ? node19999 : node19994;
														assign node19994 = (inp[10]) ? 16'b0000000111111111 : node19995;
															assign node19995 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19999 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20002 = (inp[4]) ? node20008 : node20003;
													assign node20003 = (inp[14]) ? node20005 : 16'b0000001111111111;
														assign node20005 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20008 = (inp[5]) ? 16'b0000000011111111 : node20009;
														assign node20009 = (inp[8]) ? node20011 : 16'b0000000111111111;
															assign node20011 = (inp[14]) ? 16'b0000000011111111 : node20012;
																assign node20012 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node20017 = (inp[10]) ? node20029 : node20018;
												assign node20018 = (inp[4]) ? node20024 : node20019;
													assign node20019 = (inp[5]) ? node20021 : 16'b0000001111111111;
														assign node20021 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20024 = (inp[15]) ? 16'b0000000001111111 : node20025;
														assign node20025 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20029 = (inp[4]) ? node20039 : node20030;
													assign node20030 = (inp[15]) ? node20036 : node20031;
														assign node20031 = (inp[5]) ? 16'b0000000011111111 : node20032;
															assign node20032 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20036 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20039 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node20042 = (inp[4]) ? node20068 : node20043;
											assign node20043 = (inp[12]) ? node20057 : node20044;
												assign node20044 = (inp[14]) ? node20052 : node20045;
													assign node20045 = (inp[10]) ? node20047 : 16'b0000011111111111;
														assign node20047 = (inp[8]) ? 16'b0000000111111111 : node20048;
															assign node20048 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20052 = (inp[10]) ? 16'b0000000011111111 : node20053;
														assign node20053 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20057 = (inp[10]) ? 16'b0000000001111111 : node20058;
													assign node20058 = (inp[15]) ? node20062 : node20059;
														assign node20059 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20062 = (inp[14]) ? 16'b0000000001111111 : node20063;
															assign node20063 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20068 = (inp[12]) ? node20086 : node20069;
												assign node20069 = (inp[14]) ? node20075 : node20070;
													assign node20070 = (inp[10]) ? node20072 : 16'b0000000011111111;
														assign node20072 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20075 = (inp[8]) ? node20083 : node20076;
														assign node20076 = (inp[15]) ? 16'b0000000001111111 : node20077;
															assign node20077 = (inp[10]) ? node20079 : 16'b0000000011111111;
																assign node20079 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20083 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node20086 = (inp[10]) ? node20088 : 16'b0000000001111111;
													assign node20088 = (inp[5]) ? 16'b0000000000011111 : node20089;
														assign node20089 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node20093 = (inp[14]) ? node20151 : node20094;
										assign node20094 = (inp[5]) ? node20126 : node20095;
											assign node20095 = (inp[10]) ? node20115 : node20096;
												assign node20096 = (inp[8]) ? node20104 : node20097;
													assign node20097 = (inp[4]) ? 16'b0000000111111111 : node20098;
														assign node20098 = (inp[9]) ? 16'b0000000111111111 : node20099;
															assign node20099 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20104 = (inp[4]) ? node20110 : node20105;
														assign node20105 = (inp[12]) ? 16'b0000000011111111 : node20106;
															assign node20106 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20110 = (inp[15]) ? node20112 : 16'b0000000011111111;
															assign node20112 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20115 = (inp[12]) ? node20121 : node20116;
													assign node20116 = (inp[9]) ? 16'b0000000011111111 : node20117;
														assign node20117 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node20121 = (inp[15]) ? 16'b0000000001111111 : node20122;
														assign node20122 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20126 = (inp[9]) ? node20140 : node20127;
												assign node20127 = (inp[15]) ? node20135 : node20128;
													assign node20128 = (inp[10]) ? node20132 : node20129;
														assign node20129 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20132 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20135 = (inp[12]) ? node20137 : 16'b0000000001111111;
														assign node20137 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20140 = (inp[10]) ? node20146 : node20141;
													assign node20141 = (inp[4]) ? node20143 : 16'b0000000011111111;
														assign node20143 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20146 = (inp[4]) ? 16'b0000000000011111 : node20147;
														assign node20147 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20151 = (inp[12]) ? node20195 : node20152;
											assign node20152 = (inp[9]) ? node20172 : node20153;
												assign node20153 = (inp[4]) ? node20159 : node20154;
													assign node20154 = (inp[15]) ? 16'b0000000011111111 : node20155;
														assign node20155 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20159 = (inp[10]) ? node20169 : node20160;
														assign node20160 = (inp[15]) ? node20164 : node20161;
															assign node20161 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node20164 = (inp[8]) ? 16'b0000000001111111 : node20165;
																assign node20165 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20169 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20172 = (inp[10]) ? node20184 : node20173;
													assign node20173 = (inp[15]) ? node20177 : node20174;
														assign node20174 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20177 = (inp[4]) ? 16'b0000000000111111 : node20178;
															assign node20178 = (inp[5]) ? node20180 : 16'b0000000001111111;
																assign node20180 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20184 = (inp[5]) ? node20190 : node20185;
														assign node20185 = (inp[8]) ? 16'b0000000000111111 : node20186;
															assign node20186 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node20190 = (inp[4]) ? node20192 : 16'b0000000000111111;
															assign node20192 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node20195 = (inp[10]) ? node20215 : node20196;
												assign node20196 = (inp[4]) ? node20206 : node20197;
													assign node20197 = (inp[8]) ? node20199 : 16'b0000000011111111;
														assign node20199 = (inp[15]) ? 16'b0000000000111111 : node20200;
															assign node20200 = (inp[9]) ? node20202 : 16'b0000000001111111;
																assign node20202 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20206 = (inp[5]) ? node20212 : node20207;
														assign node20207 = (inp[15]) ? 16'b0000000000111111 : node20208;
															assign node20208 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20212 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20215 = (inp[15]) ? node20227 : node20216;
													assign node20216 = (inp[9]) ? node20220 : node20217;
														assign node20217 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20220 = (inp[5]) ? node20222 : 16'b0000000000111111;
															assign node20222 = (inp[8]) ? 16'b0000000000011111 : node20223;
																assign node20223 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20227 = (inp[9]) ? 16'b0000000000011111 : node20228;
														assign node20228 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node20232 = (inp[4]) ? node20510 : node20233;
								assign node20233 = (inp[14]) ? node20361 : node20234;
									assign node20234 = (inp[5]) ? node20304 : node20235;
										assign node20235 = (inp[12]) ? node20273 : node20236;
											assign node20236 = (inp[8]) ? node20254 : node20237;
												assign node20237 = (inp[2]) ? node20243 : node20238;
													assign node20238 = (inp[10]) ? 16'b0000001111111111 : node20239;
														assign node20239 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20243 = (inp[15]) ? node20251 : node20244;
														assign node20244 = (inp[9]) ? node20246 : 16'b0000001111111111;
															assign node20246 = (inp[11]) ? 16'b0000000111111111 : node20247;
																assign node20247 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20251 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20254 = (inp[9]) ? node20266 : node20255;
													assign node20255 = (inp[11]) ? node20261 : node20256;
														assign node20256 = (inp[15]) ? 16'b0000000111111111 : node20257;
															assign node20257 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20261 = (inp[10]) ? node20263 : 16'b0000000111111111;
															assign node20263 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20266 = (inp[2]) ? node20270 : node20267;
														assign node20267 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20270 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20273 = (inp[2]) ? node20289 : node20274;
												assign node20274 = (inp[10]) ? node20278 : node20275;
													assign node20275 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20278 = (inp[11]) ? node20284 : node20279;
														assign node20279 = (inp[8]) ? node20281 : 16'b0000001111111111;
															assign node20281 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20284 = (inp[8]) ? node20286 : 16'b0000000011111111;
															assign node20286 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20289 = (inp[9]) ? node20297 : node20290;
													assign node20290 = (inp[8]) ? node20294 : node20291;
														assign node20291 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20294 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20297 = (inp[8]) ? node20301 : node20298;
														assign node20298 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20301 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20304 = (inp[11]) ? node20332 : node20305;
											assign node20305 = (inp[2]) ? node20315 : node20306;
												assign node20306 = (inp[15]) ? node20308 : 16'b0000000111111111;
													assign node20308 = (inp[10]) ? 16'b0000000011111111 : node20309;
														assign node20309 = (inp[8]) ? node20311 : 16'b0000000111111111;
															assign node20311 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node20315 = (inp[9]) ? node20323 : node20316;
													assign node20316 = (inp[12]) ? node20320 : node20317;
														assign node20317 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20320 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20323 = (inp[12]) ? node20329 : node20324;
														assign node20324 = (inp[8]) ? 16'b0000000001111111 : node20325;
															assign node20325 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20329 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node20332 = (inp[10]) ? node20346 : node20333;
												assign node20333 = (inp[8]) ? node20339 : node20334;
													assign node20334 = (inp[12]) ? node20336 : 16'b0000000011111111;
														assign node20336 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node20339 = (inp[9]) ? node20343 : node20340;
														assign node20340 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20343 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20346 = (inp[9]) ? node20356 : node20347;
													assign node20347 = (inp[12]) ? node20353 : node20348;
														assign node20348 = (inp[15]) ? 16'b0000000001111111 : node20349;
															assign node20349 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20353 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20356 = (inp[8]) ? node20358 : 16'b0000000000111111;
														assign node20358 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node20361 = (inp[11]) ? node20439 : node20362;
										assign node20362 = (inp[8]) ? node20408 : node20363;
											assign node20363 = (inp[10]) ? node20393 : node20364;
												assign node20364 = (inp[5]) ? node20380 : node20365;
													assign node20365 = (inp[12]) ? node20375 : node20366;
														assign node20366 = (inp[15]) ? node20370 : node20367;
															assign node20367 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node20370 = (inp[2]) ? 16'b0000000111111111 : node20371;
																assign node20371 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20375 = (inp[9]) ? node20377 : 16'b0000000111111111;
															assign node20377 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20380 = (inp[2]) ? node20388 : node20381;
														assign node20381 = (inp[12]) ? 16'b0000000011111111 : node20382;
															assign node20382 = (inp[9]) ? node20384 : 16'b0000000111111111;
																assign node20384 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20388 = (inp[9]) ? 16'b0000000001111111 : node20389;
															assign node20389 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20393 = (inp[9]) ? node20399 : node20394;
													assign node20394 = (inp[2]) ? 16'b0000000011111111 : node20395;
														assign node20395 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node20399 = (inp[12]) ? node20403 : node20400;
														assign node20400 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20403 = (inp[15]) ? 16'b0000000000111111 : node20404;
															assign node20404 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20408 = (inp[15]) ? node20422 : node20409;
												assign node20409 = (inp[10]) ? node20415 : node20410;
													assign node20410 = (inp[5]) ? node20412 : 16'b0000000011111111;
														assign node20412 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20415 = (inp[9]) ? node20419 : node20416;
														assign node20416 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20419 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20422 = (inp[2]) ? node20428 : node20423;
													assign node20423 = (inp[9]) ? node20425 : 16'b0000000011111111;
														assign node20425 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20428 = (inp[9]) ? node20432 : node20429;
														assign node20429 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20432 = (inp[12]) ? node20434 : 16'b0000000000111111;
															assign node20434 = (inp[5]) ? node20436 : 16'b0000000000011111;
																assign node20436 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node20439 = (inp[12]) ? node20471 : node20440;
											assign node20440 = (inp[2]) ? node20454 : node20441;
												assign node20441 = (inp[15]) ? node20447 : node20442;
													assign node20442 = (inp[10]) ? 16'b0000000011111111 : node20443;
														assign node20443 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20447 = (inp[8]) ? node20451 : node20448;
														assign node20448 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20451 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20454 = (inp[10]) ? node20460 : node20455;
													assign node20455 = (inp[9]) ? 16'b0000000001111111 : node20456;
														assign node20456 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20460 = (inp[5]) ? node20462 : 16'b0000000001111111;
														assign node20462 = (inp[8]) ? node20468 : node20463;
															assign node20463 = (inp[9]) ? 16'b0000000000111111 : node20464;
																assign node20464 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node20468 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node20471 = (inp[5]) ? node20491 : node20472;
												assign node20472 = (inp[8]) ? node20486 : node20473;
													assign node20473 = (inp[9]) ? node20477 : node20474;
														assign node20474 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20477 = (inp[15]) ? node20483 : node20478;
															assign node20478 = (inp[2]) ? node20480 : 16'b0000000001111111;
																assign node20480 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node20483 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20486 = (inp[15]) ? 16'b0000000000111111 : node20487;
														assign node20487 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20491 = (inp[2]) ? node20501 : node20492;
													assign node20492 = (inp[10]) ? node20498 : node20493;
														assign node20493 = (inp[15]) ? 16'b0000000000111111 : node20494;
															assign node20494 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20498 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20501 = (inp[10]) ? node20505 : node20502;
														assign node20502 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node20505 = (inp[9]) ? node20507 : 16'b0000000000011111;
															assign node20507 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node20510 = (inp[2]) ? node20630 : node20511;
									assign node20511 = (inp[12]) ? node20575 : node20512;
										assign node20512 = (inp[15]) ? node20536 : node20513;
											assign node20513 = (inp[9]) ? node20521 : node20514;
												assign node20514 = (inp[14]) ? node20516 : 16'b0000000111111111;
													assign node20516 = (inp[8]) ? 16'b0000000001111111 : node20517;
														assign node20517 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20521 = (inp[10]) ? node20531 : node20522;
													assign node20522 = (inp[14]) ? node20526 : node20523;
														assign node20523 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20526 = (inp[11]) ? node20528 : 16'b0000000011111111;
															assign node20528 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20531 = (inp[14]) ? 16'b0000000000111111 : node20532;
														assign node20532 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20536 = (inp[11]) ? node20554 : node20537;
												assign node20537 = (inp[14]) ? node20549 : node20538;
													assign node20538 = (inp[8]) ? node20542 : node20539;
														assign node20539 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20542 = (inp[5]) ? node20544 : 16'b0000000011111111;
															assign node20544 = (inp[10]) ? 16'b0000000001111111 : node20545;
																assign node20545 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20549 = (inp[10]) ? node20551 : 16'b0000000001111111;
														assign node20551 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20554 = (inp[10]) ? node20564 : node20555;
													assign node20555 = (inp[9]) ? node20557 : 16'b0000000011111111;
														assign node20557 = (inp[5]) ? 16'b0000000000111111 : node20558;
															assign node20558 = (inp[14]) ? node20560 : 16'b0000000001111111;
																assign node20560 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20564 = (inp[5]) ? node20568 : node20565;
														assign node20565 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20568 = (inp[14]) ? 16'b0000000000011111 : node20569;
															assign node20569 = (inp[9]) ? node20571 : 16'b0000000000111111;
																assign node20571 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node20575 = (inp[5]) ? node20603 : node20576;
											assign node20576 = (inp[8]) ? node20586 : node20577;
												assign node20577 = (inp[15]) ? node20581 : node20578;
													assign node20578 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20581 = (inp[11]) ? 16'b0000000001111111 : node20582;
														assign node20582 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20586 = (inp[11]) ? node20594 : node20587;
													assign node20587 = (inp[14]) ? node20589 : 16'b0000000001111111;
														assign node20589 = (inp[9]) ? node20591 : 16'b0000000001111111;
															assign node20591 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20594 = (inp[14]) ? node20600 : node20595;
														assign node20595 = (inp[9]) ? node20597 : 16'b0000000001111111;
															assign node20597 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20600 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node20603 = (inp[8]) ? node20615 : node20604;
												assign node20604 = (inp[10]) ? node20606 : 16'b0000000001111111;
													assign node20606 = (inp[11]) ? node20612 : node20607;
														assign node20607 = (inp[15]) ? node20609 : 16'b0000000001111111;
															assign node20609 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20612 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20615 = (inp[10]) ? node20623 : node20616;
													assign node20616 = (inp[9]) ? node20618 : 16'b0000000000111111;
														assign node20618 = (inp[14]) ? node20620 : 16'b0000000000111111;
															assign node20620 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20623 = (inp[14]) ? 16'b0000000000011111 : node20624;
														assign node20624 = (inp[15]) ? 16'b0000000000011111 : node20625;
															assign node20625 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node20630 = (inp[5]) ? node20694 : node20631;
										assign node20631 = (inp[9]) ? node20663 : node20632;
											assign node20632 = (inp[14]) ? node20650 : node20633;
												assign node20633 = (inp[12]) ? node20643 : node20634;
													assign node20634 = (inp[8]) ? node20638 : node20635;
														assign node20635 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20638 = (inp[15]) ? 16'b0000000000111111 : node20639;
															assign node20639 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20643 = (inp[10]) ? node20647 : node20644;
														assign node20644 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20647 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20650 = (inp[8]) ? node20658 : node20651;
													assign node20651 = (inp[11]) ? node20655 : node20652;
														assign node20652 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20655 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20658 = (inp[10]) ? node20660 : 16'b0000000000111111;
														assign node20660 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node20663 = (inp[10]) ? node20683 : node20664;
												assign node20664 = (inp[11]) ? node20674 : node20665;
													assign node20665 = (inp[8]) ? node20667 : 16'b0000000111111111;
														assign node20667 = (inp[15]) ? node20669 : 16'b0000000001111111;
															assign node20669 = (inp[14]) ? 16'b0000000000111111 : node20670;
																assign node20670 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20674 = (inp[15]) ? node20676 : 16'b0000000000111111;
														assign node20676 = (inp[12]) ? 16'b0000000000011111 : node20677;
															assign node20677 = (inp[8]) ? node20679 : 16'b0000000000111111;
																assign node20679 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20683 = (inp[11]) ? node20691 : node20684;
													assign node20684 = (inp[8]) ? node20686 : 16'b0000000000111111;
														assign node20686 = (inp[12]) ? 16'b0000000000011111 : node20687;
															assign node20687 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20691 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node20694 = (inp[11]) ? node20732 : node20695;
											assign node20695 = (inp[10]) ? node20711 : node20696;
												assign node20696 = (inp[15]) ? node20702 : node20697;
													assign node20697 = (inp[8]) ? node20699 : 16'b0000000001111111;
														assign node20699 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20702 = (inp[14]) ? node20704 : 16'b0000000001111111;
														assign node20704 = (inp[12]) ? node20706 : 16'b0000000000111111;
															assign node20706 = (inp[8]) ? 16'b0000000000011111 : node20707;
																assign node20707 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20711 = (inp[9]) ? node20723 : node20712;
													assign node20712 = (inp[8]) ? node20716 : node20713;
														assign node20713 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20716 = (inp[15]) ? 16'b0000000000011111 : node20717;
															assign node20717 = (inp[14]) ? node20719 : 16'b0000000000111111;
																assign node20719 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20723 = (inp[15]) ? node20729 : node20724;
														assign node20724 = (inp[12]) ? 16'b0000000000011111 : node20725;
															assign node20725 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node20729 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node20732 = (inp[8]) ? node20750 : node20733;
												assign node20733 = (inp[15]) ? node20745 : node20734;
													assign node20734 = (inp[12]) ? node20738 : node20735;
														assign node20735 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20738 = (inp[9]) ? node20740 : 16'b0000000000111111;
															assign node20740 = (inp[14]) ? node20742 : 16'b0000000000011111;
																assign node20742 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node20745 = (inp[12]) ? node20747 : 16'b0000000000011111;
														assign node20747 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node20750 = (inp[10]) ? node20758 : node20751;
													assign node20751 = (inp[12]) ? node20753 : 16'b0000000000011111;
														assign node20753 = (inp[9]) ? node20755 : 16'b0000000000011111;
															assign node20755 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node20758 = (inp[15]) ? node20764 : node20759;
														assign node20759 = (inp[12]) ? node20761 : 16'b0000000000001111;
															assign node20761 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node20764 = (inp[12]) ? node20766 : 16'b0000000000000111;
															assign node20766 = (inp[14]) ? node20768 : 16'b0000000000000111;
																assign node20768 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
				assign node20771 = (inp[5]) ? node22889 : node20772;
					assign node20772 = (inp[11]) ? node21786 : node20773;
						assign node20773 = (inp[9]) ? node21307 : node20774;
							assign node20774 = (inp[8]) ? node21060 : node20775;
								assign node20775 = (inp[4]) ? node20917 : node20776;
									assign node20776 = (inp[1]) ? node20842 : node20777;
										assign node20777 = (inp[13]) ? node20817 : node20778;
											assign node20778 = (inp[14]) ? node20802 : node20779;
												assign node20779 = (inp[15]) ? node20793 : node20780;
													assign node20780 = (inp[12]) ? node20786 : node20781;
														assign node20781 = (inp[10]) ? 16'b0000111111111111 : node20782;
															assign node20782 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node20786 = (inp[10]) ? node20788 : 16'b0000111111111111;
															assign node20788 = (inp[7]) ? node20790 : 16'b0000011111111111;
																assign node20790 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20793 = (inp[12]) ? node20799 : node20794;
														assign node20794 = (inp[7]) ? 16'b0000011111111111 : node20795;
															assign node20795 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node20799 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node20802 = (inp[2]) ? node20808 : node20803;
													assign node20803 = (inp[12]) ? node20805 : 16'b0000011111111111;
														assign node20805 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20808 = (inp[15]) ? node20814 : node20809;
														assign node20809 = (inp[10]) ? node20811 : 16'b0000011111111111;
															assign node20811 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20814 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node20817 = (inp[14]) ? node20833 : node20818;
												assign node20818 = (inp[2]) ? node20826 : node20819;
													assign node20819 = (inp[7]) ? node20821 : 16'b0000011111111111;
														assign node20821 = (inp[10]) ? node20823 : 16'b0000011111111111;
															assign node20823 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20826 = (inp[10]) ? 16'b0000001111111111 : node20827;
														assign node20827 = (inp[12]) ? 16'b0000001111111111 : node20828;
															assign node20828 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node20833 = (inp[15]) ? node20835 : 16'b0000001111111111;
													assign node20835 = (inp[2]) ? 16'b0000000011111111 : node20836;
														assign node20836 = (inp[10]) ? node20838 : 16'b0000000111111111;
															assign node20838 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node20842 = (inp[7]) ? node20892 : node20843;
											assign node20843 = (inp[13]) ? node20869 : node20844;
												assign node20844 = (inp[12]) ? node20856 : node20845;
													assign node20845 = (inp[14]) ? node20851 : node20846;
														assign node20846 = (inp[10]) ? node20848 : 16'b0000111111111111;
															assign node20848 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20851 = (inp[10]) ? 16'b0000001111111111 : node20852;
															assign node20852 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20856 = (inp[14]) ? node20862 : node20857;
														assign node20857 = (inp[15]) ? 16'b0000001111111111 : node20858;
															assign node20858 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20862 = (inp[10]) ? node20864 : 16'b0000001111111111;
															assign node20864 = (inp[15]) ? 16'b0000000111111111 : node20865;
																assign node20865 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node20869 = (inp[2]) ? node20879 : node20870;
													assign node20870 = (inp[15]) ? node20874 : node20871;
														assign node20871 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20874 = (inp[14]) ? node20876 : 16'b0000001111111111;
															assign node20876 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20879 = (inp[15]) ? node20885 : node20880;
														assign node20880 = (inp[10]) ? node20882 : 16'b0000001111111111;
															assign node20882 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node20885 = (inp[10]) ? node20887 : 16'b0000000111111111;
															assign node20887 = (inp[14]) ? node20889 : 16'b0000000111111111;
																assign node20889 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20892 = (inp[15]) ? node20904 : node20893;
												assign node20893 = (inp[2]) ? node20899 : node20894;
													assign node20894 = (inp[12]) ? 16'b0000001111111111 : node20895;
														assign node20895 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20899 = (inp[10]) ? 16'b0000000011111111 : node20900;
														assign node20900 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node20904 = (inp[14]) ? node20912 : node20905;
													assign node20905 = (inp[10]) ? node20909 : node20906;
														assign node20906 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20909 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20912 = (inp[2]) ? node20914 : 16'b0000000011111111;
														assign node20914 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node20917 = (inp[13]) ? node20995 : node20918;
										assign node20918 = (inp[15]) ? node20950 : node20919;
											assign node20919 = (inp[12]) ? node20933 : node20920;
												assign node20920 = (inp[10]) ? node20930 : node20921;
													assign node20921 = (inp[2]) ? node20923 : 16'b0000111111111111;
														assign node20923 = (inp[14]) ? 16'b0000001111111111 : node20924;
															assign node20924 = (inp[7]) ? 16'b0000011111111111 : node20925;
																assign node20925 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node20930 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node20933 = (inp[14]) ? node20943 : node20934;
													assign node20934 = (inp[7]) ? node20940 : node20935;
														assign node20935 = (inp[2]) ? node20937 : 16'b0000001111111111;
															assign node20937 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20940 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20943 = (inp[2]) ? 16'b0000000111111111 : node20944;
														assign node20944 = (inp[1]) ? node20946 : 16'b0000001111111111;
															assign node20946 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node20950 = (inp[12]) ? node20976 : node20951;
												assign node20951 = (inp[1]) ? node20965 : node20952;
													assign node20952 = (inp[10]) ? node20958 : node20953;
														assign node20953 = (inp[2]) ? 16'b0000001111111111 : node20954;
															assign node20954 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node20958 = (inp[14]) ? 16'b0000000111111111 : node20959;
															assign node20959 = (inp[2]) ? node20961 : 16'b0000001111111111;
																assign node20961 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20965 = (inp[10]) ? node20969 : node20966;
														assign node20966 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20969 = (inp[14]) ? 16'b0000000111111111 : node20970;
															assign node20970 = (inp[7]) ? 16'b0000000111111111 : node20971;
																assign node20971 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node20976 = (inp[1]) ? node20986 : node20977;
													assign node20977 = (inp[7]) ? node20983 : node20978;
														assign node20978 = (inp[2]) ? 16'b0000000111111111 : node20979;
															assign node20979 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20983 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node20986 = (inp[2]) ? node20988 : 16'b0000000111111111;
														assign node20988 = (inp[7]) ? node20990 : 16'b0000000011111111;
															assign node20990 = (inp[10]) ? node20992 : 16'b0000000001111111;
																assign node20992 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20995 = (inp[10]) ? node21019 : node20996;
											assign node20996 = (inp[15]) ? node21008 : node20997;
												assign node20997 = (inp[12]) ? 16'b0000000111111111 : node20998;
													assign node20998 = (inp[14]) ? node21004 : node20999;
														assign node20999 = (inp[7]) ? 16'b0000001111111111 : node21000;
															assign node21000 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node21004 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21008 = (inp[7]) ? node21010 : 16'b0000001111111111;
													assign node21010 = (inp[1]) ? node21012 : 16'b0000000111111111;
														assign node21012 = (inp[14]) ? 16'b0000000001111111 : node21013;
															assign node21013 = (inp[2]) ? 16'b0000000011111111 : node21014;
																assign node21014 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node21019 = (inp[1]) ? node21037 : node21020;
												assign node21020 = (inp[7]) ? node21028 : node21021;
													assign node21021 = (inp[15]) ? node21025 : node21022;
														assign node21022 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21025 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21028 = (inp[14]) ? node21032 : node21029;
														assign node21029 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node21032 = (inp[2]) ? 16'b0000000001111111 : node21033;
															assign node21033 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21037 = (inp[15]) ? node21045 : node21038;
													assign node21038 = (inp[7]) ? 16'b0000000001111111 : node21039;
														assign node21039 = (inp[12]) ? 16'b0000000011111111 : node21040;
															assign node21040 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21045 = (inp[2]) ? node21053 : node21046;
														assign node21046 = (inp[7]) ? 16'b0000000001111111 : node21047;
															assign node21047 = (inp[14]) ? node21049 : 16'b0000000011111111;
																assign node21049 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21053 = (inp[12]) ? node21055 : 16'b0000000001111111;
															assign node21055 = (inp[14]) ? 16'b0000000000111111 : node21056;
																assign node21056 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node21060 = (inp[7]) ? node21170 : node21061;
									assign node21061 = (inp[1]) ? node21111 : node21062;
										assign node21062 = (inp[14]) ? node21090 : node21063;
											assign node21063 = (inp[4]) ? node21077 : node21064;
												assign node21064 = (inp[10]) ? node21072 : node21065;
													assign node21065 = (inp[15]) ? 16'b0000011111111111 : node21066;
														assign node21066 = (inp[12]) ? node21068 : 16'b0000111111111111;
															assign node21068 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node21072 = (inp[12]) ? node21074 : 16'b0000011111111111;
														assign node21074 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21077 = (inp[13]) ? node21085 : node21078;
													assign node21078 = (inp[15]) ? node21082 : node21079;
														assign node21079 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21082 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21085 = (inp[15]) ? node21087 : 16'b0000000111111111;
														assign node21087 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node21090 = (inp[4]) ? node21100 : node21091;
												assign node21091 = (inp[13]) ? 16'b0000000111111111 : node21092;
													assign node21092 = (inp[12]) ? node21094 : 16'b0000001111111111;
														assign node21094 = (inp[10]) ? node21096 : 16'b0000001111111111;
															assign node21096 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21100 = (inp[10]) ? node21106 : node21101;
													assign node21101 = (inp[15]) ? 16'b0000000111111111 : node21102;
														assign node21102 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21106 = (inp[13]) ? 16'b0000000001111111 : node21107;
														assign node21107 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node21111 = (inp[4]) ? node21141 : node21112;
											assign node21112 = (inp[15]) ? node21134 : node21113;
												assign node21113 = (inp[12]) ? node21125 : node21114;
													assign node21114 = (inp[10]) ? node21122 : node21115;
														assign node21115 = (inp[13]) ? 16'b0000001111111111 : node21116;
															assign node21116 = (inp[14]) ? node21118 : 16'b0000011111111111;
																assign node21118 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21122 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21125 = (inp[2]) ? node21131 : node21126;
														assign node21126 = (inp[14]) ? 16'b0000000111111111 : node21127;
															assign node21127 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21131 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21134 = (inp[10]) ? node21136 : 16'b0000000111111111;
													assign node21136 = (inp[13]) ? node21138 : 16'b0000000111111111;
														assign node21138 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21141 = (inp[10]) ? node21155 : node21142;
												assign node21142 = (inp[12]) ? node21144 : 16'b0000000111111111;
													assign node21144 = (inp[2]) ? node21152 : node21145;
														assign node21145 = (inp[13]) ? node21147 : 16'b0000000111111111;
															assign node21147 = (inp[14]) ? 16'b0000000011111111 : node21148;
																assign node21148 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21152 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node21155 = (inp[12]) ? node21165 : node21156;
													assign node21156 = (inp[14]) ? node21160 : node21157;
														assign node21157 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21160 = (inp[13]) ? 16'b0000000001111111 : node21161;
															assign node21161 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21165 = (inp[13]) ? 16'b0000000000111111 : node21166;
														assign node21166 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node21170 = (inp[13]) ? node21246 : node21171;
										assign node21171 = (inp[14]) ? node21205 : node21172;
											assign node21172 = (inp[2]) ? node21188 : node21173;
												assign node21173 = (inp[10]) ? node21181 : node21174;
													assign node21174 = (inp[12]) ? node21178 : node21175;
														assign node21175 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21178 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21181 = (inp[12]) ? 16'b0000000111111111 : node21182;
														assign node21182 = (inp[4]) ? 16'b0000000111111111 : node21183;
															assign node21183 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21188 = (inp[1]) ? node21196 : node21189;
													assign node21189 = (inp[15]) ? node21191 : 16'b0000000111111111;
														assign node21191 = (inp[4]) ? 16'b0000000111111111 : node21192;
															assign node21192 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21196 = (inp[12]) ? node21198 : 16'b0000000111111111;
														assign node21198 = (inp[15]) ? node21200 : 16'b0000000011111111;
															assign node21200 = (inp[10]) ? node21202 : 16'b0000000011111111;
																assign node21202 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21205 = (inp[15]) ? node21219 : node21206;
												assign node21206 = (inp[1]) ? node21214 : node21207;
													assign node21207 = (inp[10]) ? node21211 : node21208;
														assign node21208 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21211 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21214 = (inp[2]) ? 16'b0000000001111111 : node21215;
														assign node21215 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21219 = (inp[12]) ? node21235 : node21220;
													assign node21220 = (inp[10]) ? node21226 : node21221;
														assign node21221 = (inp[2]) ? 16'b0000000011111111 : node21222;
															assign node21222 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21226 = (inp[4]) ? 16'b0000000001111111 : node21227;
															assign node21227 = (inp[2]) ? node21231 : node21228;
																assign node21228 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node21231 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21235 = (inp[1]) ? node21241 : node21236;
														assign node21236 = (inp[10]) ? node21238 : 16'b0000000011111111;
															assign node21238 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21241 = (inp[4]) ? 16'b0000000000111111 : node21242;
															assign node21242 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21246 = (inp[10]) ? node21280 : node21247;
											assign node21247 = (inp[2]) ? node21263 : node21248;
												assign node21248 = (inp[12]) ? node21256 : node21249;
													assign node21249 = (inp[4]) ? node21253 : node21250;
														assign node21250 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21253 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21256 = (inp[1]) ? node21260 : node21257;
														assign node21257 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21260 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21263 = (inp[12]) ? node21275 : node21264;
													assign node21264 = (inp[1]) ? node21270 : node21265;
														assign node21265 = (inp[15]) ? 16'b0000000011111111 : node21266;
															assign node21266 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21270 = (inp[15]) ? 16'b0000000001111111 : node21271;
															assign node21271 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21275 = (inp[14]) ? node21277 : 16'b0000000001111111;
														assign node21277 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21280 = (inp[4]) ? node21294 : node21281;
												assign node21281 = (inp[15]) ? 16'b0000000001111111 : node21282;
													assign node21282 = (inp[1]) ? node21288 : node21283;
														assign node21283 = (inp[2]) ? node21285 : 16'b0000000011111111;
															assign node21285 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21288 = (inp[2]) ? 16'b0000000001111111 : node21289;
															assign node21289 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21294 = (inp[15]) ? node21298 : node21295;
													assign node21295 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21298 = (inp[12]) ? node21300 : 16'b0000000000111111;
														assign node21300 = (inp[14]) ? node21302 : 16'b0000000000111111;
															assign node21302 = (inp[2]) ? node21304 : 16'b0000000000011111;
																assign node21304 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node21307 = (inp[15]) ? node21539 : node21308;
								assign node21308 = (inp[12]) ? node21414 : node21309;
									assign node21309 = (inp[1]) ? node21357 : node21310;
										assign node21310 = (inp[8]) ? node21336 : node21311;
											assign node21311 = (inp[14]) ? node21319 : node21312;
												assign node21312 = (inp[7]) ? node21314 : 16'b0000011111111111;
													assign node21314 = (inp[4]) ? 16'b0000001111111111 : node21315;
														assign node21315 = (inp[13]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node21319 = (inp[2]) ? 16'b0000000111111111 : node21320;
													assign node21320 = (inp[7]) ? node21328 : node21321;
														assign node21321 = (inp[13]) ? node21323 : 16'b0000011111111111;
															assign node21323 = (inp[10]) ? 16'b0000001111111111 : node21324;
																assign node21324 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21328 = (inp[10]) ? 16'b0000000111111111 : node21329;
															assign node21329 = (inp[4]) ? node21331 : 16'b0000001111111111;
																assign node21331 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node21336 = (inp[14]) ? node21344 : node21337;
												assign node21337 = (inp[10]) ? node21339 : 16'b0000001111111111;
													assign node21339 = (inp[2]) ? 16'b0000000111111111 : node21340;
														assign node21340 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21344 = (inp[7]) ? node21354 : node21345;
													assign node21345 = (inp[2]) ? node21351 : node21346;
														assign node21346 = (inp[4]) ? node21348 : 16'b0000001111111111;
															assign node21348 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node21351 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21354 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21357 = (inp[7]) ? node21385 : node21358;
											assign node21358 = (inp[14]) ? node21376 : node21359;
												assign node21359 = (inp[2]) ? node21367 : node21360;
													assign node21360 = (inp[13]) ? node21364 : node21361;
														assign node21361 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21364 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21367 = (inp[10]) ? node21369 : 16'b0000001111111111;
														assign node21369 = (inp[8]) ? 16'b0000000011111111 : node21370;
															assign node21370 = (inp[13]) ? node21372 : 16'b0000000111111111;
																assign node21372 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21376 = (inp[8]) ? node21378 : 16'b0000000111111111;
													assign node21378 = (inp[2]) ? 16'b0000000011111111 : node21379;
														assign node21379 = (inp[10]) ? node21381 : 16'b0000000111111111;
															assign node21381 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node21385 = (inp[13]) ? node21403 : node21386;
												assign node21386 = (inp[2]) ? node21394 : node21387;
													assign node21387 = (inp[8]) ? node21389 : 16'b0000001111111111;
														assign node21389 = (inp[14]) ? node21391 : 16'b0000000111111111;
															assign node21391 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21394 = (inp[10]) ? node21396 : 16'b0000000001111111;
														assign node21396 = (inp[14]) ? 16'b0000000011111111 : node21397;
															assign node21397 = (inp[4]) ? 16'b0000000011111111 : node21398;
																assign node21398 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21403 = (inp[10]) ? node21409 : node21404;
													assign node21404 = (inp[2]) ? 16'b0000000001111111 : node21405;
														assign node21405 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21409 = (inp[8]) ? node21411 : 16'b0000000001111111;
														assign node21411 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node21414 = (inp[14]) ? node21470 : node21415;
										assign node21415 = (inp[1]) ? node21441 : node21416;
											assign node21416 = (inp[10]) ? node21428 : node21417;
												assign node21417 = (inp[7]) ? node21421 : node21418;
													assign node21418 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node21421 = (inp[8]) ? 16'b0000000111111111 : node21422;
														assign node21422 = (inp[4]) ? node21424 : 16'b0000001111111111;
															assign node21424 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21428 = (inp[7]) ? node21432 : node21429;
													assign node21429 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21432 = (inp[2]) ? node21438 : node21433;
														assign node21433 = (inp[4]) ? 16'b0000000011111111 : node21434;
															assign node21434 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21438 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21441 = (inp[8]) ? node21457 : node21442;
												assign node21442 = (inp[7]) ? node21448 : node21443;
													assign node21443 = (inp[10]) ? node21445 : 16'b0000000111111111;
														assign node21445 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21448 = (inp[4]) ? node21452 : node21449;
														assign node21449 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21452 = (inp[13]) ? node21454 : 16'b0000000011111111;
															assign node21454 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21457 = (inp[7]) ? node21465 : node21458;
													assign node21458 = (inp[4]) ? node21462 : node21459;
														assign node21459 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21462 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21465 = (inp[13]) ? node21467 : 16'b0000000001111111;
														assign node21467 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21470 = (inp[7]) ? node21502 : node21471;
											assign node21471 = (inp[8]) ? node21487 : node21472;
												assign node21472 = (inp[1]) ? 16'b0000000011111111 : node21473;
													assign node21473 = (inp[4]) ? node21479 : node21474;
														assign node21474 = (inp[2]) ? 16'b0000000111111111 : node21475;
															assign node21475 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21479 = (inp[13]) ? node21481 : 16'b0000000111111111;
															assign node21481 = (inp[2]) ? 16'b0000000011111111 : node21482;
																assign node21482 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21487 = (inp[2]) ? node21495 : node21488;
													assign node21488 = (inp[1]) ? node21490 : 16'b0000000011111111;
														assign node21490 = (inp[10]) ? node21492 : 16'b0000000011111111;
															assign node21492 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21495 = (inp[13]) ? 16'b0000000000011111 : node21496;
														assign node21496 = (inp[4]) ? 16'b0000000001111111 : node21497;
															assign node21497 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21502 = (inp[2]) ? node21518 : node21503;
												assign node21503 = (inp[13]) ? node21511 : node21504;
													assign node21504 = (inp[8]) ? node21508 : node21505;
														assign node21505 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21508 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21511 = (inp[8]) ? node21515 : node21512;
														assign node21512 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21515 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21518 = (inp[4]) ? node21528 : node21519;
													assign node21519 = (inp[1]) ? node21525 : node21520;
														assign node21520 = (inp[8]) ? 16'b0000000001111111 : node21521;
															assign node21521 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21525 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21528 = (inp[8]) ? node21536 : node21529;
														assign node21529 = (inp[10]) ? node21531 : 16'b0000000001111111;
															assign node21531 = (inp[13]) ? 16'b0000000000111111 : node21532;
																assign node21532 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21536 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
								assign node21539 = (inp[14]) ? node21657 : node21540;
									assign node21540 = (inp[10]) ? node21592 : node21541;
										assign node21541 = (inp[2]) ? node21573 : node21542;
											assign node21542 = (inp[12]) ? node21556 : node21543;
												assign node21543 = (inp[13]) ? node21551 : node21544;
													assign node21544 = (inp[8]) ? node21546 : 16'b0000011111111111;
														assign node21546 = (inp[7]) ? node21548 : 16'b0000011111111111;
															assign node21548 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21551 = (inp[1]) ? 16'b0000000011111111 : node21552;
														assign node21552 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21556 = (inp[4]) ? node21562 : node21557;
													assign node21557 = (inp[8]) ? 16'b0000000111111111 : node21558;
														assign node21558 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21562 = (inp[7]) ? node21570 : node21563;
														assign node21563 = (inp[8]) ? node21565 : 16'b0000000111111111;
															assign node21565 = (inp[1]) ? 16'b0000000011111111 : node21566;
																assign node21566 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21570 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21573 = (inp[8]) ? node21585 : node21574;
												assign node21574 = (inp[7]) ? 16'b0000000011111111 : node21575;
													assign node21575 = (inp[4]) ? node21577 : 16'b0000000111111111;
														assign node21577 = (inp[13]) ? 16'b0000000011111111 : node21578;
															assign node21578 = (inp[1]) ? node21580 : 16'b0000000111111111;
																assign node21580 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21585 = (inp[12]) ? node21589 : node21586;
													assign node21586 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21589 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node21592 = (inp[2]) ? node21634 : node21593;
											assign node21593 = (inp[12]) ? node21615 : node21594;
												assign node21594 = (inp[8]) ? node21602 : node21595;
													assign node21595 = (inp[7]) ? 16'b0000000011111111 : node21596;
														assign node21596 = (inp[13]) ? node21598 : 16'b0000001111111111;
															assign node21598 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21602 = (inp[13]) ? node21610 : node21603;
														assign node21603 = (inp[1]) ? node21605 : 16'b0000000111111111;
															assign node21605 = (inp[4]) ? 16'b0000000001111111 : node21606;
																assign node21606 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21610 = (inp[1]) ? node21612 : 16'b0000000011111111;
															assign node21612 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21615 = (inp[13]) ? node21629 : node21616;
													assign node21616 = (inp[7]) ? node21624 : node21617;
														assign node21617 = (inp[8]) ? 16'b0000000011111111 : node21618;
															assign node21618 = (inp[1]) ? node21620 : 16'b0000000111111111;
																assign node21620 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21624 = (inp[1]) ? node21626 : 16'b0000000011111111;
															assign node21626 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21629 = (inp[4]) ? node21631 : 16'b0000000001111111;
														assign node21631 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21634 = (inp[1]) ? node21642 : node21635;
												assign node21635 = (inp[7]) ? 16'b0000000001111111 : node21636;
													assign node21636 = (inp[12]) ? 16'b0000000001111111 : node21637;
														assign node21637 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21642 = (inp[8]) ? node21652 : node21643;
													assign node21643 = (inp[4]) ? node21645 : 16'b0000000001111111;
														assign node21645 = (inp[13]) ? 16'b0000000000111111 : node21646;
															assign node21646 = (inp[7]) ? node21648 : 16'b0000000001111111;
																assign node21648 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21652 = (inp[13]) ? node21654 : 16'b0000000001111111;
														assign node21654 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node21657 = (inp[1]) ? node21735 : node21658;
										assign node21658 = (inp[10]) ? node21694 : node21659;
											assign node21659 = (inp[12]) ? node21679 : node21660;
												assign node21660 = (inp[7]) ? node21672 : node21661;
													assign node21661 = (inp[4]) ? node21665 : node21662;
														assign node21662 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21665 = (inp[2]) ? node21667 : 16'b0000000111111111;
															assign node21667 = (inp[13]) ? 16'b0000000011111111 : node21668;
																assign node21668 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21672 = (inp[8]) ? 16'b0000000001111111 : node21673;
														assign node21673 = (inp[13]) ? 16'b0000000011111111 : node21674;
															assign node21674 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21679 = (inp[2]) ? node21685 : node21680;
													assign node21680 = (inp[7]) ? 16'b0000000001111111 : node21681;
														assign node21681 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21685 = (inp[8]) ? node21691 : node21686;
														assign node21686 = (inp[13]) ? 16'b0000000001111111 : node21687;
															assign node21687 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21691 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node21694 = (inp[12]) ? node21720 : node21695;
												assign node21695 = (inp[4]) ? node21707 : node21696;
													assign node21696 = (inp[8]) ? node21700 : node21697;
														assign node21697 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21700 = (inp[13]) ? node21702 : 16'b0000000011111111;
															assign node21702 = (inp[2]) ? 16'b0000000001111111 : node21703;
																assign node21703 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21707 = (inp[13]) ? node21711 : node21708;
														assign node21708 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21711 = (inp[8]) ? node21717 : node21712;
															assign node21712 = (inp[7]) ? node21714 : 16'b0000000001111111;
																assign node21714 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node21717 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21720 = (inp[2]) ? node21726 : node21721;
													assign node21721 = (inp[7]) ? 16'b0000000001111111 : node21722;
														assign node21722 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21726 = (inp[7]) ? node21732 : node21727;
														assign node21727 = (inp[4]) ? 16'b0000000000111111 : node21728;
															assign node21728 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21732 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21735 = (inp[12]) ? node21765 : node21736;
											assign node21736 = (inp[4]) ? node21748 : node21737;
												assign node21737 = (inp[10]) ? node21743 : node21738;
													assign node21738 = (inp[8]) ? node21740 : 16'b0000001111111111;
														assign node21740 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21743 = (inp[2]) ? node21745 : 16'b0000000001111111;
														assign node21745 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21748 = (inp[7]) ? node21758 : node21749;
													assign node21749 = (inp[10]) ? node21753 : node21750;
														assign node21750 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21753 = (inp[8]) ? 16'b0000000001111111 : node21754;
															assign node21754 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21758 = (inp[8]) ? node21762 : node21759;
														assign node21759 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node21762 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21765 = (inp[8]) ? node21775 : node21766;
												assign node21766 = (inp[13]) ? node21772 : node21767;
													assign node21767 = (inp[10]) ? node21769 : 16'b0000000011111111;
														assign node21769 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21772 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21775 = (inp[7]) ? node21781 : node21776;
													assign node21776 = (inp[13]) ? node21778 : 16'b0000000000111111;
														assign node21778 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21781 = (inp[4]) ? node21783 : 16'b0000000000111111;
														assign node21783 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node21786 = (inp[10]) ? node22326 : node21787;
							assign node21787 = (inp[13]) ? node22061 : node21788;
								assign node21788 = (inp[8]) ? node21922 : node21789;
									assign node21789 = (inp[7]) ? node21863 : node21790;
										assign node21790 = (inp[9]) ? node21836 : node21791;
											assign node21791 = (inp[4]) ? node21815 : node21792;
												assign node21792 = (inp[1]) ? node21800 : node21793;
													assign node21793 = (inp[12]) ? node21795 : 16'b0000111111111111;
														assign node21795 = (inp[2]) ? 16'b0000011111111111 : node21796;
															assign node21796 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node21800 = (inp[2]) ? node21808 : node21801;
														assign node21801 = (inp[12]) ? 16'b0000011111111111 : node21802;
															assign node21802 = (inp[14]) ? 16'b0000011111111111 : node21803;
																assign node21803 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node21808 = (inp[15]) ? 16'b0000001111111111 : node21809;
															assign node21809 = (inp[14]) ? 16'b0000001111111111 : node21810;
																assign node21810 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21815 = (inp[2]) ? node21827 : node21816;
													assign node21816 = (inp[14]) ? node21824 : node21817;
														assign node21817 = (inp[1]) ? node21819 : 16'b0000011111111111;
															assign node21819 = (inp[15]) ? 16'b0000001111111111 : node21820;
																assign node21820 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21824 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21827 = (inp[1]) ? 16'b0000000111111111 : node21828;
														assign node21828 = (inp[12]) ? node21830 : 16'b0000011111111111;
															assign node21830 = (inp[14]) ? 16'b0000000111111111 : node21831;
																assign node21831 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node21836 = (inp[15]) ? node21850 : node21837;
												assign node21837 = (inp[1]) ? node21841 : node21838;
													assign node21838 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node21841 = (inp[14]) ? 16'b0000000111111111 : node21842;
														assign node21842 = (inp[4]) ? node21846 : node21843;
															assign node21843 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node21846 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21850 = (inp[1]) ? node21860 : node21851;
													assign node21851 = (inp[14]) ? 16'b0000000111111111 : node21852;
														assign node21852 = (inp[12]) ? node21854 : 16'b0000011111111111;
															assign node21854 = (inp[4]) ? 16'b0000000111111111 : node21855;
																assign node21855 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21860 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node21863 = (inp[4]) ? node21895 : node21864;
											assign node21864 = (inp[14]) ? node21876 : node21865;
												assign node21865 = (inp[2]) ? node21867 : 16'b0000001111111111;
													assign node21867 = (inp[1]) ? 16'b0000000111111111 : node21868;
														assign node21868 = (inp[12]) ? node21872 : node21869;
															assign node21869 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node21872 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21876 = (inp[9]) ? node21884 : node21877;
													assign node21877 = (inp[15]) ? node21881 : node21878;
														assign node21878 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21881 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21884 = (inp[1]) ? node21892 : node21885;
														assign node21885 = (inp[12]) ? node21887 : 16'b0000000111111111;
															assign node21887 = (inp[15]) ? 16'b0000000011111111 : node21888;
																assign node21888 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21892 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21895 = (inp[1]) ? node21911 : node21896;
												assign node21896 = (inp[12]) ? node21904 : node21897;
													assign node21897 = (inp[2]) ? node21899 : 16'b0000001111111111;
														assign node21899 = (inp[9]) ? 16'b0000000111111111 : node21900;
															assign node21900 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21904 = (inp[15]) ? node21908 : node21905;
														assign node21905 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21908 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node21911 = (inp[12]) ? node21917 : node21912;
													assign node21912 = (inp[15]) ? node21914 : 16'b0000000011111111;
														assign node21914 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21917 = (inp[2]) ? 16'b0000000000111111 : node21918;
														assign node21918 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node21922 = (inp[7]) ? node21986 : node21923;
										assign node21923 = (inp[9]) ? node21959 : node21924;
											assign node21924 = (inp[1]) ? node21944 : node21925;
												assign node21925 = (inp[15]) ? node21939 : node21926;
													assign node21926 = (inp[12]) ? node21930 : node21927;
														assign node21927 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node21930 = (inp[2]) ? node21936 : node21931;
															assign node21931 = (inp[4]) ? 16'b0000001111111111 : node21932;
																assign node21932 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node21936 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21939 = (inp[14]) ? node21941 : 16'b0000000011111111;
														assign node21941 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21944 = (inp[12]) ? node21952 : node21945;
													assign node21945 = (inp[2]) ? node21949 : node21946;
														assign node21946 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21949 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node21952 = (inp[4]) ? 16'b0000000011111111 : node21953;
														assign node21953 = (inp[15]) ? node21955 : 16'b0000000111111111;
															assign node21955 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21959 = (inp[12]) ? node21971 : node21960;
												assign node21960 = (inp[4]) ? node21966 : node21961;
													assign node21961 = (inp[2]) ? node21963 : 16'b0000000111111111;
														assign node21963 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21966 = (inp[2]) ? 16'b0000000011111111 : node21967;
														assign node21967 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21971 = (inp[15]) ? node21979 : node21972;
													assign node21972 = (inp[4]) ? 16'b0000000011111111 : node21973;
														assign node21973 = (inp[1]) ? 16'b0000000011111111 : node21974;
															assign node21974 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node21979 = (inp[1]) ? 16'b0000000000111111 : node21980;
														assign node21980 = (inp[14]) ? 16'b0000000001111111 : node21981;
															assign node21981 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21986 = (inp[15]) ? node22020 : node21987;
											assign node21987 = (inp[4]) ? node22005 : node21988;
												assign node21988 = (inp[2]) ? node21998 : node21989;
													assign node21989 = (inp[9]) ? node21993 : node21990;
														assign node21990 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node21993 = (inp[14]) ? node21995 : 16'b0000000111111111;
															assign node21995 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21998 = (inp[9]) ? 16'b0000000011111111 : node21999;
														assign node21999 = (inp[1]) ? 16'b0000000011111111 : node22000;
															assign node22000 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22005 = (inp[1]) ? node22015 : node22006;
													assign node22006 = (inp[2]) ? node22012 : node22007;
														assign node22007 = (inp[12]) ? 16'b0000000011111111 : node22008;
															assign node22008 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22012 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22015 = (inp[14]) ? node22017 : 16'b0000000011111111;
														assign node22017 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22020 = (inp[12]) ? node22034 : node22021;
												assign node22021 = (inp[14]) ? node22029 : node22022;
													assign node22022 = (inp[1]) ? 16'b0000000011111111 : node22023;
														assign node22023 = (inp[2]) ? node22025 : 16'b0000000111111111;
															assign node22025 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22029 = (inp[4]) ? node22031 : 16'b0000000111111111;
														assign node22031 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22034 = (inp[1]) ? node22050 : node22035;
													assign node22035 = (inp[4]) ? node22041 : node22036;
														assign node22036 = (inp[14]) ? 16'b0000000001111111 : node22037;
															assign node22037 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22041 = (inp[9]) ? 16'b0000000000111111 : node22042;
															assign node22042 = (inp[14]) ? node22046 : node22043;
																assign node22043 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
																assign node22046 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22050 = (inp[4]) ? node22054 : node22051;
														assign node22051 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22054 = (inp[9]) ? 16'b0000000000011111 : node22055;
															assign node22055 = (inp[2]) ? node22057 : 16'b0000000000111111;
																assign node22057 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node22061 = (inp[4]) ? node22183 : node22062;
									assign node22062 = (inp[12]) ? node22126 : node22063;
										assign node22063 = (inp[2]) ? node22095 : node22064;
											assign node22064 = (inp[14]) ? node22076 : node22065;
												assign node22065 = (inp[9]) ? 16'b0000000111111111 : node22066;
													assign node22066 = (inp[8]) ? node22072 : node22067;
														assign node22067 = (inp[1]) ? 16'b0000011111111111 : node22068;
															assign node22068 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node22072 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node22076 = (inp[15]) ? node22086 : node22077;
													assign node22077 = (inp[8]) ? node22083 : node22078;
														assign node22078 = (inp[9]) ? node22080 : 16'b0000001111111111;
															assign node22080 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22083 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node22086 = (inp[1]) ? node22090 : node22087;
														assign node22087 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22090 = (inp[9]) ? node22092 : 16'b0000000011111111;
															assign node22092 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22095 = (inp[8]) ? node22107 : node22096;
												assign node22096 = (inp[14]) ? 16'b0000000011111111 : node22097;
													assign node22097 = (inp[9]) ? node22101 : node22098;
														assign node22098 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22101 = (inp[15]) ? 16'b0000000011111111 : node22102;
															assign node22102 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22107 = (inp[1]) ? node22119 : node22108;
													assign node22108 = (inp[14]) ? node22114 : node22109;
														assign node22109 = (inp[15]) ? node22111 : 16'b0000001111111111;
															assign node22111 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22114 = (inp[15]) ? 16'b0000000001111111 : node22115;
															assign node22115 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22119 = (inp[9]) ? node22123 : node22120;
														assign node22120 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22123 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node22126 = (inp[9]) ? node22154 : node22127;
											assign node22127 = (inp[15]) ? node22139 : node22128;
												assign node22128 = (inp[8]) ? node22134 : node22129;
													assign node22129 = (inp[7]) ? 16'b0000000111111111 : node22130;
														assign node22130 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22134 = (inp[2]) ? 16'b0000000011111111 : node22135;
														assign node22135 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22139 = (inp[2]) ? node22149 : node22140;
													assign node22140 = (inp[14]) ? node22142 : 16'b0000000111111111;
														assign node22142 = (inp[1]) ? 16'b0000000001111111 : node22143;
															assign node22143 = (inp[8]) ? 16'b0000000001111111 : node22144;
																assign node22144 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22149 = (inp[1]) ? node22151 : 16'b0000000001111111;
														assign node22151 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22154 = (inp[15]) ? node22164 : node22155;
												assign node22155 = (inp[2]) ? node22157 : 16'b0000000011111111;
													assign node22157 = (inp[14]) ? node22161 : node22158;
														assign node22158 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22161 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22164 = (inp[2]) ? node22174 : node22165;
													assign node22165 = (inp[1]) ? node22169 : node22166;
														assign node22166 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22169 = (inp[14]) ? 16'b0000000000111111 : node22170;
															assign node22170 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22174 = (inp[7]) ? node22178 : node22175;
														assign node22175 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22178 = (inp[1]) ? 16'b0000000000011111 : node22179;
															assign node22179 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22183 = (inp[1]) ? node22241 : node22184;
										assign node22184 = (inp[7]) ? node22212 : node22185;
											assign node22185 = (inp[8]) ? node22201 : node22186;
												assign node22186 = (inp[9]) ? node22194 : node22187;
													assign node22187 = (inp[15]) ? node22189 : 16'b0000001111111111;
														assign node22189 = (inp[12]) ? 16'b0000000111111111 : node22190;
															assign node22190 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22194 = (inp[2]) ? 16'b0000000011111111 : node22195;
														assign node22195 = (inp[12]) ? node22197 : 16'b0000000111111111;
															assign node22197 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22201 = (inp[9]) ? 16'b0000000001111111 : node22202;
													assign node22202 = (inp[12]) ? node22206 : node22203;
														assign node22203 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22206 = (inp[2]) ? 16'b0000000001111111 : node22207;
															assign node22207 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22212 = (inp[2]) ? node22230 : node22213;
												assign node22213 = (inp[9]) ? node22227 : node22214;
													assign node22214 = (inp[8]) ? node22220 : node22215;
														assign node22215 = (inp[14]) ? node22217 : 16'b0000000111111111;
															assign node22217 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22220 = (inp[15]) ? 16'b0000000001111111 : node22221;
															assign node22221 = (inp[12]) ? node22223 : 16'b0000000011111111;
																assign node22223 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22227 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22230 = (inp[12]) ? node22238 : node22231;
													assign node22231 = (inp[8]) ? node22235 : node22232;
														assign node22232 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22235 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22238 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22241 = (inp[12]) ? node22281 : node22242;
											assign node22242 = (inp[8]) ? node22266 : node22243;
												assign node22243 = (inp[9]) ? node22257 : node22244;
													assign node22244 = (inp[15]) ? node22250 : node22245;
														assign node22245 = (inp[2]) ? node22247 : 16'b0000000111111111;
															assign node22247 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22250 = (inp[7]) ? 16'b0000000001111111 : node22251;
															assign node22251 = (inp[14]) ? node22253 : 16'b0000000011111111;
																assign node22253 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22257 = (inp[15]) ? node22261 : node22258;
														assign node22258 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22261 = (inp[7]) ? 16'b0000000000111111 : node22262;
															assign node22262 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22266 = (inp[2]) ? node22268 : 16'b0000000001111111;
													assign node22268 = (inp[14]) ? node22278 : node22269;
														assign node22269 = (inp[15]) ? node22273 : node22270;
															assign node22270 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node22273 = (inp[9]) ? 16'b0000000000111111 : node22274;
																assign node22274 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22278 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22281 = (inp[15]) ? node22299 : node22282;
												assign node22282 = (inp[7]) ? 16'b0000000000111111 : node22283;
													assign node22283 = (inp[2]) ? node22287 : node22284;
														assign node22284 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22287 = (inp[9]) ? node22293 : node22288;
															assign node22288 = (inp[8]) ? node22290 : 16'b0000000001111111;
																assign node22290 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node22293 = (inp[14]) ? 16'b0000000000111111 : node22294;
																assign node22294 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22299 = (inp[2]) ? node22315 : node22300;
													assign node22300 = (inp[7]) ? node22310 : node22301;
														assign node22301 = (inp[8]) ? node22305 : node22302;
															assign node22302 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node22305 = (inp[14]) ? 16'b0000000000111111 : node22306;
																assign node22306 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22310 = (inp[8]) ? 16'b0000000000011111 : node22311;
															assign node22311 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22315 = (inp[9]) ? node22319 : node22316;
														assign node22316 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22319 = (inp[8]) ? node22321 : 16'b0000000000011111;
															assign node22321 = (inp[14]) ? 16'b0000000000001111 : node22322;
																assign node22322 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node22326 = (inp[14]) ? node22590 : node22327;
								assign node22327 = (inp[2]) ? node22453 : node22328;
									assign node22328 = (inp[7]) ? node22388 : node22329;
										assign node22329 = (inp[4]) ? node22365 : node22330;
											assign node22330 = (inp[9]) ? node22348 : node22331;
												assign node22331 = (inp[15]) ? node22341 : node22332;
													assign node22332 = (inp[13]) ? node22336 : node22333;
														assign node22333 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node22336 = (inp[12]) ? node22338 : 16'b0000001111111111;
															assign node22338 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22341 = (inp[13]) ? node22345 : node22342;
														assign node22342 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22345 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22348 = (inp[15]) ? node22360 : node22349;
													assign node22349 = (inp[8]) ? node22357 : node22350;
														assign node22350 = (inp[12]) ? 16'b0000000111111111 : node22351;
															assign node22351 = (inp[1]) ? node22353 : 16'b0000001111111111;
																assign node22353 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22357 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22360 = (inp[13]) ? 16'b0000000011111111 : node22361;
														assign node22361 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node22365 = (inp[12]) ? node22377 : node22366;
												assign node22366 = (inp[13]) ? node22368 : 16'b0000000111111111;
													assign node22368 = (inp[8]) ? node22372 : node22369;
														assign node22369 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22372 = (inp[15]) ? node22374 : 16'b0000000011111111;
															assign node22374 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22377 = (inp[13]) ? 16'b0000000001111111 : node22378;
													assign node22378 = (inp[15]) ? node22382 : node22379;
														assign node22379 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22382 = (inp[8]) ? node22384 : 16'b0000000011111111;
															assign node22384 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node22388 = (inp[1]) ? node22430 : node22389;
											assign node22389 = (inp[9]) ? node22413 : node22390;
												assign node22390 = (inp[12]) ? node22400 : node22391;
													assign node22391 = (inp[8]) ? node22397 : node22392;
														assign node22392 = (inp[15]) ? 16'b0000000111111111 : node22393;
															assign node22393 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22397 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node22400 = (inp[8]) ? node22408 : node22401;
														assign node22401 = (inp[15]) ? 16'b0000000011111111 : node22402;
															assign node22402 = (inp[4]) ? node22404 : 16'b0000000111111111;
																assign node22404 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22408 = (inp[15]) ? node22410 : 16'b0000000011111111;
															assign node22410 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22413 = (inp[13]) ? node22421 : node22414;
													assign node22414 = (inp[8]) ? node22418 : node22415;
														assign node22415 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node22418 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22421 = (inp[12]) ? 16'b0000000001111111 : node22422;
														assign node22422 = (inp[8]) ? node22424 : 16'b0000000011111111;
															assign node22424 = (inp[4]) ? 16'b0000000000111111 : node22425;
																assign node22425 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node22430 = (inp[12]) ? node22440 : node22431;
												assign node22431 = (inp[15]) ? 16'b0000000011111111 : node22432;
													assign node22432 = (inp[9]) ? node22436 : node22433;
														assign node22433 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22436 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22440 = (inp[8]) ? node22446 : node22441;
													assign node22441 = (inp[9]) ? node22443 : 16'b0000000001111111;
														assign node22443 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node22446 = (inp[15]) ? node22450 : node22447;
														assign node22447 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node22450 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22453 = (inp[9]) ? node22535 : node22454;
										assign node22454 = (inp[7]) ? node22490 : node22455;
											assign node22455 = (inp[13]) ? node22469 : node22456;
												assign node22456 = (inp[1]) ? node22460 : node22457;
													assign node22457 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22460 = (inp[12]) ? node22466 : node22461;
														assign node22461 = (inp[15]) ? node22463 : 16'b0000000111111111;
															assign node22463 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22466 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22469 = (inp[1]) ? node22479 : node22470;
													assign node22470 = (inp[8]) ? 16'b0000000011111111 : node22471;
														assign node22471 = (inp[4]) ? 16'b0000000011111111 : node22472;
															assign node22472 = (inp[12]) ? node22474 : 16'b0000000111111111;
																assign node22474 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22479 = (inp[8]) ? node22487 : node22480;
														assign node22480 = (inp[4]) ? node22482 : 16'b0000000011111111;
															assign node22482 = (inp[15]) ? 16'b0000000001111111 : node22483;
																assign node22483 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22487 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22490 = (inp[12]) ? node22512 : node22491;
												assign node22491 = (inp[15]) ? node22503 : node22492;
													assign node22492 = (inp[13]) ? node22498 : node22493;
														assign node22493 = (inp[1]) ? 16'b0000000111111111 : node22494;
															assign node22494 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22498 = (inp[8]) ? node22500 : 16'b0000000011111111;
															assign node22500 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22503 = (inp[8]) ? node22507 : node22504;
														assign node22504 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22507 = (inp[13]) ? node22509 : 16'b0000000001111111;
															assign node22509 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22512 = (inp[1]) ? node22520 : node22513;
													assign node22513 = (inp[13]) ? node22515 : 16'b0000000011111111;
														assign node22515 = (inp[15]) ? node22517 : 16'b0000000001111111;
															assign node22517 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22520 = (inp[8]) ? node22528 : node22521;
														assign node22521 = (inp[13]) ? 16'b0000000000111111 : node22522;
															assign node22522 = (inp[15]) ? node22524 : 16'b0000000001111111;
																assign node22524 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22528 = (inp[13]) ? node22530 : 16'b0000000000111111;
															assign node22530 = (inp[4]) ? 16'b0000000000001111 : node22531;
																assign node22531 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22535 = (inp[4]) ? node22563 : node22536;
											assign node22536 = (inp[15]) ? node22546 : node22537;
												assign node22537 = (inp[8]) ? node22539 : 16'b0000000011111111;
													assign node22539 = (inp[12]) ? node22541 : 16'b0000000011111111;
														assign node22541 = (inp[7]) ? 16'b0000000000111111 : node22542;
															assign node22542 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22546 = (inp[1]) ? node22556 : node22547;
													assign node22547 = (inp[12]) ? node22549 : 16'b0000000011111111;
														assign node22549 = (inp[8]) ? 16'b0000000000111111 : node22550;
															assign node22550 = (inp[7]) ? node22552 : 16'b0000000001111111;
																assign node22552 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22556 = (inp[13]) ? node22558 : 16'b0000000001111111;
														assign node22558 = (inp[8]) ? node22560 : 16'b0000000000111111;
															assign node22560 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22563 = (inp[15]) ? node22575 : node22564;
												assign node22564 = (inp[1]) ? node22568 : node22565;
													assign node22565 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22568 = (inp[8]) ? 16'b0000000000001111 : node22569;
														assign node22569 = (inp[7]) ? node22571 : 16'b0000000000111111;
															assign node22571 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22575 = (inp[1]) ? node22583 : node22576;
													assign node22576 = (inp[8]) ? 16'b0000000000011111 : node22577;
														assign node22577 = (inp[7]) ? node22579 : 16'b0000000000111111;
															assign node22579 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22583 = (inp[8]) ? node22585 : 16'b0000000000011111;
														assign node22585 = (inp[12]) ? node22587 : 16'b0000000000011111;
															assign node22587 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node22590 = (inp[9]) ? node22734 : node22591;
									assign node22591 = (inp[4]) ? node22657 : node22592;
										assign node22592 = (inp[1]) ? node22626 : node22593;
											assign node22593 = (inp[13]) ? node22611 : node22594;
												assign node22594 = (inp[7]) ? node22606 : node22595;
													assign node22595 = (inp[12]) ? node22603 : node22596;
														assign node22596 = (inp[8]) ? 16'b0000000111111111 : node22597;
															assign node22597 = (inp[15]) ? 16'b0000000111111111 : node22598;
																assign node22598 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node22603 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node22606 = (inp[8]) ? 16'b0000000011111111 : node22607;
														assign node22607 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node22611 = (inp[2]) ? node22617 : node22612;
													assign node22612 = (inp[15]) ? 16'b0000000011111111 : node22613;
														assign node22613 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22617 = (inp[8]) ? node22623 : node22618;
														assign node22618 = (inp[7]) ? node22620 : 16'b0000000011111111;
															assign node22620 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22623 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22626 = (inp[7]) ? node22644 : node22627;
												assign node22627 = (inp[15]) ? node22633 : node22628;
													assign node22628 = (inp[12]) ? 16'b0000000011111111 : node22629;
														assign node22629 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22633 = (inp[13]) ? node22641 : node22634;
														assign node22634 = (inp[12]) ? 16'b0000000001111111 : node22635;
															assign node22635 = (inp[2]) ? node22637 : 16'b0000000011111111;
																assign node22637 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22641 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node22644 = (inp[15]) ? node22650 : node22645;
													assign node22645 = (inp[13]) ? node22647 : 16'b0000000011111111;
														assign node22647 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22650 = (inp[12]) ? node22652 : 16'b0000000000111111;
														assign node22652 = (inp[8]) ? node22654 : 16'b0000000000111111;
															assign node22654 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22657 = (inp[12]) ? node22699 : node22658;
											assign node22658 = (inp[8]) ? node22680 : node22659;
												assign node22659 = (inp[1]) ? node22667 : node22660;
													assign node22660 = (inp[15]) ? node22664 : node22661;
														assign node22661 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22664 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22667 = (inp[15]) ? node22675 : node22668;
														assign node22668 = (inp[2]) ? node22670 : 16'b0000000011111111;
															assign node22670 = (inp[13]) ? node22672 : 16'b0000000001111111;
																assign node22672 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22675 = (inp[7]) ? 16'b0000000000111111 : node22676;
															assign node22676 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22680 = (inp[7]) ? node22686 : node22681;
													assign node22681 = (inp[2]) ? node22683 : 16'b0000000001111111;
														assign node22683 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22686 = (inp[1]) ? 16'b0000000000111111 : node22687;
														assign node22687 = (inp[2]) ? node22693 : node22688;
															assign node22688 = (inp[13]) ? node22690 : 16'b0000000001111111;
																assign node22690 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node22693 = (inp[15]) ? 16'b0000000000111111 : node22694;
																assign node22694 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22699 = (inp[2]) ? node22721 : node22700;
												assign node22700 = (inp[15]) ? node22708 : node22701;
													assign node22701 = (inp[13]) ? node22703 : 16'b0000000001111111;
														assign node22703 = (inp[1]) ? node22705 : 16'b0000000001111111;
															assign node22705 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22708 = (inp[13]) ? node22714 : node22709;
														assign node22709 = (inp[1]) ? node22711 : 16'b0000000001111111;
															assign node22711 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22714 = (inp[7]) ? node22716 : 16'b0000000000111111;
															assign node22716 = (inp[8]) ? 16'b0000000000011111 : node22717;
																assign node22717 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22721 = (inp[1]) ? node22727 : node22722;
													assign node22722 = (inp[15]) ? 16'b0000000000111111 : node22723;
														assign node22723 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22727 = (inp[7]) ? 16'b0000000000001111 : node22728;
														assign node22728 = (inp[13]) ? node22730 : 16'b0000000000111111;
															assign node22730 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22734 = (inp[7]) ? node22808 : node22735;
										assign node22735 = (inp[2]) ? node22777 : node22736;
											assign node22736 = (inp[15]) ? node22758 : node22737;
												assign node22737 = (inp[4]) ? node22747 : node22738;
													assign node22738 = (inp[13]) ? node22742 : node22739;
														assign node22739 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22742 = (inp[1]) ? node22744 : 16'b0000000011111111;
															assign node22744 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22747 = (inp[1]) ? node22753 : node22748;
														assign node22748 = (inp[12]) ? 16'b0000000001111111 : node22749;
															assign node22749 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22753 = (inp[12]) ? 16'b0000000000011111 : node22754;
															assign node22754 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22758 = (inp[4]) ? node22772 : node22759;
													assign node22759 = (inp[13]) ? node22763 : node22760;
														assign node22760 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22763 = (inp[1]) ? node22769 : node22764;
															assign node22764 = (inp[12]) ? node22766 : 16'b0000000001111111;
																assign node22766 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node22769 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22772 = (inp[12]) ? node22774 : 16'b0000000000111111;
														assign node22774 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22777 = (inp[4]) ? node22791 : node22778;
												assign node22778 = (inp[12]) ? node22786 : node22779;
													assign node22779 = (inp[15]) ? node22781 : 16'b0000000111111111;
														assign node22781 = (inp[1]) ? 16'b0000000000111111 : node22782;
															assign node22782 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22786 = (inp[15]) ? node22788 : 16'b0000000000111111;
														assign node22788 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22791 = (inp[8]) ? node22801 : node22792;
													assign node22792 = (inp[15]) ? node22798 : node22793;
														assign node22793 = (inp[12]) ? 16'b0000000000111111 : node22794;
															assign node22794 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22798 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22801 = (inp[15]) ? node22805 : node22802;
														assign node22802 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22805 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node22808 = (inp[15]) ? node22860 : node22809;
											assign node22809 = (inp[12]) ? node22837 : node22810;
												assign node22810 = (inp[8]) ? node22822 : node22811;
													assign node22811 = (inp[2]) ? node22817 : node22812;
														assign node22812 = (inp[4]) ? 16'b0000000001111111 : node22813;
															assign node22813 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22817 = (inp[1]) ? node22819 : 16'b0000000001111111;
															assign node22819 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22822 = (inp[4]) ? node22830 : node22823;
														assign node22823 = (inp[13]) ? 16'b0000000000111111 : node22824;
															assign node22824 = (inp[2]) ? node22826 : 16'b0000000001111111;
																assign node22826 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22830 = (inp[1]) ? 16'b0000000000011111 : node22831;
															assign node22831 = (inp[2]) ? node22833 : 16'b0000000000111111;
																assign node22833 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22837 = (inp[4]) ? node22851 : node22838;
													assign node22838 = (inp[13]) ? node22846 : node22839;
														assign node22839 = (inp[8]) ? node22841 : 16'b0000000000111111;
															assign node22841 = (inp[1]) ? node22843 : 16'b0000000000111111;
																assign node22843 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22846 = (inp[2]) ? 16'b0000000000011111 : node22847;
															assign node22847 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22851 = (inp[13]) ? 16'b0000000000001111 : node22852;
														assign node22852 = (inp[8]) ? node22854 : 16'b0000000000111111;
															assign node22854 = (inp[1]) ? node22856 : 16'b0000000000011111;
																assign node22856 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node22860 = (inp[2]) ? node22870 : node22861;
												assign node22861 = (inp[1]) ? 16'b0000000000011111 : node22862;
													assign node22862 = (inp[4]) ? node22864 : 16'b0000000000111111;
														assign node22864 = (inp[8]) ? 16'b0000000000011111 : node22865;
															assign node22865 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22870 = (inp[13]) ? node22876 : node22871;
													assign node22871 = (inp[1]) ? node22873 : 16'b0000000000011111;
														assign node22873 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22876 = (inp[8]) ? node22884 : node22877;
														assign node22877 = (inp[4]) ? 16'b0000000000001111 : node22878;
															assign node22878 = (inp[1]) ? node22880 : 16'b0000000000011111;
																assign node22880 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node22884 = (inp[4]) ? 16'b0000000000000111 : node22885;
															assign node22885 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node22889 = (inp[1]) ? node23981 : node22890;
						assign node22890 = (inp[11]) ? node23434 : node22891;
							assign node22891 = (inp[9]) ? node23153 : node22892;
								assign node22892 = (inp[2]) ? node23020 : node22893;
									assign node22893 = (inp[15]) ? node22963 : node22894;
										assign node22894 = (inp[10]) ? node22932 : node22895;
											assign node22895 = (inp[13]) ? node22917 : node22896;
												assign node22896 = (inp[7]) ? node22908 : node22897;
													assign node22897 = (inp[12]) ? node22901 : node22898;
														assign node22898 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node22901 = (inp[14]) ? node22903 : 16'b0000011111111111;
															assign node22903 = (inp[8]) ? 16'b0000001111111111 : node22904;
																assign node22904 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node22908 = (inp[12]) ? node22914 : node22909;
														assign node22909 = (inp[14]) ? node22911 : 16'b0000011111111111;
															assign node22911 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node22914 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node22917 = (inp[12]) ? node22923 : node22918;
													assign node22918 = (inp[7]) ? node22920 : 16'b0000011111111111;
														assign node22920 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22923 = (inp[7]) ? 16'b0000000111111111 : node22924;
														assign node22924 = (inp[14]) ? 16'b0000000111111111 : node22925;
															assign node22925 = (inp[4]) ? node22927 : 16'b0000001111111111;
																assign node22927 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node22932 = (inp[4]) ? node22946 : node22933;
												assign node22933 = (inp[8]) ? 16'b0000000111111111 : node22934;
													assign node22934 = (inp[12]) ? node22940 : node22935;
														assign node22935 = (inp[7]) ? node22937 : 16'b0000001111111111;
															assign node22937 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22940 = (inp[13]) ? 16'b0000001111111111 : node22941;
															assign node22941 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node22946 = (inp[14]) ? node22956 : node22947;
													assign node22947 = (inp[12]) ? node22953 : node22948;
														assign node22948 = (inp[8]) ? node22950 : 16'b0000011111111111;
															assign node22950 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22953 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22956 = (inp[12]) ? node22960 : node22957;
														assign node22957 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22960 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node22963 = (inp[14]) ? node22997 : node22964;
											assign node22964 = (inp[8]) ? node22984 : node22965;
												assign node22965 = (inp[12]) ? node22971 : node22966;
													assign node22966 = (inp[7]) ? 16'b0000001111111111 : node22967;
														assign node22967 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node22971 = (inp[10]) ? node22979 : node22972;
														assign node22972 = (inp[7]) ? node22974 : 16'b0000001111111111;
															assign node22974 = (inp[4]) ? 16'b0000000111111111 : node22975;
																assign node22975 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22979 = (inp[7]) ? node22981 : 16'b0000000111111111;
															assign node22981 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22984 = (inp[7]) ? node22990 : node22985;
													assign node22985 = (inp[4]) ? 16'b0000000111111111 : node22986;
														assign node22986 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22990 = (inp[13]) ? node22992 : 16'b0000000111111111;
														assign node22992 = (inp[4]) ? 16'b0000000011111111 : node22993;
															assign node22993 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node22997 = (inp[13]) ? node23007 : node22998;
												assign node22998 = (inp[8]) ? node23004 : node22999;
													assign node22999 = (inp[10]) ? node23001 : 16'b0000000111111111;
														assign node23001 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23004 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node23007 = (inp[7]) ? node23015 : node23008;
													assign node23008 = (inp[10]) ? node23012 : node23009;
														assign node23009 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node23012 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23015 = (inp[4]) ? node23017 : 16'b0000000011111111;
														assign node23017 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node23020 = (inp[8]) ? node23088 : node23021;
										assign node23021 = (inp[14]) ? node23061 : node23022;
											assign node23022 = (inp[4]) ? node23044 : node23023;
												assign node23023 = (inp[10]) ? node23037 : node23024;
													assign node23024 = (inp[12]) ? node23032 : node23025;
														assign node23025 = (inp[13]) ? node23029 : node23026;
															assign node23026 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node23029 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23032 = (inp[13]) ? 16'b0000001111111111 : node23033;
															assign node23033 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23037 = (inp[7]) ? 16'b0000001111111111 : node23038;
														assign node23038 = (inp[13]) ? 16'b0000000111111111 : node23039;
															assign node23039 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23044 = (inp[12]) ? node23054 : node23045;
													assign node23045 = (inp[15]) ? 16'b0000000111111111 : node23046;
														assign node23046 = (inp[13]) ? node23048 : 16'b0000001111111111;
															assign node23048 = (inp[10]) ? node23050 : 16'b0000001111111111;
																assign node23050 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23054 = (inp[7]) ? node23056 : 16'b0000000011111111;
														assign node23056 = (inp[13]) ? 16'b0000000011111111 : node23057;
															assign node23057 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node23061 = (inp[12]) ? node23075 : node23062;
												assign node23062 = (inp[13]) ? node23072 : node23063;
													assign node23063 = (inp[7]) ? node23069 : node23064;
														assign node23064 = (inp[15]) ? 16'b0000000111111111 : node23065;
															assign node23065 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23069 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23072 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23075 = (inp[13]) ? node23081 : node23076;
													assign node23076 = (inp[7]) ? 16'b0000000011111111 : node23077;
														assign node23077 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node23081 = (inp[4]) ? node23085 : node23082;
														assign node23082 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23085 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node23088 = (inp[12]) ? node23122 : node23089;
											assign node23089 = (inp[4]) ? node23103 : node23090;
												assign node23090 = (inp[14]) ? node23096 : node23091;
													assign node23091 = (inp[15]) ? node23093 : 16'b0000000111111111;
														assign node23093 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23096 = (inp[7]) ? 16'b0000000011111111 : node23097;
														assign node23097 = (inp[15]) ? node23099 : 16'b0000000111111111;
															assign node23099 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23103 = (inp[15]) ? node23111 : node23104;
													assign node23104 = (inp[10]) ? node23106 : 16'b0000000111111111;
														assign node23106 = (inp[14]) ? node23108 : 16'b0000000011111111;
															assign node23108 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23111 = (inp[14]) ? node23117 : node23112;
														assign node23112 = (inp[10]) ? 16'b0000000001111111 : node23113;
															assign node23113 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23117 = (inp[7]) ? node23119 : 16'b0000000001111111;
															assign node23119 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23122 = (inp[14]) ? node23140 : node23123;
												assign node23123 = (inp[7]) ? node23131 : node23124;
													assign node23124 = (inp[10]) ? node23128 : node23125;
														assign node23125 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23128 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23131 = (inp[4]) ? 16'b0000000001111111 : node23132;
														assign node23132 = (inp[13]) ? node23134 : 16'b0000000011111111;
															assign node23134 = (inp[10]) ? 16'b0000000001111111 : node23135;
																assign node23135 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23140 = (inp[13]) ? node23146 : node23141;
													assign node23141 = (inp[15]) ? 16'b0000000001111111 : node23142;
														assign node23142 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23146 = (inp[7]) ? 16'b0000000000111111 : node23147;
														assign node23147 = (inp[4]) ? 16'b0000000000111111 : node23148;
															assign node23148 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node23153 = (inp[4]) ? node23285 : node23154;
									assign node23154 = (inp[13]) ? node23232 : node23155;
										assign node23155 = (inp[8]) ? node23189 : node23156;
											assign node23156 = (inp[14]) ? node23178 : node23157;
												assign node23157 = (inp[7]) ? node23167 : node23158;
													assign node23158 = (inp[2]) ? 16'b0000001111111111 : node23159;
														assign node23159 = (inp[12]) ? 16'b0000001111111111 : node23160;
															assign node23160 = (inp[15]) ? node23162 : 16'b0000011111111111;
																assign node23162 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23167 = (inp[12]) ? node23173 : node23168;
														assign node23168 = (inp[10]) ? node23170 : 16'b0000001111111111;
															assign node23170 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23173 = (inp[2]) ? node23175 : 16'b0000000111111111;
															assign node23175 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23178 = (inp[10]) ? node23182 : node23179;
													assign node23179 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23182 = (inp[2]) ? 16'b0000000001111111 : node23183;
														assign node23183 = (inp[12]) ? node23185 : 16'b0000000111111111;
															assign node23185 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node23189 = (inp[14]) ? node23215 : node23190;
												assign node23190 = (inp[7]) ? node23202 : node23191;
													assign node23191 = (inp[2]) ? node23197 : node23192;
														assign node23192 = (inp[15]) ? 16'b0000000111111111 : node23193;
															assign node23193 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23197 = (inp[12]) ? node23199 : 16'b0000000111111111;
															assign node23199 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23202 = (inp[12]) ? node23208 : node23203;
														assign node23203 = (inp[10]) ? 16'b0000000011111111 : node23204;
															assign node23204 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23208 = (inp[15]) ? 16'b0000000001111111 : node23209;
															assign node23209 = (inp[2]) ? node23211 : 16'b0000000011111111;
																assign node23211 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23215 = (inp[2]) ? node23223 : node23216;
													assign node23216 = (inp[15]) ? node23220 : node23217;
														assign node23217 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23220 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23223 = (inp[12]) ? node23227 : node23224;
														assign node23224 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23227 = (inp[7]) ? node23229 : 16'b0000000001111111;
															assign node23229 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23232 = (inp[7]) ? node23252 : node23233;
											assign node23233 = (inp[15]) ? node23241 : node23234;
												assign node23234 = (inp[8]) ? node23238 : node23235;
													assign node23235 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23238 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23241 = (inp[14]) ? node23247 : node23242;
													assign node23242 = (inp[8]) ? node23244 : 16'b0000000111111111;
														assign node23244 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node23247 = (inp[8]) ? node23249 : 16'b0000000001111111;
														assign node23249 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node23252 = (inp[8]) ? node23268 : node23253;
												assign node23253 = (inp[15]) ? node23261 : node23254;
													assign node23254 = (inp[10]) ? node23258 : node23255;
														assign node23255 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23258 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23261 = (inp[12]) ? node23265 : node23262;
														assign node23262 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23265 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23268 = (inp[12]) ? node23278 : node23269;
													assign node23269 = (inp[14]) ? node23271 : 16'b0000000001111111;
														assign node23271 = (inp[2]) ? 16'b0000000000111111 : node23272;
															assign node23272 = (inp[15]) ? node23274 : 16'b0000000001111111;
																assign node23274 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23278 = (inp[14]) ? node23280 : 16'b0000000000111111;
														assign node23280 = (inp[10]) ? 16'b0000000000011111 : node23281;
															assign node23281 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node23285 = (inp[7]) ? node23353 : node23286;
										assign node23286 = (inp[10]) ? node23314 : node23287;
											assign node23287 = (inp[15]) ? node23297 : node23288;
												assign node23288 = (inp[8]) ? 16'b0000000011111111 : node23289;
													assign node23289 = (inp[13]) ? node23291 : 16'b0000001111111111;
														assign node23291 = (inp[14]) ? 16'b0000000111111111 : node23292;
															assign node23292 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23297 = (inp[2]) ? node23305 : node23298;
													assign node23298 = (inp[12]) ? node23300 : 16'b0000000011111111;
														assign node23300 = (inp[8]) ? node23302 : 16'b0000000011111111;
															assign node23302 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23305 = (inp[8]) ? node23311 : node23306;
														assign node23306 = (inp[12]) ? node23308 : 16'b0000000011111111;
															assign node23308 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23311 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23314 = (inp[15]) ? node23336 : node23315;
												assign node23315 = (inp[14]) ? node23323 : node23316;
													assign node23316 = (inp[13]) ? 16'b0000000001111111 : node23317;
														assign node23317 = (inp[2]) ? node23319 : 16'b0000000111111111;
															assign node23319 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23323 = (inp[2]) ? node23331 : node23324;
														assign node23324 = (inp[8]) ? node23326 : 16'b0000000011111111;
															assign node23326 = (inp[12]) ? 16'b0000000001111111 : node23327;
																assign node23327 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23331 = (inp[8]) ? 16'b0000000000111111 : node23332;
															assign node23332 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23336 = (inp[2]) ? node23348 : node23337;
													assign node23337 = (inp[14]) ? node23341 : node23338;
														assign node23338 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23341 = (inp[8]) ? node23343 : 16'b0000000001111111;
															assign node23343 = (inp[12]) ? 16'b0000000000111111 : node23344;
																assign node23344 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23348 = (inp[12]) ? 16'b0000000000111111 : node23349;
														assign node23349 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node23353 = (inp[13]) ? node23397 : node23354;
											assign node23354 = (inp[2]) ? node23376 : node23355;
												assign node23355 = (inp[12]) ? node23369 : node23356;
													assign node23356 = (inp[14]) ? node23362 : node23357;
														assign node23357 = (inp[10]) ? 16'b0000000111111111 : node23358;
															assign node23358 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23362 = (inp[10]) ? 16'b0000000001111111 : node23363;
															assign node23363 = (inp[15]) ? node23365 : 16'b0000000011111111;
																assign node23365 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23369 = (inp[14]) ? node23371 : 16'b0000000001111111;
														assign node23371 = (inp[8]) ? 16'b0000000000111111 : node23372;
															assign node23372 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23376 = (inp[14]) ? node23390 : node23377;
													assign node23377 = (inp[10]) ? node23383 : node23378;
														assign node23378 = (inp[8]) ? 16'b0000000001111111 : node23379;
															assign node23379 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23383 = (inp[8]) ? 16'b0000000000111111 : node23384;
															assign node23384 = (inp[12]) ? node23386 : 16'b0000000001111111;
																assign node23386 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23390 = (inp[15]) ? node23394 : node23391;
														assign node23391 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23394 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23397 = (inp[12]) ? node23417 : node23398;
												assign node23398 = (inp[14]) ? node23410 : node23399;
													assign node23399 = (inp[10]) ? node23403 : node23400;
														assign node23400 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23403 = (inp[8]) ? 16'b0000000000111111 : node23404;
															assign node23404 = (inp[2]) ? node23406 : 16'b0000000001111111;
																assign node23406 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23410 = (inp[8]) ? node23414 : node23411;
														assign node23411 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23414 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23417 = (inp[2]) ? 16'b0000000000011111 : node23418;
													assign node23418 = (inp[10]) ? node23422 : node23419;
														assign node23419 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23422 = (inp[15]) ? node23428 : node23423;
															assign node23423 = (inp[14]) ? node23425 : 16'b0000000000111111;
																assign node23425 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node23428 = (inp[8]) ? node23430 : 16'b0000000000011111;
																assign node23430 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node23434 = (inp[13]) ? node23706 : node23435;
								assign node23435 = (inp[8]) ? node23553 : node23436;
									assign node23436 = (inp[4]) ? node23496 : node23437;
										assign node23437 = (inp[10]) ? node23471 : node23438;
											assign node23438 = (inp[9]) ? node23458 : node23439;
												assign node23439 = (inp[7]) ? node23447 : node23440;
													assign node23440 = (inp[2]) ? 16'b0000000111111111 : node23441;
														assign node23441 = (inp[14]) ? node23443 : 16'b0000011111111111;
															assign node23443 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23447 = (inp[14]) ? node23453 : node23448;
														assign node23448 = (inp[15]) ? 16'b0000000111111111 : node23449;
															assign node23449 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23453 = (inp[15]) ? 16'b0000000011111111 : node23454;
															assign node23454 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23458 = (inp[14]) ? node23462 : node23459;
													assign node23459 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23462 = (inp[7]) ? node23466 : node23463;
														assign node23463 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23466 = (inp[15]) ? node23468 : 16'b0000000011111111;
															assign node23468 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23471 = (inp[2]) ? node23485 : node23472;
												assign node23472 = (inp[15]) ? node23480 : node23473;
													assign node23473 = (inp[12]) ? node23475 : 16'b0000000111111111;
														assign node23475 = (inp[9]) ? 16'b0000000011111111 : node23476;
															assign node23476 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23480 = (inp[9]) ? 16'b0000000011111111 : node23481;
														assign node23481 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23485 = (inp[7]) ? node23491 : node23486;
													assign node23486 = (inp[14]) ? node23488 : 16'b0000000011111111;
														assign node23488 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23491 = (inp[15]) ? 16'b0000000000011111 : node23492;
														assign node23492 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node23496 = (inp[9]) ? node23520 : node23497;
											assign node23497 = (inp[15]) ? node23511 : node23498;
												assign node23498 = (inp[2]) ? node23502 : node23499;
													assign node23499 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23502 = (inp[7]) ? node23506 : node23503;
														assign node23503 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23506 = (inp[10]) ? node23508 : 16'b0000000011111111;
															assign node23508 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23511 = (inp[14]) ? node23513 : 16'b0000000011111111;
													assign node23513 = (inp[12]) ? 16'b0000000001111111 : node23514;
														assign node23514 = (inp[7]) ? node23516 : 16'b0000000011111111;
															assign node23516 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23520 = (inp[7]) ? node23538 : node23521;
												assign node23521 = (inp[2]) ? node23529 : node23522;
													assign node23522 = (inp[14]) ? node23524 : 16'b0000000111111111;
														assign node23524 = (inp[10]) ? 16'b0000000011111111 : node23525;
															assign node23525 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23529 = (inp[14]) ? 16'b0000000000111111 : node23530;
														assign node23530 = (inp[12]) ? 16'b0000000001111111 : node23531;
															assign node23531 = (inp[15]) ? node23533 : 16'b0000000111111111;
																assign node23533 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23538 = (inp[2]) ? node23546 : node23539;
													assign node23539 = (inp[12]) ? node23543 : node23540;
														assign node23540 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23543 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23546 = (inp[12]) ? node23550 : node23547;
														assign node23547 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23550 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node23553 = (inp[7]) ? node23637 : node23554;
										assign node23554 = (inp[4]) ? node23592 : node23555;
											assign node23555 = (inp[2]) ? node23573 : node23556;
												assign node23556 = (inp[10]) ? node23564 : node23557;
													assign node23557 = (inp[14]) ? 16'b0000000111111111 : node23558;
														assign node23558 = (inp[12]) ? 16'b0000001111111111 : node23559;
															assign node23559 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23564 = (inp[14]) ? 16'b0000000011111111 : node23565;
														assign node23565 = (inp[15]) ? 16'b0000000011111111 : node23566;
															assign node23566 = (inp[12]) ? node23568 : 16'b0000000111111111;
																assign node23568 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23573 = (inp[12]) ? node23581 : node23574;
													assign node23574 = (inp[15]) ? node23576 : 16'b0000001111111111;
														assign node23576 = (inp[9]) ? node23578 : 16'b0000000011111111;
															assign node23578 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23581 = (inp[15]) ? node23589 : node23582;
														assign node23582 = (inp[14]) ? node23584 : 16'b0000000111111111;
															assign node23584 = (inp[9]) ? 16'b0000000001111111 : node23585;
																assign node23585 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23589 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23592 = (inp[14]) ? node23618 : node23593;
												assign node23593 = (inp[9]) ? node23609 : node23594;
													assign node23594 = (inp[10]) ? node23598 : node23595;
														assign node23595 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23598 = (inp[12]) ? node23604 : node23599;
															assign node23599 = (inp[15]) ? node23601 : 16'b0000000011111111;
																assign node23601 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node23604 = (inp[15]) ? 16'b0000000001111111 : node23605;
																assign node23605 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23609 = (inp[12]) ? node23613 : node23610;
														assign node23610 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23613 = (inp[10]) ? node23615 : 16'b0000000001111111;
															assign node23615 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node23618 = (inp[2]) ? node23628 : node23619;
													assign node23619 = (inp[10]) ? node23623 : node23620;
														assign node23620 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node23623 = (inp[12]) ? node23625 : 16'b0000000001111111;
															assign node23625 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23628 = (inp[9]) ? node23634 : node23629;
														assign node23629 = (inp[15]) ? 16'b0000000000111111 : node23630;
															assign node23630 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23634 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23637 = (inp[2]) ? node23675 : node23638;
											assign node23638 = (inp[15]) ? node23660 : node23639;
												assign node23639 = (inp[4]) ? node23645 : node23640;
													assign node23640 = (inp[10]) ? node23642 : 16'b0000000011111111;
														assign node23642 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23645 = (inp[14]) ? node23657 : node23646;
														assign node23646 = (inp[10]) ? node23652 : node23647;
															assign node23647 = (inp[12]) ? node23649 : 16'b0000000011111111;
																assign node23649 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node23652 = (inp[12]) ? node23654 : 16'b0000000001111111;
																assign node23654 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23657 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23660 = (inp[9]) ? node23670 : node23661;
													assign node23661 = (inp[14]) ? 16'b0000000000111111 : node23662;
														assign node23662 = (inp[10]) ? node23666 : node23663;
															assign node23663 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node23666 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23670 = (inp[14]) ? node23672 : 16'b0000000000111111;
														assign node23672 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23675 = (inp[9]) ? node23687 : node23676;
												assign node23676 = (inp[14]) ? node23680 : node23677;
													assign node23677 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23680 = (inp[4]) ? node23684 : node23681;
														assign node23681 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23684 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23687 = (inp[15]) ? node23693 : node23688;
													assign node23688 = (inp[12]) ? node23690 : 16'b0000000000111111;
														assign node23690 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23693 = (inp[14]) ? node23701 : node23694;
														assign node23694 = (inp[12]) ? node23696 : 16'b0000000001111111;
															assign node23696 = (inp[4]) ? 16'b0000000000011111 : node23697;
																assign node23697 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23701 = (inp[4]) ? node23703 : 16'b0000000000011111;
															assign node23703 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node23706 = (inp[14]) ? node23848 : node23707;
									assign node23707 = (inp[2]) ? node23767 : node23708;
										assign node23708 = (inp[4]) ? node23738 : node23709;
											assign node23709 = (inp[15]) ? node23725 : node23710;
												assign node23710 = (inp[12]) ? node23718 : node23711;
													assign node23711 = (inp[9]) ? 16'b0000000111111111 : node23712;
														assign node23712 = (inp[8]) ? node23714 : 16'b0000001111111111;
															assign node23714 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23718 = (inp[10]) ? 16'b0000000011111111 : node23719;
														assign node23719 = (inp[7]) ? 16'b0000000011111111 : node23720;
															assign node23720 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23725 = (inp[8]) ? node23731 : node23726;
													assign node23726 = (inp[9]) ? 16'b0000000011111111 : node23727;
														assign node23727 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23731 = (inp[9]) ? node23733 : 16'b0000000011111111;
														assign node23733 = (inp[10]) ? node23735 : 16'b0000000001111111;
															assign node23735 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23738 = (inp[15]) ? node23756 : node23739;
												assign node23739 = (inp[9]) ? node23747 : node23740;
													assign node23740 = (inp[12]) ? node23742 : 16'b0000000111111111;
														assign node23742 = (inp[7]) ? 16'b0000000001111111 : node23743;
															assign node23743 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23747 = (inp[10]) ? node23753 : node23748;
														assign node23748 = (inp[8]) ? 16'b0000000001111111 : node23749;
															assign node23749 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23753 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23756 = (inp[8]) ? node23762 : node23757;
													assign node23757 = (inp[12]) ? node23759 : 16'b0000000001111111;
														assign node23759 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23762 = (inp[9]) ? node23764 : 16'b0000000000111111;
														assign node23764 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node23767 = (inp[9]) ? node23803 : node23768;
											assign node23768 = (inp[12]) ? node23788 : node23769;
												assign node23769 = (inp[10]) ? node23777 : node23770;
													assign node23770 = (inp[7]) ? node23772 : 16'b0000000111111111;
														assign node23772 = (inp[15]) ? 16'b0000000001111111 : node23773;
															assign node23773 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23777 = (inp[4]) ? node23783 : node23778;
														assign node23778 = (inp[7]) ? 16'b0000000001111111 : node23779;
															assign node23779 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23783 = (inp[15]) ? 16'b0000000000111111 : node23784;
															assign node23784 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23788 = (inp[8]) ? node23794 : node23789;
													assign node23789 = (inp[4]) ? 16'b0000000001111111 : node23790;
														assign node23790 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000111111111;
													assign node23794 = (inp[10]) ? 16'b0000000000011111 : node23795;
														assign node23795 = (inp[7]) ? node23797 : 16'b0000000000111111;
															assign node23797 = (inp[4]) ? node23799 : 16'b0000000000111111;
																assign node23799 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23803 = (inp[7]) ? node23827 : node23804;
												assign node23804 = (inp[10]) ? node23812 : node23805;
													assign node23805 = (inp[4]) ? node23809 : node23806;
														assign node23806 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23809 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23812 = (inp[8]) ? node23820 : node23813;
														assign node23813 = (inp[15]) ? 16'b0000000000111111 : node23814;
															assign node23814 = (inp[4]) ? node23816 : 16'b0000000001111111;
																assign node23816 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23820 = (inp[4]) ? 16'b0000000000011111 : node23821;
															assign node23821 = (inp[15]) ? node23823 : 16'b0000000000111111;
																assign node23823 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23827 = (inp[4]) ? node23837 : node23828;
													assign node23828 = (inp[10]) ? 16'b0000000000011111 : node23829;
														assign node23829 = (inp[12]) ? node23831 : 16'b0000000001111111;
															assign node23831 = (inp[8]) ? node23833 : 16'b0000000000111111;
																assign node23833 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23837 = (inp[15]) ? node23841 : node23838;
														assign node23838 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23841 = (inp[10]) ? node23843 : 16'b0000000000011111;
															assign node23843 = (inp[12]) ? 16'b0000000000001111 : node23844;
																assign node23844 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node23848 = (inp[7]) ? node23908 : node23849;
										assign node23849 = (inp[12]) ? node23879 : node23850;
											assign node23850 = (inp[9]) ? node23862 : node23851;
												assign node23851 = (inp[10]) ? node23857 : node23852;
													assign node23852 = (inp[8]) ? 16'b0000000001111111 : node23853;
														assign node23853 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23857 = (inp[4]) ? 16'b0000000001111111 : node23858;
														assign node23858 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node23862 = (inp[2]) ? node23874 : node23863;
													assign node23863 = (inp[10]) ? node23869 : node23864;
														assign node23864 = (inp[4]) ? 16'b0000000001111111 : node23865;
															assign node23865 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23869 = (inp[8]) ? 16'b0000000000011111 : node23870;
															assign node23870 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23874 = (inp[8]) ? node23876 : 16'b0000000000111111;
														assign node23876 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23879 = (inp[10]) ? node23895 : node23880;
												assign node23880 = (inp[9]) ? node23890 : node23881;
													assign node23881 = (inp[4]) ? node23883 : 16'b0000000001111111;
														assign node23883 = (inp[15]) ? node23885 : 16'b0000000001111111;
															assign node23885 = (inp[8]) ? 16'b0000000000111111 : node23886;
																assign node23886 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23890 = (inp[15]) ? node23892 : 16'b0000000000111111;
														assign node23892 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23895 = (inp[9]) ? node23899 : node23896;
													assign node23896 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23899 = (inp[4]) ? node23901 : 16'b0000000000111111;
														assign node23901 = (inp[15]) ? node23903 : 16'b0000000000011111;
															assign node23903 = (inp[2]) ? 16'b0000000000001111 : node23904;
																assign node23904 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23908 = (inp[15]) ? node23938 : node23909;
											assign node23909 = (inp[8]) ? node23923 : node23910;
												assign node23910 = (inp[10]) ? node23916 : node23911;
													assign node23911 = (inp[2]) ? node23913 : 16'b0000000111111111;
														assign node23913 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23916 = (inp[9]) ? node23920 : node23917;
														assign node23917 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23920 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23923 = (inp[2]) ? node23931 : node23924;
													assign node23924 = (inp[9]) ? node23926 : 16'b0000000000111111;
														assign node23926 = (inp[4]) ? 16'b0000000000011111 : node23927;
															assign node23927 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23931 = (inp[12]) ? 16'b0000000000001111 : node23932;
														assign node23932 = (inp[9]) ? 16'b0000000000011111 : node23933;
															assign node23933 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23938 = (inp[4]) ? node23960 : node23939;
												assign node23939 = (inp[12]) ? node23953 : node23940;
													assign node23940 = (inp[9]) ? node23950 : node23941;
														assign node23941 = (inp[8]) ? node23945 : node23942;
															assign node23942 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node23945 = (inp[2]) ? 16'b0000000000111111 : node23946;
																assign node23946 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23950 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23953 = (inp[8]) ? node23955 : 16'b0000000000011111;
														assign node23955 = (inp[2]) ? 16'b0000000000001111 : node23956;
															assign node23956 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23960 = (inp[2]) ? node23968 : node23961;
													assign node23961 = (inp[8]) ? node23963 : 16'b0000000000011111;
														assign node23963 = (inp[12]) ? 16'b0000000000001111 : node23964;
															assign node23964 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23968 = (inp[9]) ? node23970 : 16'b0000000000001111;
														assign node23970 = (inp[10]) ? node23976 : node23971;
															assign node23971 = (inp[12]) ? node23973 : 16'b0000000000001111;
																assign node23973 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node23976 = (inp[8]) ? 16'b0000000000000111 : node23977;
																assign node23977 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node23981 = (inp[8]) ? node24475 : node23982;
							assign node23982 = (inp[11]) ? node24230 : node23983;
								assign node23983 = (inp[4]) ? node24083 : node23984;
									assign node23984 = (inp[15]) ? node24026 : node23985;
										assign node23985 = (inp[7]) ? node24001 : node23986;
											assign node23986 = (inp[10]) ? node23996 : node23987;
												assign node23987 = (inp[9]) ? node23993 : node23988;
													assign node23988 = (inp[12]) ? 16'b0000001111111111 : node23989;
														assign node23989 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23993 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23996 = (inp[13]) ? node23998 : 16'b0000000111111111;
													assign node23998 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node24001 = (inp[10]) ? node24015 : node24002;
												assign node24002 = (inp[12]) ? node24010 : node24003;
													assign node24003 = (inp[14]) ? 16'b0000000111111111 : node24004;
														assign node24004 = (inp[13]) ? node24006 : 16'b0000001111111111;
															assign node24006 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24010 = (inp[2]) ? 16'b0000000011111111 : node24011;
														assign node24011 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24015 = (inp[13]) ? node24017 : 16'b0000000011111111;
													assign node24017 = (inp[14]) ? node24021 : node24018;
														assign node24018 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24021 = (inp[2]) ? node24023 : 16'b0000000001111111;
															assign node24023 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node24026 = (inp[12]) ? node24060 : node24027;
											assign node24027 = (inp[2]) ? node24041 : node24028;
												assign node24028 = (inp[7]) ? node24038 : node24029;
													assign node24029 = (inp[10]) ? node24033 : node24030;
														assign node24030 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24033 = (inp[14]) ? node24035 : 16'b0000000111111111;
															assign node24035 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24038 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24041 = (inp[7]) ? node24051 : node24042;
													assign node24042 = (inp[13]) ? node24048 : node24043;
														assign node24043 = (inp[14]) ? 16'b0000000011111111 : node24044;
															assign node24044 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24048 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24051 = (inp[14]) ? node24055 : node24052;
														assign node24052 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24055 = (inp[10]) ? node24057 : 16'b0000000001111111;
															assign node24057 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24060 = (inp[13]) ? node24066 : node24061;
												assign node24061 = (inp[7]) ? node24063 : 16'b0000000111111111;
													assign node24063 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24066 = (inp[7]) ? node24074 : node24067;
													assign node24067 = (inp[10]) ? node24071 : node24068;
														assign node24068 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24071 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24074 = (inp[2]) ? node24080 : node24075;
														assign node24075 = (inp[14]) ? 16'b0000000000111111 : node24076;
															assign node24076 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24080 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node24083 = (inp[15]) ? node24161 : node24084;
										assign node24084 = (inp[14]) ? node24116 : node24085;
											assign node24085 = (inp[12]) ? node24099 : node24086;
												assign node24086 = (inp[7]) ? node24090 : node24087;
													assign node24087 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24090 = (inp[10]) ? 16'b0000000011111111 : node24091;
														assign node24091 = (inp[2]) ? node24093 : 16'b0000000111111111;
															assign node24093 = (inp[13]) ? 16'b0000000011111111 : node24094;
																assign node24094 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24099 = (inp[13]) ? node24109 : node24100;
													assign node24100 = (inp[10]) ? node24102 : 16'b0000001111111111;
														assign node24102 = (inp[7]) ? 16'b0000000001111111 : node24103;
															assign node24103 = (inp[2]) ? 16'b0000000011111111 : node24104;
																assign node24104 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24109 = (inp[7]) ? 16'b0000000001111111 : node24110;
														assign node24110 = (inp[9]) ? 16'b0000000001111111 : node24111;
															assign node24111 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24116 = (inp[13]) ? node24144 : node24117;
												assign node24117 = (inp[10]) ? node24133 : node24118;
													assign node24118 = (inp[9]) ? node24128 : node24119;
														assign node24119 = (inp[7]) ? node24125 : node24120;
															assign node24120 = (inp[12]) ? node24122 : 16'b0000000111111111;
																assign node24122 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node24125 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24128 = (inp[12]) ? node24130 : 16'b0000000011111111;
															assign node24130 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24133 = (inp[2]) ? node24139 : node24134;
														assign node24134 = (inp[12]) ? node24136 : 16'b0000000111111111;
															assign node24136 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24139 = (inp[7]) ? 16'b0000000000111111 : node24140;
															assign node24140 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24144 = (inp[7]) ? node24152 : node24145;
													assign node24145 = (inp[2]) ? node24147 : 16'b0000000001111111;
														assign node24147 = (inp[10]) ? node24149 : 16'b0000000001111111;
															assign node24149 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24152 = (inp[12]) ? node24158 : node24153;
														assign node24153 = (inp[9]) ? node24155 : 16'b0000000001111111;
															assign node24155 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24158 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node24161 = (inp[14]) ? node24201 : node24162;
											assign node24162 = (inp[7]) ? node24186 : node24163;
												assign node24163 = (inp[9]) ? node24175 : node24164;
													assign node24164 = (inp[2]) ? node24170 : node24165;
														assign node24165 = (inp[12]) ? node24167 : 16'b0000000111111111;
															assign node24167 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24170 = (inp[12]) ? node24172 : 16'b0000000011111111;
															assign node24172 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24175 = (inp[12]) ? node24179 : node24176;
														assign node24176 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node24179 = (inp[10]) ? 16'b0000000000111111 : node24180;
															assign node24180 = (inp[2]) ? node24182 : 16'b0000000001111111;
																assign node24182 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24186 = (inp[12]) ? node24192 : node24187;
													assign node24187 = (inp[9]) ? node24189 : 16'b0000000001111111;
														assign node24189 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node24192 = (inp[9]) ? node24198 : node24193;
														assign node24193 = (inp[10]) ? 16'b0000000000111111 : node24194;
															assign node24194 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24198 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node24201 = (inp[13]) ? node24217 : node24202;
												assign node24202 = (inp[7]) ? node24210 : node24203;
													assign node24203 = (inp[2]) ? node24207 : node24204;
														assign node24204 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24207 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node24210 = (inp[10]) ? node24214 : node24211;
														assign node24211 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24214 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24217 = (inp[12]) ? node24227 : node24218;
													assign node24218 = (inp[7]) ? 16'b0000000000011111 : node24219;
														assign node24219 = (inp[2]) ? node24223 : node24220;
															assign node24220 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node24223 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24227 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node24230 = (inp[4]) ? node24368 : node24231;
									assign node24231 = (inp[2]) ? node24295 : node24232;
										assign node24232 = (inp[12]) ? node24256 : node24233;
											assign node24233 = (inp[13]) ? node24247 : node24234;
												assign node24234 = (inp[10]) ? node24242 : node24235;
													assign node24235 = (inp[15]) ? 16'b0000000011111111 : node24236;
														assign node24236 = (inp[14]) ? 16'b0000000111111111 : node24237;
															assign node24237 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node24242 = (inp[14]) ? node24244 : 16'b0000000011111111;
														assign node24244 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24247 = (inp[9]) ? node24249 : 16'b0000000011111111;
													assign node24249 = (inp[15]) ? 16'b0000000001111111 : node24250;
														assign node24250 = (inp[7]) ? node24252 : 16'b0000000011111111;
															assign node24252 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24256 = (inp[9]) ? node24278 : node24257;
												assign node24257 = (inp[7]) ? node24267 : node24258;
													assign node24258 = (inp[13]) ? node24262 : node24259;
														assign node24259 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24262 = (inp[15]) ? node24264 : 16'b0000000011111111;
															assign node24264 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24267 = (inp[10]) ? node24275 : node24268;
														assign node24268 = (inp[15]) ? 16'b0000000001111111 : node24269;
															assign node24269 = (inp[14]) ? node24271 : 16'b0000000011111111;
																assign node24271 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24275 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24278 = (inp[15]) ? node24290 : node24279;
													assign node24279 = (inp[14]) ? node24283 : node24280;
														assign node24280 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24283 = (inp[7]) ? node24285 : 16'b0000000001111111;
															assign node24285 = (inp[10]) ? 16'b0000000000111111 : node24286;
																assign node24286 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24290 = (inp[10]) ? node24292 : 16'b0000000000111111;
														assign node24292 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node24295 = (inp[13]) ? node24335 : node24296;
											assign node24296 = (inp[14]) ? node24318 : node24297;
												assign node24297 = (inp[9]) ? node24309 : node24298;
													assign node24298 = (inp[7]) ? node24306 : node24299;
														assign node24299 = (inp[15]) ? node24301 : 16'b0000000111111111;
															assign node24301 = (inp[10]) ? 16'b0000000011111111 : node24302;
																assign node24302 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24306 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24309 = (inp[15]) ? node24313 : node24310;
														assign node24310 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24313 = (inp[7]) ? node24315 : 16'b0000000001111111;
															assign node24315 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24318 = (inp[15]) ? node24326 : node24319;
													assign node24319 = (inp[12]) ? node24321 : 16'b0000000001111111;
														assign node24321 = (inp[10]) ? 16'b0000000000111111 : node24322;
															assign node24322 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24326 = (inp[9]) ? node24330 : node24327;
														assign node24327 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24330 = (inp[12]) ? node24332 : 16'b0000000000111111;
															assign node24332 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24335 = (inp[10]) ? node24353 : node24336;
												assign node24336 = (inp[14]) ? node24344 : node24337;
													assign node24337 = (inp[9]) ? node24341 : node24338;
														assign node24338 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24341 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24344 = (inp[12]) ? node24346 : 16'b0000000000111111;
														assign node24346 = (inp[7]) ? 16'b0000000000011111 : node24347;
															assign node24347 = (inp[9]) ? node24349 : 16'b0000000000111111;
																assign node24349 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24353 = (inp[9]) ? node24359 : node24354;
													assign node24354 = (inp[15]) ? node24356 : 16'b0000000000111111;
														assign node24356 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24359 = (inp[14]) ? node24363 : node24360;
														assign node24360 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24363 = (inp[7]) ? node24365 : 16'b0000000000011111;
															assign node24365 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node24368 = (inp[7]) ? node24406 : node24369;
										assign node24369 = (inp[10]) ? node24385 : node24370;
											assign node24370 = (inp[9]) ? node24380 : node24371;
												assign node24371 = (inp[15]) ? node24375 : node24372;
													assign node24372 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24375 = (inp[14]) ? 16'b0000000001111111 : node24376;
														assign node24376 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node24380 = (inp[14]) ? node24382 : 16'b0000000001111111;
													assign node24382 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24385 = (inp[15]) ? node24393 : node24386;
												assign node24386 = (inp[13]) ? 16'b0000000000111111 : node24387;
													assign node24387 = (inp[14]) ? node24389 : 16'b0000000001111111;
														assign node24389 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24393 = (inp[14]) ? node24399 : node24394;
													assign node24394 = (inp[12]) ? 16'b0000000000111111 : node24395;
														assign node24395 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24399 = (inp[9]) ? node24401 : 16'b0000000000111111;
														assign node24401 = (inp[12]) ? 16'b0000000000001111 : node24402;
															assign node24402 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node24406 = (inp[15]) ? node24442 : node24407;
											assign node24407 = (inp[12]) ? node24425 : node24408;
												assign node24408 = (inp[13]) ? node24416 : node24409;
													assign node24409 = (inp[9]) ? 16'b0000000011111111 : node24410;
														assign node24410 = (inp[14]) ? 16'b0000000001111111 : node24411;
															assign node24411 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24416 = (inp[10]) ? node24420 : node24417;
														assign node24417 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24420 = (inp[9]) ? node24422 : 16'b0000000000111111;
															assign node24422 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24425 = (inp[2]) ? node24433 : node24426;
													assign node24426 = (inp[10]) ? 16'b0000000000011111 : node24427;
														assign node24427 = (inp[9]) ? 16'b0000000000111111 : node24428;
															assign node24428 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24433 = (inp[9]) ? node24437 : node24434;
														assign node24434 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24437 = (inp[14]) ? node24439 : 16'b0000000000001111;
															assign node24439 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node24442 = (inp[13]) ? node24452 : node24443;
												assign node24443 = (inp[9]) ? node24447 : node24444;
													assign node24444 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node24447 = (inp[10]) ? node24449 : 16'b0000000000011111;
														assign node24449 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node24452 = (inp[14]) ? node24462 : node24453;
													assign node24453 = (inp[2]) ? node24457 : node24454;
														assign node24454 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24457 = (inp[10]) ? node24459 : 16'b0000000000011111;
															assign node24459 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node24462 = (inp[9]) ? node24470 : node24463;
														assign node24463 = (inp[12]) ? node24465 : 16'b0000000000001111;
															assign node24465 = (inp[2]) ? node24467 : 16'b0000000000001111;
																assign node24467 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node24470 = (inp[10]) ? 16'b0000000000000111 : node24471;
															assign node24471 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node24475 = (inp[9]) ? node24753 : node24476;
								assign node24476 = (inp[4]) ? node24622 : node24477;
									assign node24477 = (inp[2]) ? node24543 : node24478;
										assign node24478 = (inp[12]) ? node24508 : node24479;
											assign node24479 = (inp[10]) ? node24491 : node24480;
												assign node24480 = (inp[11]) ? node24486 : node24481;
													assign node24481 = (inp[15]) ? 16'b0000000111111111 : node24482;
														assign node24482 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24486 = (inp[13]) ? 16'b0000000001111111 : node24487;
														assign node24487 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24491 = (inp[11]) ? node24501 : node24492;
													assign node24492 = (inp[15]) ? node24496 : node24493;
														assign node24493 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24496 = (inp[7]) ? 16'b0000000001111111 : node24497;
															assign node24497 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24501 = (inp[13]) ? 16'b0000000000111111 : node24502;
														assign node24502 = (inp[7]) ? 16'b0000000001111111 : node24503;
															assign node24503 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24508 = (inp[15]) ? node24532 : node24509;
												assign node24509 = (inp[7]) ? node24523 : node24510;
													assign node24510 = (inp[13]) ? node24518 : node24511;
														assign node24511 = (inp[14]) ? node24513 : 16'b0000000011111111;
															assign node24513 = (inp[10]) ? node24515 : 16'b0000000011111111;
																assign node24515 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24518 = (inp[14]) ? 16'b0000000001111111 : node24519;
															assign node24519 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24523 = (inp[13]) ? node24527 : node24524;
														assign node24524 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node24527 = (inp[10]) ? node24529 : 16'b0000000001111111;
															assign node24529 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24532 = (inp[14]) ? node24540 : node24533;
													assign node24533 = (inp[11]) ? 16'b0000000000111111 : node24534;
														assign node24534 = (inp[10]) ? 16'b0000000001111111 : node24535;
															assign node24535 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24540 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node24543 = (inp[10]) ? node24589 : node24544;
											assign node24544 = (inp[15]) ? node24568 : node24545;
												assign node24545 = (inp[14]) ? node24551 : node24546;
													assign node24546 = (inp[7]) ? 16'b0000000011111111 : node24547;
														assign node24547 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24551 = (inp[12]) ? node24561 : node24552;
														assign node24552 = (inp[13]) ? node24556 : node24553;
															assign node24553 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node24556 = (inp[7]) ? 16'b0000000001111111 : node24557;
																assign node24557 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24561 = (inp[7]) ? node24563 : 16'b0000000001111111;
															assign node24563 = (inp[13]) ? 16'b0000000000111111 : node24564;
																assign node24564 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24568 = (inp[12]) ? node24582 : node24569;
													assign node24569 = (inp[14]) ? node24575 : node24570;
														assign node24570 = (inp[13]) ? 16'b0000000001111111 : node24571;
															assign node24571 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24575 = (inp[11]) ? node24577 : 16'b0000000001111111;
															assign node24577 = (inp[7]) ? node24579 : 16'b0000000000111111;
																assign node24579 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24582 = (inp[11]) ? 16'b0000000000011111 : node24583;
														assign node24583 = (inp[13]) ? node24585 : 16'b0000000001111111;
															assign node24585 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24589 = (inp[14]) ? node24611 : node24590;
												assign node24590 = (inp[11]) ? node24600 : node24591;
													assign node24591 = (inp[12]) ? node24593 : 16'b0000000011111111;
														assign node24593 = (inp[13]) ? node24595 : 16'b0000000001111111;
															assign node24595 = (inp[7]) ? 16'b0000000000111111 : node24596;
																assign node24596 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24600 = (inp[12]) ? node24604 : node24601;
														assign node24601 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24604 = (inp[13]) ? node24606 : 16'b0000000000111111;
															assign node24606 = (inp[15]) ? 16'b0000000000011111 : node24607;
																assign node24607 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24611 = (inp[15]) ? node24613 : 16'b0000000000111111;
													assign node24613 = (inp[7]) ? node24615 : 16'b0000000000111111;
														assign node24615 = (inp[11]) ? 16'b0000000000001111 : node24616;
															assign node24616 = (inp[12]) ? node24618 : 16'b0000000000011111;
																assign node24618 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node24622 = (inp[14]) ? node24692 : node24623;
										assign node24623 = (inp[7]) ? node24653 : node24624;
											assign node24624 = (inp[12]) ? node24638 : node24625;
												assign node24625 = (inp[15]) ? node24633 : node24626;
													assign node24626 = (inp[10]) ? node24630 : node24627;
														assign node24627 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24630 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24633 = (inp[11]) ? 16'b0000000001111111 : node24634;
														assign node24634 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24638 = (inp[15]) ? 16'b0000000000111111 : node24639;
													assign node24639 = (inp[2]) ? node24647 : node24640;
														assign node24640 = (inp[10]) ? node24642 : 16'b0000000011111111;
															assign node24642 = (inp[11]) ? node24644 : 16'b0000000011111111;
																assign node24644 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24647 = (inp[11]) ? 16'b0000000000111111 : node24648;
															assign node24648 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24653 = (inp[12]) ? node24669 : node24654;
												assign node24654 = (inp[13]) ? node24664 : node24655;
													assign node24655 = (inp[15]) ? 16'b0000000000111111 : node24656;
														assign node24656 = (inp[2]) ? node24658 : 16'b0000000001111111;
															assign node24658 = (inp[11]) ? node24660 : 16'b0000000001111111;
																assign node24660 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24664 = (inp[11]) ? 16'b0000000000011111 : node24665;
														assign node24665 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24669 = (inp[11]) ? node24681 : node24670;
													assign node24670 = (inp[2]) ? node24678 : node24671;
														assign node24671 = (inp[10]) ? node24673 : 16'b0000000001111111;
															assign node24673 = (inp[15]) ? node24675 : 16'b0000000000111111;
																assign node24675 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24678 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24681 = (inp[10]) ? node24687 : node24682;
														assign node24682 = (inp[13]) ? 16'b0000000000011111 : node24683;
															assign node24683 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24687 = (inp[2]) ? 16'b0000000000001111 : node24688;
															assign node24688 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node24692 = (inp[13]) ? node24716 : node24693;
											assign node24693 = (inp[10]) ? node24703 : node24694;
												assign node24694 = (inp[12]) ? 16'b0000000000111111 : node24695;
													assign node24695 = (inp[15]) ? node24697 : 16'b0000000001111111;
														assign node24697 = (inp[2]) ? 16'b0000000000111111 : node24698;
															assign node24698 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24703 = (inp[15]) ? node24711 : node24704;
													assign node24704 = (inp[11]) ? node24708 : node24705;
														assign node24705 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24708 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24711 = (inp[7]) ? node24713 : 16'b0000000000011111;
														assign node24713 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node24716 = (inp[11]) ? node24730 : node24717;
												assign node24717 = (inp[2]) ? node24725 : node24718;
													assign node24718 = (inp[7]) ? node24722 : node24719;
														assign node24719 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24722 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24725 = (inp[10]) ? 16'b0000000000011111 : node24726;
														assign node24726 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24730 = (inp[12]) ? node24740 : node24731;
													assign node24731 = (inp[7]) ? node24733 : 16'b0000000000011111;
														assign node24733 = (inp[15]) ? 16'b0000000000001111 : node24734;
															assign node24734 = (inp[10]) ? node24736 : 16'b0000000000011111;
																assign node24736 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24740 = (inp[15]) ? node24744 : node24741;
														assign node24741 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24744 = (inp[10]) ? node24750 : node24745;
															assign node24745 = (inp[2]) ? node24747 : 16'b0000000000001111;
																assign node24747 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node24750 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
								assign node24753 = (inp[10]) ? node24853 : node24754;
									assign node24754 = (inp[14]) ? node24802 : node24755;
										assign node24755 = (inp[15]) ? node24779 : node24756;
											assign node24756 = (inp[7]) ? node24772 : node24757;
												assign node24757 = (inp[4]) ? node24763 : node24758;
													assign node24758 = (inp[13]) ? 16'b0000000011111111 : node24759;
														assign node24759 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24763 = (inp[11]) ? node24769 : node24764;
														assign node24764 = (inp[12]) ? 16'b0000000001111111 : node24765;
															assign node24765 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24769 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24772 = (inp[4]) ? 16'b0000000000111111 : node24773;
													assign node24773 = (inp[12]) ? 16'b0000000000111111 : node24774;
														assign node24774 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24779 = (inp[13]) ? node24789 : node24780;
												assign node24780 = (inp[2]) ? 16'b0000000000111111 : node24781;
													assign node24781 = (inp[11]) ? node24783 : 16'b0000000011111111;
														assign node24783 = (inp[7]) ? node24785 : 16'b0000000001111111;
															assign node24785 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24789 = (inp[7]) ? node24795 : node24790;
													assign node24790 = (inp[11]) ? 16'b0000000000011111 : node24791;
														assign node24791 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24795 = (inp[12]) ? node24799 : node24796;
														assign node24796 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node24799 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node24802 = (inp[11]) ? node24834 : node24803;
											assign node24803 = (inp[4]) ? node24825 : node24804;
												assign node24804 = (inp[15]) ? node24814 : node24805;
													assign node24805 = (inp[12]) ? 16'b0000000001111111 : node24806;
														assign node24806 = (inp[13]) ? 16'b0000000001111111 : node24807;
															assign node24807 = (inp[7]) ? node24809 : 16'b0000000011111111;
																assign node24809 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24814 = (inp[12]) ? node24820 : node24815;
														assign node24815 = (inp[13]) ? 16'b0000000000111111 : node24816;
															assign node24816 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24820 = (inp[13]) ? node24822 : 16'b0000000000111111;
															assign node24822 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24825 = (inp[13]) ? 16'b0000000000011111 : node24826;
													assign node24826 = (inp[2]) ? node24828 : 16'b0000000000111111;
														assign node24828 = (inp[7]) ? 16'b0000000000011111 : node24829;
															assign node24829 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24834 = (inp[7]) ? node24836 : 16'b0000000000011111;
												assign node24836 = (inp[2]) ? node24844 : node24837;
													assign node24837 = (inp[4]) ? node24841 : node24838;
														assign node24838 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24841 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24844 = (inp[15]) ? node24848 : node24845;
														assign node24845 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node24848 = (inp[13]) ? 16'b0000000000000111 : node24849;
															assign node24849 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node24853 = (inp[12]) ? node24929 : node24854;
										assign node24854 = (inp[2]) ? node24898 : node24855;
											assign node24855 = (inp[11]) ? node24875 : node24856;
												assign node24856 = (inp[4]) ? node24864 : node24857;
													assign node24857 = (inp[13]) ? node24861 : node24858;
														assign node24858 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24861 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24864 = (inp[14]) ? node24868 : node24865;
														assign node24865 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24868 = (inp[13]) ? 16'b0000000000011111 : node24869;
															assign node24869 = (inp[15]) ? node24871 : 16'b0000000000111111;
																assign node24871 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24875 = (inp[7]) ? node24887 : node24876;
													assign node24876 = (inp[14]) ? node24882 : node24877;
														assign node24877 = (inp[4]) ? node24879 : 16'b0000000001111111;
															assign node24879 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24882 = (inp[15]) ? 16'b0000000000011111 : node24883;
															assign node24883 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24887 = (inp[13]) ? node24891 : node24888;
														assign node24888 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24891 = (inp[14]) ? node24893 : 16'b0000000000011111;
															assign node24893 = (inp[4]) ? 16'b0000000000001111 : node24894;
																assign node24894 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node24898 = (inp[7]) ? node24914 : node24899;
												assign node24899 = (inp[4]) ? node24905 : node24900;
													assign node24900 = (inp[15]) ? 16'b0000000000011111 : node24901;
														assign node24901 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24905 = (inp[11]) ? node24909 : node24906;
														assign node24906 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24909 = (inp[14]) ? node24911 : 16'b0000000000011111;
															assign node24911 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node24914 = (inp[4]) ? node24922 : node24915;
													assign node24915 = (inp[11]) ? node24919 : node24916;
														assign node24916 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24919 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24922 = (inp[13]) ? 16'b0000000000000111 : node24923;
														assign node24923 = (inp[14]) ? 16'b0000000000001111 : node24924;
															assign node24924 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node24929 = (inp[4]) ? node24949 : node24930;
											assign node24930 = (inp[14]) ? node24936 : node24931;
												assign node24931 = (inp[15]) ? node24933 : 16'b0000000011111111;
													assign node24933 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24936 = (inp[15]) ? node24946 : node24937;
													assign node24937 = (inp[13]) ? 16'b0000000000001111 : node24938;
														assign node24938 = (inp[7]) ? node24940 : 16'b0000000000011111;
															assign node24940 = (inp[2]) ? node24942 : 16'b0000000000011111;
																assign node24942 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24946 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node24949 = (inp[7]) ? node24959 : node24950;
												assign node24950 = (inp[13]) ? node24954 : node24951;
													assign node24951 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node24954 = (inp[11]) ? node24956 : 16'b0000000000011111;
														assign node24956 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node24959 = (inp[2]) ? node24969 : node24960;
													assign node24960 = (inp[15]) ? node24966 : node24961;
														assign node24961 = (inp[14]) ? node24963 : 16'b0000000000011111;
															assign node24963 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node24966 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node24969 = (inp[15]) ? node24971 : 16'b0000000000000111;
														assign node24971 = (inp[14]) ? 16'b0000000000000011 : node24972;
															assign node24972 = (inp[11]) ? node24976 : node24973;
																assign node24973 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
																assign node24976 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;
			assign node24980 = (inp[5]) ? node29082 : node24981;
				assign node24981 = (inp[13]) ? node26989 : node24982;
					assign node24982 = (inp[1]) ? node25972 : node24983;
						assign node24983 = (inp[15]) ? node25505 : node24984;
							assign node24984 = (inp[11]) ? node25236 : node24985;
								assign node24985 = (inp[7]) ? node25119 : node24986;
									assign node24986 = (inp[14]) ? node25048 : node24987;
										assign node24987 = (inp[2]) ? node25017 : node24988;
											assign node24988 = (inp[8]) ? node24998 : node24989;
												assign node24989 = (inp[10]) ? node24995 : node24990;
													assign node24990 = (inp[4]) ? 16'b0000111111111111 : node24991;
														assign node24991 = (inp[6]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node24995 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node24998 = (inp[6]) ? node25006 : node24999;
													assign node24999 = (inp[4]) ? 16'b0000011111111111 : node25000;
														assign node25000 = (inp[9]) ? node25002 : 16'b0001111111111111;
															assign node25002 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node25006 = (inp[9]) ? node25012 : node25007;
														assign node25007 = (inp[12]) ? 16'b0000011111111111 : node25008;
															assign node25008 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node25012 = (inp[4]) ? 16'b0000001111111111 : node25013;
															assign node25013 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node25017 = (inp[6]) ? node25033 : node25018;
												assign node25018 = (inp[9]) ? node25024 : node25019;
													assign node25019 = (inp[12]) ? 16'b0000011111111111 : node25020;
														assign node25020 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node25024 = (inp[10]) ? node25028 : node25025;
														assign node25025 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25028 = (inp[8]) ? node25030 : 16'b0000001111111111;
															assign node25030 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25033 = (inp[10]) ? node25043 : node25034;
													assign node25034 = (inp[12]) ? 16'b0000000111111111 : node25035;
														assign node25035 = (inp[4]) ? node25037 : 16'b0000011111111111;
															assign node25037 = (inp[9]) ? 16'b0000001111111111 : node25038;
																assign node25038 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25043 = (inp[4]) ? 16'b0000000011111111 : node25044;
														assign node25044 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node25048 = (inp[2]) ? node25092 : node25049;
											assign node25049 = (inp[8]) ? node25071 : node25050;
												assign node25050 = (inp[4]) ? node25058 : node25051;
													assign node25051 = (inp[6]) ? node25053 : 16'b0000111111111111;
														assign node25053 = (inp[10]) ? 16'b0000001111111111 : node25054;
															assign node25054 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node25058 = (inp[9]) ? node25064 : node25059;
														assign node25059 = (inp[6]) ? 16'b0000001111111111 : node25060;
															assign node25060 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node25064 = (inp[12]) ? node25066 : 16'b0000001111111111;
															assign node25066 = (inp[6]) ? 16'b0000000111111111 : node25067;
																assign node25067 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25071 = (inp[4]) ? node25079 : node25072;
													assign node25072 = (inp[6]) ? node25076 : node25073;
														assign node25073 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25076 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25079 = (inp[10]) ? 16'b0000000011111111 : node25080;
														assign node25080 = (inp[12]) ? node25086 : node25081;
															assign node25081 = (inp[6]) ? node25083 : 16'b0000001111111111;
																assign node25083 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node25086 = (inp[9]) ? node25088 : 16'b0000000111111111;
																assign node25088 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node25092 = (inp[10]) ? node25108 : node25093;
												assign node25093 = (inp[9]) ? node25099 : node25094;
													assign node25094 = (inp[8]) ? node25096 : 16'b0000001111111111;
														assign node25096 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25099 = (inp[8]) ? node25105 : node25100;
														assign node25100 = (inp[6]) ? 16'b0000000111111111 : node25101;
															assign node25101 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25105 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25108 = (inp[8]) ? 16'b0000000011111111 : node25109;
													assign node25109 = (inp[12]) ? node25111 : 16'b0000001111111111;
														assign node25111 = (inp[6]) ? 16'b0000000011111111 : node25112;
															assign node25112 = (inp[9]) ? node25114 : 16'b0000000111111111;
																assign node25114 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node25119 = (inp[8]) ? node25175 : node25120;
										assign node25120 = (inp[6]) ? node25144 : node25121;
											assign node25121 = (inp[2]) ? node25137 : node25122;
												assign node25122 = (inp[10]) ? node25132 : node25123;
													assign node25123 = (inp[12]) ? node25129 : node25124;
														assign node25124 = (inp[14]) ? 16'b0000111111111111 : node25125;
															assign node25125 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node25129 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25132 = (inp[12]) ? 16'b0000001111111111 : node25133;
														assign node25133 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node25137 = (inp[12]) ? node25139 : 16'b0000001111111111;
													assign node25139 = (inp[14]) ? 16'b0000000111111111 : node25140;
														assign node25140 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node25144 = (inp[9]) ? node25166 : node25145;
												assign node25145 = (inp[4]) ? node25157 : node25146;
													assign node25146 = (inp[10]) ? node25152 : node25147;
														assign node25147 = (inp[2]) ? node25149 : 16'b0000011111111111;
															assign node25149 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25152 = (inp[2]) ? 16'b0000000111111111 : node25153;
															assign node25153 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25157 = (inp[14]) ? node25161 : node25158;
														assign node25158 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25161 = (inp[10]) ? node25163 : 16'b0000000111111111;
															assign node25163 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25166 = (inp[2]) ? node25170 : node25167;
													assign node25167 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25170 = (inp[4]) ? node25172 : 16'b0000000011111111;
														assign node25172 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node25175 = (inp[12]) ? node25199 : node25176;
											assign node25176 = (inp[2]) ? node25180 : node25177;
												assign node25177 = (inp[6]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node25180 = (inp[4]) ? node25190 : node25181;
													assign node25181 = (inp[6]) ? node25185 : node25182;
														assign node25182 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25185 = (inp[9]) ? node25187 : 16'b0000000111111111;
															assign node25187 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25190 = (inp[14]) ? 16'b0000000011111111 : node25191;
														assign node25191 = (inp[10]) ? node25193 : 16'b0000000111111111;
															assign node25193 = (inp[6]) ? 16'b0000000011111111 : node25194;
																assign node25194 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node25199 = (inp[9]) ? node25217 : node25200;
												assign node25200 = (inp[6]) ? node25206 : node25201;
													assign node25201 = (inp[2]) ? 16'b0000000011111111 : node25202;
														assign node25202 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25206 = (inp[4]) ? node25214 : node25207;
														assign node25207 = (inp[14]) ? 16'b0000000011111111 : node25208;
															assign node25208 = (inp[2]) ? node25210 : 16'b0000000111111111;
																assign node25210 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25214 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25217 = (inp[14]) ? node25229 : node25218;
													assign node25218 = (inp[6]) ? node25224 : node25219;
														assign node25219 = (inp[10]) ? 16'b0000000011111111 : node25220;
															assign node25220 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25224 = (inp[10]) ? node25226 : 16'b0000000011111111;
															assign node25226 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25229 = (inp[10]) ? node25231 : 16'b0000000001111111;
														assign node25231 = (inp[2]) ? 16'b0000000000111111 : node25232;
															assign node25232 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node25236 = (inp[6]) ? node25384 : node25237;
									assign node25237 = (inp[7]) ? node25325 : node25238;
										assign node25238 = (inp[9]) ? node25280 : node25239;
											assign node25239 = (inp[8]) ? node25257 : node25240;
												assign node25240 = (inp[2]) ? node25248 : node25241;
													assign node25241 = (inp[10]) ? node25245 : node25242;
														assign node25242 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node25245 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25248 = (inp[10]) ? node25254 : node25249;
														assign node25249 = (inp[12]) ? 16'b0000001111111111 : node25250;
															assign node25250 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25254 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25257 = (inp[12]) ? node25275 : node25258;
													assign node25258 = (inp[14]) ? node25270 : node25259;
														assign node25259 = (inp[2]) ? node25265 : node25260;
															assign node25260 = (inp[10]) ? node25262 : 16'b0000011111111111;
																assign node25262 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node25265 = (inp[10]) ? node25267 : 16'b0000001111111111;
																assign node25267 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25270 = (inp[2]) ? 16'b0000000111111111 : node25271;
															assign node25271 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25275 = (inp[4]) ? 16'b0000000011111111 : node25276;
														assign node25276 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node25280 = (inp[4]) ? node25304 : node25281;
												assign node25281 = (inp[10]) ? node25293 : node25282;
													assign node25282 = (inp[14]) ? node25290 : node25283;
														assign node25283 = (inp[8]) ? node25285 : 16'b0000011111111111;
															assign node25285 = (inp[2]) ? 16'b0000001111111111 : node25286;
																assign node25286 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25290 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node25293 = (inp[2]) ? node25301 : node25294;
														assign node25294 = (inp[14]) ? 16'b0000000111111111 : node25295;
															assign node25295 = (inp[12]) ? node25297 : 16'b0000001111111111;
																assign node25297 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25301 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25304 = (inp[8]) ? node25314 : node25305;
													assign node25305 = (inp[10]) ? node25309 : node25306;
														assign node25306 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25309 = (inp[14]) ? node25311 : 16'b0000000111111111;
															assign node25311 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25314 = (inp[10]) ? node25322 : node25315;
														assign node25315 = (inp[12]) ? 16'b0000000011111111 : node25316;
															assign node25316 = (inp[14]) ? node25318 : 16'b0000000111111111;
																assign node25318 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25322 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node25325 = (inp[8]) ? node25355 : node25326;
											assign node25326 = (inp[10]) ? node25346 : node25327;
												assign node25327 = (inp[14]) ? node25337 : node25328;
													assign node25328 = (inp[9]) ? node25334 : node25329;
														assign node25329 = (inp[4]) ? 16'b0000001111111111 : node25330;
															assign node25330 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25334 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25337 = (inp[12]) ? node25343 : node25338;
														assign node25338 = (inp[2]) ? 16'b0000000111111111 : node25339;
															assign node25339 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25343 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node25346 = (inp[4]) ? node25348 : 16'b0000000111111111;
													assign node25348 = (inp[14]) ? node25352 : node25349;
														assign node25349 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25352 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25355 = (inp[2]) ? node25367 : node25356;
												assign node25356 = (inp[4]) ? node25358 : 16'b0000001111111111;
													assign node25358 = (inp[9]) ? 16'b0000000001111111 : node25359;
														assign node25359 = (inp[10]) ? 16'b0000000011111111 : node25360;
															assign node25360 = (inp[14]) ? node25362 : 16'b0000000111111111;
																assign node25362 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25367 = (inp[12]) ? node25375 : node25368;
													assign node25368 = (inp[4]) ? node25370 : 16'b0000000011111111;
														assign node25370 = (inp[10]) ? node25372 : 16'b0000000011111111;
															assign node25372 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25375 = (inp[4]) ? 16'b0000000001111111 : node25376;
														assign node25376 = (inp[9]) ? node25378 : 16'b0000000011111111;
															assign node25378 = (inp[14]) ? 16'b0000000001111111 : node25379;
																assign node25379 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node25384 = (inp[2]) ? node25450 : node25385;
										assign node25385 = (inp[12]) ? node25421 : node25386;
											assign node25386 = (inp[10]) ? node25408 : node25387;
												assign node25387 = (inp[4]) ? node25399 : node25388;
													assign node25388 = (inp[9]) ? node25396 : node25389;
														assign node25389 = (inp[8]) ? node25391 : 16'b0000011111111111;
															assign node25391 = (inp[14]) ? 16'b0000001111111111 : node25392;
																assign node25392 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25396 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25399 = (inp[7]) ? node25405 : node25400;
														assign node25400 = (inp[8]) ? 16'b0000000111111111 : node25401;
															assign node25401 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25405 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node25408 = (inp[4]) ? node25414 : node25409;
													assign node25409 = (inp[9]) ? 16'b0000000011111111 : node25410;
														assign node25410 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25414 = (inp[9]) ? node25416 : 16'b0000000011111111;
														assign node25416 = (inp[8]) ? 16'b0000000001111111 : node25417;
															assign node25417 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25421 = (inp[8]) ? node25437 : node25422;
												assign node25422 = (inp[10]) ? node25430 : node25423;
													assign node25423 = (inp[4]) ? node25425 : 16'b0000000111111111;
														assign node25425 = (inp[9]) ? 16'b0000000011111111 : node25426;
															assign node25426 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25430 = (inp[9]) ? 16'b0000000011111111 : node25431;
														assign node25431 = (inp[4]) ? 16'b0000000011111111 : node25432;
															assign node25432 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25437 = (inp[9]) ? node25443 : node25438;
													assign node25438 = (inp[10]) ? 16'b0000000001111111 : node25439;
														assign node25439 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25443 = (inp[14]) ? node25447 : node25444;
														assign node25444 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node25447 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node25450 = (inp[9]) ? node25476 : node25451;
											assign node25451 = (inp[12]) ? node25459 : node25452;
												assign node25452 = (inp[7]) ? 16'b0000000011111111 : node25453;
													assign node25453 = (inp[8]) ? 16'b0000000111111111 : node25454;
														assign node25454 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25459 = (inp[4]) ? node25467 : node25460;
													assign node25460 = (inp[8]) ? node25464 : node25461;
														assign node25461 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25464 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25467 = (inp[10]) ? node25471 : node25468;
														assign node25468 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node25471 = (inp[8]) ? node25473 : 16'b0000000001111111;
															assign node25473 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node25476 = (inp[14]) ? node25484 : node25477;
												assign node25477 = (inp[8]) ? node25479 : 16'b0000000011111111;
													assign node25479 = (inp[4]) ? 16'b0000000000111111 : node25480;
														assign node25480 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25484 = (inp[7]) ? node25498 : node25485;
													assign node25485 = (inp[4]) ? node25491 : node25486;
														assign node25486 = (inp[12]) ? 16'b0000000001111111 : node25487;
															assign node25487 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25491 = (inp[8]) ? node25493 : 16'b0000000001111111;
															assign node25493 = (inp[12]) ? node25495 : 16'b0000000000111111;
																assign node25495 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25498 = (inp[8]) ? node25500 : 16'b0000000000111111;
														assign node25500 = (inp[4]) ? node25502 : 16'b0000000000011111;
															assign node25502 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node25505 = (inp[2]) ? node25733 : node25506;
								assign node25506 = (inp[8]) ? node25610 : node25507;
									assign node25507 = (inp[7]) ? node25559 : node25508;
										assign node25508 = (inp[6]) ? node25534 : node25509;
											assign node25509 = (inp[14]) ? node25525 : node25510;
												assign node25510 = (inp[10]) ? node25522 : node25511;
													assign node25511 = (inp[9]) ? node25513 : 16'b0000111111111111;
														assign node25513 = (inp[12]) ? node25517 : node25514;
															assign node25514 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node25517 = (inp[4]) ? 16'b0000001111111111 : node25518;
																assign node25518 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25522 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25525 = (inp[11]) ? node25531 : node25526;
													assign node25526 = (inp[9]) ? node25528 : 16'b0000001111111111;
														assign node25528 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25531 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node25534 = (inp[11]) ? node25546 : node25535;
												assign node25535 = (inp[12]) ? node25541 : node25536;
													assign node25536 = (inp[10]) ? node25538 : 16'b0000001111111111;
														assign node25538 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25541 = (inp[14]) ? 16'b0000000111111111 : node25542;
														assign node25542 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25546 = (inp[12]) ? node25552 : node25547;
													assign node25547 = (inp[9]) ? 16'b0000000111111111 : node25548;
														assign node25548 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node25552 = (inp[10]) ? node25556 : node25553;
														assign node25553 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node25556 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node25559 = (inp[14]) ? node25583 : node25560;
											assign node25560 = (inp[4]) ? node25570 : node25561;
												assign node25561 = (inp[12]) ? node25563 : 16'b0000001111111111;
													assign node25563 = (inp[6]) ? node25567 : node25564;
														assign node25564 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25567 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25570 = (inp[9]) ? node25576 : node25571;
													assign node25571 = (inp[6]) ? 16'b0000000111111111 : node25572;
														assign node25572 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25576 = (inp[11]) ? node25580 : node25577;
														assign node25577 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25580 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25583 = (inp[4]) ? node25603 : node25584;
												assign node25584 = (inp[12]) ? node25598 : node25585;
													assign node25585 = (inp[6]) ? node25593 : node25586;
														assign node25586 = (inp[9]) ? node25588 : 16'b0000001111111111;
															assign node25588 = (inp[11]) ? 16'b0000000111111111 : node25589;
																assign node25589 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25593 = (inp[11]) ? 16'b0000000011111111 : node25594;
															assign node25594 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25598 = (inp[9]) ? node25600 : 16'b0000000111111111;
														assign node25600 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25603 = (inp[9]) ? node25605 : 16'b0000000011111111;
													assign node25605 = (inp[6]) ? 16'b0000000001111111 : node25606;
														assign node25606 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node25610 = (inp[12]) ? node25672 : node25611;
										assign node25611 = (inp[14]) ? node25637 : node25612;
											assign node25612 = (inp[9]) ? node25628 : node25613;
												assign node25613 = (inp[6]) ? node25619 : node25614;
													assign node25614 = (inp[4]) ? 16'b0000001111111111 : node25615;
														assign node25615 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25619 = (inp[10]) ? 16'b0000000111111111 : node25620;
														assign node25620 = (inp[7]) ? node25622 : 16'b0000001111111111;
															assign node25622 = (inp[4]) ? 16'b0000000111111111 : node25623;
																assign node25623 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25628 = (inp[6]) ? node25634 : node25629;
													assign node25629 = (inp[4]) ? node25631 : 16'b0000001111111111;
														assign node25631 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25634 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node25637 = (inp[11]) ? node25657 : node25638;
												assign node25638 = (inp[7]) ? node25652 : node25639;
													assign node25639 = (inp[4]) ? node25649 : node25640;
														assign node25640 = (inp[10]) ? node25646 : node25641;
															assign node25641 = (inp[6]) ? 16'b0000001111111111 : node25642;
																assign node25642 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node25646 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25649 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25652 = (inp[10]) ? node25654 : 16'b0000000011111111;
														assign node25654 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node25657 = (inp[6]) ? node25665 : node25658;
													assign node25658 = (inp[10]) ? 16'b0000000011111111 : node25659;
														assign node25659 = (inp[4]) ? 16'b0000000011111111 : node25660;
															assign node25660 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25665 = (inp[10]) ? node25669 : node25666;
														assign node25666 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25669 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node25672 = (inp[9]) ? node25698 : node25673;
											assign node25673 = (inp[6]) ? node25681 : node25674;
												assign node25674 = (inp[14]) ? node25676 : 16'b0000000111111111;
													assign node25676 = (inp[4]) ? 16'b0000000011111111 : node25677;
														assign node25677 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25681 = (inp[4]) ? 16'b0000000001111111 : node25682;
													assign node25682 = (inp[11]) ? node25690 : node25683;
														assign node25683 = (inp[7]) ? 16'b0000000011111111 : node25684;
															assign node25684 = (inp[10]) ? node25686 : 16'b0000000111111111;
																assign node25686 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25690 = (inp[7]) ? node25692 : 16'b0000000011111111;
															assign node25692 = (inp[10]) ? 16'b0000000001111111 : node25693;
																assign node25693 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25698 = (inp[14]) ? node25718 : node25699;
												assign node25699 = (inp[11]) ? node25711 : node25700;
													assign node25700 = (inp[6]) ? node25704 : node25701;
														assign node25701 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25704 = (inp[4]) ? node25706 : 16'b0000000011111111;
															assign node25706 = (inp[7]) ? 16'b0000000001111111 : node25707;
																assign node25707 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25711 = (inp[7]) ? 16'b0000000001111111 : node25712;
														assign node25712 = (inp[6]) ? node25714 : 16'b0000000011111111;
															assign node25714 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25718 = (inp[11]) ? node25722 : node25719;
													assign node25719 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25722 = (inp[7]) ? node25726 : node25723;
														assign node25723 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25726 = (inp[4]) ? node25728 : 16'b0000000000111111;
															assign node25728 = (inp[6]) ? node25730 : 16'b0000000000011111;
																assign node25730 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node25733 = (inp[6]) ? node25859 : node25734;
									assign node25734 = (inp[12]) ? node25806 : node25735;
										assign node25735 = (inp[10]) ? node25775 : node25736;
											assign node25736 = (inp[14]) ? node25752 : node25737;
												assign node25737 = (inp[7]) ? node25745 : node25738;
													assign node25738 = (inp[4]) ? 16'b0000001111111111 : node25739;
														assign node25739 = (inp[9]) ? 16'b0000001111111111 : node25740;
															assign node25740 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node25745 = (inp[4]) ? node25747 : 16'b0000001111111111;
														assign node25747 = (inp[8]) ? node25749 : 16'b0000000111111111;
															assign node25749 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25752 = (inp[8]) ? node25764 : node25753;
													assign node25753 = (inp[11]) ? node25757 : node25754;
														assign node25754 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25757 = (inp[7]) ? node25759 : 16'b0000000111111111;
															assign node25759 = (inp[4]) ? 16'b0000000011111111 : node25760;
																assign node25760 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25764 = (inp[7]) ? node25768 : node25765;
														assign node25765 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25768 = (inp[11]) ? node25772 : node25769;
															assign node25769 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node25772 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25775 = (inp[4]) ? node25791 : node25776;
												assign node25776 = (inp[14]) ? node25784 : node25777;
													assign node25777 = (inp[8]) ? node25779 : 16'b0000001111111111;
														assign node25779 = (inp[9]) ? node25781 : 16'b0000000111111111;
															assign node25781 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25784 = (inp[8]) ? node25788 : node25785;
														assign node25785 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25788 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25791 = (inp[11]) ? node25795 : node25792;
													assign node25792 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node25795 = (inp[8]) ? node25803 : node25796;
														assign node25796 = (inp[9]) ? node25798 : 16'b0000000001111111;
															assign node25798 = (inp[14]) ? node25800 : 16'b0000000001111111;
																assign node25800 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25803 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node25806 = (inp[9]) ? node25846 : node25807;
											assign node25807 = (inp[14]) ? node25823 : node25808;
												assign node25808 = (inp[4]) ? node25816 : node25809;
													assign node25809 = (inp[11]) ? 16'b0000000011111111 : node25810;
														assign node25810 = (inp[10]) ? node25812 : 16'b0000001111111111;
															assign node25812 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25816 = (inp[8]) ? 16'b0000000011111111 : node25817;
														assign node25817 = (inp[10]) ? 16'b0000000011111111 : node25818;
															assign node25818 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25823 = (inp[4]) ? node25833 : node25824;
													assign node25824 = (inp[8]) ? node25830 : node25825;
														assign node25825 = (inp[7]) ? node25827 : 16'b0000000111111111;
															assign node25827 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25830 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25833 = (inp[7]) ? node25841 : node25834;
														assign node25834 = (inp[8]) ? 16'b0000000001111111 : node25835;
															assign node25835 = (inp[10]) ? node25837 : 16'b0000000011111111;
																assign node25837 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25841 = (inp[11]) ? node25843 : 16'b0000000001111111;
															assign node25843 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node25846 = (inp[8]) ? node25854 : node25847;
												assign node25847 = (inp[14]) ? node25849 : 16'b0000000011111111;
													assign node25849 = (inp[7]) ? 16'b0000000000111111 : node25850;
														assign node25850 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25854 = (inp[7]) ? 16'b0000000000011111 : node25855;
													assign node25855 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node25859 = (inp[4]) ? node25921 : node25860;
										assign node25860 = (inp[7]) ? node25894 : node25861;
											assign node25861 = (inp[9]) ? node25875 : node25862;
												assign node25862 = (inp[12]) ? node25868 : node25863;
													assign node25863 = (inp[8]) ? node25865 : 16'b0000000111111111;
														assign node25865 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25868 = (inp[10]) ? node25872 : node25869;
														assign node25869 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25872 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25875 = (inp[8]) ? node25889 : node25876;
													assign node25876 = (inp[10]) ? node25886 : node25877;
														assign node25877 = (inp[14]) ? node25881 : node25878;
															assign node25878 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node25881 = (inp[12]) ? 16'b0000000011111111 : node25882;
																assign node25882 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25886 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node25889 = (inp[11]) ? 16'b0000000001111111 : node25890;
														assign node25890 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25894 = (inp[14]) ? node25908 : node25895;
												assign node25895 = (inp[8]) ? node25901 : node25896;
													assign node25896 = (inp[9]) ? 16'b0000000011111111 : node25897;
														assign node25897 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25901 = (inp[9]) ? node25903 : 16'b0000000011111111;
														assign node25903 = (inp[10]) ? node25905 : 16'b0000000001111111;
															assign node25905 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25908 = (inp[8]) ? node25914 : node25909;
													assign node25909 = (inp[12]) ? node25911 : 16'b0000000001111111;
														assign node25911 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25914 = (inp[10]) ? 16'b0000000000111111 : node25915;
														assign node25915 = (inp[9]) ? 16'b0000000000111111 : node25916;
															assign node25916 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node25921 = (inp[14]) ? node25939 : node25922;
											assign node25922 = (inp[9]) ? node25932 : node25923;
												assign node25923 = (inp[10]) ? node25925 : 16'b0000000111111111;
													assign node25925 = (inp[11]) ? node25929 : node25926;
														assign node25926 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25929 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25932 = (inp[8]) ? node25934 : 16'b0000000001111111;
													assign node25934 = (inp[11]) ? node25936 : 16'b0000000001111111;
														assign node25936 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node25939 = (inp[12]) ? node25957 : node25940;
												assign node25940 = (inp[8]) ? node25948 : node25941;
													assign node25941 = (inp[11]) ? 16'b0000000000111111 : node25942;
														assign node25942 = (inp[10]) ? 16'b0000000001111111 : node25943;
															assign node25943 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25948 = (inp[9]) ? node25950 : 16'b0000000001111111;
														assign node25950 = (inp[7]) ? 16'b0000000000011111 : node25951;
															assign node25951 = (inp[11]) ? node25953 : 16'b0000000000111111;
																assign node25953 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node25957 = (inp[9]) ? node25963 : node25958;
													assign node25958 = (inp[10]) ? node25960 : 16'b0000000000111111;
														assign node25960 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25963 = (inp[11]) ? node25967 : node25964;
														assign node25964 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node25967 = (inp[8]) ? node25969 : 16'b0000000000011111;
															assign node25969 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node25972 = (inp[14]) ? node26486 : node25973;
							assign node25973 = (inp[12]) ? node26227 : node25974;
								assign node25974 = (inp[9]) ? node26108 : node25975;
									assign node25975 = (inp[15]) ? node26045 : node25976;
										assign node25976 = (inp[10]) ? node26012 : node25977;
											assign node25977 = (inp[4]) ? node26005 : node25978;
												assign node25978 = (inp[8]) ? node25994 : node25979;
													assign node25979 = (inp[11]) ? node25987 : node25980;
														assign node25980 = (inp[2]) ? node25982 : 16'b0000111111111111;
															assign node25982 = (inp[6]) ? 16'b0000011111111111 : node25983;
																assign node25983 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node25987 = (inp[2]) ? 16'b0000000111111111 : node25988;
															assign node25988 = (inp[6]) ? node25990 : 16'b0000011111111111;
																assign node25990 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25994 = (inp[2]) ? node25998 : node25995;
														assign node25995 = (inp[6]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25998 = (inp[11]) ? 16'b0000000111111111 : node25999;
															assign node25999 = (inp[7]) ? node26001 : 16'b0000001111111111;
																assign node26001 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node26005 = (inp[8]) ? 16'b0000000111111111 : node26006;
													assign node26006 = (inp[7]) ? node26008 : 16'b0000001111111111;
														assign node26008 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node26012 = (inp[11]) ? node26028 : node26013;
												assign node26013 = (inp[2]) ? node26021 : node26014;
													assign node26014 = (inp[8]) ? node26018 : node26015;
														assign node26015 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node26018 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26021 = (inp[8]) ? node26025 : node26022;
														assign node26022 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26025 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26028 = (inp[4]) ? node26038 : node26029;
													assign node26029 = (inp[2]) ? node26031 : 16'b0000000111111111;
														assign node26031 = (inp[8]) ? 16'b0000000011111111 : node26032;
															assign node26032 = (inp[7]) ? node26034 : 16'b0000000111111111;
																assign node26034 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26038 = (inp[6]) ? node26042 : node26039;
														assign node26039 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26042 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node26045 = (inp[10]) ? node26079 : node26046;
											assign node26046 = (inp[2]) ? node26060 : node26047;
												assign node26047 = (inp[7]) ? node26055 : node26048;
													assign node26048 = (inp[8]) ? node26050 : 16'b0000011111111111;
														assign node26050 = (inp[11]) ? 16'b0000000111111111 : node26051;
															assign node26051 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26055 = (inp[6]) ? node26057 : 16'b0000000111111111;
														assign node26057 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26060 = (inp[6]) ? node26074 : node26061;
													assign node26061 = (inp[7]) ? node26069 : node26062;
														assign node26062 = (inp[11]) ? node26064 : 16'b0000000111111111;
															assign node26064 = (inp[8]) ? node26066 : 16'b0000000111111111;
																assign node26066 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26069 = (inp[4]) ? 16'b0000000011111111 : node26070;
															assign node26070 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26074 = (inp[8]) ? 16'b0000000011111111 : node26075;
														assign node26075 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node26079 = (inp[7]) ? node26093 : node26080;
												assign node26080 = (inp[6]) ? node26088 : node26081;
													assign node26081 = (inp[4]) ? node26083 : 16'b0000001111111111;
														assign node26083 = (inp[11]) ? 16'b0000000111111111 : node26084;
															assign node26084 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26088 = (inp[8]) ? 16'b0000000000111111 : node26089;
														assign node26089 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26093 = (inp[2]) ? node26095 : 16'b0000000011111111;
													assign node26095 = (inp[8]) ? node26101 : node26096;
														assign node26096 = (inp[4]) ? node26098 : 16'b0000000011111111;
															assign node26098 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26101 = (inp[6]) ? 16'b0000000001111111 : node26102;
															assign node26102 = (inp[4]) ? 16'b0000000001111111 : node26103;
																assign node26103 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node26108 = (inp[6]) ? node26168 : node26109;
										assign node26109 = (inp[10]) ? node26137 : node26110;
											assign node26110 = (inp[11]) ? node26122 : node26111;
												assign node26111 = (inp[15]) ? node26117 : node26112;
													assign node26112 = (inp[8]) ? 16'b0000001111111111 : node26113;
														assign node26113 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node26117 = (inp[2]) ? node26119 : 16'b0000001111111111;
														assign node26119 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26122 = (inp[7]) ? node26132 : node26123;
													assign node26123 = (inp[4]) ? node26127 : node26124;
														assign node26124 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26127 = (inp[8]) ? node26129 : 16'b0000000111111111;
															assign node26129 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26132 = (inp[8]) ? 16'b0000000011111111 : node26133;
														assign node26133 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node26137 = (inp[7]) ? node26157 : node26138;
												assign node26138 = (inp[15]) ? node26148 : node26139;
													assign node26139 = (inp[8]) ? node26145 : node26140;
														assign node26140 = (inp[4]) ? 16'b0000000111111111 : node26141;
															assign node26141 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node26145 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26148 = (inp[11]) ? node26154 : node26149;
														assign node26149 = (inp[2]) ? 16'b0000000011111111 : node26150;
															assign node26150 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26154 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26157 = (inp[4]) ? 16'b0000000001111111 : node26158;
													assign node26158 = (inp[2]) ? node26162 : node26159;
														assign node26159 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node26162 = (inp[11]) ? node26164 : 16'b0000000011111111;
															assign node26164 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node26168 = (inp[2]) ? node26202 : node26169;
											assign node26169 = (inp[11]) ? node26183 : node26170;
												assign node26170 = (inp[10]) ? node26178 : node26171;
													assign node26171 = (inp[7]) ? node26173 : 16'b0000000111111111;
														assign node26173 = (inp[4]) ? node26175 : 16'b0000000111111111;
															assign node26175 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26178 = (inp[4]) ? 16'b0000000011111111 : node26179;
														assign node26179 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26183 = (inp[8]) ? node26195 : node26184;
													assign node26184 = (inp[4]) ? node26190 : node26185;
														assign node26185 = (inp[7]) ? node26187 : 16'b0000000111111111;
															assign node26187 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26190 = (inp[7]) ? 16'b0000000001111111 : node26191;
															assign node26191 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26195 = (inp[4]) ? node26199 : node26196;
														assign node26196 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26199 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node26202 = (inp[8]) ? node26218 : node26203;
												assign node26203 = (inp[7]) ? node26209 : node26204;
													assign node26204 = (inp[10]) ? node26206 : 16'b0000000111111111;
														assign node26206 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node26209 = (inp[4]) ? node26213 : node26210;
														assign node26210 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26213 = (inp[11]) ? node26215 : 16'b0000000001111111;
															assign node26215 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26218 = (inp[10]) ? node26224 : node26219;
													assign node26219 = (inp[4]) ? node26221 : 16'b0000000001111111;
														assign node26221 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26224 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node26227 = (inp[8]) ? node26361 : node26228;
									assign node26228 = (inp[6]) ? node26290 : node26229;
										assign node26229 = (inp[10]) ? node26265 : node26230;
											assign node26230 = (inp[4]) ? node26248 : node26231;
												assign node26231 = (inp[15]) ? node26241 : node26232;
													assign node26232 = (inp[7]) ? node26236 : node26233;
														assign node26233 = (inp[11]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node26236 = (inp[11]) ? 16'b0000000111111111 : node26237;
															assign node26237 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26241 = (inp[11]) ? node26245 : node26242;
														assign node26242 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26245 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26248 = (inp[11]) ? node26258 : node26249;
													assign node26249 = (inp[9]) ? node26255 : node26250;
														assign node26250 = (inp[7]) ? 16'b0000000111111111 : node26251;
															assign node26251 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26255 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26258 = (inp[15]) ? 16'b0000000001111111 : node26259;
														assign node26259 = (inp[7]) ? 16'b0000000011111111 : node26260;
															assign node26260 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node26265 = (inp[7]) ? node26281 : node26266;
												assign node26266 = (inp[4]) ? node26274 : node26267;
													assign node26267 = (inp[9]) ? node26271 : node26268;
														assign node26268 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26271 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26274 = (inp[11]) ? node26278 : node26275;
														assign node26275 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26278 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26281 = (inp[9]) ? node26287 : node26282;
													assign node26282 = (inp[2]) ? node26284 : 16'b0000000011111111;
														assign node26284 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26287 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node26290 = (inp[11]) ? node26318 : node26291;
											assign node26291 = (inp[15]) ? node26307 : node26292;
												assign node26292 = (inp[4]) ? node26300 : node26293;
													assign node26293 = (inp[10]) ? node26295 : 16'b0000001111111111;
														assign node26295 = (inp[2]) ? 16'b0000000011111111 : node26296;
															assign node26296 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26300 = (inp[9]) ? node26304 : node26301;
														assign node26301 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26304 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26307 = (inp[2]) ? node26313 : node26308;
													assign node26308 = (inp[7]) ? 16'b0000000011111111 : node26309;
														assign node26309 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26313 = (inp[9]) ? 16'b0000000001111111 : node26314;
														assign node26314 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node26318 = (inp[9]) ? node26340 : node26319;
												assign node26319 = (inp[4]) ? node26327 : node26320;
													assign node26320 = (inp[2]) ? node26324 : node26321;
														assign node26321 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26324 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26327 = (inp[15]) ? node26335 : node26328;
														assign node26328 = (inp[2]) ? node26330 : 16'b0000000011111111;
															assign node26330 = (inp[10]) ? 16'b0000000001111111 : node26331;
																assign node26331 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26335 = (inp[10]) ? node26337 : 16'b0000000001111111;
															assign node26337 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26340 = (inp[10]) ? node26350 : node26341;
													assign node26341 = (inp[7]) ? node26343 : 16'b0000000011111111;
														assign node26343 = (inp[2]) ? 16'b0000000000111111 : node26344;
															assign node26344 = (inp[4]) ? 16'b0000000001111111 : node26345;
																assign node26345 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26350 = (inp[2]) ? node26358 : node26351;
														assign node26351 = (inp[15]) ? node26353 : 16'b0000000001111111;
															assign node26353 = (inp[7]) ? 16'b0000000000111111 : node26354;
																assign node26354 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26358 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node26361 = (inp[7]) ? node26423 : node26362;
										assign node26362 = (inp[4]) ? node26394 : node26363;
											assign node26363 = (inp[11]) ? node26375 : node26364;
												assign node26364 = (inp[10]) ? node26370 : node26365;
													assign node26365 = (inp[9]) ? 16'b0000000111111111 : node26366;
														assign node26366 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26370 = (inp[15]) ? 16'b0000000011111111 : node26371;
														assign node26371 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26375 = (inp[9]) ? node26387 : node26376;
													assign node26376 = (inp[15]) ? node26382 : node26377;
														assign node26377 = (inp[10]) ? node26379 : 16'b0000000111111111;
															assign node26379 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26382 = (inp[10]) ? 16'b0000000001111111 : node26383;
															assign node26383 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26387 = (inp[6]) ? node26389 : 16'b0000000001111111;
														assign node26389 = (inp[2]) ? 16'b0000000000111111 : node26390;
															assign node26390 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26394 = (inp[11]) ? node26410 : node26395;
												assign node26395 = (inp[2]) ? node26405 : node26396;
													assign node26396 = (inp[15]) ? node26398 : 16'b0000000011111111;
														assign node26398 = (inp[6]) ? 16'b0000000001111111 : node26399;
															assign node26399 = (inp[9]) ? node26401 : 16'b0000000011111111;
																assign node26401 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26405 = (inp[9]) ? 16'b0000000000111111 : node26406;
														assign node26406 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26410 = (inp[10]) ? node26414 : node26411;
													assign node26411 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26414 = (inp[15]) ? node26416 : 16'b0000000000111111;
														assign node26416 = (inp[6]) ? 16'b0000000000011111 : node26417;
															assign node26417 = (inp[2]) ? node26419 : 16'b0000000001111111;
																assign node26419 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node26423 = (inp[11]) ? node26451 : node26424;
											assign node26424 = (inp[2]) ? node26436 : node26425;
												assign node26425 = (inp[10]) ? node26433 : node26426;
													assign node26426 = (inp[6]) ? 16'b0000000001111111 : node26427;
														assign node26427 = (inp[4]) ? 16'b0000000011111111 : node26428;
															assign node26428 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26433 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26436 = (inp[10]) ? node26444 : node26437;
													assign node26437 = (inp[6]) ? node26439 : 16'b0000000001111111;
														assign node26439 = (inp[4]) ? 16'b0000000000011111 : node26440;
															assign node26440 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26444 = (inp[4]) ? node26446 : 16'b0000000000111111;
														assign node26446 = (inp[6]) ? 16'b0000000000011111 : node26447;
															assign node26447 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26451 = (inp[2]) ? node26469 : node26452;
												assign node26452 = (inp[9]) ? node26462 : node26453;
													assign node26453 = (inp[10]) ? node26455 : 16'b0000000001111111;
														assign node26455 = (inp[4]) ? 16'b0000000000111111 : node26456;
															assign node26456 = (inp[15]) ? node26458 : 16'b0000000001111111;
																assign node26458 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26462 = (inp[15]) ? node26464 : 16'b0000000000111111;
														assign node26464 = (inp[4]) ? node26466 : 16'b0000000000111111;
															assign node26466 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node26469 = (inp[10]) ? node26479 : node26470;
													assign node26470 = (inp[4]) ? node26476 : node26471;
														assign node26471 = (inp[6]) ? 16'b0000000000111111 : node26472;
															assign node26472 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26476 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26479 = (inp[9]) ? node26483 : node26480;
														assign node26480 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26483 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node26486 = (inp[4]) ? node26728 : node26487;
								assign node26487 = (inp[2]) ? node26611 : node26488;
									assign node26488 = (inp[8]) ? node26558 : node26489;
										assign node26489 = (inp[7]) ? node26529 : node26490;
											assign node26490 = (inp[11]) ? node26510 : node26491;
												assign node26491 = (inp[15]) ? node26501 : node26492;
													assign node26492 = (inp[9]) ? node26498 : node26493;
														assign node26493 = (inp[12]) ? 16'b0000001111111111 : node26494;
															assign node26494 = (inp[6]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node26498 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26501 = (inp[10]) ? node26505 : node26502;
														assign node26502 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26505 = (inp[6]) ? node26507 : 16'b0000000111111111;
															assign node26507 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26510 = (inp[10]) ? node26524 : node26511;
													assign node26511 = (inp[6]) ? node26519 : node26512;
														assign node26512 = (inp[9]) ? 16'b0000000111111111 : node26513;
															assign node26513 = (inp[12]) ? node26515 : 16'b0000001111111111;
																assign node26515 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26519 = (inp[12]) ? node26521 : 16'b0000000111111111;
															assign node26521 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26524 = (inp[12]) ? 16'b0000000011111111 : node26525;
														assign node26525 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node26529 = (inp[15]) ? node26545 : node26530;
												assign node26530 = (inp[9]) ? node26536 : node26531;
													assign node26531 = (inp[6]) ? 16'b0000000111111111 : node26532;
														assign node26532 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26536 = (inp[12]) ? node26542 : node26537;
														assign node26537 = (inp[6]) ? node26539 : 16'b0000000111111111;
															assign node26539 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26542 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node26545 = (inp[6]) ? node26553 : node26546;
													assign node26546 = (inp[9]) ? node26548 : 16'b0000000011111111;
														assign node26548 = (inp[10]) ? node26550 : 16'b0000000011111111;
															assign node26550 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26553 = (inp[9]) ? 16'b0000000000111111 : node26554;
														assign node26554 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node26558 = (inp[9]) ? node26586 : node26559;
											assign node26559 = (inp[6]) ? node26573 : node26560;
												assign node26560 = (inp[15]) ? node26562 : 16'b0000000111111111;
													assign node26562 = (inp[11]) ? node26570 : node26563;
														assign node26563 = (inp[7]) ? 16'b0000000011111111 : node26564;
															assign node26564 = (inp[10]) ? 16'b0000000111111111 : node26565;
																assign node26565 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26570 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26573 = (inp[15]) ? node26581 : node26574;
													assign node26574 = (inp[10]) ? 16'b0000000011111111 : node26575;
														assign node26575 = (inp[7]) ? 16'b0000000011111111 : node26576;
															assign node26576 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26581 = (inp[10]) ? node26583 : 16'b0000000011111111;
														assign node26583 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26586 = (inp[11]) ? node26600 : node26587;
												assign node26587 = (inp[12]) ? node26593 : node26588;
													assign node26588 = (inp[7]) ? node26590 : 16'b0000000011111111;
														assign node26590 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26593 = (inp[10]) ? node26597 : node26594;
														assign node26594 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node26597 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26600 = (inp[12]) ? node26608 : node26601;
													assign node26601 = (inp[10]) ? node26605 : node26602;
														assign node26602 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26605 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26608 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node26611 = (inp[9]) ? node26675 : node26612;
										assign node26612 = (inp[15]) ? node26638 : node26613;
											assign node26613 = (inp[6]) ? node26621 : node26614;
												assign node26614 = (inp[12]) ? 16'b0000000011111111 : node26615;
													assign node26615 = (inp[7]) ? 16'b0000000011111111 : node26616;
														assign node26616 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node26621 = (inp[10]) ? node26631 : node26622;
													assign node26622 = (inp[11]) ? node26626 : node26623;
														assign node26623 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26626 = (inp[7]) ? node26628 : 16'b0000000011111111;
															assign node26628 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26631 = (inp[11]) ? node26635 : node26632;
														assign node26632 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26635 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26638 = (inp[7]) ? node26658 : node26639;
												assign node26639 = (inp[12]) ? node26647 : node26640;
													assign node26640 = (inp[6]) ? 16'b0000000011111111 : node26641;
														assign node26641 = (inp[11]) ? node26643 : 16'b0000000111111111;
															assign node26643 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26647 = (inp[6]) ? node26653 : node26648;
														assign node26648 = (inp[10]) ? 16'b0000000001111111 : node26649;
															assign node26649 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26653 = (inp[8]) ? 16'b0000000000111111 : node26654;
															assign node26654 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26658 = (inp[12]) ? 16'b0000000000111111 : node26659;
													assign node26659 = (inp[10]) ? node26665 : node26660;
														assign node26660 = (inp[11]) ? 16'b0000000001111111 : node26661;
															assign node26661 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26665 = (inp[11]) ? node26667 : 16'b0000000001111111;
															assign node26667 = (inp[6]) ? node26671 : node26668;
																assign node26668 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
																assign node26671 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node26675 = (inp[10]) ? node26695 : node26676;
											assign node26676 = (inp[7]) ? node26680 : node26677;
												assign node26677 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26680 = (inp[6]) ? node26686 : node26681;
													assign node26681 = (inp[11]) ? 16'b0000000001111111 : node26682;
														assign node26682 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26686 = (inp[8]) ? node26692 : node26687;
														assign node26687 = (inp[15]) ? node26689 : 16'b0000000001111111;
															assign node26689 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26692 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26695 = (inp[12]) ? node26713 : node26696;
												assign node26696 = (inp[15]) ? node26704 : node26697;
													assign node26697 = (inp[11]) ? 16'b0000000000111111 : node26698;
														assign node26698 = (inp[7]) ? 16'b0000000001111111 : node26699;
															assign node26699 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26704 = (inp[6]) ? node26710 : node26705;
														assign node26705 = (inp[7]) ? 16'b0000000000111111 : node26706;
															assign node26706 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26710 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26713 = (inp[6]) ? node26719 : node26714;
													assign node26714 = (inp[15]) ? 16'b0000000000111111 : node26715;
														assign node26715 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26719 = (inp[11]) ? 16'b0000000000001111 : node26720;
														assign node26720 = (inp[7]) ? node26724 : node26721;
															assign node26721 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node26724 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node26728 = (inp[7]) ? node26850 : node26729;
									assign node26729 = (inp[8]) ? node26799 : node26730;
										assign node26730 = (inp[9]) ? node26760 : node26731;
											assign node26731 = (inp[2]) ? node26749 : node26732;
												assign node26732 = (inp[6]) ? node26738 : node26733;
													assign node26733 = (inp[11]) ? 16'b0000000111111111 : node26734;
														assign node26734 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node26738 = (inp[12]) ? node26742 : node26739;
														assign node26739 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26742 = (inp[11]) ? 16'b0000000001111111 : node26743;
															assign node26743 = (inp[10]) ? node26745 : 16'b0000000011111111;
																assign node26745 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26749 = (inp[15]) ? 16'b0000000001111111 : node26750;
													assign node26750 = (inp[6]) ? node26752 : 16'b0000000011111111;
														assign node26752 = (inp[10]) ? node26754 : 16'b0000000011111111;
															assign node26754 = (inp[12]) ? 16'b0000000001111111 : node26755;
																assign node26755 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node26760 = (inp[12]) ? node26782 : node26761;
												assign node26761 = (inp[2]) ? node26769 : node26762;
													assign node26762 = (inp[6]) ? node26766 : node26763;
														assign node26763 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26766 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26769 = (inp[15]) ? 16'b0000000000111111 : node26770;
														assign node26770 = (inp[6]) ? node26776 : node26771;
															assign node26771 = (inp[10]) ? node26773 : 16'b0000000011111111;
																assign node26773 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node26776 = (inp[11]) ? node26778 : 16'b0000000001111111;
																assign node26778 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26782 = (inp[15]) ? node26790 : node26783;
													assign node26783 = (inp[11]) ? node26787 : node26784;
														assign node26784 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26787 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26790 = (inp[2]) ? node26796 : node26791;
														assign node26791 = (inp[10]) ? 16'b0000000000111111 : node26792;
															assign node26792 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26796 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node26799 = (inp[12]) ? node26825 : node26800;
											assign node26800 = (inp[10]) ? node26814 : node26801;
												assign node26801 = (inp[2]) ? node26809 : node26802;
													assign node26802 = (inp[15]) ? node26806 : node26803;
														assign node26803 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node26806 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26809 = (inp[15]) ? node26811 : 16'b0000000001111111;
														assign node26811 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node26814 = (inp[15]) ? node26816 : 16'b0000000001111111;
													assign node26816 = (inp[6]) ? 16'b0000000000111111 : node26817;
														assign node26817 = (inp[11]) ? 16'b0000000000111111 : node26818;
															assign node26818 = (inp[9]) ? node26820 : 16'b0000000001111111;
																assign node26820 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26825 = (inp[11]) ? node26831 : node26826;
												assign node26826 = (inp[10]) ? node26828 : 16'b0000000001111111;
													assign node26828 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26831 = (inp[10]) ? node26843 : node26832;
													assign node26832 = (inp[6]) ? node26840 : node26833;
														assign node26833 = (inp[2]) ? node26835 : 16'b0000000001111111;
															assign node26835 = (inp[15]) ? 16'b0000000000111111 : node26836;
																assign node26836 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26840 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26843 = (inp[15]) ? node26845 : 16'b0000000000011111;
														assign node26845 = (inp[6]) ? node26847 : 16'b0000000000011111;
															assign node26847 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node26850 = (inp[6]) ? node26922 : node26851;
										assign node26851 = (inp[15]) ? node26877 : node26852;
											assign node26852 = (inp[10]) ? node26866 : node26853;
												assign node26853 = (inp[11]) ? node26861 : node26854;
													assign node26854 = (inp[2]) ? 16'b0000000011111111 : node26855;
														assign node26855 = (inp[12]) ? node26857 : 16'b0000000111111111;
															assign node26857 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26861 = (inp[8]) ? 16'b0000000000111111 : node26862;
														assign node26862 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26866 = (inp[2]) ? 16'b0000000000111111 : node26867;
													assign node26867 = (inp[8]) ? node26869 : 16'b0000000001111111;
														assign node26869 = (inp[12]) ? 16'b0000000000111111 : node26870;
															assign node26870 = (inp[9]) ? node26872 : 16'b0000000001111111;
																assign node26872 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26877 = (inp[9]) ? node26897 : node26878;
												assign node26878 = (inp[10]) ? node26884 : node26879;
													assign node26879 = (inp[8]) ? node26881 : 16'b0000000001111111;
														assign node26881 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26884 = (inp[11]) ? node26894 : node26885;
														assign node26885 = (inp[2]) ? node26889 : node26886;
															assign node26886 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node26889 = (inp[8]) ? 16'b0000000000111111 : node26890;
																assign node26890 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26894 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26897 = (inp[11]) ? node26905 : node26898;
													assign node26898 = (inp[12]) ? node26902 : node26899;
														assign node26899 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26902 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26905 = (inp[12]) ? node26917 : node26906;
														assign node26906 = (inp[8]) ? node26912 : node26907;
															assign node26907 = (inp[2]) ? node26909 : 16'b0000000000111111;
																assign node26909 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node26912 = (inp[10]) ? 16'b0000000000011111 : node26913;
																assign node26913 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26917 = (inp[10]) ? node26919 : 16'b0000000000011111;
															assign node26919 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node26922 = (inp[12]) ? node26958 : node26923;
											assign node26923 = (inp[11]) ? node26939 : node26924;
												assign node26924 = (inp[9]) ? node26930 : node26925;
													assign node26925 = (inp[10]) ? node26927 : 16'b0000000011111111;
														assign node26927 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26930 = (inp[8]) ? node26936 : node26931;
														assign node26931 = (inp[10]) ? node26933 : 16'b0000000001111111;
															assign node26933 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26936 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26939 = (inp[9]) ? node26951 : node26940;
													assign node26940 = (inp[10]) ? node26944 : node26941;
														assign node26941 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26944 = (inp[15]) ? node26946 : 16'b0000000000111111;
															assign node26946 = (inp[8]) ? node26948 : 16'b0000000000111111;
																assign node26948 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node26951 = (inp[15]) ? node26953 : 16'b0000000000011111;
														assign node26953 = (inp[2]) ? node26955 : 16'b0000000000011111;
															assign node26955 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node26958 = (inp[2]) ? node26974 : node26959;
												assign node26959 = (inp[8]) ? node26969 : node26960;
													assign node26960 = (inp[9]) ? node26964 : node26961;
														assign node26961 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26964 = (inp[15]) ? 16'b0000000000011111 : node26965;
															assign node26965 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26969 = (inp[9]) ? 16'b0000000000011111 : node26970;
														assign node26970 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node26974 = (inp[11]) ? node26982 : node26975;
													assign node26975 = (inp[15]) ? node26977 : 16'b0000000000011111;
														assign node26977 = (inp[10]) ? node26979 : 16'b0000000000011111;
															assign node26979 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node26982 = (inp[15]) ? node26984 : 16'b0000000000001111;
														assign node26984 = (inp[10]) ? 16'b0000000000000011 : node26985;
															assign node26985 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node26989 = (inp[15]) ? node28017 : node26990;
						assign node26990 = (inp[7]) ? node27486 : node26991;
							assign node26991 = (inp[4]) ? node27245 : node26992;
								assign node26992 = (inp[6]) ? node27116 : node26993;
									assign node26993 = (inp[12]) ? node27063 : node26994;
										assign node26994 = (inp[2]) ? node27032 : node26995;
											assign node26995 = (inp[10]) ? node27015 : node26996;
												assign node26996 = (inp[14]) ? node27008 : node26997;
													assign node26997 = (inp[1]) ? node27001 : node26998;
														assign node26998 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node27001 = (inp[11]) ? 16'b0000001111111111 : node27002;
															assign node27002 = (inp[9]) ? node27004 : 16'b0000011111111111;
																assign node27004 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node27008 = (inp[9]) ? node27012 : node27009;
														assign node27009 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27012 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node27015 = (inp[9]) ? node27023 : node27016;
													assign node27016 = (inp[1]) ? node27020 : node27017;
														assign node27017 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node27020 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27023 = (inp[11]) ? node27027 : node27024;
														assign node27024 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27027 = (inp[14]) ? node27029 : 16'b0000000111111111;
															assign node27029 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27032 = (inp[11]) ? node27046 : node27033;
												assign node27033 = (inp[8]) ? node27039 : node27034;
													assign node27034 = (inp[1]) ? 16'b0000001111111111 : node27035;
														assign node27035 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node27039 = (inp[9]) ? node27043 : node27040;
														assign node27040 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27043 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27046 = (inp[10]) ? node27054 : node27047;
													assign node27047 = (inp[14]) ? node27051 : node27048;
														assign node27048 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27051 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node27054 = (inp[8]) ? node27060 : node27055;
														assign node27055 = (inp[9]) ? 16'b0000000011111111 : node27056;
															assign node27056 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27060 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node27063 = (inp[9]) ? node27089 : node27064;
											assign node27064 = (inp[10]) ? node27076 : node27065;
												assign node27065 = (inp[14]) ? node27071 : node27066;
													assign node27066 = (inp[1]) ? 16'b0000001111111111 : node27067;
														assign node27067 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node27071 = (inp[11]) ? node27073 : 16'b0000001111111111;
														assign node27073 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27076 = (inp[11]) ? node27078 : 16'b0000000111111111;
													assign node27078 = (inp[14]) ? node27082 : node27079;
														assign node27079 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27082 = (inp[1]) ? 16'b0000000001111111 : node27083;
															assign node27083 = (inp[8]) ? 16'b0000000011111111 : node27084;
																assign node27084 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27089 = (inp[2]) ? node27101 : node27090;
												assign node27090 = (inp[10]) ? node27096 : node27091;
													assign node27091 = (inp[1]) ? node27093 : 16'b0000001111111111;
														assign node27093 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27096 = (inp[14]) ? 16'b0000000011111111 : node27097;
														assign node27097 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27101 = (inp[14]) ? node27109 : node27102;
													assign node27102 = (inp[11]) ? node27106 : node27103;
														assign node27103 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27106 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27109 = (inp[1]) ? node27113 : node27110;
														assign node27110 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27113 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node27116 = (inp[8]) ? node27178 : node27117;
										assign node27117 = (inp[9]) ? node27149 : node27118;
											assign node27118 = (inp[2]) ? node27130 : node27119;
												assign node27119 = (inp[14]) ? node27121 : 16'b0000001111111111;
													assign node27121 = (inp[1]) ? node27125 : node27122;
														assign node27122 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27125 = (inp[11]) ? node27127 : 16'b0000000111111111;
															assign node27127 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27130 = (inp[14]) ? node27142 : node27131;
													assign node27131 = (inp[10]) ? node27137 : node27132;
														assign node27132 = (inp[11]) ? 16'b0000000111111111 : node27133;
															assign node27133 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27137 = (inp[11]) ? node27139 : 16'b0000000111111111;
															assign node27139 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27142 = (inp[12]) ? 16'b0000000001111111 : node27143;
														assign node27143 = (inp[11]) ? node27145 : 16'b0000000111111111;
															assign node27145 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27149 = (inp[10]) ? node27163 : node27150;
												assign node27150 = (inp[12]) ? node27154 : node27151;
													assign node27151 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27154 = (inp[1]) ? 16'b0000000011111111 : node27155;
														assign node27155 = (inp[11]) ? 16'b0000000011111111 : node27156;
															assign node27156 = (inp[14]) ? node27158 : 16'b0000000111111111;
																assign node27158 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27163 = (inp[14]) ? node27171 : node27164;
													assign node27164 = (inp[2]) ? node27166 : 16'b0000001111111111;
														assign node27166 = (inp[1]) ? 16'b0000000011111111 : node27167;
															assign node27167 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27171 = (inp[12]) ? 16'b0000000001111111 : node27172;
														assign node27172 = (inp[1]) ? node27174 : 16'b0000000011111111;
															assign node27174 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node27178 = (inp[12]) ? node27212 : node27179;
											assign node27179 = (inp[2]) ? node27199 : node27180;
												assign node27180 = (inp[14]) ? node27188 : node27181;
													assign node27181 = (inp[9]) ? 16'b0000000111111111 : node27182;
														assign node27182 = (inp[1]) ? node27184 : 16'b0000001111111111;
															assign node27184 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27188 = (inp[9]) ? node27194 : node27189;
														assign node27189 = (inp[10]) ? node27191 : 16'b0000000111111111;
															assign node27191 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27194 = (inp[11]) ? node27196 : 16'b0000000011111111;
															assign node27196 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27199 = (inp[11]) ? node27201 : 16'b0000000011111111;
													assign node27201 = (inp[9]) ? node27207 : node27202;
														assign node27202 = (inp[1]) ? 16'b0000000001111111 : node27203;
															assign node27203 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27207 = (inp[14]) ? 16'b0000000000111111 : node27208;
															assign node27208 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27212 = (inp[1]) ? node27232 : node27213;
												assign node27213 = (inp[14]) ? node27221 : node27214;
													assign node27214 = (inp[2]) ? node27218 : node27215;
														assign node27215 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27218 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27221 = (inp[10]) ? node27229 : node27222;
														assign node27222 = (inp[2]) ? node27224 : 16'b0000000011111111;
															assign node27224 = (inp[9]) ? 16'b0000000001111111 : node27225;
																assign node27225 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27229 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27232 = (inp[14]) ? node27240 : node27233;
													assign node27233 = (inp[2]) ? node27235 : 16'b0000000001111111;
														assign node27235 = (inp[11]) ? node27237 : 16'b0000000001111111;
															assign node27237 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27240 = (inp[9]) ? node27242 : 16'b0000000000111111;
														assign node27242 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node27245 = (inp[9]) ? node27365 : node27246;
									assign node27246 = (inp[14]) ? node27302 : node27247;
										assign node27247 = (inp[10]) ? node27273 : node27248;
											assign node27248 = (inp[12]) ? node27264 : node27249;
												assign node27249 = (inp[11]) ? node27257 : node27250;
													assign node27250 = (inp[6]) ? node27254 : node27251;
														assign node27251 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node27254 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27257 = (inp[8]) ? node27261 : node27258;
														assign node27258 = (inp[6]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node27261 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27264 = (inp[8]) ? node27266 : 16'b0000000111111111;
													assign node27266 = (inp[2]) ? node27268 : 16'b0000000111111111;
														assign node27268 = (inp[1]) ? 16'b0000000011111111 : node27269;
															assign node27269 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27273 = (inp[12]) ? node27283 : node27274;
												assign node27274 = (inp[2]) ? node27280 : node27275;
													assign node27275 = (inp[1]) ? node27277 : 16'b0000000111111111;
														assign node27277 = (inp[6]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node27280 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27283 = (inp[11]) ? node27291 : node27284;
													assign node27284 = (inp[6]) ? node27288 : node27285;
														assign node27285 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27288 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27291 = (inp[1]) ? node27295 : node27292;
														assign node27292 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node27295 = (inp[6]) ? 16'b0000000000011111 : node27296;
															assign node27296 = (inp[8]) ? node27298 : 16'b0000000001111111;
																assign node27298 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node27302 = (inp[2]) ? node27332 : node27303;
											assign node27303 = (inp[12]) ? node27321 : node27304;
												assign node27304 = (inp[8]) ? node27312 : node27305;
													assign node27305 = (inp[1]) ? 16'b0000000111111111 : node27306;
														assign node27306 = (inp[11]) ? 16'b0000000111111111 : node27307;
															assign node27307 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node27312 = (inp[11]) ? node27318 : node27313;
														assign node27313 = (inp[6]) ? 16'b0000000011111111 : node27314;
															assign node27314 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27318 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27321 = (inp[1]) ? node27323 : 16'b0000000011111111;
													assign node27323 = (inp[10]) ? node27327 : node27324;
														assign node27324 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node27327 = (inp[11]) ? node27329 : 16'b0000000001111111;
															assign node27329 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27332 = (inp[6]) ? node27348 : node27333;
												assign node27333 = (inp[12]) ? node27345 : node27334;
													assign node27334 = (inp[1]) ? node27340 : node27335;
														assign node27335 = (inp[10]) ? 16'b0000000011111111 : node27336;
															assign node27336 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27340 = (inp[11]) ? 16'b0000000001111111 : node27341;
															assign node27341 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node27345 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node27348 = (inp[8]) ? node27350 : 16'b0000000001111111;
													assign node27350 = (inp[1]) ? node27362 : node27351;
														assign node27351 = (inp[12]) ? node27357 : node27352;
															assign node27352 = (inp[11]) ? node27354 : 16'b0000000001111111;
																assign node27354 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node27357 = (inp[10]) ? 16'b0000000000111111 : node27358;
																assign node27358 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27362 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node27365 = (inp[2]) ? node27437 : node27366;
										assign node27366 = (inp[12]) ? node27394 : node27367;
											assign node27367 = (inp[6]) ? node27379 : node27368;
												assign node27368 = (inp[8]) ? node27374 : node27369;
													assign node27369 = (inp[11]) ? node27371 : 16'b0000001111111111;
														assign node27371 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27374 = (inp[1]) ? node27376 : 16'b0000000011111111;
														assign node27376 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27379 = (inp[11]) ? 16'b0000000001111111 : node27380;
													assign node27380 = (inp[14]) ? node27386 : node27381;
														assign node27381 = (inp[1]) ? 16'b0000000011111111 : node27382;
															assign node27382 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27386 = (inp[10]) ? node27388 : 16'b0000000011111111;
															assign node27388 = (inp[1]) ? 16'b0000000001111111 : node27389;
																assign node27389 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node27394 = (inp[11]) ? node27418 : node27395;
												assign node27395 = (inp[14]) ? node27411 : node27396;
													assign node27396 = (inp[8]) ? node27400 : node27397;
														assign node27397 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27400 = (inp[6]) ? node27406 : node27401;
															assign node27401 = (inp[10]) ? node27403 : 16'b0000000011111111;
																assign node27403 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node27406 = (inp[10]) ? 16'b0000000001111111 : node27407;
																assign node27407 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27411 = (inp[10]) ? 16'b0000000000111111 : node27412;
														assign node27412 = (inp[1]) ? 16'b0000000001111111 : node27413;
															assign node27413 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27418 = (inp[1]) ? node27430 : node27419;
													assign node27419 = (inp[14]) ? node27425 : node27420;
														assign node27420 = (inp[10]) ? node27422 : 16'b0000000011111111;
															assign node27422 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27425 = (inp[8]) ? 16'b0000000000111111 : node27426;
															assign node27426 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27430 = (inp[10]) ? node27432 : 16'b0000000000111111;
														assign node27432 = (inp[8]) ? node27434 : 16'b0000000000111111;
															assign node27434 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node27437 = (inp[10]) ? node27459 : node27438;
											assign node27438 = (inp[1]) ? node27450 : node27439;
												assign node27439 = (inp[14]) ? node27443 : node27440;
													assign node27440 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27443 = (inp[11]) ? node27445 : 16'b0000000011111111;
														assign node27445 = (inp[8]) ? node27447 : 16'b0000000001111111;
															assign node27447 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27450 = (inp[12]) ? 16'b0000000000111111 : node27451;
													assign node27451 = (inp[6]) ? node27455 : node27452;
														assign node27452 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27455 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27459 = (inp[1]) ? node27475 : node27460;
												assign node27460 = (inp[6]) ? node27466 : node27461;
													assign node27461 = (inp[11]) ? node27463 : 16'b0000000001111111;
														assign node27463 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27466 = (inp[11]) ? node27470 : node27467;
														assign node27467 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node27470 = (inp[14]) ? node27472 : 16'b0000000000111111;
															assign node27472 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node27475 = (inp[14]) ? node27479 : node27476;
													assign node27476 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27479 = (inp[6]) ? node27481 : 16'b0000000000011111;
														assign node27481 = (inp[8]) ? 16'b0000000000001111 : node27482;
															assign node27482 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node27486 = (inp[12]) ? node27750 : node27487;
								assign node27487 = (inp[8]) ? node27629 : node27488;
									assign node27488 = (inp[9]) ? node27562 : node27489;
										assign node27489 = (inp[2]) ? node27527 : node27490;
											assign node27490 = (inp[6]) ? node27510 : node27491;
												assign node27491 = (inp[1]) ? node27505 : node27492;
													assign node27492 = (inp[10]) ? node27498 : node27493;
														assign node27493 = (inp[4]) ? node27495 : 16'b0000111111111111;
															assign node27495 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27498 = (inp[4]) ? 16'b0000000111111111 : node27499;
															assign node27499 = (inp[14]) ? 16'b0000001111111111 : node27500;
																assign node27500 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node27505 = (inp[4]) ? node27507 : 16'b0000000111111111;
														assign node27507 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27510 = (inp[11]) ? node27520 : node27511;
													assign node27511 = (inp[1]) ? node27513 : 16'b0000001111111111;
														assign node27513 = (inp[4]) ? 16'b0000000011111111 : node27514;
															assign node27514 = (inp[14]) ? 16'b0000000111111111 : node27515;
																assign node27515 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27520 = (inp[10]) ? 16'b0000000011111111 : node27521;
														assign node27521 = (inp[4]) ? 16'b0000000011111111 : node27522;
															assign node27522 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27527 = (inp[10]) ? node27549 : node27528;
												assign node27528 = (inp[4]) ? node27542 : node27529;
													assign node27529 = (inp[6]) ? node27537 : node27530;
														assign node27530 = (inp[11]) ? node27532 : 16'b0000000111111111;
															assign node27532 = (inp[1]) ? node27534 : 16'b0000000111111111;
																assign node27534 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27537 = (inp[1]) ? 16'b0000000111111111 : node27538;
															assign node27538 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27542 = (inp[11]) ? 16'b0000000001111111 : node27543;
														assign node27543 = (inp[1]) ? 16'b0000000001111111 : node27544;
															assign node27544 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node27549 = (inp[14]) ? node27555 : node27550;
													assign node27550 = (inp[1]) ? node27552 : 16'b0000000011111111;
														assign node27552 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27555 = (inp[11]) ? 16'b0000000001111111 : node27556;
														assign node27556 = (inp[6]) ? 16'b0000000001111111 : node27557;
															assign node27557 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node27562 = (inp[10]) ? node27598 : node27563;
											assign node27563 = (inp[2]) ? node27579 : node27564;
												assign node27564 = (inp[14]) ? node27574 : node27565;
													assign node27565 = (inp[6]) ? node27567 : 16'b0000000111111111;
														assign node27567 = (inp[11]) ? node27569 : 16'b0000000111111111;
															assign node27569 = (inp[4]) ? 16'b0000000011111111 : node27570;
																assign node27570 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27574 = (inp[6]) ? 16'b0000000001111111 : node27575;
														assign node27575 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node27579 = (inp[11]) ? node27589 : node27580;
													assign node27580 = (inp[6]) ? node27582 : 16'b0000000111111111;
														assign node27582 = (inp[4]) ? node27584 : 16'b0000000011111111;
															assign node27584 = (inp[1]) ? 16'b0000000001111111 : node27585;
																assign node27585 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27589 = (inp[1]) ? node27593 : node27590;
														assign node27590 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27593 = (inp[14]) ? node27595 : 16'b0000000001111111;
															assign node27595 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27598 = (inp[1]) ? node27614 : node27599;
												assign node27599 = (inp[6]) ? node27607 : node27600;
													assign node27600 = (inp[2]) ? node27604 : node27601;
														assign node27601 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27604 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27607 = (inp[4]) ? node27611 : node27608;
														assign node27608 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27611 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27614 = (inp[14]) ? node27624 : node27615;
													assign node27615 = (inp[11]) ? node27619 : node27616;
														assign node27616 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node27619 = (inp[4]) ? node27621 : 16'b0000000001111111;
															assign node27621 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27624 = (inp[6]) ? node27626 : 16'b0000000000111111;
														assign node27626 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node27629 = (inp[6]) ? node27685 : node27630;
										assign node27630 = (inp[14]) ? node27660 : node27631;
											assign node27631 = (inp[4]) ? node27645 : node27632;
												assign node27632 = (inp[1]) ? node27638 : node27633;
													assign node27633 = (inp[10]) ? 16'b0000000011111111 : node27634;
														assign node27634 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27638 = (inp[9]) ? node27642 : node27639;
														assign node27639 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27642 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27645 = (inp[10]) ? node27655 : node27646;
													assign node27646 = (inp[11]) ? node27652 : node27647;
														assign node27647 = (inp[1]) ? 16'b0000000011111111 : node27648;
															assign node27648 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27652 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27655 = (inp[1]) ? 16'b0000000001111111 : node27656;
														assign node27656 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node27660 = (inp[1]) ? node27666 : node27661;
												assign node27661 = (inp[11]) ? node27663 : 16'b0000000011111111;
													assign node27663 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node27666 = (inp[10]) ? node27678 : node27667;
													assign node27667 = (inp[11]) ? node27675 : node27668;
														assign node27668 = (inp[9]) ? node27670 : 16'b0000000001111111;
															assign node27670 = (inp[2]) ? node27672 : 16'b0000000001111111;
																assign node27672 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27675 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27678 = (inp[4]) ? node27682 : node27679;
														assign node27679 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27682 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node27685 = (inp[11]) ? node27715 : node27686;
											assign node27686 = (inp[2]) ? node27704 : node27687;
												assign node27687 = (inp[9]) ? node27697 : node27688;
													assign node27688 = (inp[10]) ? 16'b0000000111111111 : node27689;
														assign node27689 = (inp[4]) ? node27691 : 16'b0000000011111111;
															assign node27691 = (inp[1]) ? node27693 : 16'b0000000011111111;
																assign node27693 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27697 = (inp[4]) ? node27701 : node27698;
														assign node27698 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27701 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27704 = (inp[9]) ? 16'b0000000000111111 : node27705;
													assign node27705 = (inp[14]) ? node27709 : node27706;
														assign node27706 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27709 = (inp[4]) ? 16'b0000000000111111 : node27710;
															assign node27710 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27715 = (inp[4]) ? node27735 : node27716;
												assign node27716 = (inp[2]) ? node27726 : node27717;
													assign node27717 = (inp[9]) ? node27723 : node27718;
														assign node27718 = (inp[14]) ? 16'b0000000001111111 : node27719;
															assign node27719 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27723 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node27726 = (inp[14]) ? node27732 : node27727;
														assign node27727 = (inp[9]) ? 16'b0000000000111111 : node27728;
															assign node27728 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27732 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node27735 = (inp[2]) ? node27743 : node27736;
													assign node27736 = (inp[9]) ? node27738 : 16'b0000000000111111;
														assign node27738 = (inp[10]) ? 16'b0000000000011111 : node27739;
															assign node27739 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27743 = (inp[14]) ? node27745 : 16'b0000000000011111;
														assign node27745 = (inp[10]) ? node27747 : 16'b0000000000011111;
															assign node27747 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node27750 = (inp[11]) ? node27900 : node27751;
									assign node27751 = (inp[6]) ? node27815 : node27752;
										assign node27752 = (inp[2]) ? node27788 : node27753;
											assign node27753 = (inp[10]) ? node27769 : node27754;
												assign node27754 = (inp[9]) ? node27760 : node27755;
													assign node27755 = (inp[1]) ? node27757 : 16'b0000001111111111;
														assign node27757 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27760 = (inp[14]) ? node27766 : node27761;
														assign node27761 = (inp[4]) ? node27763 : 16'b0000000011111111;
															assign node27763 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27766 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27769 = (inp[1]) ? node27777 : node27770;
													assign node27770 = (inp[8]) ? node27772 : 16'b0000000111111111;
														assign node27772 = (inp[9]) ? node27774 : 16'b0000000011111111;
															assign node27774 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27777 = (inp[4]) ? node27785 : node27778;
														assign node27778 = (inp[8]) ? node27780 : 16'b0000000011111111;
															assign node27780 = (inp[9]) ? 16'b0000000001111111 : node27781;
																assign node27781 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27785 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27788 = (inp[14]) ? node27804 : node27789;
												assign node27789 = (inp[1]) ? node27797 : node27790;
													assign node27790 = (inp[8]) ? node27792 : 16'b0000000111111111;
														assign node27792 = (inp[10]) ? node27794 : 16'b0000000011111111;
															assign node27794 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27797 = (inp[4]) ? node27801 : node27798;
														assign node27798 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27801 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node27804 = (inp[1]) ? node27812 : node27805;
													assign node27805 = (inp[10]) ? node27807 : 16'b0000000001111111;
														assign node27807 = (inp[9]) ? 16'b0000000000111111 : node27808;
															assign node27808 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27812 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node27815 = (inp[10]) ? node27857 : node27816;
											assign node27816 = (inp[9]) ? node27838 : node27817;
												assign node27817 = (inp[1]) ? node27827 : node27818;
													assign node27818 = (inp[2]) ? node27824 : node27819;
														assign node27819 = (inp[14]) ? 16'b0000000011111111 : node27820;
															assign node27820 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27824 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27827 = (inp[14]) ? node27835 : node27828;
														assign node27828 = (inp[8]) ? 16'b0000000001111111 : node27829;
															assign node27829 = (inp[4]) ? node27831 : 16'b0000000011111111;
																assign node27831 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27835 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27838 = (inp[1]) ? node27850 : node27839;
													assign node27839 = (inp[14]) ? node27847 : node27840;
														assign node27840 = (inp[4]) ? 16'b0000000001111111 : node27841;
															assign node27841 = (inp[8]) ? node27843 : 16'b0000000011111111;
																assign node27843 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27847 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27850 = (inp[2]) ? 16'b0000000000011111 : node27851;
														assign node27851 = (inp[4]) ? 16'b0000000000111111 : node27852;
															assign node27852 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27857 = (inp[2]) ? node27885 : node27858;
												assign node27858 = (inp[4]) ? node27868 : node27859;
													assign node27859 = (inp[8]) ? node27865 : node27860;
														assign node27860 = (inp[1]) ? 16'b0000000011111111 : node27861;
															assign node27861 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27865 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27868 = (inp[14]) ? node27876 : node27869;
														assign node27869 = (inp[8]) ? node27871 : 16'b0000000001111111;
															assign node27871 = (inp[1]) ? 16'b0000000000111111 : node27872;
																assign node27872 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27876 = (inp[1]) ? node27880 : node27877;
															assign node27877 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node27880 = (inp[8]) ? 16'b0000000000011111 : node27881;
																assign node27881 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node27885 = (inp[9]) ? node27891 : node27886;
													assign node27886 = (inp[1]) ? 16'b0000000000111111 : node27887;
														assign node27887 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27891 = (inp[8]) ? node27895 : node27892;
														assign node27892 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27895 = (inp[14]) ? node27897 : 16'b0000000000011111;
															assign node27897 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node27900 = (inp[14]) ? node27956 : node27901;
										assign node27901 = (inp[10]) ? node27925 : node27902;
											assign node27902 = (inp[1]) ? node27912 : node27903;
												assign node27903 = (inp[8]) ? node27905 : 16'b0000000011111111;
													assign node27905 = (inp[9]) ? node27909 : node27906;
														assign node27906 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27909 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27912 = (inp[2]) ? node27918 : node27913;
													assign node27913 = (inp[8]) ? node27915 : 16'b0000000001111111;
														assign node27915 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27918 = (inp[9]) ? node27922 : node27919;
														assign node27919 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node27922 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node27925 = (inp[4]) ? node27939 : node27926;
												assign node27926 = (inp[9]) ? node27934 : node27927;
													assign node27927 = (inp[8]) ? node27929 : 16'b0000000001111111;
														assign node27929 = (inp[2]) ? node27931 : 16'b0000000001111111;
															assign node27931 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27934 = (inp[2]) ? node27936 : 16'b0000000000111111;
														assign node27936 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node27939 = (inp[6]) ? node27947 : node27940;
													assign node27940 = (inp[1]) ? node27942 : 16'b0000000000111111;
														assign node27942 = (inp[9]) ? 16'b0000000000011111 : node27943;
															assign node27943 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27947 = (inp[2]) ? node27949 : 16'b0000000000111111;
														assign node27949 = (inp[1]) ? 16'b0000000000000111 : node27950;
															assign node27950 = (inp[8]) ? node27952 : 16'b0000000000011111;
																assign node27952 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node27956 = (inp[10]) ? node27990 : node27957;
											assign node27957 = (inp[4]) ? node27975 : node27958;
												assign node27958 = (inp[1]) ? node27960 : 16'b0000000001111111;
													assign node27960 = (inp[9]) ? node27968 : node27961;
														assign node27961 = (inp[8]) ? 16'b0000000000111111 : node27962;
															assign node27962 = (inp[6]) ? node27964 : 16'b0000000001111111;
																assign node27964 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27968 = (inp[2]) ? node27970 : 16'b0000000000111111;
															assign node27970 = (inp[6]) ? node27972 : 16'b0000000000111111;
																assign node27972 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node27975 = (inp[6]) ? node27983 : node27976;
													assign node27976 = (inp[8]) ? 16'b0000000000011111 : node27977;
														assign node27977 = (inp[9]) ? node27979 : 16'b0000000000111111;
															assign node27979 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27983 = (inp[9]) ? node27985 : 16'b0000000000011111;
														assign node27985 = (inp[2]) ? 16'b0000000000001111 : node27986;
															assign node27986 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node27990 = (inp[8]) ? node28002 : node27991;
												assign node27991 = (inp[9]) ? node27999 : node27992;
													assign node27992 = (inp[2]) ? 16'b0000000000011111 : node27993;
														assign node27993 = (inp[1]) ? node27995 : 16'b0000000000111111;
															assign node27995 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27999 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node28002 = (inp[2]) ? node28008 : node28003;
													assign node28003 = (inp[6]) ? 16'b0000000000001111 : node28004;
														assign node28004 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28008 = (inp[9]) ? node28010 : 16'b0000000000001111;
														assign node28010 = (inp[1]) ? node28014 : node28011;
															assign node28011 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node28014 = (inp[4]) ? 16'b0000000000000011 : 16'b0000000000000111;
						assign node28017 = (inp[1]) ? node28565 : node28018;
							assign node28018 = (inp[9]) ? node28278 : node28019;
								assign node28019 = (inp[8]) ? node28155 : node28020;
									assign node28020 = (inp[14]) ? node28090 : node28021;
										assign node28021 = (inp[10]) ? node28057 : node28022;
											assign node28022 = (inp[7]) ? node28036 : node28023;
												assign node28023 = (inp[11]) ? node28029 : node28024;
													assign node28024 = (inp[6]) ? 16'b0000001111111111 : node28025;
														assign node28025 = (inp[12]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node28029 = (inp[6]) ? node28033 : node28030;
														assign node28030 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28033 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node28036 = (inp[4]) ? node28044 : node28037;
													assign node28037 = (inp[2]) ? node28039 : 16'b0000000111111111;
														assign node28039 = (inp[12]) ? node28041 : 16'b0000000111111111;
															assign node28041 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28044 = (inp[2]) ? node28052 : node28045;
														assign node28045 = (inp[6]) ? node28047 : 16'b0000000111111111;
															assign node28047 = (inp[11]) ? 16'b0000000011111111 : node28048;
																assign node28048 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28052 = (inp[12]) ? node28054 : 16'b0000000011111111;
															assign node28054 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node28057 = (inp[6]) ? node28075 : node28058;
												assign node28058 = (inp[12]) ? node28070 : node28059;
													assign node28059 = (inp[2]) ? node28065 : node28060;
														assign node28060 = (inp[11]) ? node28062 : 16'b0000001111111111;
															assign node28062 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28065 = (inp[4]) ? node28067 : 16'b0000000111111111;
															assign node28067 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28070 = (inp[2]) ? 16'b0000000011111111 : node28071;
														assign node28071 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node28075 = (inp[11]) ? node28085 : node28076;
													assign node28076 = (inp[12]) ? node28082 : node28077;
														assign node28077 = (inp[7]) ? 16'b0000000011111111 : node28078;
															assign node28078 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28082 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28085 = (inp[2]) ? 16'b0000000001111111 : node28086;
														assign node28086 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node28090 = (inp[2]) ? node28116 : node28091;
											assign node28091 = (inp[7]) ? node28107 : node28092;
												assign node28092 = (inp[11]) ? node28100 : node28093;
													assign node28093 = (inp[10]) ? node28097 : node28094;
														assign node28094 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28097 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28100 = (inp[12]) ? node28104 : node28101;
														assign node28101 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28104 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28107 = (inp[6]) ? node28109 : 16'b0000000011111111;
													assign node28109 = (inp[10]) ? 16'b0000000001111111 : node28110;
														assign node28110 = (inp[12]) ? 16'b0000000001111111 : node28111;
															assign node28111 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node28116 = (inp[4]) ? node28138 : node28117;
												assign node28117 = (inp[11]) ? node28131 : node28118;
													assign node28118 = (inp[6]) ? node28124 : node28119;
														assign node28119 = (inp[12]) ? 16'b0000000011111111 : node28120;
															assign node28120 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28124 = (inp[7]) ? node28126 : 16'b0000000111111111;
															assign node28126 = (inp[10]) ? 16'b0000000001111111 : node28127;
																assign node28127 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28131 = (inp[7]) ? node28135 : node28132;
														assign node28132 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28135 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28138 = (inp[10]) ? node28144 : node28139;
													assign node28139 = (inp[6]) ? 16'b0000000001111111 : node28140;
														assign node28140 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28144 = (inp[7]) ? node28148 : node28145;
														assign node28145 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node28148 = (inp[6]) ? node28150 : 16'b0000000000111111;
															assign node28150 = (inp[11]) ? 16'b0000000000011111 : node28151;
																assign node28151 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node28155 = (inp[7]) ? node28209 : node28156;
										assign node28156 = (inp[2]) ? node28182 : node28157;
											assign node28157 = (inp[6]) ? node28171 : node28158;
												assign node28158 = (inp[10]) ? node28164 : node28159;
													assign node28159 = (inp[11]) ? 16'b0000000111111111 : node28160;
														assign node28160 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node28164 = (inp[4]) ? node28168 : node28165;
														assign node28165 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28168 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28171 = (inp[14]) ? node28177 : node28172;
													assign node28172 = (inp[11]) ? 16'b0000000011111111 : node28173;
														assign node28173 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28177 = (inp[11]) ? 16'b0000000001111111 : node28178;
														assign node28178 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node28182 = (inp[4]) ? node28198 : node28183;
												assign node28183 = (inp[6]) ? node28191 : node28184;
													assign node28184 = (inp[10]) ? 16'b0000000011111111 : node28185;
														assign node28185 = (inp[14]) ? 16'b0000000011111111 : node28186;
															assign node28186 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node28191 = (inp[10]) ? node28195 : node28192;
														assign node28192 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28195 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28198 = (inp[10]) ? node28204 : node28199;
													assign node28199 = (inp[6]) ? node28201 : 16'b0000000001111111;
														assign node28201 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28204 = (inp[12]) ? 16'b0000000000011111 : node28205;
														assign node28205 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node28209 = (inp[4]) ? node28241 : node28210;
											assign node28210 = (inp[11]) ? node28226 : node28211;
												assign node28211 = (inp[14]) ? node28219 : node28212;
													assign node28212 = (inp[2]) ? node28216 : node28213;
														assign node28213 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node28216 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28219 = (inp[12]) ? 16'b0000000000111111 : node28220;
														assign node28220 = (inp[6]) ? 16'b0000000001111111 : node28221;
															assign node28221 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28226 = (inp[12]) ? node28234 : node28227;
													assign node28227 = (inp[2]) ? node28231 : node28228;
														assign node28228 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28231 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28234 = (inp[6]) ? 16'b0000000000111111 : node28235;
														assign node28235 = (inp[14]) ? node28237 : 16'b0000000001111111;
															assign node28237 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28241 = (inp[2]) ? node28261 : node28242;
												assign node28242 = (inp[14]) ? node28254 : node28243;
													assign node28243 = (inp[11]) ? node28247 : node28244;
														assign node28244 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28247 = (inp[10]) ? 16'b0000000000111111 : node28248;
															assign node28248 = (inp[12]) ? node28250 : 16'b0000000001111111;
																assign node28250 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28254 = (inp[6]) ? 16'b0000000000011111 : node28255;
														assign node28255 = (inp[12]) ? node28257 : 16'b0000000001111111;
															assign node28257 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28261 = (inp[11]) ? node28267 : node28262;
													assign node28262 = (inp[10]) ? node28264 : 16'b0000000000111111;
														assign node28264 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28267 = (inp[14]) ? 16'b0000000000001111 : node28268;
														assign node28268 = (inp[10]) ? node28272 : node28269;
															assign node28269 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node28272 = (inp[6]) ? node28274 : 16'b0000000000011111;
																assign node28274 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node28278 = (inp[2]) ? node28418 : node28279;
									assign node28279 = (inp[8]) ? node28351 : node28280;
										assign node28280 = (inp[14]) ? node28320 : node28281;
											assign node28281 = (inp[12]) ? node28297 : node28282;
												assign node28282 = (inp[11]) ? node28290 : node28283;
													assign node28283 = (inp[7]) ? node28285 : 16'b0000001111111111;
														assign node28285 = (inp[10]) ? node28287 : 16'b0000000111111111;
															assign node28287 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28290 = (inp[7]) ? 16'b0000000001111111 : node28291;
														assign node28291 = (inp[6]) ? 16'b0000000011111111 : node28292;
															assign node28292 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node28297 = (inp[4]) ? node28313 : node28298;
													assign node28298 = (inp[10]) ? node28302 : node28299;
														assign node28299 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28302 = (inp[7]) ? node28308 : node28303;
															assign node28303 = (inp[6]) ? 16'b0000000011111111 : node28304;
																assign node28304 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node28308 = (inp[6]) ? 16'b0000000001111111 : node28309;
																assign node28309 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28313 = (inp[10]) ? node28317 : node28314;
														assign node28314 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28317 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28320 = (inp[4]) ? node28336 : node28321;
												assign node28321 = (inp[12]) ? node28327 : node28322;
													assign node28322 = (inp[7]) ? 16'b0000000011111111 : node28323;
														assign node28323 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node28327 = (inp[11]) ? 16'b0000000000111111 : node28328;
														assign node28328 = (inp[6]) ? 16'b0000000000111111 : node28329;
															assign node28329 = (inp[7]) ? node28331 : 16'b0000000011111111;
																assign node28331 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28336 = (inp[10]) ? node28344 : node28337;
													assign node28337 = (inp[12]) ? node28341 : node28338;
														assign node28338 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28341 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28344 = (inp[7]) ? node28346 : 16'b0000000000111111;
														assign node28346 = (inp[12]) ? 16'b0000000000011111 : node28347;
															assign node28347 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node28351 = (inp[12]) ? node28385 : node28352;
											assign node28352 = (inp[11]) ? node28372 : node28353;
												assign node28353 = (inp[4]) ? node28359 : node28354;
													assign node28354 = (inp[10]) ? 16'b0000000011111111 : node28355;
														assign node28355 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28359 = (inp[10]) ? node28363 : node28360;
														assign node28360 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28363 = (inp[14]) ? node28367 : node28364;
															assign node28364 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node28367 = (inp[7]) ? 16'b0000000000111111 : node28368;
																assign node28368 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28372 = (inp[4]) ? node28378 : node28373;
													assign node28373 = (inp[6]) ? node28375 : 16'b0000000001111111;
														assign node28375 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28378 = (inp[14]) ? node28382 : node28379;
														assign node28379 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28382 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28385 = (inp[14]) ? node28407 : node28386;
												assign node28386 = (inp[4]) ? node28398 : node28387;
													assign node28387 = (inp[11]) ? node28393 : node28388;
														assign node28388 = (inp[7]) ? node28390 : 16'b0000000011111111;
															assign node28390 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28393 = (inp[10]) ? node28395 : 16'b0000000001111111;
															assign node28395 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28398 = (inp[7]) ? node28404 : node28399;
														assign node28399 = (inp[10]) ? 16'b0000000000111111 : node28400;
															assign node28400 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28404 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28407 = (inp[6]) ? node28411 : node28408;
													assign node28408 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28411 = (inp[11]) ? node28415 : node28412;
														assign node28412 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28415 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000001111;
									assign node28418 = (inp[11]) ? node28496 : node28419;
										assign node28419 = (inp[6]) ? node28465 : node28420;
											assign node28420 = (inp[8]) ? node28442 : node28421;
												assign node28421 = (inp[7]) ? node28433 : node28422;
													assign node28422 = (inp[14]) ? node28428 : node28423;
														assign node28423 = (inp[10]) ? node28425 : 16'b0000000111111111;
															assign node28425 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28428 = (inp[4]) ? 16'b0000000001111111 : node28429;
															assign node28429 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28433 = (inp[4]) ? node28437 : node28434;
														assign node28434 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28437 = (inp[14]) ? 16'b0000000001111111 : node28438;
															assign node28438 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28442 = (inp[12]) ? node28458 : node28443;
													assign node28443 = (inp[7]) ? node28451 : node28444;
														assign node28444 = (inp[14]) ? 16'b0000000001111111 : node28445;
															assign node28445 = (inp[10]) ? node28447 : 16'b0000000011111111;
																assign node28447 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28451 = (inp[14]) ? 16'b0000000000011111 : node28452;
															assign node28452 = (inp[4]) ? node28454 : 16'b0000000001111111;
																assign node28454 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28458 = (inp[14]) ? 16'b0000000000111111 : node28459;
														assign node28459 = (inp[4]) ? node28461 : 16'b0000000000111111;
															assign node28461 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28465 = (inp[4]) ? node28475 : node28466;
												assign node28466 = (inp[14]) ? node28468 : 16'b0000000001111111;
													assign node28468 = (inp[12]) ? 16'b0000000000111111 : node28469;
														assign node28469 = (inp[8]) ? node28471 : 16'b0000000001111111;
															assign node28471 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28475 = (inp[14]) ? node28485 : node28476;
													assign node28476 = (inp[10]) ? node28482 : node28477;
														assign node28477 = (inp[7]) ? 16'b0000000000111111 : node28478;
															assign node28478 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28482 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28485 = (inp[12]) ? node28489 : node28486;
														assign node28486 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28489 = (inp[7]) ? node28491 : 16'b0000000000011111;
															assign node28491 = (inp[10]) ? 16'b0000000000001111 : node28492;
																assign node28492 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28496 = (inp[8]) ? node28534 : node28497;
											assign node28497 = (inp[4]) ? node28515 : node28498;
												assign node28498 = (inp[7]) ? node28510 : node28499;
													assign node28499 = (inp[12]) ? node28505 : node28500;
														assign node28500 = (inp[14]) ? 16'b0000000001111111 : node28501;
															assign node28501 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28505 = (inp[14]) ? 16'b0000000000111111 : node28506;
															assign node28506 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28510 = (inp[12]) ? 16'b0000000000011111 : node28511;
														assign node28511 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28515 = (inp[6]) ? node28525 : node28516;
													assign node28516 = (inp[12]) ? node28520 : node28517;
														assign node28517 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28520 = (inp[10]) ? node28522 : 16'b0000000000111111;
															assign node28522 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28525 = (inp[7]) ? node28527 : 16'b0000000000011111;
														assign node28527 = (inp[10]) ? node28529 : 16'b0000000000011111;
															assign node28529 = (inp[12]) ? 16'b0000000000001111 : node28530;
																assign node28530 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28534 = (inp[14]) ? node28548 : node28535;
												assign node28535 = (inp[6]) ? node28543 : node28536;
													assign node28536 = (inp[10]) ? node28540 : node28537;
														assign node28537 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28540 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28543 = (inp[10]) ? node28545 : 16'b0000000000011111;
														assign node28545 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000001111;
												assign node28548 = (inp[12]) ? node28556 : node28549;
													assign node28549 = (inp[4]) ? node28553 : node28550;
														assign node28550 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28553 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28556 = (inp[6]) ? 16'b0000000000000111 : node28557;
														assign node28557 = (inp[4]) ? node28559 : 16'b0000000000011111;
															assign node28559 = (inp[10]) ? node28561 : 16'b0000000000001111;
																assign node28561 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node28565 = (inp[10]) ? node28817 : node28566;
								assign node28566 = (inp[14]) ? node28682 : node28567;
									assign node28567 = (inp[8]) ? node28627 : node28568;
										assign node28568 = (inp[9]) ? node28604 : node28569;
											assign node28569 = (inp[7]) ? node28583 : node28570;
												assign node28570 = (inp[4]) ? node28576 : node28571;
													assign node28571 = (inp[2]) ? 16'b0000000111111111 : node28572;
														assign node28572 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node28576 = (inp[2]) ? node28578 : 16'b0000000111111111;
														assign node28578 = (inp[12]) ? node28580 : 16'b0000000011111111;
															assign node28580 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28583 = (inp[4]) ? node28599 : node28584;
													assign node28584 = (inp[12]) ? node28586 : 16'b0000000111111111;
														assign node28586 = (inp[11]) ? node28594 : node28587;
															assign node28587 = (inp[6]) ? node28591 : node28588;
																assign node28588 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
																assign node28591 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node28594 = (inp[2]) ? 16'b0000000001111111 : node28595;
																assign node28595 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28599 = (inp[12]) ? 16'b0000000001111111 : node28600;
														assign node28600 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node28604 = (inp[7]) ? node28608 : node28605;
												assign node28605 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28608 = (inp[4]) ? node28618 : node28609;
													assign node28609 = (inp[2]) ? node28613 : node28610;
														assign node28610 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node28613 = (inp[11]) ? node28615 : 16'b0000000001111111;
															assign node28615 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28618 = (inp[12]) ? node28622 : node28619;
														assign node28619 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28622 = (inp[2]) ? node28624 : 16'b0000000000111111;
															assign node28624 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28627 = (inp[4]) ? node28659 : node28628;
											assign node28628 = (inp[12]) ? node28642 : node28629;
												assign node28629 = (inp[6]) ? node28635 : node28630;
													assign node28630 = (inp[9]) ? node28632 : 16'b0000000011111111;
														assign node28632 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28635 = (inp[2]) ? node28639 : node28636;
														assign node28636 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28639 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28642 = (inp[11]) ? node28654 : node28643;
													assign node28643 = (inp[7]) ? node28651 : node28644;
														assign node28644 = (inp[2]) ? 16'b0000000001111111 : node28645;
															assign node28645 = (inp[6]) ? node28647 : 16'b0000000011111111;
																assign node28647 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28651 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28654 = (inp[9]) ? node28656 : 16'b0000000000111111;
														assign node28656 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28659 = (inp[12]) ? node28669 : node28660;
												assign node28660 = (inp[2]) ? 16'b0000000000111111 : node28661;
													assign node28661 = (inp[11]) ? node28665 : node28662;
														assign node28662 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node28665 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node28669 = (inp[9]) ? node28677 : node28670;
													assign node28670 = (inp[11]) ? 16'b0000000000001111 : node28671;
														assign node28671 = (inp[2]) ? node28673 : 16'b0000000000111111;
															assign node28673 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28677 = (inp[6]) ? 16'b0000000000011111 : node28678;
														assign node28678 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node28682 = (inp[12]) ? node28752 : node28683;
										assign node28683 = (inp[8]) ? node28717 : node28684;
											assign node28684 = (inp[11]) ? node28702 : node28685;
												assign node28685 = (inp[2]) ? node28691 : node28686;
													assign node28686 = (inp[9]) ? node28688 : 16'b0000000011111111;
														assign node28688 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28691 = (inp[6]) ? node28695 : node28692;
														assign node28692 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28695 = (inp[7]) ? node28697 : 16'b0000000001111111;
															assign node28697 = (inp[4]) ? 16'b0000000000111111 : node28698;
																assign node28698 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28702 = (inp[4]) ? node28710 : node28703;
													assign node28703 = (inp[6]) ? node28707 : node28704;
														assign node28704 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node28707 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28710 = (inp[7]) ? node28712 : 16'b0000000000111111;
														assign node28712 = (inp[6]) ? node28714 : 16'b0000000000111111;
															assign node28714 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28717 = (inp[7]) ? node28727 : node28718;
												assign node28718 = (inp[11]) ? node28720 : 16'b0000000001111111;
													assign node28720 = (inp[4]) ? 16'b0000000000111111 : node28721;
														assign node28721 = (inp[2]) ? node28723 : 16'b0000000001111111;
															assign node28723 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28727 = (inp[11]) ? node28743 : node28728;
													assign node28728 = (inp[6]) ? node28734 : node28729;
														assign node28729 = (inp[2]) ? 16'b0000000000111111 : node28730;
															assign node28730 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28734 = (inp[4]) ? node28738 : node28735;
															assign node28735 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node28738 = (inp[2]) ? 16'b0000000000011111 : node28739;
																assign node28739 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28743 = (inp[6]) ? 16'b0000000000011111 : node28744;
														assign node28744 = (inp[2]) ? 16'b0000000000011111 : node28745;
															assign node28745 = (inp[4]) ? node28747 : 16'b0000000000111111;
																assign node28747 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node28752 = (inp[4]) ? node28782 : node28753;
											assign node28753 = (inp[6]) ? node28773 : node28754;
												assign node28754 = (inp[11]) ? node28764 : node28755;
													assign node28755 = (inp[9]) ? node28761 : node28756;
														assign node28756 = (inp[7]) ? 16'b0000000001111111 : node28757;
															assign node28757 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28761 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28764 = (inp[7]) ? node28768 : node28765;
														assign node28765 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28768 = (inp[9]) ? node28770 : 16'b0000000000111111;
															assign node28770 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28773 = (inp[9]) ? node28775 : 16'b0000000000111111;
													assign node28775 = (inp[2]) ? node28779 : node28776;
														assign node28776 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node28779 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28782 = (inp[7]) ? node28798 : node28783;
												assign node28783 = (inp[11]) ? node28789 : node28784;
													assign node28784 = (inp[2]) ? 16'b0000000000111111 : node28785;
														assign node28785 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node28789 = (inp[8]) ? node28791 : 16'b0000000000111111;
														assign node28791 = (inp[6]) ? node28793 : 16'b0000000000011111;
															assign node28793 = (inp[2]) ? node28795 : 16'b0000000000001111;
																assign node28795 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node28798 = (inp[9]) ? node28804 : node28799;
													assign node28799 = (inp[6]) ? node28801 : 16'b0000000000011111;
														assign node28801 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28804 = (inp[6]) ? node28812 : node28805;
														assign node28805 = (inp[8]) ? node28807 : 16'b0000000000011111;
															assign node28807 = (inp[2]) ? node28809 : 16'b0000000000001111;
																assign node28809 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node28812 = (inp[8]) ? 16'b0000000000000111 : node28813;
															assign node28813 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node28817 = (inp[2]) ? node28963 : node28818;
									assign node28818 = (inp[8]) ? node28880 : node28819;
										assign node28819 = (inp[12]) ? node28851 : node28820;
											assign node28820 = (inp[9]) ? node28844 : node28821;
												assign node28821 = (inp[4]) ? node28831 : node28822;
													assign node28822 = (inp[14]) ? node28826 : node28823;
														assign node28823 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node28826 = (inp[6]) ? node28828 : 16'b0000000011111111;
															assign node28828 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28831 = (inp[6]) ? node28839 : node28832;
														assign node28832 = (inp[7]) ? 16'b0000000001111111 : node28833;
															assign node28833 = (inp[14]) ? node28835 : 16'b0000000011111111;
																assign node28835 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28839 = (inp[11]) ? 16'b0000000000111111 : node28840;
															assign node28840 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28844 = (inp[11]) ? node28848 : node28845;
													assign node28845 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28848 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28851 = (inp[4]) ? node28865 : node28852;
												assign node28852 = (inp[7]) ? node28860 : node28853;
													assign node28853 = (inp[6]) ? node28857 : node28854;
														assign node28854 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28857 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28860 = (inp[11]) ? 16'b0000000000111111 : node28861;
														assign node28861 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28865 = (inp[9]) ? node28875 : node28866;
													assign node28866 = (inp[7]) ? node28868 : 16'b0000000000111111;
														assign node28868 = (inp[6]) ? 16'b0000000000011111 : node28869;
															assign node28869 = (inp[14]) ? 16'b0000000000011111 : node28870;
																assign node28870 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28875 = (inp[7]) ? node28877 : 16'b0000000000011111;
														assign node28877 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28880 = (inp[7]) ? node28926 : node28881;
											assign node28881 = (inp[14]) ? node28901 : node28882;
												assign node28882 = (inp[6]) ? node28894 : node28883;
													assign node28883 = (inp[12]) ? node28887 : node28884;
														assign node28884 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28887 = (inp[4]) ? 16'b0000000000111111 : node28888;
															assign node28888 = (inp[11]) ? node28890 : 16'b0000000001111111;
																assign node28890 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28894 = (inp[12]) ? 16'b0000000000011111 : node28895;
														assign node28895 = (inp[4]) ? 16'b0000000000111111 : node28896;
															assign node28896 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28901 = (inp[12]) ? node28913 : node28902;
													assign node28902 = (inp[9]) ? node28910 : node28903;
														assign node28903 = (inp[4]) ? 16'b0000000000111111 : node28904;
															assign node28904 = (inp[11]) ? node28906 : 16'b0000000001111111;
																assign node28906 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28910 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28913 = (inp[9]) ? node28917 : node28914;
														assign node28914 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28917 = (inp[4]) ? node28921 : node28918;
															assign node28918 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node28921 = (inp[6]) ? node28923 : 16'b0000000000001111;
																assign node28923 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node28926 = (inp[14]) ? node28948 : node28927;
												assign node28927 = (inp[9]) ? node28939 : node28928;
													assign node28928 = (inp[4]) ? node28932 : node28929;
														assign node28929 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28932 = (inp[11]) ? 16'b0000000000011111 : node28933;
															assign node28933 = (inp[6]) ? node28935 : 16'b0000000000111111;
																assign node28935 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28939 = (inp[4]) ? node28945 : node28940;
														assign node28940 = (inp[12]) ? 16'b0000000000011111 : node28941;
															assign node28941 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28945 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node28948 = (inp[4]) ? node28950 : 16'b0000000000011111;
													assign node28950 = (inp[6]) ? node28954 : node28951;
														assign node28951 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node28954 = (inp[11]) ? node28958 : node28955;
															assign node28955 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node28958 = (inp[12]) ? 16'b0000000000000111 : node28959;
																assign node28959 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node28963 = (inp[7]) ? node29013 : node28964;
										assign node28964 = (inp[14]) ? node28986 : node28965;
											assign node28965 = (inp[11]) ? node28971 : node28966;
												assign node28966 = (inp[4]) ? 16'b0000000000111111 : node28967;
													assign node28967 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28971 = (inp[9]) ? node28979 : node28972;
													assign node28972 = (inp[6]) ? node28976 : node28973;
														assign node28973 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28976 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28979 = (inp[12]) ? node28981 : 16'b0000000000011111;
														assign node28981 = (inp[4]) ? node28983 : 16'b0000000000011111;
															assign node28983 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28986 = (inp[9]) ? node29004 : node28987;
												assign node28987 = (inp[8]) ? node28993 : node28988;
													assign node28988 = (inp[6]) ? node28990 : 16'b0000000001111111;
														assign node28990 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28993 = (inp[6]) ? node28997 : node28994;
														assign node28994 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28997 = (inp[12]) ? node28999 : 16'b0000000000011111;
															assign node28999 = (inp[11]) ? 16'b0000000000001111 : node29000;
																assign node29000 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29004 = (inp[6]) ? node29006 : 16'b0000000000011111;
													assign node29006 = (inp[12]) ? node29008 : 16'b0000000000001111;
														assign node29008 = (inp[4]) ? 16'b0000000000000111 : node29009;
															assign node29009 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node29013 = (inp[8]) ? node29051 : node29014;
											assign node29014 = (inp[12]) ? node29036 : node29015;
												assign node29015 = (inp[14]) ? node29025 : node29016;
													assign node29016 = (inp[9]) ? node29018 : 16'b0000000001111111;
														assign node29018 = (inp[4]) ? 16'b0000000000011111 : node29019;
															assign node29019 = (inp[6]) ? node29021 : 16'b0000000000111111;
																assign node29021 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29025 = (inp[9]) ? node29033 : node29026;
														assign node29026 = (inp[11]) ? 16'b0000000000001111 : node29027;
															assign node29027 = (inp[4]) ? node29029 : 16'b0000000000111111;
																assign node29029 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29033 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29036 = (inp[11]) ? node29046 : node29037;
													assign node29037 = (inp[9]) ? node29041 : node29038;
														assign node29038 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29041 = (inp[4]) ? 16'b0000000000001111 : node29042;
															assign node29042 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29046 = (inp[6]) ? node29048 : 16'b0000000000001111;
														assign node29048 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node29051 = (inp[14]) ? node29061 : node29052;
												assign node29052 = (inp[11]) ? node29054 : 16'b0000000000011111;
													assign node29054 = (inp[6]) ? node29056 : 16'b0000000000011111;
														assign node29056 = (inp[9]) ? node29058 : 16'b0000000000001111;
															assign node29058 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000001111;
												assign node29061 = (inp[11]) ? node29073 : node29062;
													assign node29062 = (inp[12]) ? node29066 : node29063;
														assign node29063 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node29066 = (inp[4]) ? 16'b0000000000000111 : node29067;
															assign node29067 = (inp[9]) ? node29069 : 16'b0000000000001111;
																assign node29069 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node29073 = (inp[6]) ? node29077 : node29074;
														assign node29074 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node29077 = (inp[4]) ? node29079 : 16'b0000000000000111;
															assign node29079 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000000111;
				assign node29082 = (inp[7]) ? node31218 : node29083;
					assign node29083 = (inp[6]) ? node30165 : node29084;
						assign node29084 = (inp[9]) ? node29618 : node29085;
							assign node29085 = (inp[2]) ? node29349 : node29086;
								assign node29086 = (inp[11]) ? node29224 : node29087;
									assign node29087 = (inp[12]) ? node29171 : node29088;
										assign node29088 = (inp[15]) ? node29136 : node29089;
											assign node29089 = (inp[10]) ? node29109 : node29090;
												assign node29090 = (inp[4]) ? node29100 : node29091;
													assign node29091 = (inp[8]) ? node29093 : 16'b0000011111111111;
														assign node29093 = (inp[13]) ? 16'b0000001111111111 : node29094;
															assign node29094 = (inp[1]) ? node29096 : 16'b0000011111111111;
																assign node29096 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node29100 = (inp[8]) ? 16'b0000000111111111 : node29101;
														assign node29101 = (inp[1]) ? 16'b0000001111111111 : node29102;
															assign node29102 = (inp[14]) ? node29104 : 16'b0000011111111111;
																assign node29104 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node29109 = (inp[14]) ? node29123 : node29110;
													assign node29110 = (inp[1]) ? node29118 : node29111;
														assign node29111 = (inp[4]) ? 16'b0000001111111111 : node29112;
															assign node29112 = (inp[13]) ? node29114 : 16'b0000011111111111;
																assign node29114 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node29118 = (inp[4]) ? node29120 : 16'b0000001111111111;
															assign node29120 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node29123 = (inp[8]) ? node29131 : node29124;
														assign node29124 = (inp[1]) ? 16'b0000000111111111 : node29125;
															assign node29125 = (inp[13]) ? 16'b0000001111111111 : node29126;
																assign node29126 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node29131 = (inp[4]) ? 16'b0000000011111111 : node29132;
															assign node29132 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node29136 = (inp[1]) ? node29152 : node29137;
												assign node29137 = (inp[8]) ? node29143 : node29138;
													assign node29138 = (inp[4]) ? 16'b0000001111111111 : node29139;
														assign node29139 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node29143 = (inp[13]) ? 16'b0000000111111111 : node29144;
														assign node29144 = (inp[10]) ? node29146 : 16'b0000001111111111;
															assign node29146 = (inp[14]) ? 16'b0000000111111111 : node29147;
																assign node29147 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node29152 = (inp[10]) ? node29164 : node29153;
													assign node29153 = (inp[14]) ? node29159 : node29154;
														assign node29154 = (inp[13]) ? 16'b0000000111111111 : node29155;
															assign node29155 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29159 = (inp[4]) ? node29161 : 16'b0000000111111111;
															assign node29161 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29164 = (inp[14]) ? node29168 : node29165;
														assign node29165 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29168 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node29171 = (inp[15]) ? node29195 : node29172;
											assign node29172 = (inp[10]) ? node29184 : node29173;
												assign node29173 = (inp[1]) ? node29175 : 16'b0000001111111111;
													assign node29175 = (inp[4]) ? node29179 : node29176;
														assign node29176 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29179 = (inp[13]) ? node29181 : 16'b0000000111111111;
															assign node29181 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29184 = (inp[1]) ? node29190 : node29185;
													assign node29185 = (inp[14]) ? node29187 : 16'b0000000111111111;
														assign node29187 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29190 = (inp[13]) ? 16'b0000000011111111 : node29191;
														assign node29191 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node29195 = (inp[1]) ? node29207 : node29196;
												assign node29196 = (inp[10]) ? node29202 : node29197;
													assign node29197 = (inp[13]) ? node29199 : 16'b0000000111111111;
														assign node29199 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29202 = (inp[13]) ? node29204 : 16'b0000000011111111;
														assign node29204 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29207 = (inp[8]) ? node29217 : node29208;
													assign node29208 = (inp[4]) ? node29212 : node29209;
														assign node29209 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node29212 = (inp[13]) ? node29214 : 16'b0000000011111111;
															assign node29214 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29217 = (inp[13]) ? 16'b0000000001111111 : node29218;
														assign node29218 = (inp[10]) ? 16'b0000000001111111 : node29219;
															assign node29219 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node29224 = (inp[15]) ? node29286 : node29225;
										assign node29225 = (inp[10]) ? node29249 : node29226;
											assign node29226 = (inp[14]) ? node29238 : node29227;
												assign node29227 = (inp[8]) ? node29233 : node29228;
													assign node29228 = (inp[13]) ? 16'b0000001111111111 : node29229;
														assign node29229 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node29233 = (inp[13]) ? node29235 : 16'b0000001111111111;
														assign node29235 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29238 = (inp[1]) ? node29246 : node29239;
													assign node29239 = (inp[13]) ? node29241 : 16'b0000001111111111;
														assign node29241 = (inp[8]) ? node29243 : 16'b0000000111111111;
															assign node29243 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29246 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node29249 = (inp[1]) ? node29275 : node29250;
												assign node29250 = (inp[12]) ? node29264 : node29251;
													assign node29251 = (inp[4]) ? node29257 : node29252;
														assign node29252 = (inp[8]) ? node29254 : 16'b0000011111111111;
															assign node29254 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29257 = (inp[8]) ? node29259 : 16'b0000000111111111;
															assign node29259 = (inp[13]) ? 16'b0000000011111111 : node29260;
																assign node29260 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29264 = (inp[14]) ? node29268 : node29265;
														assign node29265 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29268 = (inp[8]) ? node29270 : 16'b0000000011111111;
															assign node29270 = (inp[13]) ? 16'b0000000001111111 : node29271;
																assign node29271 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29275 = (inp[13]) ? node29279 : node29276;
													assign node29276 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29279 = (inp[4]) ? node29281 : 16'b0000000001111111;
														assign node29281 = (inp[14]) ? 16'b0000000000011111 : node29282;
															assign node29282 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node29286 = (inp[4]) ? node29316 : node29287;
											assign node29287 = (inp[13]) ? node29303 : node29288;
												assign node29288 = (inp[12]) ? node29298 : node29289;
													assign node29289 = (inp[8]) ? node29295 : node29290;
														assign node29290 = (inp[1]) ? 16'b0000000111111111 : node29291;
															assign node29291 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29295 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29298 = (inp[8]) ? 16'b0000000011111111 : node29299;
														assign node29299 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29303 = (inp[12]) ? node29313 : node29304;
													assign node29304 = (inp[14]) ? node29310 : node29305;
														assign node29305 = (inp[1]) ? 16'b0000000011111111 : node29306;
															assign node29306 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29310 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29313 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node29316 = (inp[14]) ? node29328 : node29317;
												assign node29317 = (inp[10]) ? node29323 : node29318;
													assign node29318 = (inp[8]) ? node29320 : 16'b0000000111111111;
														assign node29320 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node29323 = (inp[13]) ? 16'b0000000001111111 : node29324;
														assign node29324 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29328 = (inp[12]) ? node29338 : node29329;
													assign node29329 = (inp[10]) ? node29333 : node29330;
														assign node29330 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29333 = (inp[1]) ? 16'b0000000000111111 : node29334;
															assign node29334 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29338 = (inp[10]) ? node29340 : 16'b0000000000111111;
														assign node29340 = (inp[1]) ? node29346 : node29341;
															assign node29341 = (inp[13]) ? node29343 : 16'b0000000000111111;
																assign node29343 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node29346 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node29349 = (inp[1]) ? node29475 : node29350;
									assign node29350 = (inp[14]) ? node29414 : node29351;
										assign node29351 = (inp[15]) ? node29385 : node29352;
											assign node29352 = (inp[13]) ? node29364 : node29353;
												assign node29353 = (inp[11]) ? 16'b0000000111111111 : node29354;
													assign node29354 = (inp[4]) ? node29356 : 16'b0000011111111111;
														assign node29356 = (inp[10]) ? 16'b0000001111111111 : node29357;
															assign node29357 = (inp[12]) ? 16'b0000001111111111 : node29358;
																assign node29358 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node29364 = (inp[4]) ? node29380 : node29365;
													assign node29365 = (inp[8]) ? node29373 : node29366;
														assign node29366 = (inp[10]) ? node29368 : 16'b0000001111111111;
															assign node29368 = (inp[11]) ? 16'b0000000111111111 : node29369;
																assign node29369 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29373 = (inp[12]) ? node29375 : 16'b0000000111111111;
															assign node29375 = (inp[10]) ? 16'b0000000011111111 : node29376;
																assign node29376 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29380 = (inp[12]) ? node29382 : 16'b0000000011111111;
														assign node29382 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node29385 = (inp[10]) ? node29399 : node29386;
												assign node29386 = (inp[11]) ? node29394 : node29387;
													assign node29387 = (inp[13]) ? node29391 : node29388;
														assign node29388 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node29391 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29394 = (inp[4]) ? 16'b0000000001111111 : node29395;
														assign node29395 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29399 = (inp[12]) ? node29401 : 16'b0000000011111111;
													assign node29401 = (inp[8]) ? node29409 : node29402;
														assign node29402 = (inp[4]) ? node29404 : 16'b0000000011111111;
															assign node29404 = (inp[13]) ? 16'b0000000001111111 : node29405;
																assign node29405 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29409 = (inp[13]) ? node29411 : 16'b0000000001111111;
															assign node29411 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node29414 = (inp[13]) ? node29446 : node29415;
											assign node29415 = (inp[10]) ? node29433 : node29416;
												assign node29416 = (inp[11]) ? node29424 : node29417;
													assign node29417 = (inp[12]) ? node29419 : 16'b0000000111111111;
														assign node29419 = (inp[15]) ? node29421 : 16'b0000000111111111;
															assign node29421 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29424 = (inp[4]) ? node29430 : node29425;
														assign node29425 = (inp[15]) ? 16'b0000000011111111 : node29426;
															assign node29426 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29430 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29433 = (inp[15]) ? node29441 : node29434;
													assign node29434 = (inp[8]) ? node29436 : 16'b0000000111111111;
														assign node29436 = (inp[12]) ? 16'b0000000001111111 : node29437;
															assign node29437 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29441 = (inp[4]) ? node29443 : 16'b0000000001111111;
														assign node29443 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node29446 = (inp[11]) ? node29464 : node29447;
												assign node29447 = (inp[15]) ? node29457 : node29448;
													assign node29448 = (inp[8]) ? node29450 : 16'b0000000011111111;
														assign node29450 = (inp[4]) ? 16'b0000000001111111 : node29451;
															assign node29451 = (inp[10]) ? node29453 : 16'b0000000011111111;
																assign node29453 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29457 = (inp[4]) ? 16'b0000000000111111 : node29458;
														assign node29458 = (inp[8]) ? 16'b0000000001111111 : node29459;
															assign node29459 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29464 = (inp[12]) ? node29466 : 16'b0000000001111111;
													assign node29466 = (inp[10]) ? 16'b0000000000011111 : node29467;
														assign node29467 = (inp[4]) ? node29469 : 16'b0000000001111111;
															assign node29469 = (inp[8]) ? 16'b0000000000111111 : node29470;
																assign node29470 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node29475 = (inp[4]) ? node29545 : node29476;
										assign node29476 = (inp[12]) ? node29512 : node29477;
											assign node29477 = (inp[11]) ? node29495 : node29478;
												assign node29478 = (inp[10]) ? node29486 : node29479;
													assign node29479 = (inp[14]) ? node29483 : node29480;
														assign node29480 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29483 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29486 = (inp[13]) ? node29488 : 16'b0000000001111111;
														assign node29488 = (inp[15]) ? 16'b0000000011111111 : node29489;
															assign node29489 = (inp[14]) ? 16'b0000000011111111 : node29490;
																assign node29490 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29495 = (inp[14]) ? node29497 : 16'b0000000011111111;
													assign node29497 = (inp[15]) ? node29507 : node29498;
														assign node29498 = (inp[8]) ? node29504 : node29499;
															assign node29499 = (inp[13]) ? 16'b0000000011111111 : node29500;
																assign node29500 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node29504 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29507 = (inp[10]) ? 16'b0000000000111111 : node29508;
															assign node29508 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node29512 = (inp[13]) ? node29528 : node29513;
												assign node29513 = (inp[15]) ? node29521 : node29514;
													assign node29514 = (inp[10]) ? node29518 : node29515;
														assign node29515 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node29518 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29521 = (inp[10]) ? node29525 : node29522;
														assign node29522 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29525 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node29528 = (inp[8]) ? node29538 : node29529;
													assign node29529 = (inp[11]) ? node29535 : node29530;
														assign node29530 = (inp[15]) ? 16'b0000000001111111 : node29531;
															assign node29531 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29535 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29538 = (inp[14]) ? node29542 : node29539;
														assign node29539 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29542 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node29545 = (inp[14]) ? node29577 : node29546;
											assign node29546 = (inp[10]) ? node29558 : node29547;
												assign node29547 = (inp[11]) ? node29551 : node29548;
													assign node29548 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node29551 = (inp[12]) ? 16'b0000000001111111 : node29552;
														assign node29552 = (inp[8]) ? 16'b0000000001111111 : node29553;
															assign node29553 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29558 = (inp[12]) ? node29566 : node29559;
													assign node29559 = (inp[13]) ? node29563 : node29560;
														assign node29560 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29563 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node29566 = (inp[8]) ? node29574 : node29567;
														assign node29567 = (inp[15]) ? node29569 : 16'b0000000001111111;
															assign node29569 = (inp[13]) ? 16'b0000000000111111 : node29570;
																assign node29570 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29574 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29577 = (inp[12]) ? node29599 : node29578;
												assign node29578 = (inp[10]) ? node29590 : node29579;
													assign node29579 = (inp[15]) ? node29583 : node29580;
														assign node29580 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node29583 = (inp[8]) ? node29585 : 16'b0000000001111111;
															assign node29585 = (inp[13]) ? 16'b0000000000111111 : node29586;
																assign node29586 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29590 = (inp[8]) ? node29594 : node29591;
														assign node29591 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29594 = (inp[11]) ? 16'b0000000000011111 : node29595;
															assign node29595 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29599 = (inp[13]) ? node29609 : node29600;
													assign node29600 = (inp[11]) ? node29602 : 16'b0000000001111111;
														assign node29602 = (inp[10]) ? node29604 : 16'b0000000000111111;
															assign node29604 = (inp[15]) ? 16'b0000000000011111 : node29605;
																assign node29605 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29609 = (inp[15]) ? node29615 : node29610;
														assign node29610 = (inp[10]) ? 16'b0000000000011111 : node29611;
															assign node29611 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29615 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node29618 = (inp[4]) ? node29908 : node29619;
								assign node29619 = (inp[14]) ? node29761 : node29620;
									assign node29620 = (inp[15]) ? node29702 : node29621;
										assign node29621 = (inp[12]) ? node29661 : node29622;
											assign node29622 = (inp[8]) ? node29646 : node29623;
												assign node29623 = (inp[10]) ? node29635 : node29624;
													assign node29624 = (inp[1]) ? node29628 : node29625;
														assign node29625 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node29628 = (inp[11]) ? node29630 : 16'b0000001111111111;
															assign node29630 = (inp[2]) ? 16'b0000000111111111 : node29631;
																assign node29631 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node29635 = (inp[2]) ? node29639 : node29636;
														assign node29636 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29639 = (inp[13]) ? node29641 : 16'b0000000111111111;
															assign node29641 = (inp[1]) ? 16'b0000000011111111 : node29642;
																assign node29642 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29646 = (inp[11]) ? node29654 : node29647;
													assign node29647 = (inp[1]) ? 16'b0000000111111111 : node29648;
														assign node29648 = (inp[2]) ? 16'b0000000111111111 : node29649;
															assign node29649 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node29654 = (inp[13]) ? node29658 : node29655;
														assign node29655 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29658 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node29661 = (inp[2]) ? node29685 : node29662;
												assign node29662 = (inp[10]) ? node29676 : node29663;
													assign node29663 = (inp[1]) ? node29671 : node29664;
														assign node29664 = (inp[11]) ? node29666 : 16'b0000011111111111;
															assign node29666 = (inp[13]) ? 16'b0000000111111111 : node29667;
																assign node29667 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29671 = (inp[13]) ? node29673 : 16'b0000000111111111;
															assign node29673 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29676 = (inp[11]) ? node29680 : node29677;
														assign node29677 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29680 = (inp[13]) ? node29682 : 16'b0000000011111111;
															assign node29682 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29685 = (inp[11]) ? node29689 : node29686;
													assign node29686 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node29689 = (inp[10]) ? node29699 : node29690;
														assign node29690 = (inp[13]) ? node29696 : node29691;
															assign node29691 = (inp[8]) ? node29693 : 16'b0000000011111111;
																assign node29693 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node29696 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29699 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node29702 = (inp[13]) ? node29732 : node29703;
											assign node29703 = (inp[10]) ? node29717 : node29704;
												assign node29704 = (inp[1]) ? node29710 : node29705;
													assign node29705 = (inp[11]) ? 16'b0000000111111111 : node29706;
														assign node29706 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node29710 = (inp[8]) ? node29712 : 16'b0000001111111111;
														assign node29712 = (inp[2]) ? 16'b0000000001111111 : node29713;
															assign node29713 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29717 = (inp[11]) ? node29727 : node29718;
													assign node29718 = (inp[2]) ? node29722 : node29719;
														assign node29719 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29722 = (inp[1]) ? node29724 : 16'b0000000011111111;
															assign node29724 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29727 = (inp[1]) ? 16'b0000000000111111 : node29728;
														assign node29728 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node29732 = (inp[10]) ? node29746 : node29733;
												assign node29733 = (inp[12]) ? node29739 : node29734;
													assign node29734 = (inp[11]) ? node29736 : 16'b0000000011111111;
														assign node29736 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29739 = (inp[11]) ? 16'b0000000000111111 : node29740;
														assign node29740 = (inp[8]) ? 16'b0000000001111111 : node29741;
															assign node29741 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29746 = (inp[1]) ? node29754 : node29747;
													assign node29747 = (inp[8]) ? node29751 : node29748;
														assign node29748 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29751 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29754 = (inp[12]) ? node29758 : node29755;
														assign node29755 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29758 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node29761 = (inp[12]) ? node29831 : node29762;
										assign node29762 = (inp[10]) ? node29800 : node29763;
											assign node29763 = (inp[13]) ? node29773 : node29764;
												assign node29764 = (inp[2]) ? 16'b0000000011111111 : node29765;
													assign node29765 = (inp[11]) ? node29767 : 16'b0000001111111111;
														assign node29767 = (inp[1]) ? 16'b0000000111111111 : node29768;
															assign node29768 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node29773 = (inp[15]) ? node29789 : node29774;
													assign node29774 = (inp[2]) ? node29786 : node29775;
														assign node29775 = (inp[1]) ? node29781 : node29776;
															assign node29776 = (inp[11]) ? node29778 : 16'b0000000111111111;
																assign node29778 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node29781 = (inp[11]) ? 16'b0000000011111111 : node29782;
																assign node29782 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29786 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29789 = (inp[11]) ? node29795 : node29790;
														assign node29790 = (inp[1]) ? node29792 : 16'b0000000011111111;
															assign node29792 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29795 = (inp[1]) ? 16'b0000000000111111 : node29796;
															assign node29796 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node29800 = (inp[2]) ? node29820 : node29801;
												assign node29801 = (inp[13]) ? node29813 : node29802;
													assign node29802 = (inp[8]) ? node29806 : node29803;
														assign node29803 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29806 = (inp[1]) ? 16'b0000000001111111 : node29807;
															assign node29807 = (inp[15]) ? node29809 : 16'b0000000011111111;
																assign node29809 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29813 = (inp[15]) ? 16'b0000000000011111 : node29814;
														assign node29814 = (inp[11]) ? node29816 : 16'b0000000001111111;
															assign node29816 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29820 = (inp[8]) ? node29828 : node29821;
													assign node29821 = (inp[15]) ? 16'b0000000000111111 : node29822;
														assign node29822 = (inp[11]) ? 16'b0000000001111111 : node29823;
															assign node29823 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29828 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node29831 = (inp[1]) ? node29875 : node29832;
											assign node29832 = (inp[2]) ? node29860 : node29833;
												assign node29833 = (inp[13]) ? node29845 : node29834;
													assign node29834 = (inp[11]) ? node29838 : node29835;
														assign node29835 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node29838 = (inp[8]) ? 16'b0000000001111111 : node29839;
															assign node29839 = (inp[10]) ? node29841 : 16'b0000000011111111;
																assign node29841 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29845 = (inp[11]) ? node29855 : node29846;
														assign node29846 = (inp[10]) ? node29852 : node29847;
															assign node29847 = (inp[15]) ? node29849 : 16'b0000000011111111;
																assign node29849 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
															assign node29852 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29855 = (inp[8]) ? node29857 : 16'b0000000001111111;
															assign node29857 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29860 = (inp[13]) ? node29870 : node29861;
													assign node29861 = (inp[15]) ? node29865 : node29862;
														assign node29862 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29865 = (inp[8]) ? 16'b0000000000111111 : node29866;
															assign node29866 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29870 = (inp[15]) ? node29872 : 16'b0000000000111111;
														assign node29872 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29875 = (inp[13]) ? node29887 : node29876;
												assign node29876 = (inp[2]) ? node29880 : node29877;
													assign node29877 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29880 = (inp[8]) ? node29882 : 16'b0000000001111111;
														assign node29882 = (inp[10]) ? node29884 : 16'b0000000000111111;
															assign node29884 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node29887 = (inp[10]) ? node29893 : node29888;
													assign node29888 = (inp[11]) ? node29890 : 16'b0000000000111111;
														assign node29890 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29893 = (inp[11]) ? node29897 : node29894;
														assign node29894 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29897 = (inp[2]) ? node29903 : node29898;
															assign node29898 = (inp[8]) ? node29900 : 16'b0000000000011111;
																assign node29900 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node29903 = (inp[8]) ? node29905 : 16'b0000000000001111;
																assign node29905 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node29908 = (inp[1]) ? node30034 : node29909;
									assign node29909 = (inp[12]) ? node29963 : node29910;
										assign node29910 = (inp[2]) ? node29942 : node29911;
											assign node29911 = (inp[13]) ? node29925 : node29912;
												assign node29912 = (inp[10]) ? node29920 : node29913;
													assign node29913 = (inp[8]) ? 16'b0000000111111111 : node29914;
														assign node29914 = (inp[15]) ? node29916 : 16'b0000000111111111;
															assign node29916 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29920 = (inp[11]) ? node29922 : 16'b0000000011111111;
														assign node29922 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29925 = (inp[15]) ? node29937 : node29926;
													assign node29926 = (inp[14]) ? node29930 : node29927;
														assign node29927 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29930 = (inp[10]) ? node29932 : 16'b0000000011111111;
															assign node29932 = (inp[8]) ? 16'b0000000001111111 : node29933;
																assign node29933 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29937 = (inp[14]) ? node29939 : 16'b0000000001111111;
														assign node29939 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node29942 = (inp[10]) ? node29952 : node29943;
												assign node29943 = (inp[13]) ? 16'b0000000001111111 : node29944;
													assign node29944 = (inp[14]) ? node29946 : 16'b0000001111111111;
														assign node29946 = (inp[15]) ? node29948 : 16'b0000000011111111;
															assign node29948 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29952 = (inp[14]) ? node29958 : node29953;
													assign node29953 = (inp[11]) ? node29955 : 16'b0000000001111111;
														assign node29955 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29958 = (inp[15]) ? node29960 : 16'b0000000001111111;
														assign node29960 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node29963 = (inp[11]) ? node30007 : node29964;
											assign node29964 = (inp[10]) ? node29984 : node29965;
												assign node29965 = (inp[13]) ? node29971 : node29966;
													assign node29966 = (inp[2]) ? 16'b0000000011111111 : node29967;
														assign node29967 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29971 = (inp[14]) ? node29979 : node29972;
														assign node29972 = (inp[2]) ? 16'b0000000001111111 : node29973;
															assign node29973 = (inp[15]) ? node29975 : 16'b0000000011111111;
																assign node29975 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29979 = (inp[2]) ? node29981 : 16'b0000000001111111;
															assign node29981 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29984 = (inp[2]) ? node30002 : node29985;
													assign node29985 = (inp[15]) ? node29991 : node29986;
														assign node29986 = (inp[8]) ? node29988 : 16'b0000000111111111;
															assign node29988 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29991 = (inp[14]) ? node29997 : node29992;
															assign node29992 = (inp[13]) ? node29994 : 16'b0000000001111111;
																assign node29994 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node29997 = (inp[13]) ? 16'b0000000000111111 : node29998;
																assign node29998 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30002 = (inp[13]) ? 16'b0000000000011111 : node30003;
														assign node30003 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30007 = (inp[14]) ? node30019 : node30008;
												assign node30008 = (inp[10]) ? node30012 : node30009;
													assign node30009 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30012 = (inp[2]) ? node30016 : node30013;
														assign node30013 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30016 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30019 = (inp[2]) ? node30029 : node30020;
													assign node30020 = (inp[13]) ? node30026 : node30021;
														assign node30021 = (inp[15]) ? 16'b0000000000111111 : node30022;
															assign node30022 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30026 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30029 = (inp[10]) ? 16'b0000000000001111 : node30030;
														assign node30030 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node30034 = (inp[8]) ? node30086 : node30035;
										assign node30035 = (inp[11]) ? node30059 : node30036;
											assign node30036 = (inp[13]) ? node30046 : node30037;
												assign node30037 = (inp[14]) ? node30041 : node30038;
													assign node30038 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30041 = (inp[10]) ? node30043 : 16'b0000000011111111;
														assign node30043 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30046 = (inp[12]) ? node30050 : node30047;
													assign node30047 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30050 = (inp[2]) ? 16'b0000000000011111 : node30051;
														assign node30051 = (inp[14]) ? node30053 : 16'b0000000001111111;
															assign node30053 = (inp[15]) ? 16'b0000000000111111 : node30054;
																assign node30054 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30059 = (inp[10]) ? node30077 : node30060;
												assign node30060 = (inp[14]) ? node30072 : node30061;
													assign node30061 = (inp[15]) ? node30067 : node30062;
														assign node30062 = (inp[12]) ? 16'b0000000001111111 : node30063;
															assign node30063 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30067 = (inp[2]) ? node30069 : 16'b0000000001111111;
															assign node30069 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30072 = (inp[2]) ? 16'b0000000000111111 : node30073;
														assign node30073 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30077 = (inp[14]) ? node30081 : node30078;
													assign node30078 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30081 = (inp[12]) ? node30083 : 16'b0000000000011111;
														assign node30083 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node30086 = (inp[13]) ? node30124 : node30087;
											assign node30087 = (inp[2]) ? node30107 : node30088;
												assign node30088 = (inp[12]) ? node30100 : node30089;
													assign node30089 = (inp[14]) ? node30093 : node30090;
														assign node30090 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30093 = (inp[11]) ? node30095 : 16'b0000000001111111;
															assign node30095 = (inp[15]) ? node30097 : 16'b0000000001111111;
																assign node30097 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30100 = (inp[15]) ? node30104 : node30101;
														assign node30101 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30104 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30107 = (inp[12]) ? node30117 : node30108;
													assign node30108 = (inp[14]) ? node30114 : node30109;
														assign node30109 = (inp[15]) ? node30111 : 16'b0000000001111111;
															assign node30111 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30114 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30117 = (inp[14]) ? 16'b0000000000001111 : node30118;
														assign node30118 = (inp[11]) ? 16'b0000000000011111 : node30119;
															assign node30119 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30124 = (inp[14]) ? node30140 : node30125;
												assign node30125 = (inp[15]) ? node30135 : node30126;
													assign node30126 = (inp[11]) ? node30128 : 16'b0000000000111111;
														assign node30128 = (inp[10]) ? node30130 : 16'b0000000000111111;
															assign node30130 = (inp[12]) ? 16'b0000000000011111 : node30131;
																assign node30131 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30135 = (inp[12]) ? 16'b0000000000011111 : node30136;
														assign node30136 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30140 = (inp[2]) ? node30154 : node30141;
													assign node30141 = (inp[15]) ? node30149 : node30142;
														assign node30142 = (inp[12]) ? node30144 : 16'b0000000000111111;
															assign node30144 = (inp[10]) ? 16'b0000000000011111 : node30145;
																assign node30145 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30149 = (inp[12]) ? node30151 : 16'b0000000000011111;
															assign node30151 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node30154 = (inp[11]) ? node30158 : node30155;
														assign node30155 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30158 = (inp[10]) ? 16'b0000000000000111 : node30159;
															assign node30159 = (inp[15]) ? node30161 : 16'b0000000000001111;
																assign node30161 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node30165 = (inp[8]) ? node30673 : node30166;
							assign node30166 = (inp[14]) ? node30412 : node30167;
								assign node30167 = (inp[9]) ? node30301 : node30168;
									assign node30168 = (inp[1]) ? node30238 : node30169;
										assign node30169 = (inp[11]) ? node30193 : node30170;
											assign node30170 = (inp[13]) ? node30184 : node30171;
												assign node30171 = (inp[10]) ? 16'b0000000111111111 : node30172;
													assign node30172 = (inp[12]) ? node30180 : node30173;
														assign node30173 = (inp[4]) ? node30175 : 16'b0000011111111111;
															assign node30175 = (inp[2]) ? 16'b0000001111111111 : node30176;
																assign node30176 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node30180 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node30184 = (inp[4]) ? node30186 : 16'b0000000111111111;
													assign node30186 = (inp[15]) ? 16'b0000000001111111 : node30187;
														assign node30187 = (inp[10]) ? 16'b0000000011111111 : node30188;
															assign node30188 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node30193 = (inp[15]) ? node30215 : node30194;
												assign node30194 = (inp[10]) ? node30204 : node30195;
													assign node30195 = (inp[12]) ? node30199 : node30196;
														assign node30196 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node30199 = (inp[4]) ? node30201 : 16'b0000000111111111;
															assign node30201 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30204 = (inp[13]) ? 16'b0000000001111111 : node30205;
														assign node30205 = (inp[12]) ? node30211 : node30206;
															assign node30206 = (inp[4]) ? node30208 : 16'b0000000111111111;
																assign node30208 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node30211 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30215 = (inp[4]) ? node30227 : node30216;
													assign node30216 = (inp[13]) ? node30220 : node30217;
														assign node30217 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30220 = (inp[10]) ? node30222 : 16'b0000000011111111;
															assign node30222 = (inp[12]) ? 16'b0000000001111111 : node30223;
																assign node30223 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30227 = (inp[12]) ? node30231 : node30228;
														assign node30228 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30231 = (inp[10]) ? node30233 : 16'b0000000001111111;
															assign node30233 = (inp[13]) ? 16'b0000000000111111 : node30234;
																assign node30234 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node30238 = (inp[10]) ? node30268 : node30239;
											assign node30239 = (inp[11]) ? node30247 : node30240;
												assign node30240 = (inp[4]) ? 16'b0000000011111111 : node30241;
													assign node30241 = (inp[12]) ? 16'b0000000011111111 : node30242;
														assign node30242 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node30247 = (inp[4]) ? node30261 : node30248;
													assign node30248 = (inp[2]) ? node30254 : node30249;
														assign node30249 = (inp[13]) ? 16'b0000000011111111 : node30250;
															assign node30250 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30254 = (inp[15]) ? 16'b0000000001111111 : node30255;
															assign node30255 = (inp[13]) ? node30257 : 16'b0000000011111111;
																assign node30257 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30261 = (inp[12]) ? 16'b0000000000111111 : node30262;
														assign node30262 = (inp[2]) ? 16'b0000000001111111 : node30263;
															assign node30263 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node30268 = (inp[2]) ? node30284 : node30269;
												assign node30269 = (inp[12]) ? node30279 : node30270;
													assign node30270 = (inp[4]) ? node30276 : node30271;
														assign node30271 = (inp[15]) ? node30273 : 16'b0000000111111111;
															assign node30273 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30276 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30279 = (inp[15]) ? node30281 : 16'b0000000011111111;
														assign node30281 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30284 = (inp[15]) ? node30290 : node30285;
													assign node30285 = (inp[13]) ? 16'b0000000001111111 : node30286;
														assign node30286 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30290 = (inp[13]) ? node30294 : node30291;
														assign node30291 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30294 = (inp[11]) ? node30296 : 16'b0000000001111111;
															assign node30296 = (inp[12]) ? 16'b0000000000011111 : node30297;
																assign node30297 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node30301 = (inp[11]) ? node30359 : node30302;
										assign node30302 = (inp[15]) ? node30334 : node30303;
											assign node30303 = (inp[4]) ? node30321 : node30304;
												assign node30304 = (inp[12]) ? node30314 : node30305;
													assign node30305 = (inp[13]) ? node30311 : node30306;
														assign node30306 = (inp[2]) ? node30308 : 16'b0000001111111111;
															assign node30308 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node30311 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node30314 = (inp[1]) ? 16'b0000000011111111 : node30315;
														assign node30315 = (inp[2]) ? node30317 : 16'b0000000111111111;
															assign node30317 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node30321 = (inp[10]) ? node30327 : node30322;
													assign node30322 = (inp[13]) ? 16'b0000000011111111 : node30323;
														assign node30323 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node30327 = (inp[13]) ? node30331 : node30328;
														assign node30328 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30331 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30334 = (inp[2]) ? node30348 : node30335;
												assign node30335 = (inp[13]) ? node30341 : node30336;
													assign node30336 = (inp[1]) ? node30338 : 16'b0000000011111111;
														assign node30338 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30341 = (inp[10]) ? 16'b0000000001111111 : node30342;
														assign node30342 = (inp[4]) ? 16'b0000000001111111 : node30343;
															assign node30343 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30348 = (inp[13]) ? node30354 : node30349;
													assign node30349 = (inp[1]) ? 16'b0000000001111111 : node30350;
														assign node30350 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30354 = (inp[10]) ? node30356 : 16'b0000000000111111;
														assign node30356 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node30359 = (inp[15]) ? node30385 : node30360;
											assign node30360 = (inp[13]) ? node30378 : node30361;
												assign node30361 = (inp[1]) ? node30367 : node30362;
													assign node30362 = (inp[12]) ? 16'b0000000011111111 : node30363;
														assign node30363 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node30367 = (inp[12]) ? node30371 : node30368;
														assign node30368 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30371 = (inp[4]) ? 16'b0000000000111111 : node30372;
															assign node30372 = (inp[2]) ? node30374 : 16'b0000000001111111;
																assign node30374 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30378 = (inp[10]) ? 16'b0000000000111111 : node30379;
													assign node30379 = (inp[12]) ? node30381 : 16'b0000000001111111;
														assign node30381 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30385 = (inp[4]) ? node30395 : node30386;
												assign node30386 = (inp[12]) ? node30388 : 16'b0000000011111111;
													assign node30388 = (inp[2]) ? node30392 : node30389;
														assign node30389 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30392 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30395 = (inp[10]) ? node30407 : node30396;
													assign node30396 = (inp[2]) ? node30400 : node30397;
														assign node30397 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30400 = (inp[13]) ? node30402 : 16'b0000000000111111;
															assign node30402 = (inp[12]) ? node30404 : 16'b0000000000011111;
																assign node30404 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30407 = (inp[2]) ? node30409 : 16'b0000000000011111;
														assign node30409 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node30412 = (inp[2]) ? node30574 : node30413;
									assign node30413 = (inp[4]) ? node30485 : node30414;
										assign node30414 = (inp[12]) ? node30452 : node30415;
											assign node30415 = (inp[11]) ? node30443 : node30416;
												assign node30416 = (inp[15]) ? node30426 : node30417;
													assign node30417 = (inp[10]) ? node30423 : node30418;
														assign node30418 = (inp[9]) ? 16'b0000001111111111 : node30419;
															assign node30419 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node30423 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30426 = (inp[9]) ? node30432 : node30427;
														assign node30427 = (inp[10]) ? node30429 : 16'b0000000111111111;
															assign node30429 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30432 = (inp[13]) ? node30438 : node30433;
															assign node30433 = (inp[1]) ? 16'b0000000011111111 : node30434;
																assign node30434 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node30438 = (inp[10]) ? 16'b0000000001111111 : node30439;
																assign node30439 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30443 = (inp[9]) ? node30445 : 16'b0000000011111111;
													assign node30445 = (inp[1]) ? node30449 : node30446;
														assign node30446 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30449 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30452 = (inp[10]) ? node30470 : node30453;
												assign node30453 = (inp[1]) ? node30463 : node30454;
													assign node30454 = (inp[13]) ? node30456 : 16'b0000000111111111;
														assign node30456 = (inp[11]) ? node30458 : 16'b0000000011111111;
															assign node30458 = (inp[15]) ? 16'b0000000001111111 : node30459;
																assign node30459 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30463 = (inp[9]) ? node30467 : node30464;
														assign node30464 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30467 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30470 = (inp[15]) ? node30476 : node30471;
													assign node30471 = (inp[11]) ? node30473 : 16'b0000000001111111;
														assign node30473 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node30476 = (inp[11]) ? node30482 : node30477;
														assign node30477 = (inp[13]) ? 16'b0000000000111111 : node30478;
															assign node30478 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30482 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node30485 = (inp[9]) ? node30521 : node30486;
											assign node30486 = (inp[12]) ? node30504 : node30487;
												assign node30487 = (inp[1]) ? node30499 : node30488;
													assign node30488 = (inp[11]) ? node30492 : node30489;
														assign node30489 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30492 = (inp[13]) ? node30494 : 16'b0000000011111111;
															assign node30494 = (inp[10]) ? 16'b0000000001111111 : node30495;
																assign node30495 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30499 = (inp[15]) ? node30501 : 16'b0000000011111111;
														assign node30501 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30504 = (inp[13]) ? node30514 : node30505;
													assign node30505 = (inp[10]) ? 16'b0000000000111111 : node30506;
														assign node30506 = (inp[15]) ? 16'b0000000001111111 : node30507;
															assign node30507 = (inp[1]) ? node30509 : 16'b0000000011111111;
																assign node30509 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30514 = (inp[1]) ? node30518 : node30515;
														assign node30515 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30518 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30521 = (inp[10]) ? node30547 : node30522;
												assign node30522 = (inp[11]) ? node30534 : node30523;
													assign node30523 = (inp[12]) ? node30525 : 16'b0000000001111111;
														assign node30525 = (inp[13]) ? 16'b0000000000111111 : node30526;
															assign node30526 = (inp[1]) ? node30530 : node30527;
																assign node30527 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
																assign node30530 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30534 = (inp[13]) ? node30542 : node30535;
														assign node30535 = (inp[15]) ? node30537 : 16'b0000000001111111;
															assign node30537 = (inp[1]) ? 16'b0000000000111111 : node30538;
																assign node30538 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30542 = (inp[12]) ? node30544 : 16'b0000000000111111;
															assign node30544 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30547 = (inp[11]) ? node30561 : node30548;
													assign node30548 = (inp[12]) ? node30554 : node30549;
														assign node30549 = (inp[13]) ? node30551 : 16'b0000000001111111;
															assign node30551 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node30554 = (inp[1]) ? node30556 : 16'b0000000000111111;
															assign node30556 = (inp[15]) ? node30558 : 16'b0000000000111111;
																assign node30558 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30561 = (inp[1]) ? 16'b0000000000011111 : node30562;
														assign node30562 = (inp[12]) ? node30568 : node30563;
															assign node30563 = (inp[13]) ? node30565 : 16'b0000000000111111;
																assign node30565 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node30568 = (inp[13]) ? 16'b0000000000011111 : node30569;
																assign node30569 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node30574 = (inp[1]) ? node30630 : node30575;
										assign node30575 = (inp[4]) ? node30603 : node30576;
											assign node30576 = (inp[15]) ? node30590 : node30577;
												assign node30577 = (inp[10]) ? node30585 : node30578;
													assign node30578 = (inp[12]) ? node30582 : node30579;
														assign node30579 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30582 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node30585 = (inp[9]) ? node30587 : 16'b0000000001111111;
														assign node30587 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30590 = (inp[12]) ? node30598 : node30591;
													assign node30591 = (inp[11]) ? node30595 : node30592;
														assign node30592 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30595 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30598 = (inp[13]) ? node30600 : 16'b0000000000111111;
														assign node30600 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30603 = (inp[12]) ? node30621 : node30604;
												assign node30604 = (inp[9]) ? node30612 : node30605;
													assign node30605 = (inp[11]) ? node30609 : node30606;
														assign node30606 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30609 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30612 = (inp[15]) ? node30616 : node30613;
														assign node30613 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30616 = (inp[10]) ? 16'b0000000000011111 : node30617;
															assign node30617 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30621 = (inp[15]) ? node30625 : node30622;
													assign node30622 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30625 = (inp[11]) ? node30627 : 16'b0000000000011111;
														assign node30627 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node30630 = (inp[13]) ? node30650 : node30631;
											assign node30631 = (inp[9]) ? node30639 : node30632;
												assign node30632 = (inp[10]) ? 16'b0000000000111111 : node30633;
													assign node30633 = (inp[12]) ? 16'b0000000000111111 : node30634;
														assign node30634 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30639 = (inp[12]) ? node30645 : node30640;
													assign node30640 = (inp[4]) ? node30642 : 16'b0000000000111111;
														assign node30642 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30645 = (inp[15]) ? 16'b0000000000011111 : node30646;
														assign node30646 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30650 = (inp[9]) ? node30666 : node30651;
												assign node30651 = (inp[15]) ? node30659 : node30652;
													assign node30652 = (inp[11]) ? node30656 : node30653;
														assign node30653 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30656 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30659 = (inp[10]) ? node30663 : node30660;
														assign node30660 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30663 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30666 = (inp[10]) ? 16'b0000000000001111 : node30667;
													assign node30667 = (inp[11]) ? node30669 : 16'b0000000000011111;
														assign node30669 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node30673 = (inp[2]) ? node30933 : node30674;
								assign node30674 = (inp[13]) ? node30800 : node30675;
									assign node30675 = (inp[4]) ? node30727 : node30676;
										assign node30676 = (inp[12]) ? node30700 : node30677;
											assign node30677 = (inp[9]) ? node30689 : node30678;
												assign node30678 = (inp[10]) ? node30682 : node30679;
													assign node30679 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node30682 = (inp[11]) ? 16'b0000000011111111 : node30683;
														assign node30683 = (inp[1]) ? node30685 : 16'b0000001111111111;
															assign node30685 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node30689 = (inp[10]) ? node30693 : node30690;
													assign node30690 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30693 = (inp[11]) ? 16'b0000000011111111 : node30694;
														assign node30694 = (inp[15]) ? node30696 : 16'b0000000001111111;
															assign node30696 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30700 = (inp[1]) ? node30714 : node30701;
												assign node30701 = (inp[15]) ? node30709 : node30702;
													assign node30702 = (inp[10]) ? node30706 : node30703;
														assign node30703 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30706 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30709 = (inp[14]) ? 16'b0000000000111111 : node30710;
														assign node30710 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30714 = (inp[10]) ? node30722 : node30715;
													assign node30715 = (inp[9]) ? node30717 : 16'b0000000011111111;
														assign node30717 = (inp[14]) ? node30719 : 16'b0000000001111111;
															assign node30719 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30722 = (inp[9]) ? 16'b0000000000111111 : node30723;
														assign node30723 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node30727 = (inp[1]) ? node30765 : node30728;
											assign node30728 = (inp[9]) ? node30750 : node30729;
												assign node30729 = (inp[15]) ? node30739 : node30730;
													assign node30730 = (inp[14]) ? node30734 : node30731;
														assign node30731 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node30734 = (inp[10]) ? node30736 : 16'b0000000011111111;
															assign node30736 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30739 = (inp[10]) ? node30747 : node30740;
														assign node30740 = (inp[12]) ? node30742 : 16'b0000000011111111;
															assign node30742 = (inp[14]) ? 16'b0000000001111111 : node30743;
																assign node30743 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30747 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node30750 = (inp[14]) ? node30758 : node30751;
													assign node30751 = (inp[15]) ? node30755 : node30752;
														assign node30752 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30755 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30758 = (inp[11]) ? node30762 : node30759;
														assign node30759 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30762 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30765 = (inp[14]) ? node30787 : node30766;
												assign node30766 = (inp[9]) ? node30776 : node30767;
													assign node30767 = (inp[11]) ? node30769 : 16'b0000000001111111;
														assign node30769 = (inp[12]) ? 16'b0000000000011111 : node30770;
															assign node30770 = (inp[10]) ? node30772 : 16'b0000000001111111;
																assign node30772 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30776 = (inp[12]) ? node30782 : node30777;
														assign node30777 = (inp[15]) ? 16'b0000000000111111 : node30778;
															assign node30778 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30782 = (inp[11]) ? node30784 : 16'b0000000000111111;
															assign node30784 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30787 = (inp[10]) ? node30793 : node30788;
													assign node30788 = (inp[15]) ? node30790 : 16'b0000000001111111;
														assign node30790 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30793 = (inp[9]) ? node30797 : node30794;
														assign node30794 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30797 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node30800 = (inp[10]) ? node30876 : node30801;
										assign node30801 = (inp[1]) ? node30839 : node30802;
											assign node30802 = (inp[4]) ? node30824 : node30803;
												assign node30803 = (inp[15]) ? node30813 : node30804;
													assign node30804 = (inp[9]) ? node30808 : node30805;
														assign node30805 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30808 = (inp[14]) ? 16'b0000000001111111 : node30809;
															assign node30809 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30813 = (inp[14]) ? node30817 : node30814;
														assign node30814 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node30817 = (inp[12]) ? node30819 : 16'b0000000001111111;
															assign node30819 = (inp[11]) ? 16'b0000000000111111 : node30820;
																assign node30820 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30824 = (inp[9]) ? node30832 : node30825;
													assign node30825 = (inp[14]) ? node30829 : node30826;
														assign node30826 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30829 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30832 = (inp[11]) ? node30836 : node30833;
														assign node30833 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30836 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30839 = (inp[9]) ? node30861 : node30840;
												assign node30840 = (inp[11]) ? node30850 : node30841;
													assign node30841 = (inp[15]) ? node30845 : node30842;
														assign node30842 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30845 = (inp[12]) ? node30847 : 16'b0000000001111111;
															assign node30847 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30850 = (inp[4]) ? node30858 : node30851;
														assign node30851 = (inp[15]) ? node30853 : 16'b0000000001111111;
															assign node30853 = (inp[14]) ? 16'b0000000000111111 : node30854;
																assign node30854 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30858 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node30861 = (inp[14]) ? node30867 : node30862;
													assign node30862 = (inp[15]) ? node30864 : 16'b0000000001111111;
														assign node30864 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30867 = (inp[11]) ? node30871 : node30868;
														assign node30868 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000011111;
														assign node30871 = (inp[12]) ? 16'b0000000000001111 : node30872;
															assign node30872 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node30876 = (inp[12]) ? node30902 : node30877;
											assign node30877 = (inp[15]) ? node30889 : node30878;
												assign node30878 = (inp[4]) ? node30884 : node30879;
													assign node30879 = (inp[11]) ? 16'b0000000001111111 : node30880;
														assign node30880 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30884 = (inp[11]) ? 16'b0000000000111111 : node30885;
														assign node30885 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30889 = (inp[4]) ? node30893 : node30890;
													assign node30890 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node30893 = (inp[14]) ? node30897 : node30894;
														assign node30894 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30897 = (inp[1]) ? node30899 : 16'b0000000000011111;
															assign node30899 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30902 = (inp[11]) ? node30924 : node30903;
												assign node30903 = (inp[4]) ? node30909 : node30904;
													assign node30904 = (inp[1]) ? node30906 : 16'b0000000000111111;
														assign node30906 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30909 = (inp[1]) ? node30921 : node30910;
														assign node30910 = (inp[9]) ? node30916 : node30911;
															assign node30911 = (inp[14]) ? node30913 : 16'b0000000000111111;
																assign node30913 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node30916 = (inp[15]) ? node30918 : 16'b0000000000011111;
																assign node30918 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30921 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30924 = (inp[9]) ? node30926 : 16'b0000000000011111;
													assign node30926 = (inp[1]) ? node30930 : node30927;
														assign node30927 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30930 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node30933 = (inp[9]) ? node31081 : node30934;
									assign node30934 = (inp[13]) ? node31010 : node30935;
										assign node30935 = (inp[4]) ? node30969 : node30936;
											assign node30936 = (inp[12]) ? node30952 : node30937;
												assign node30937 = (inp[10]) ? node30947 : node30938;
													assign node30938 = (inp[14]) ? node30944 : node30939;
														assign node30939 = (inp[11]) ? node30941 : 16'b0000000111111111;
															assign node30941 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30944 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30947 = (inp[11]) ? 16'b0000000001111111 : node30948;
														assign node30948 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node30952 = (inp[14]) ? node30958 : node30953;
													assign node30953 = (inp[1]) ? 16'b0000000001111111 : node30954;
														assign node30954 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30958 = (inp[10]) ? node30962 : node30959;
														assign node30959 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30962 = (inp[15]) ? 16'b0000000000011111 : node30963;
															assign node30963 = (inp[1]) ? node30965 : 16'b0000000000111111;
																assign node30965 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30969 = (inp[1]) ? node30993 : node30970;
												assign node30970 = (inp[15]) ? node30980 : node30971;
													assign node30971 = (inp[12]) ? node30977 : node30972;
														assign node30972 = (inp[14]) ? 16'b0000000001111111 : node30973;
															assign node30973 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30977 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30980 = (inp[11]) ? node30986 : node30981;
														assign node30981 = (inp[10]) ? node30983 : 16'b0000000001111111;
															assign node30983 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30986 = (inp[14]) ? 16'b0000000000011111 : node30987;
															assign node30987 = (inp[12]) ? 16'b0000000000111111 : node30988;
																assign node30988 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30993 = (inp[11]) ? node30999 : node30994;
													assign node30994 = (inp[12]) ? 16'b0000000000111111 : node30995;
														assign node30995 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30999 = (inp[14]) ? node31005 : node31000;
														assign node31000 = (inp[15]) ? node31002 : 16'b0000000000111111;
															assign node31002 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node31005 = (inp[10]) ? 16'b0000000000000111 : node31006;
															assign node31006 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node31010 = (inp[10]) ? node31046 : node31011;
											assign node31011 = (inp[4]) ? node31025 : node31012;
												assign node31012 = (inp[14]) ? 16'b0000000000111111 : node31013;
													assign node31013 = (inp[1]) ? node31017 : node31014;
														assign node31014 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31017 = (inp[11]) ? node31019 : 16'b0000000001111111;
															assign node31019 = (inp[15]) ? 16'b0000000000111111 : node31020;
																assign node31020 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31025 = (inp[12]) ? node31033 : node31026;
													assign node31026 = (inp[1]) ? node31030 : node31027;
														assign node31027 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31030 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31033 = (inp[15]) ? node31037 : node31034;
														assign node31034 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node31037 = (inp[14]) ? node31043 : node31038;
															assign node31038 = (inp[1]) ? node31040 : 16'b0000000000011111;
																assign node31040 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node31043 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node31046 = (inp[14]) ? node31058 : node31047;
												assign node31047 = (inp[1]) ? node31053 : node31048;
													assign node31048 = (inp[12]) ? node31050 : 16'b0000000000111111;
														assign node31050 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node31053 = (inp[4]) ? node31055 : 16'b0000000000011111;
														assign node31055 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node31058 = (inp[4]) ? node31062 : node31059;
													assign node31059 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000001111;
													assign node31062 = (inp[12]) ? node31072 : node31063;
														assign node31063 = (inp[1]) ? node31067 : node31064;
															assign node31064 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node31067 = (inp[15]) ? node31069 : 16'b0000000000001111;
																assign node31069 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node31072 = (inp[15]) ? node31078 : node31073;
															assign node31073 = (inp[11]) ? node31075 : 16'b0000000000001111;
																assign node31075 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node31078 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node31081 = (inp[15]) ? node31145 : node31082;
										assign node31082 = (inp[11]) ? node31114 : node31083;
											assign node31083 = (inp[14]) ? node31101 : node31084;
												assign node31084 = (inp[10]) ? node31098 : node31085;
													assign node31085 = (inp[13]) ? node31091 : node31086;
														assign node31086 = (inp[4]) ? 16'b0000000001111111 : node31087;
															assign node31087 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node31091 = (inp[4]) ? 16'b0000000000111111 : node31092;
															assign node31092 = (inp[1]) ? node31094 : 16'b0000000001111111;
																assign node31094 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31098 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node31101 = (inp[13]) ? node31109 : node31102;
													assign node31102 = (inp[4]) ? node31106 : node31103;
														assign node31103 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31106 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31109 = (inp[1]) ? node31111 : 16'b0000000000011111;
														assign node31111 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node31114 = (inp[4]) ? node31128 : node31115;
												assign node31115 = (inp[10]) ? node31123 : node31116;
													assign node31116 = (inp[13]) ? node31120 : node31117;
														assign node31117 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31120 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31123 = (inp[12]) ? node31125 : 16'b0000000000011111;
														assign node31125 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node31128 = (inp[10]) ? node31140 : node31129;
													assign node31129 = (inp[1]) ? node31131 : 16'b0000000000011111;
														assign node31131 = (inp[14]) ? node31135 : node31132;
															assign node31132 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node31135 = (inp[13]) ? node31137 : 16'b0000000000001111;
																assign node31137 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node31140 = (inp[1]) ? node31142 : 16'b0000000000001111;
														assign node31142 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node31145 = (inp[12]) ? node31173 : node31146;
											assign node31146 = (inp[13]) ? node31152 : node31147;
												assign node31147 = (inp[14]) ? 16'b0000000000011111 : node31148;
													assign node31148 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node31152 = (inp[1]) ? node31166 : node31153;
													assign node31153 = (inp[14]) ? node31159 : node31154;
														assign node31154 = (inp[11]) ? 16'b0000000000011111 : node31155;
															assign node31155 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31159 = (inp[11]) ? node31161 : 16'b0000000000011111;
															assign node31161 = (inp[10]) ? node31163 : 16'b0000000000001111;
																assign node31163 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node31166 = (inp[14]) ? 16'b0000000000000111 : node31167;
														assign node31167 = (inp[10]) ? node31169 : 16'b0000000000001111;
															assign node31169 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node31173 = (inp[13]) ? node31195 : node31174;
												assign node31174 = (inp[4]) ? node31182 : node31175;
													assign node31175 = (inp[1]) ? node31177 : 16'b0000000000011111;
														assign node31177 = (inp[11]) ? 16'b0000000000001111 : node31178;
															assign node31178 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node31182 = (inp[10]) ? node31190 : node31183;
														assign node31183 = (inp[14]) ? node31185 : 16'b0000000000001111;
															assign node31185 = (inp[1]) ? node31187 : 16'b0000000000001111;
																assign node31187 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node31190 = (inp[14]) ? 16'b0000000000000111 : node31191;
															assign node31191 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node31195 = (inp[11]) ? node31201 : node31196;
													assign node31196 = (inp[10]) ? 16'b0000000000000111 : node31197;
														assign node31197 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000001111;
													assign node31201 = (inp[4]) ? node31211 : node31202;
														assign node31202 = (inp[1]) ? node31206 : node31203;
															assign node31203 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node31206 = (inp[14]) ? node31208 : 16'b0000000000000111;
																assign node31208 = (inp[10]) ? 16'b0000000000000011 : 16'b0000000000000111;
														assign node31211 = (inp[10]) ? node31213 : 16'b0000000000000011;
															assign node31213 = (inp[14]) ? node31215 : 16'b0000000000000011;
																assign node31215 = (inp[1]) ? 16'b0000000000000001 : 16'b0000000000000011;
					assign node31218 = (inp[11]) ? node32276 : node31219;
						assign node31219 = (inp[13]) ? node31767 : node31220;
							assign node31220 = (inp[12]) ? node31508 : node31221;
								assign node31221 = (inp[4]) ? node31359 : node31222;
									assign node31222 = (inp[2]) ? node31294 : node31223;
										assign node31223 = (inp[10]) ? node31263 : node31224;
											assign node31224 = (inp[8]) ? node31246 : node31225;
												assign node31225 = (inp[6]) ? node31235 : node31226;
													assign node31226 = (inp[15]) ? 16'b0000001111111111 : node31227;
														assign node31227 = (inp[9]) ? node31231 : node31228;
															assign node31228 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
															assign node31231 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node31235 = (inp[9]) ? node31243 : node31236;
														assign node31236 = (inp[14]) ? node31240 : node31237;
															assign node31237 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
															assign node31240 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node31243 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node31246 = (inp[6]) ? node31256 : node31247;
													assign node31247 = (inp[1]) ? node31253 : node31248;
														assign node31248 = (inp[14]) ? 16'b0000000111111111 : node31249;
															assign node31249 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node31253 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node31256 = (inp[15]) ? node31258 : 16'b0000001111111111;
														assign node31258 = (inp[1]) ? 16'b0000000001111111 : node31259;
															assign node31259 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node31263 = (inp[14]) ? node31277 : node31264;
												assign node31264 = (inp[9]) ? 16'b0000000001111111 : node31265;
													assign node31265 = (inp[15]) ? node31267 : 16'b0000001111111111;
														assign node31267 = (inp[8]) ? node31271 : node31268;
															assign node31268 = (inp[6]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node31271 = (inp[1]) ? 16'b0000000011111111 : node31272;
																assign node31272 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node31277 = (inp[8]) ? node31289 : node31278;
													assign node31278 = (inp[1]) ? node31284 : node31279;
														assign node31279 = (inp[15]) ? node31281 : 16'b0000000111111111;
															assign node31281 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31284 = (inp[15]) ? node31286 : 16'b0000000011111111;
															assign node31286 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31289 = (inp[9]) ? node31291 : 16'b0000000011111111;
														assign node31291 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node31294 = (inp[10]) ? node31326 : node31295;
											assign node31295 = (inp[15]) ? node31317 : node31296;
												assign node31296 = (inp[14]) ? node31310 : node31297;
													assign node31297 = (inp[9]) ? node31305 : node31298;
														assign node31298 = (inp[6]) ? node31300 : 16'b0000001111111111;
															assign node31300 = (inp[8]) ? 16'b0000000111111111 : node31301;
																assign node31301 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node31305 = (inp[1]) ? 16'b0000000011111111 : node31306;
															assign node31306 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31310 = (inp[8]) ? node31312 : 16'b0000000011111111;
														assign node31312 = (inp[1]) ? 16'b0000000001111111 : node31313;
															assign node31313 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31317 = (inp[1]) ? 16'b0000000001111111 : node31318;
													assign node31318 = (inp[9]) ? node31322 : node31319;
														assign node31319 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31322 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node31326 = (inp[9]) ? node31338 : node31327;
												assign node31327 = (inp[8]) ? node31331 : node31328;
													assign node31328 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31331 = (inp[14]) ? node31333 : 16'b0000000011111111;
														assign node31333 = (inp[1]) ? node31335 : 16'b0000000001111111;
															assign node31335 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31338 = (inp[1]) ? node31350 : node31339;
													assign node31339 = (inp[14]) ? node31343 : node31340;
														assign node31340 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31343 = (inp[6]) ? 16'b0000000000111111 : node31344;
															assign node31344 = (inp[15]) ? node31346 : 16'b0000000001111111;
																assign node31346 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31350 = (inp[15]) ? node31354 : node31351;
														assign node31351 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31354 = (inp[14]) ? node31356 : 16'b0000000000111111;
															assign node31356 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node31359 = (inp[8]) ? node31435 : node31360;
										assign node31360 = (inp[10]) ? node31400 : node31361;
											assign node31361 = (inp[9]) ? node31381 : node31362;
												assign node31362 = (inp[6]) ? node31376 : node31363;
													assign node31363 = (inp[14]) ? node31373 : node31364;
														assign node31364 = (inp[1]) ? node31366 : 16'b0000001111111111;
															assign node31366 = (inp[2]) ? node31370 : node31367;
																assign node31367 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
																assign node31370 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31373 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31376 = (inp[14]) ? 16'b0000000011111111 : node31377;
														assign node31377 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31381 = (inp[1]) ? node31395 : node31382;
													assign node31382 = (inp[15]) ? node31388 : node31383;
														assign node31383 = (inp[14]) ? 16'b0000000011111111 : node31384;
															assign node31384 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31388 = (inp[14]) ? node31390 : 16'b0000000011111111;
															assign node31390 = (inp[6]) ? 16'b0000000001111111 : node31391;
																assign node31391 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31395 = (inp[6]) ? node31397 : 16'b0000000001111111;
														assign node31397 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node31400 = (inp[1]) ? node31422 : node31401;
												assign node31401 = (inp[14]) ? node31417 : node31402;
													assign node31402 = (inp[2]) ? node31412 : node31403;
														assign node31403 = (inp[6]) ? node31409 : node31404;
															assign node31404 = (inp[9]) ? node31406 : 16'b0000000111111111;
																assign node31406 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
															assign node31409 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31412 = (inp[9]) ? node31414 : 16'b0000000011111111;
															assign node31414 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31417 = (inp[15]) ? node31419 : 16'b0000000001111111;
														assign node31419 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31422 = (inp[6]) ? node31424 : 16'b0000000001111111;
													assign node31424 = (inp[9]) ? node31428 : node31425;
														assign node31425 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31428 = (inp[2]) ? 16'b0000000000011111 : node31429;
															assign node31429 = (inp[15]) ? 16'b0000000000111111 : node31430;
																assign node31430 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node31435 = (inp[1]) ? node31473 : node31436;
											assign node31436 = (inp[2]) ? node31452 : node31437;
												assign node31437 = (inp[6]) ? node31443 : node31438;
													assign node31438 = (inp[14]) ? 16'b0000000011111111 : node31439;
														assign node31439 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31443 = (inp[10]) ? node31447 : node31444;
														assign node31444 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node31447 = (inp[15]) ? node31449 : 16'b0000000001111111;
															assign node31449 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31452 = (inp[10]) ? node31464 : node31453;
													assign node31453 = (inp[9]) ? node31457 : node31454;
														assign node31454 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31457 = (inp[6]) ? node31459 : 16'b0000000001111111;
															assign node31459 = (inp[14]) ? 16'b0000000000111111 : node31460;
																assign node31460 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31464 = (inp[9]) ? 16'b0000000000011111 : node31465;
														assign node31465 = (inp[14]) ? node31467 : 16'b0000000001111111;
															assign node31467 = (inp[6]) ? 16'b0000000000111111 : node31468;
																assign node31468 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node31473 = (inp[9]) ? node31491 : node31474;
												assign node31474 = (inp[6]) ? node31484 : node31475;
													assign node31475 = (inp[2]) ? 16'b0000000001111111 : node31476;
														assign node31476 = (inp[14]) ? node31478 : 16'b0000000011111111;
															assign node31478 = (inp[10]) ? 16'b0000000001111111 : node31479;
																assign node31479 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31484 = (inp[15]) ? 16'b0000000000111111 : node31485;
														assign node31485 = (inp[14]) ? 16'b0000000000111111 : node31486;
															assign node31486 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31491 = (inp[15]) ? node31501 : node31492;
													assign node31492 = (inp[6]) ? 16'b0000000000011111 : node31493;
														assign node31493 = (inp[2]) ? node31495 : 16'b0000000001111111;
															assign node31495 = (inp[10]) ? 16'b0000000000111111 : node31496;
																assign node31496 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31501 = (inp[10]) ? node31503 : 16'b0000000000011111;
														assign node31503 = (inp[14]) ? node31505 : 16'b0000000000011111;
															assign node31505 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node31508 = (inp[10]) ? node31640 : node31509;
									assign node31509 = (inp[2]) ? node31571 : node31510;
										assign node31510 = (inp[1]) ? node31540 : node31511;
											assign node31511 = (inp[8]) ? node31525 : node31512;
												assign node31512 = (inp[4]) ? node31520 : node31513;
													assign node31513 = (inp[15]) ? node31517 : node31514;
														assign node31514 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node31517 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31520 = (inp[9]) ? node31522 : 16'b0000000111111111;
														assign node31522 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31525 = (inp[6]) ? node31533 : node31526;
													assign node31526 = (inp[9]) ? node31530 : node31527;
														assign node31527 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31530 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31533 = (inp[14]) ? node31537 : node31534;
														assign node31534 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31537 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node31540 = (inp[14]) ? node31556 : node31541;
												assign node31541 = (inp[15]) ? node31549 : node31542;
													assign node31542 = (inp[9]) ? node31546 : node31543;
														assign node31543 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31546 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31549 = (inp[8]) ? node31553 : node31550;
														assign node31550 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31553 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31556 = (inp[9]) ? node31564 : node31557;
													assign node31557 = (inp[15]) ? node31561 : node31558;
														assign node31558 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node31561 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31564 = (inp[8]) ? node31568 : node31565;
														assign node31565 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31568 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node31571 = (inp[9]) ? node31599 : node31572;
											assign node31572 = (inp[4]) ? node31584 : node31573;
												assign node31573 = (inp[15]) ? node31579 : node31574;
													assign node31574 = (inp[6]) ? 16'b0000000011111111 : node31575;
														assign node31575 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node31579 = (inp[8]) ? node31581 : 16'b0000000001111111;
														assign node31581 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31584 = (inp[1]) ? node31592 : node31585;
													assign node31585 = (inp[8]) ? node31589 : node31586;
														assign node31586 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31589 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31592 = (inp[6]) ? node31596 : node31593;
														assign node31593 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31596 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node31599 = (inp[15]) ? node31615 : node31600;
												assign node31600 = (inp[4]) ? node31606 : node31601;
													assign node31601 = (inp[14]) ? node31603 : 16'b0000000011111111;
														assign node31603 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31606 = (inp[8]) ? node31612 : node31607;
														assign node31607 = (inp[6]) ? 16'b0000000000111111 : node31608;
															assign node31608 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31612 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node31615 = (inp[1]) ? node31627 : node31616;
													assign node31616 = (inp[6]) ? node31620 : node31617;
														assign node31617 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31620 = (inp[4]) ? 16'b0000000000011111 : node31621;
															assign node31621 = (inp[8]) ? node31623 : 16'b0000000000111111;
																assign node31623 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31627 = (inp[8]) ? node31635 : node31628;
														assign node31628 = (inp[6]) ? node31630 : 16'b0000000000111111;
															assign node31630 = (inp[4]) ? node31632 : 16'b0000000000011111;
																assign node31632 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node31635 = (inp[6]) ? node31637 : 16'b0000000000001111;
															assign node31637 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node31640 = (inp[8]) ? node31702 : node31641;
										assign node31641 = (inp[4]) ? node31671 : node31642;
											assign node31642 = (inp[14]) ? node31654 : node31643;
												assign node31643 = (inp[1]) ? node31647 : node31644;
													assign node31644 = (inp[6]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31647 = (inp[15]) ? node31651 : node31648;
														assign node31648 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node31651 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31654 = (inp[15]) ? node31660 : node31655;
													assign node31655 = (inp[9]) ? node31657 : 16'b0000000011111111;
														assign node31657 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31660 = (inp[6]) ? node31666 : node31661;
														assign node31661 = (inp[9]) ? 16'b0000000000111111 : node31662;
															assign node31662 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31666 = (inp[2]) ? node31668 : 16'b0000000000111111;
															assign node31668 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node31671 = (inp[15]) ? node31689 : node31672;
												assign node31672 = (inp[14]) ? node31678 : node31673;
													assign node31673 = (inp[1]) ? node31675 : 16'b0000000001111111;
														assign node31675 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31678 = (inp[1]) ? node31682 : node31679;
														assign node31679 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31682 = (inp[6]) ? node31684 : 16'b0000000000111111;
															assign node31684 = (inp[2]) ? 16'b0000000000011111 : node31685;
																assign node31685 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node31689 = (inp[6]) ? node31697 : node31690;
													assign node31690 = (inp[1]) ? node31692 : 16'b0000000000111111;
														assign node31692 = (inp[14]) ? node31694 : 16'b0000000000111111;
															assign node31694 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31697 = (inp[2]) ? node31699 : 16'b0000000000111111;
														assign node31699 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node31702 = (inp[14]) ? node31738 : node31703;
											assign node31703 = (inp[4]) ? node31715 : node31704;
												assign node31704 = (inp[9]) ? node31708 : node31705;
													assign node31705 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31708 = (inp[6]) ? node31710 : 16'b0000000001111111;
														assign node31710 = (inp[15]) ? 16'b0000000000011111 : node31711;
															assign node31711 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31715 = (inp[9]) ? node31729 : node31716;
													assign node31716 = (inp[6]) ? node31718 : 16'b0000000001111111;
														assign node31718 = (inp[15]) ? node31724 : node31719;
															assign node31719 = (inp[1]) ? 16'b0000000000111111 : node31720;
																assign node31720 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node31724 = (inp[1]) ? 16'b0000000000011111 : node31725;
																assign node31725 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31729 = (inp[15]) ? 16'b0000000000011111 : node31730;
														assign node31730 = (inp[1]) ? 16'b0000000000011111 : node31731;
															assign node31731 = (inp[6]) ? node31733 : 16'b0000000000111111;
																assign node31733 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node31738 = (inp[9]) ? node31746 : node31739;
												assign node31739 = (inp[15]) ? 16'b0000000000011111 : node31740;
													assign node31740 = (inp[6]) ? 16'b0000000000011111 : node31741;
														assign node31741 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31746 = (inp[15]) ? node31754 : node31747;
													assign node31747 = (inp[2]) ? node31749 : 16'b0000000000011111;
														assign node31749 = (inp[1]) ? node31751 : 16'b0000000000011111;
															assign node31751 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node31754 = (inp[2]) ? node31760 : node31755;
														assign node31755 = (inp[6]) ? 16'b0000000000001111 : node31756;
															assign node31756 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node31760 = (inp[6]) ? 16'b0000000000000111 : node31761;
															assign node31761 = (inp[4]) ? node31763 : 16'b0000000000001111;
																assign node31763 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node31767 = (inp[8]) ? node32021 : node31768;
								assign node31768 = (inp[2]) ? node31874 : node31769;
									assign node31769 = (inp[4]) ? node31823 : node31770;
										assign node31770 = (inp[9]) ? node31806 : node31771;
											assign node31771 = (inp[6]) ? node31791 : node31772;
												assign node31772 = (inp[1]) ? node31786 : node31773;
													assign node31773 = (inp[10]) ? node31781 : node31774;
														assign node31774 = (inp[14]) ? 16'b0000000111111111 : node31775;
															assign node31775 = (inp[12]) ? node31777 : 16'b0000001111111111;
																assign node31777 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node31781 = (inp[15]) ? node31783 : 16'b0000000111111111;
															assign node31783 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31786 = (inp[15]) ? node31788 : 16'b0000000111111111;
														assign node31788 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31791 = (inp[14]) ? node31799 : node31792;
													assign node31792 = (inp[12]) ? 16'b0000000001111111 : node31793;
														assign node31793 = (inp[15]) ? 16'b0000000011111111 : node31794;
															assign node31794 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node31799 = (inp[1]) ? 16'b0000000000111111 : node31800;
														assign node31800 = (inp[12]) ? 16'b0000000001111111 : node31801;
															assign node31801 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node31806 = (inp[10]) ? node31816 : node31807;
												assign node31807 = (inp[14]) ? node31811 : node31808;
													assign node31808 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node31811 = (inp[15]) ? 16'b0000000001111111 : node31812;
														assign node31812 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node31816 = (inp[12]) ? 16'b0000000000111111 : node31817;
													assign node31817 = (inp[14]) ? node31819 : 16'b0000000001111111;
														assign node31819 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node31823 = (inp[15]) ? node31851 : node31824;
											assign node31824 = (inp[6]) ? node31836 : node31825;
												assign node31825 = (inp[1]) ? node31833 : node31826;
													assign node31826 = (inp[14]) ? 16'b0000000011111111 : node31827;
														assign node31827 = (inp[10]) ? 16'b0000000011111111 : node31828;
															assign node31828 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node31833 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node31836 = (inp[14]) ? node31842 : node31837;
													assign node31837 = (inp[12]) ? 16'b0000000001111111 : node31838;
														assign node31838 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31842 = (inp[9]) ? node31848 : node31843;
														assign node31843 = (inp[12]) ? node31845 : 16'b0000000001111111;
															assign node31845 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31848 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node31851 = (inp[1]) ? node31859 : node31852;
												assign node31852 = (inp[10]) ? 16'b0000000000111111 : node31853;
													assign node31853 = (inp[6]) ? node31855 : 16'b0000000001111111;
														assign node31855 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31859 = (inp[12]) ? node31865 : node31860;
													assign node31860 = (inp[6]) ? 16'b0000000000111111 : node31861;
														assign node31861 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node31865 = (inp[10]) ? node31871 : node31866;
														assign node31866 = (inp[14]) ? 16'b0000000000011111 : node31867;
															assign node31867 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node31871 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node31874 = (inp[12]) ? node31946 : node31875;
										assign node31875 = (inp[9]) ? node31915 : node31876;
											assign node31876 = (inp[4]) ? node31896 : node31877;
												assign node31877 = (inp[6]) ? node31885 : node31878;
													assign node31878 = (inp[10]) ? node31882 : node31879;
														assign node31879 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node31882 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node31885 = (inp[10]) ? node31893 : node31886;
														assign node31886 = (inp[14]) ? node31888 : 16'b0000000011111111;
															assign node31888 = (inp[1]) ? 16'b0000000001111111 : node31889;
																assign node31889 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31893 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31896 = (inp[14]) ? node31910 : node31897;
													assign node31897 = (inp[6]) ? node31905 : node31898;
														assign node31898 = (inp[15]) ? node31900 : 16'b0000000011111111;
															assign node31900 = (inp[10]) ? 16'b0000000001111111 : node31901;
																assign node31901 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31905 = (inp[10]) ? 16'b0000000000111111 : node31906;
															assign node31906 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31910 = (inp[15]) ? node31912 : 16'b0000000000111111;
														assign node31912 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node31915 = (inp[10]) ? node31933 : node31916;
												assign node31916 = (inp[15]) ? node31924 : node31917;
													assign node31917 = (inp[6]) ? node31921 : node31918;
														assign node31918 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node31921 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node31924 = (inp[14]) ? 16'b0000000000111111 : node31925;
														assign node31925 = (inp[1]) ? 16'b0000000000111111 : node31926;
															assign node31926 = (inp[6]) ? node31928 : 16'b0000000001111111;
																assign node31928 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node31933 = (inp[4]) ? node31939 : node31934;
													assign node31934 = (inp[1]) ? node31936 : 16'b0000000000111111;
														assign node31936 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node31939 = (inp[1]) ? node31943 : node31940;
														assign node31940 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node31943 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node31946 = (inp[15]) ? node31978 : node31947;
											assign node31947 = (inp[6]) ? node31961 : node31948;
												assign node31948 = (inp[10]) ? node31950 : 16'b0000000001111111;
													assign node31950 = (inp[4]) ? node31958 : node31951;
														assign node31951 = (inp[14]) ? node31953 : 16'b0000000001111111;
															assign node31953 = (inp[1]) ? 16'b0000000000111111 : node31954;
																assign node31954 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31958 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node31961 = (inp[14]) ? node31969 : node31962;
													assign node31962 = (inp[9]) ? node31966 : node31963;
														assign node31963 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31966 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31969 = (inp[1]) ? node31971 : 16'b0000000000111111;
														assign node31971 = (inp[9]) ? 16'b0000000000001111 : node31972;
															assign node31972 = (inp[4]) ? 16'b0000000000011111 : node31973;
																assign node31973 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node31978 = (inp[6]) ? node32000 : node31979;
												assign node31979 = (inp[9]) ? node31991 : node31980;
													assign node31980 = (inp[10]) ? node31984 : node31981;
														assign node31981 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node31984 = (inp[14]) ? node31986 : 16'b0000000000111111;
															assign node31986 = (inp[4]) ? 16'b0000000000011111 : node31987;
																assign node31987 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node31991 = (inp[10]) ? node31995 : node31992;
														assign node31992 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node31995 = (inp[1]) ? node31997 : 16'b0000000000011111;
															assign node31997 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node32000 = (inp[4]) ? node32016 : node32001;
													assign node32001 = (inp[1]) ? node32007 : node32002;
														assign node32002 = (inp[9]) ? 16'b0000000000011111 : node32003;
															assign node32003 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32007 = (inp[10]) ? node32011 : node32008;
															assign node32008 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
															assign node32011 = (inp[14]) ? 16'b0000000000001111 : node32012;
																assign node32012 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32016 = (inp[9]) ? 16'b0000000000001111 : node32017;
														assign node32017 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node32021 = (inp[9]) ? node32139 : node32022;
									assign node32022 = (inp[4]) ? node32074 : node32023;
										assign node32023 = (inp[1]) ? node32043 : node32024;
											assign node32024 = (inp[15]) ? node32038 : node32025;
												assign node32025 = (inp[12]) ? node32031 : node32026;
													assign node32026 = (inp[6]) ? 16'b0000000011111111 : node32027;
														assign node32027 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node32031 = (inp[6]) ? node32035 : node32032;
														assign node32032 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32035 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32038 = (inp[12]) ? node32040 : 16'b0000000001111111;
													assign node32040 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node32043 = (inp[14]) ? node32055 : node32044;
												assign node32044 = (inp[15]) ? node32050 : node32045;
													assign node32045 = (inp[10]) ? 16'b0000000000111111 : node32046;
														assign node32046 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32050 = (inp[2]) ? 16'b0000000000111111 : node32051;
														assign node32051 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32055 = (inp[2]) ? node32067 : node32056;
													assign node32056 = (inp[10]) ? node32062 : node32057;
														assign node32057 = (inp[12]) ? node32059 : 16'b0000000001111111;
															assign node32059 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32062 = (inp[15]) ? node32064 : 16'b0000000000111111;
															assign node32064 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32067 = (inp[6]) ? 16'b0000000000011111 : node32068;
														assign node32068 = (inp[12]) ? node32070 : 16'b0000000000111111;
															assign node32070 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node32074 = (inp[15]) ? node32114 : node32075;
											assign node32075 = (inp[12]) ? node32097 : node32076;
												assign node32076 = (inp[2]) ? node32090 : node32077;
													assign node32077 = (inp[6]) ? node32083 : node32078;
														assign node32078 = (inp[10]) ? 16'b0000000001111111 : node32079;
															assign node32079 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32083 = (inp[1]) ? node32085 : 16'b0000000001111111;
															assign node32085 = (inp[14]) ? 16'b0000000000111111 : node32086;
																assign node32086 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32090 = (inp[1]) ? node32092 : 16'b0000000001111111;
														assign node32092 = (inp[10]) ? node32094 : 16'b0000000000111111;
															assign node32094 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32097 = (inp[1]) ? node32105 : node32098;
													assign node32098 = (inp[14]) ? node32102 : node32099;
														assign node32099 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32102 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32105 = (inp[10]) ? 16'b0000000000011111 : node32106;
														assign node32106 = (inp[14]) ? node32108 : 16'b0000000000111111;
															assign node32108 = (inp[2]) ? 16'b0000000000011111 : node32109;
																assign node32109 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node32114 = (inp[6]) ? node32134 : node32115;
												assign node32115 = (inp[2]) ? node32129 : node32116;
													assign node32116 = (inp[12]) ? node32122 : node32117;
														assign node32117 = (inp[10]) ? 16'b0000000000111111 : node32118;
															assign node32118 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32122 = (inp[14]) ? 16'b0000000000011111 : node32123;
															assign node32123 = (inp[1]) ? node32125 : 16'b0000000000111111;
																assign node32125 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32129 = (inp[12]) ? 16'b0000000000011111 : node32130;
														assign node32130 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32134 = (inp[12]) ? 16'b0000000000001111 : node32135;
													assign node32135 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node32139 = (inp[4]) ? node32213 : node32140;
										assign node32140 = (inp[15]) ? node32182 : node32141;
											assign node32141 = (inp[10]) ? node32161 : node32142;
												assign node32142 = (inp[1]) ? node32154 : node32143;
													assign node32143 = (inp[12]) ? node32149 : node32144;
														assign node32144 = (inp[2]) ? 16'b0000000001111111 : node32145;
															assign node32145 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32149 = (inp[6]) ? node32151 : 16'b0000000001111111;
															assign node32151 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32154 = (inp[14]) ? node32158 : node32155;
														assign node32155 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32158 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32161 = (inp[6]) ? node32171 : node32162;
													assign node32162 = (inp[14]) ? node32166 : node32163;
														assign node32163 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32166 = (inp[2]) ? node32168 : 16'b0000000000111111;
															assign node32168 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32171 = (inp[1]) ? node32179 : node32172;
														assign node32172 = (inp[14]) ? node32174 : 16'b0000000000111111;
															assign node32174 = (inp[12]) ? 16'b0000000000011111 : node32175;
																assign node32175 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32179 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node32182 = (inp[1]) ? node32198 : node32183;
												assign node32183 = (inp[14]) ? node32189 : node32184;
													assign node32184 = (inp[2]) ? 16'b0000000000011111 : node32185;
														assign node32185 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32189 = (inp[12]) ? node32193 : node32190;
														assign node32190 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32193 = (inp[10]) ? node32195 : 16'b0000000000011111;
															assign node32195 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32198 = (inp[14]) ? node32206 : node32199;
													assign node32199 = (inp[12]) ? node32203 : node32200;
														assign node32200 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32203 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32206 = (inp[2]) ? 16'b0000000000000111 : node32207;
														assign node32207 = (inp[10]) ? 16'b0000000000000111 : node32208;
															assign node32208 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node32213 = (inp[2]) ? node32249 : node32214;
											assign node32214 = (inp[14]) ? node32226 : node32215;
												assign node32215 = (inp[10]) ? 16'b0000000000011111 : node32216;
													assign node32216 = (inp[15]) ? node32222 : node32217;
														assign node32217 = (inp[6]) ? 16'b0000000000111111 : node32218;
															assign node32218 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32222 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32226 = (inp[1]) ? node32236 : node32227;
													assign node32227 = (inp[6]) ? node32231 : node32228;
														assign node32228 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32231 = (inp[12]) ? node32233 : 16'b0000000000011111;
															assign node32233 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32236 = (inp[12]) ? node32240 : node32237;
														assign node32237 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node32240 = (inp[6]) ? node32244 : node32241;
															assign node32241 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
															assign node32244 = (inp[15]) ? 16'b0000000000000111 : node32245;
																assign node32245 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node32249 = (inp[1]) ? node32261 : node32250;
												assign node32250 = (inp[12]) ? 16'b0000000000001111 : node32251;
													assign node32251 = (inp[10]) ? node32253 : 16'b0000000000011111;
														assign node32253 = (inp[14]) ? node32255 : 16'b0000000000011111;
															assign node32255 = (inp[6]) ? node32257 : 16'b0000000000001111;
																assign node32257 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node32261 = (inp[10]) ? node32269 : node32262;
													assign node32262 = (inp[14]) ? 16'b0000000000000111 : node32263;
														assign node32263 = (inp[12]) ? 16'b0000000000001111 : node32264;
															assign node32264 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node32269 = (inp[15]) ? node32273 : node32270;
														assign node32270 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node32273 = (inp[14]) ? 16'b0000000000000011 : 16'b0000000000000111;
						assign node32276 = (inp[13]) ? node32826 : node32277;
							assign node32277 = (inp[4]) ? node32559 : node32278;
								assign node32278 = (inp[6]) ? node32416 : node32279;
									assign node32279 = (inp[9]) ? node32357 : node32280;
										assign node32280 = (inp[1]) ? node32322 : node32281;
											assign node32281 = (inp[12]) ? node32301 : node32282;
												assign node32282 = (inp[8]) ? node32292 : node32283;
													assign node32283 = (inp[14]) ? node32289 : node32284;
														assign node32284 = (inp[10]) ? node32286 : 16'b0000000111111111;
															assign node32286 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node32289 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node32292 = (inp[2]) ? node32298 : node32293;
														assign node32293 = (inp[10]) ? node32295 : 16'b0000000111111111;
															assign node32295 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node32298 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node32301 = (inp[8]) ? node32315 : node32302;
													assign node32302 = (inp[10]) ? node32308 : node32303;
														assign node32303 = (inp[15]) ? 16'b0000000011111111 : node32304;
															assign node32304 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node32308 = (inp[14]) ? node32310 : 16'b0000000011111111;
															assign node32310 = (inp[2]) ? 16'b0000000001111111 : node32311;
																assign node32311 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32315 = (inp[10]) ? 16'b0000000000111111 : node32316;
														assign node32316 = (inp[14]) ? 16'b0000000001111111 : node32317;
															assign node32317 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node32322 = (inp[8]) ? node32334 : node32323;
												assign node32323 = (inp[15]) ? node32329 : node32324;
													assign node32324 = (inp[14]) ? 16'b0000000011111111 : node32325;
														assign node32325 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node32329 = (inp[10]) ? 16'b0000000001111111 : node32330;
														assign node32330 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node32334 = (inp[12]) ? node32348 : node32335;
													assign node32335 = (inp[2]) ? node32341 : node32336;
														assign node32336 = (inp[15]) ? 16'b0000000011111111 : node32337;
															assign node32337 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node32341 = (inp[15]) ? 16'b0000000000111111 : node32342;
															assign node32342 = (inp[10]) ? 16'b0000000001111111 : node32343;
																assign node32343 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32348 = (inp[2]) ? node32354 : node32349;
														assign node32349 = (inp[14]) ? node32351 : 16'b0000000001111111;
															assign node32351 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node32354 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node32357 = (inp[2]) ? node32387 : node32358;
											assign node32358 = (inp[10]) ? node32380 : node32359;
												assign node32359 = (inp[8]) ? node32371 : node32360;
													assign node32360 = (inp[15]) ? node32362 : 16'b0000000011111111;
														assign node32362 = (inp[12]) ? node32364 : 16'b0000000111111111;
															assign node32364 = (inp[1]) ? node32368 : node32365;
																assign node32365 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
																assign node32368 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32371 = (inp[1]) ? node32373 : 16'b0000000001111111;
														assign node32373 = (inp[14]) ? 16'b0000000000111111 : node32374;
															assign node32374 = (inp[15]) ? 16'b0000000000111111 : node32375;
																assign node32375 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node32380 = (inp[12]) ? node32382 : 16'b0000000001111111;
													assign node32382 = (inp[8]) ? 16'b0000000000111111 : node32383;
														assign node32383 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node32387 = (inp[12]) ? node32401 : node32388;
												assign node32388 = (inp[10]) ? node32394 : node32389;
													assign node32389 = (inp[15]) ? node32391 : 16'b0000000011111111;
														assign node32391 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32394 = (inp[15]) ? node32398 : node32395;
														assign node32395 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32398 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32401 = (inp[14]) ? node32411 : node32402;
													assign node32402 = (inp[10]) ? node32406 : node32403;
														assign node32403 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32406 = (inp[8]) ? 16'b0000000000011111 : node32407;
															assign node32407 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32411 = (inp[8]) ? node32413 : 16'b0000000000011111;
														assign node32413 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node32416 = (inp[14]) ? node32484 : node32417;
										assign node32417 = (inp[8]) ? node32445 : node32418;
											assign node32418 = (inp[15]) ? node32430 : node32419;
												assign node32419 = (inp[12]) ? node32425 : node32420;
													assign node32420 = (inp[2]) ? node32422 : 16'b0000000111111111;
														assign node32422 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node32425 = (inp[9]) ? 16'b0000000001111111 : node32426;
														assign node32426 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node32430 = (inp[2]) ? node32434 : node32431;
													assign node32431 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node32434 = (inp[12]) ? node32442 : node32435;
														assign node32435 = (inp[1]) ? node32437 : 16'b0000000001111111;
															assign node32437 = (inp[9]) ? 16'b0000000000111111 : node32438;
																assign node32438 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32442 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node32445 = (inp[1]) ? node32461 : node32446;
												assign node32446 = (inp[12]) ? node32456 : node32447;
													assign node32447 = (inp[10]) ? node32451 : node32448;
														assign node32448 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32451 = (inp[2]) ? node32453 : 16'b0000000001111111;
															assign node32453 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32456 = (inp[9]) ? 16'b0000000000111111 : node32457;
														assign node32457 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32461 = (inp[2]) ? node32475 : node32462;
													assign node32462 = (inp[15]) ? node32470 : node32463;
														assign node32463 = (inp[9]) ? node32465 : 16'b0000000001111111;
															assign node32465 = (inp[12]) ? 16'b0000000000111111 : node32466;
																assign node32466 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32470 = (inp[10]) ? 16'b0000000000011111 : node32471;
															assign node32471 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32475 = (inp[9]) ? 16'b0000000000001111 : node32476;
														assign node32476 = (inp[12]) ? node32478 : 16'b0000000000111111;
															assign node32478 = (inp[15]) ? 16'b0000000000011111 : node32479;
																assign node32479 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node32484 = (inp[10]) ? node32524 : node32485;
											assign node32485 = (inp[12]) ? node32503 : node32486;
												assign node32486 = (inp[1]) ? node32496 : node32487;
													assign node32487 = (inp[8]) ? node32493 : node32488;
														assign node32488 = (inp[15]) ? node32490 : 16'b0000000011111111;
															assign node32490 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32493 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32496 = (inp[9]) ? node32498 : 16'b0000000000011111;
														assign node32498 = (inp[2]) ? 16'b0000000000111111 : node32499;
															assign node32499 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32503 = (inp[2]) ? node32515 : node32504;
													assign node32504 = (inp[15]) ? node32508 : node32505;
														assign node32505 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node32508 = (inp[8]) ? node32510 : 16'b0000000000111111;
															assign node32510 = (inp[9]) ? 16'b0000000000011111 : node32511;
																assign node32511 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32515 = (inp[15]) ? node32521 : node32516;
														assign node32516 = (inp[9]) ? 16'b0000000000011111 : node32517;
															assign node32517 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32521 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node32524 = (inp[8]) ? node32538 : node32525;
												assign node32525 = (inp[1]) ? node32529 : node32526;
													assign node32526 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32529 = (inp[12]) ? node32533 : node32530;
														assign node32530 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32533 = (inp[9]) ? 16'b0000000000001111 : node32534;
															assign node32534 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32538 = (inp[1]) ? node32544 : node32539;
													assign node32539 = (inp[9]) ? node32541 : 16'b0000000000011111;
														assign node32541 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32544 = (inp[9]) ? node32550 : node32545;
														assign node32545 = (inp[12]) ? node32547 : 16'b0000000000011111;
															assign node32547 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node32550 = (inp[2]) ? node32554 : node32551;
															assign node32551 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node32554 = (inp[12]) ? node32556 : 16'b0000000000000111;
																assign node32556 = (inp[15]) ? 16'b0000000000000011 : 16'b0000000000000111;
								assign node32559 = (inp[15]) ? node32683 : node32560;
									assign node32560 = (inp[12]) ? node32616 : node32561;
										assign node32561 = (inp[6]) ? node32585 : node32562;
											assign node32562 = (inp[8]) ? node32572 : node32563;
												assign node32563 = (inp[2]) ? node32565 : 16'b0000000011111111;
													assign node32565 = (inp[9]) ? 16'b0000000001111111 : node32566;
														assign node32566 = (inp[10]) ? node32568 : 16'b0000000011111111;
															assign node32568 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node32572 = (inp[14]) ? node32578 : node32573;
													assign node32573 = (inp[2]) ? 16'b0000000001111111 : node32574;
														assign node32574 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node32578 = (inp[1]) ? 16'b0000000000111111 : node32579;
														assign node32579 = (inp[9]) ? node32581 : 16'b0000000001111111;
															assign node32581 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node32585 = (inp[10]) ? node32603 : node32586;
												assign node32586 = (inp[8]) ? node32594 : node32587;
													assign node32587 = (inp[14]) ? 16'b0000000000111111 : node32588;
														assign node32588 = (inp[2]) ? 16'b0000000001111111 : node32589;
															assign node32589 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32594 = (inp[2]) ? node32598 : node32595;
														assign node32595 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32598 = (inp[9]) ? node32600 : 16'b0000000000111111;
															assign node32600 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32603 = (inp[2]) ? node32609 : node32604;
													assign node32604 = (inp[14]) ? 16'b0000000000111111 : node32605;
														assign node32605 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node32609 = (inp[1]) ? 16'b0000000000001111 : node32610;
														assign node32610 = (inp[9]) ? 16'b0000000000001111 : node32611;
															assign node32611 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node32616 = (inp[8]) ? node32646 : node32617;
											assign node32617 = (inp[6]) ? node32627 : node32618;
												assign node32618 = (inp[2]) ? node32620 : 16'b0000000001111111;
													assign node32620 = (inp[9]) ? node32624 : node32621;
														assign node32621 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32624 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32627 = (inp[14]) ? node32639 : node32628;
													assign node32628 = (inp[2]) ? node32634 : node32629;
														assign node32629 = (inp[1]) ? 16'b0000000000111111 : node32630;
															assign node32630 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32634 = (inp[10]) ? node32636 : 16'b0000000000111111;
															assign node32636 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32639 = (inp[2]) ? node32641 : 16'b0000000000011111;
														assign node32641 = (inp[1]) ? node32643 : 16'b0000000000011111;
															assign node32643 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node32646 = (inp[9]) ? node32668 : node32647;
												assign node32647 = (inp[10]) ? node32659 : node32648;
													assign node32648 = (inp[2]) ? node32652 : node32649;
														assign node32649 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32652 = (inp[1]) ? 16'b0000000000011111 : node32653;
															assign node32653 = (inp[6]) ? node32655 : 16'b0000000000111111;
																assign node32655 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32659 = (inp[6]) ? node32665 : node32660;
														assign node32660 = (inp[14]) ? node32662 : 16'b0000000000111111;
															assign node32662 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32665 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32668 = (inp[2]) ? node32678 : node32669;
													assign node32669 = (inp[14]) ? node32675 : node32670;
														assign node32670 = (inp[10]) ? 16'b0000000000011111 : node32671;
															assign node32671 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32675 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32678 = (inp[14]) ? 16'b0000000000001111 : node32679;
														assign node32679 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000001111;
									assign node32683 = (inp[2]) ? node32761 : node32684;
										assign node32684 = (inp[6]) ? node32722 : node32685;
											assign node32685 = (inp[10]) ? node32701 : node32686;
												assign node32686 = (inp[1]) ? node32692 : node32687;
													assign node32687 = (inp[14]) ? 16'b0000000000111111 : node32688;
														assign node32688 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32692 = (inp[9]) ? node32696 : node32693;
														assign node32693 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32696 = (inp[8]) ? node32698 : 16'b0000000000111111;
															assign node32698 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32701 = (inp[12]) ? node32711 : node32702;
													assign node32702 = (inp[14]) ? node32706 : node32703;
														assign node32703 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node32706 = (inp[9]) ? node32708 : 16'b0000000000111111;
															assign node32708 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32711 = (inp[1]) ? node32715 : node32712;
														assign node32712 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32715 = (inp[8]) ? 16'b0000000000001111 : node32716;
															assign node32716 = (inp[9]) ? node32718 : 16'b0000000000011111;
																assign node32718 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node32722 = (inp[14]) ? node32744 : node32723;
												assign node32723 = (inp[12]) ? node32739 : node32724;
													assign node32724 = (inp[1]) ? node32734 : node32725;
														assign node32725 = (inp[10]) ? node32731 : node32726;
															assign node32726 = (inp[9]) ? node32728 : 16'b0000000001111111;
																assign node32728 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
															assign node32731 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32734 = (inp[8]) ? node32736 : 16'b0000000000111111;
															assign node32736 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32739 = (inp[10]) ? 16'b0000000000011111 : node32740;
														assign node32740 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32744 = (inp[9]) ? node32752 : node32745;
													assign node32745 = (inp[1]) ? 16'b0000000000000111 : node32746;
														assign node32746 = (inp[10]) ? 16'b0000000000011111 : node32747;
															assign node32747 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32752 = (inp[8]) ? node32754 : 16'b0000000000001111;
														assign node32754 = (inp[12]) ? node32756 : 16'b0000000000001111;
															assign node32756 = (inp[1]) ? node32758 : 16'b0000000000000111;
																assign node32758 = (inp[10]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node32761 = (inp[8]) ? node32785 : node32762;
											assign node32762 = (inp[6]) ? node32776 : node32763;
												assign node32763 = (inp[9]) ? node32769 : node32764;
													assign node32764 = (inp[14]) ? node32766 : 16'b0000000001111111;
														assign node32766 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32769 = (inp[12]) ? node32773 : node32770;
														assign node32770 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32773 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32776 = (inp[1]) ? node32782 : node32777;
													assign node32777 = (inp[9]) ? 16'b0000000000001111 : node32778;
														assign node32778 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32782 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node32785 = (inp[14]) ? node32811 : node32786;
												assign node32786 = (inp[12]) ? node32800 : node32787;
													assign node32787 = (inp[10]) ? node32793 : node32788;
														assign node32788 = (inp[6]) ? 16'b0000000000011111 : node32789;
															assign node32789 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32793 = (inp[1]) ? node32795 : 16'b0000000000011111;
															assign node32795 = (inp[6]) ? 16'b0000000000001111 : node32796;
																assign node32796 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32800 = (inp[1]) ? node32804 : node32801;
														assign node32801 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node32804 = (inp[6]) ? node32806 : 16'b0000000000001111;
															assign node32806 = (inp[10]) ? node32808 : 16'b0000000000000111;
																assign node32808 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
												assign node32811 = (inp[10]) ? node32817 : node32812;
													assign node32812 = (inp[9]) ? node32814 : 16'b0000000000001111;
														assign node32814 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node32817 = (inp[9]) ? node32819 : 16'b0000000000000111;
														assign node32819 = (inp[6]) ? node32821 : 16'b0000000000000111;
															assign node32821 = (inp[1]) ? node32823 : 16'b0000000000000111;
																assign node32823 = (inp[12]) ? 16'b0000000000000001 : 16'b0000000000000011;
							assign node32826 = (inp[14]) ? node33074 : node32827;
								assign node32827 = (inp[4]) ? node32939 : node32828;
									assign node32828 = (inp[2]) ? node32876 : node32829;
										assign node32829 = (inp[10]) ? node32867 : node32830;
											assign node32830 = (inp[15]) ? node32848 : node32831;
												assign node32831 = (inp[6]) ? node32839 : node32832;
													assign node32832 = (inp[9]) ? node32834 : 16'b0000000111111111;
														assign node32834 = (inp[1]) ? 16'b0000000001111111 : node32835;
															assign node32835 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32839 = (inp[8]) ? node32843 : node32840;
														assign node32840 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32843 = (inp[12]) ? 16'b0000000000111111 : node32844;
															assign node32844 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32848 = (inp[9]) ? node32858 : node32849;
													assign node32849 = (inp[12]) ? node32851 : 16'b0000000001111111;
														assign node32851 = (inp[6]) ? 16'b0000000000111111 : node32852;
															assign node32852 = (inp[8]) ? node32854 : 16'b0000000001111111;
																assign node32854 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32858 = (inp[1]) ? node32864 : node32859;
														assign node32859 = (inp[12]) ? 16'b0000000000111111 : node32860;
															assign node32860 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32864 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node32867 = (inp[15]) ? node32871 : node32868;
												assign node32868 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node32871 = (inp[9]) ? node32873 : 16'b0000000000111111;
													assign node32873 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node32876 = (inp[8]) ? node32904 : node32877;
											assign node32877 = (inp[1]) ? node32891 : node32878;
												assign node32878 = (inp[12]) ? node32886 : node32879;
													assign node32879 = (inp[15]) ? node32881 : 16'b0000000011111111;
														assign node32881 = (inp[10]) ? 16'b0000000001111111 : node32882;
															assign node32882 = (inp[6]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node32886 = (inp[9]) ? node32888 : 16'b0000000001111111;
														assign node32888 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node32891 = (inp[9]) ? node32899 : node32892;
													assign node32892 = (inp[10]) ? node32896 : node32893;
														assign node32893 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32896 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32899 = (inp[12]) ? node32901 : 16'b0000000000011111;
														assign node32901 = (inp[6]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node32904 = (inp[10]) ? node32922 : node32905;
												assign node32905 = (inp[1]) ? node32913 : node32906;
													assign node32906 = (inp[9]) ? node32910 : node32907;
														assign node32907 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32910 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32913 = (inp[6]) ? node32919 : node32914;
														assign node32914 = (inp[15]) ? 16'b0000000000011111 : node32915;
															assign node32915 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32919 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node32922 = (inp[12]) ? node32930 : node32923;
													assign node32923 = (inp[6]) ? node32927 : node32924;
														assign node32924 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node32927 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node32930 = (inp[15]) ? node32936 : node32931;
														assign node32931 = (inp[9]) ? node32933 : 16'b0000000000011111;
															assign node32933 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node32936 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node32939 = (inp[1]) ? node33017 : node32940;
										assign node32940 = (inp[9]) ? node32978 : node32941;
											assign node32941 = (inp[10]) ? node32961 : node32942;
												assign node32942 = (inp[8]) ? node32952 : node32943;
													assign node32943 = (inp[12]) ? node32947 : node32944;
														assign node32944 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node32947 = (inp[6]) ? node32949 : 16'b0000000001111111;
															assign node32949 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32952 = (inp[12]) ? node32958 : node32953;
														assign node32953 = (inp[6]) ? node32955 : 16'b0000000001111111;
															assign node32955 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32958 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32961 = (inp[6]) ? node32975 : node32962;
													assign node32962 = (inp[8]) ? node32968 : node32963;
														assign node32963 = (inp[2]) ? 16'b0000000000111111 : node32964;
															assign node32964 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node32968 = (inp[2]) ? 16'b0000000000011111 : node32969;
															assign node32969 = (inp[12]) ? 16'b0000000000011111 : node32970;
																assign node32970 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node32975 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node32978 = (inp[8]) ? node32994 : node32979;
												assign node32979 = (inp[15]) ? node32985 : node32980;
													assign node32980 = (inp[12]) ? node32982 : 16'b0000000000111111;
														assign node32982 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node32985 = (inp[6]) ? 16'b0000000000011111 : node32986;
														assign node32986 = (inp[2]) ? node32988 : 16'b0000000000111111;
															assign node32988 = (inp[10]) ? 16'b0000000000011111 : node32989;
																assign node32989 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node32994 = (inp[6]) ? node33006 : node32995;
													assign node32995 = (inp[2]) ? node33003 : node32996;
														assign node32996 = (inp[15]) ? node32998 : 16'b0000000000111111;
															assign node32998 = (inp[12]) ? 16'b0000000000011111 : node32999;
																assign node32999 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node33003 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node33006 = (inp[12]) ? node33010 : node33007;
														assign node33007 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33010 = (inp[10]) ? 16'b0000000000000111 : node33011;
															assign node33011 = (inp[15]) ? node33013 : 16'b0000000000001111;
																assign node33013 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node33017 = (inp[9]) ? node33051 : node33018;
											assign node33018 = (inp[2]) ? node33030 : node33019;
												assign node33019 = (inp[6]) ? node33025 : node33020;
													assign node33020 = (inp[12]) ? node33022 : 16'b0000000000111111;
														assign node33022 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node33025 = (inp[8]) ? node33027 : 16'b0000000000011111;
														assign node33027 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node33030 = (inp[10]) ? node33044 : node33031;
													assign node33031 = (inp[8]) ? node33035 : node33032;
														assign node33032 = (inp[6]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node33035 = (inp[6]) ? node33039 : node33036;
															assign node33036 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
															assign node33039 = (inp[12]) ? node33041 : 16'b0000000000001111;
																assign node33041 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node33044 = (inp[6]) ? node33046 : 16'b0000000000001111;
														assign node33046 = (inp[8]) ? 16'b0000000000000111 : node33047;
															assign node33047 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node33051 = (inp[15]) ? node33061 : node33052;
												assign node33052 = (inp[8]) ? node33054 : 16'b0000000000011111;
													assign node33054 = (inp[6]) ? node33058 : node33055;
														assign node33055 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33058 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node33061 = (inp[10]) ? node33069 : node33062;
													assign node33062 = (inp[2]) ? 16'b0000000000000111 : node33063;
														assign node33063 = (inp[8]) ? node33065 : 16'b0000000000001111;
															assign node33065 = (inp[6]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node33069 = (inp[6]) ? node33071 : 16'b0000000000000011;
														assign node33071 = (inp[12]) ? 16'b0000000000000001 : 16'b0000000000000011;
								assign node33074 = (inp[8]) ? node33196 : node33075;
									assign node33075 = (inp[9]) ? node33151 : node33076;
										assign node33076 = (inp[10]) ? node33106 : node33077;
											assign node33077 = (inp[12]) ? node33093 : node33078;
												assign node33078 = (inp[4]) ? node33088 : node33079;
													assign node33079 = (inp[15]) ? node33083 : node33080;
														assign node33080 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node33083 = (inp[2]) ? 16'b0000000000111111 : node33084;
															assign node33084 = (inp[6]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node33088 = (inp[15]) ? node33090 : 16'b0000000000111111;
														assign node33090 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node33093 = (inp[6]) ? node33097 : node33094;
													assign node33094 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node33097 = (inp[4]) ? node33103 : node33098;
														assign node33098 = (inp[15]) ? 16'b0000000000011111 : node33099;
															assign node33099 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node33103 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node33106 = (inp[6]) ? node33124 : node33107;
												assign node33107 = (inp[1]) ? node33113 : node33108;
													assign node33108 = (inp[15]) ? node33110 : 16'b0000000001111111;
														assign node33110 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node33113 = (inp[15]) ? node33119 : node33114;
														assign node33114 = (inp[4]) ? node33116 : 16'b0000000000111111;
															assign node33116 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node33119 = (inp[12]) ? node33121 : 16'b0000000000011111;
															assign node33121 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node33124 = (inp[1]) ? node33136 : node33125;
													assign node33125 = (inp[4]) ? node33129 : node33126;
														assign node33126 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node33129 = (inp[2]) ? node33131 : 16'b0000000000011111;
															assign node33131 = (inp[12]) ? 16'b0000000000001111 : node33132;
																assign node33132 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node33136 = (inp[12]) ? node33144 : node33137;
														assign node33137 = (inp[4]) ? node33139 : 16'b0000000000011111;
															assign node33139 = (inp[15]) ? 16'b0000000000001111 : node33140;
																assign node33140 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33144 = (inp[2]) ? node33148 : node33145;
															assign node33145 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
															assign node33148 = (inp[4]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node33151 = (inp[1]) ? node33181 : node33152;
											assign node33152 = (inp[6]) ? node33170 : node33153;
												assign node33153 = (inp[4]) ? node33157 : node33154;
													assign node33154 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node33157 = (inp[10]) ? node33163 : node33158;
														assign node33158 = (inp[15]) ? 16'b0000000000011111 : node33159;
															assign node33159 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node33163 = (inp[2]) ? node33165 : 16'b0000000000011111;
															assign node33165 = (inp[15]) ? 16'b0000000000001111 : node33166;
																assign node33166 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node33170 = (inp[4]) ? node33176 : node33171;
													assign node33171 = (inp[15]) ? node33173 : 16'b0000000000011111;
														assign node33173 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node33176 = (inp[10]) ? 16'b0000000000001111 : node33177;
														assign node33177 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node33181 = (inp[15]) ? node33191 : node33182;
												assign node33182 = (inp[2]) ? node33188 : node33183;
													assign node33183 = (inp[12]) ? node33185 : 16'b0000000000011111;
														assign node33185 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node33188 = (inp[6]) ? 16'b0000000000000011 : 16'b0000000000001111;
												assign node33191 = (inp[4]) ? node33193 : 16'b0000000000001111;
													assign node33193 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node33196 = (inp[1]) ? node33250 : node33197;
										assign node33197 = (inp[6]) ? node33217 : node33198;
											assign node33198 = (inp[9]) ? node33206 : node33199;
												assign node33199 = (inp[2]) ? 16'b0000000000011111 : node33200;
													assign node33200 = (inp[15]) ? node33202 : 16'b0000000000111111;
														assign node33202 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node33206 = (inp[4]) ? node33208 : 16'b0000000000011111;
													assign node33208 = (inp[15]) ? node33214 : node33209;
														assign node33209 = (inp[12]) ? node33211 : 16'b0000000000011111;
															assign node33211 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33214 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node33217 = (inp[15]) ? node33235 : node33218;
												assign node33218 = (inp[9]) ? node33224 : node33219;
													assign node33219 = (inp[2]) ? node33221 : 16'b0000000000011111;
														assign node33221 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node33224 = (inp[4]) ? node33230 : node33225;
														assign node33225 = (inp[12]) ? 16'b0000000000001111 : node33226;
															assign node33226 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33230 = (inp[10]) ? node33232 : 16'b0000000000001111;
															assign node33232 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node33235 = (inp[9]) ? node33243 : node33236;
													assign node33236 = (inp[2]) ? node33240 : node33237;
														assign node33237 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33240 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node33243 = (inp[10]) ? node33245 : 16'b0000000000000111;
														assign node33245 = (inp[12]) ? node33247 : 16'b0000000000000111;
															assign node33247 = (inp[4]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node33250 = (inp[10]) ? node33278 : node33251;
											assign node33251 = (inp[15]) ? node33259 : node33252;
												assign node33252 = (inp[4]) ? 16'b0000000000000111 : node33253;
													assign node33253 = (inp[6]) ? node33255 : 16'b0000000000011111;
														assign node33255 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node33259 = (inp[12]) ? node33269 : node33260;
													assign node33260 = (inp[2]) ? node33264 : node33261;
														assign node33261 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node33264 = (inp[4]) ? node33266 : 16'b0000000000001111;
															assign node33266 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node33269 = (inp[9]) ? node33273 : node33270;
														assign node33270 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node33273 = (inp[4]) ? node33275 : 16'b0000000000000111;
															assign node33275 = (inp[2]) ? 16'b0000000000000011 : 16'b0000000000000111;
											assign node33278 = (inp[6]) ? node33290 : node33279;
												assign node33279 = (inp[12]) ? node33285 : node33280;
													assign node33280 = (inp[15]) ? node33282 : 16'b0000000000011111;
														assign node33282 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node33285 = (inp[2]) ? 16'b0000000000000111 : node33286;
														assign node33286 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node33290 = (inp[4]) ? node33304 : node33291;
													assign node33291 = (inp[12]) ? node33297 : node33292;
														assign node33292 = (inp[15]) ? node33294 : 16'b0000000000001111;
															assign node33294 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000001111;
														assign node33297 = (inp[9]) ? 16'b0000000000000011 : node33298;
															assign node33298 = (inp[2]) ? node33300 : 16'b0000000000000111;
																assign node33300 = (inp[15]) ? 16'b0000000000000011 : 16'b0000000000000111;
													assign node33304 = (inp[2]) ? node33316 : node33305;
														assign node33305 = (inp[12]) ? node33311 : node33306;
															assign node33306 = (inp[15]) ? node33308 : 16'b0000000000000111;
																assign node33308 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
															assign node33311 = (inp[15]) ? 16'b0000000000000011 : node33312;
																assign node33312 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
														assign node33316 = (inp[15]) ? 16'b0000000000000001 : 16'b0000000000000011;

endmodule