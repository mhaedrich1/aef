module dtc_split25_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;

	assign outp = (inp[9]) ? node172 : node1;
		assign node1 = (inp[6]) ? node105 : node2;
			assign node2 = (inp[10]) ? node42 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[3]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[8]) ? 3'b011 : 3'b111;
					assign node11 = (inp[8]) ? node29 : node12;
						assign node12 = (inp[11]) ? node18 : node13;
							assign node13 = (inp[4]) ? node15 : 3'b111;
								assign node15 = (inp[3]) ? 3'b011 : 3'b111;
							assign node18 = (inp[3]) ? node24 : node19;
								assign node19 = (inp[4]) ? 3'b011 : node20;
									assign node20 = (inp[2]) ? 3'b011 : 3'b111;
								assign node24 = (inp[5]) ? 3'b101 : node25;
									assign node25 = (inp[0]) ? 3'b111 : 3'b011;
						assign node29 = (inp[11]) ? node35 : node30;
							assign node30 = (inp[3]) ? 3'b011 : node31;
								assign node31 = (inp[1]) ? 3'b011 : 3'b111;
							assign node35 = (inp[3]) ? 3'b101 : node36;
								assign node36 = (inp[1]) ? node38 : 3'b011;
									assign node38 = (inp[2]) ? 3'b011 : 3'b001;
				assign node42 = (inp[11]) ? node84 : node43;
					assign node43 = (inp[8]) ? node59 : node44;
						assign node44 = (inp[3]) ? node54 : node45;
							assign node45 = (inp[4]) ? node51 : node46;
								assign node46 = (inp[2]) ? 3'b111 : node47;
									assign node47 = (inp[7]) ? 3'b011 : 3'b111;
								assign node51 = (inp[7]) ? 3'b101 : 3'b111;
							assign node54 = (inp[7]) ? node56 : 3'b011;
								assign node56 = (inp[4]) ? 3'b001 : 3'b111;
						assign node59 = (inp[3]) ? node69 : node60;
							assign node60 = (inp[7]) ? node62 : 3'b011;
								assign node62 = (inp[2]) ? node64 : 3'b101;
									assign node64 = (inp[4]) ? node66 : 3'b001;
										assign node66 = (inp[1]) ? 3'b010 : 3'b001;
							assign node69 = (inp[1]) ? node71 : 3'b001;
								assign node71 = (inp[5]) ? node77 : node72;
									assign node72 = (inp[0]) ? 3'b001 : node73;
										assign node73 = (inp[7]) ? 3'b001 : 3'b101;
									assign node77 = (inp[0]) ? node81 : node78;
										assign node78 = (inp[4]) ? 3'b101 : 3'b001;
										assign node81 = (inp[7]) ? 3'b110 : 3'b101;
					assign node84 = (inp[7]) ? node94 : node85;
						assign node85 = (inp[3]) ? node89 : node86;
							assign node86 = (inp[8]) ? 3'b101 : 3'b011;
							assign node89 = (inp[8]) ? node91 : 3'b101;
								assign node91 = (inp[4]) ? 3'b001 : 3'b101;
						assign node94 = (inp[8]) ? node96 : 3'b101;
							assign node96 = (inp[3]) ? node102 : node97;
								assign node97 = (inp[1]) ? node99 : 3'b101;
									assign node99 = (inp[2]) ? 3'b101 : 3'b110;
								assign node102 = (inp[0]) ? 3'b010 : 3'b110;
			assign node105 = (inp[10]) ? node161 : node106;
				assign node106 = (inp[7]) ? node126 : node107;
					assign node107 = (inp[8]) ? node115 : node108;
						assign node108 = (inp[11]) ? 3'b001 : node109;
							assign node109 = (inp[4]) ? node111 : 3'b011;
								assign node111 = (inp[3]) ? 3'b101 : 3'b011;
						assign node115 = (inp[11]) ? 3'b110 : node116;
							assign node116 = (inp[5]) ? node120 : node117;
								assign node117 = (inp[4]) ? 3'b001 : 3'b011;
								assign node120 = (inp[2]) ? 3'b001 : node121;
									assign node121 = (inp[1]) ? 3'b001 : 3'b101;
					assign node126 = (inp[11]) ? node146 : node127;
						assign node127 = (inp[8]) ? node137 : node128;
							assign node128 = (inp[3]) ? node134 : node129;
								assign node129 = (inp[4]) ? 3'b001 : node130;
									assign node130 = (inp[2]) ? 3'b001 : 3'b101;
								assign node134 = (inp[4]) ? 3'b110 : 3'b001;
							assign node137 = (inp[4]) ? node141 : node138;
								assign node138 = (inp[3]) ? 3'b110 : 3'b001;
								assign node141 = (inp[1]) ? node143 : 3'b110;
									assign node143 = (inp[2]) ? 3'b110 : 3'b010;
						assign node146 = (inp[8]) ? node152 : node147;
							assign node147 = (inp[4]) ? node149 : 3'b110;
								assign node149 = (inp[3]) ? 3'b010 : 3'b110;
							assign node152 = (inp[1]) ? node154 : 3'b010;
								assign node154 = (inp[2]) ? node156 : 3'b010;
									assign node156 = (inp[0]) ? node158 : 3'b010;
										assign node158 = (inp[4]) ? 3'b100 : 3'b010;
				assign node161 = (inp[7]) ? node169 : node162;
					assign node162 = (inp[11]) ? node166 : node163;
						assign node163 = (inp[8]) ? 3'b010 : 3'b110;
						assign node166 = (inp[8]) ? 3'b100 : 3'b010;
					assign node169 = (inp[11]) ? 3'b000 : 3'b100;
		assign node172 = (inp[6]) ? node226 : node173;
			assign node173 = (inp[10]) ? node211 : node174;
				assign node174 = (inp[8]) ? node194 : node175;
					assign node175 = (inp[7]) ? node191 : node176;
						assign node176 = (inp[4]) ? node186 : node177;
							assign node177 = (inp[11]) ? 3'b001 : node178;
								assign node178 = (inp[3]) ? node180 : 3'b101;
									assign node180 = (inp[0]) ? node182 : 3'b101;
										assign node182 = (inp[5]) ? 3'b001 : 3'b101;
							assign node186 = (inp[11]) ? node188 : 3'b101;
								assign node188 = (inp[3]) ? 3'b110 : 3'b101;
						assign node191 = (inp[11]) ? 3'b100 : 3'b010;
					assign node194 = (inp[7]) ? node202 : node195;
						assign node195 = (inp[11]) ? node197 : 3'b000;
							assign node197 = (inp[4]) ? node199 : 3'b010;
								assign node199 = (inp[0]) ? 3'b101 : 3'b010;
						assign node202 = (inp[11]) ? node208 : node203;
							assign node203 = (inp[3]) ? node205 : 3'b010;
								assign node205 = (inp[2]) ? 3'b100 : 3'b010;
							assign node208 = (inp[4]) ? 3'b000 : 3'b100;
				assign node211 = (inp[7]) ? 3'b000 : node212;
					assign node212 = (inp[8]) ? node222 : node213;
						assign node213 = (inp[11]) ? node215 : 3'b010;
							assign node215 = (inp[0]) ? node217 : 3'b100;
								assign node217 = (inp[4]) ? node219 : 3'b100;
									assign node219 = (inp[1]) ? 3'b100 : 3'b000;
						assign node222 = (inp[11]) ? 3'b000 : 3'b100;
			assign node226 = (inp[7]) ? 3'b000 : node227;
				assign node227 = (inp[11]) ? 3'b000 : node228;
					assign node228 = (inp[10]) ? 3'b000 : node229;
						assign node229 = (inp[8]) ? 3'b000 : 3'b100;

endmodule