module dtc_split75_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node642;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node692;
	wire [3-1:0] node696;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node738;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node764;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node814;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node878;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node968;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1012;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1048;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1056;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1063;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1077;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1107;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1115;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1158;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1167;
	wire [3-1:0] node1171;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1179;
	wire [3-1:0] node1183;
	wire [3-1:0] node1185;
	wire [3-1:0] node1187;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1202;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1221;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;

	assign outp = (inp[6]) ? node384 : node1;
		assign node1 = (inp[9]) ? node343 : node2;
			assign node2 = (inp[0]) ? node256 : node3;
				assign node3 = (inp[7]) ? node109 : node4;
					assign node4 = (inp[10]) ? node84 : node5;
						assign node5 = (inp[1]) ? node55 : node6;
							assign node6 = (inp[8]) ? node34 : node7;
								assign node7 = (inp[11]) ? node19 : node8;
									assign node8 = (inp[3]) ? node16 : node9;
										assign node9 = (inp[2]) ? 3'b010 : node10;
											assign node10 = (inp[4]) ? 3'b010 : node11;
												assign node11 = (inp[5]) ? 3'b010 : 3'b110;
										assign node16 = (inp[2]) ? 3'b100 : 3'b010;
									assign node19 = (inp[4]) ? node29 : node20;
										assign node20 = (inp[5]) ? node26 : node21;
											assign node21 = (inp[2]) ? 3'b100 : node22;
												assign node22 = (inp[3]) ? 3'b100 : 3'b010;
											assign node26 = (inp[3]) ? 3'b000 : 3'b100;
										assign node29 = (inp[3]) ? node31 : 3'b100;
											assign node31 = (inp[2]) ? 3'b000 : 3'b100;
								assign node34 = (inp[11]) ? node44 : node35;
									assign node35 = (inp[2]) ? node41 : node36;
										assign node36 = (inp[4]) ? 3'b110 : node37;
											assign node37 = (inp[3]) ? 3'b110 : 3'b001;
										assign node41 = (inp[4]) ? 3'b010 : 3'b110;
									assign node44 = (inp[2]) ? node50 : node45;
										assign node45 = (inp[4]) ? 3'b010 : node46;
											assign node46 = (inp[3]) ? 3'b010 : 3'b110;
										assign node50 = (inp[4]) ? node52 : 3'b010;
											assign node52 = (inp[3]) ? 3'b100 : 3'b010;
							assign node55 = (inp[2]) ? node63 : node56;
								assign node56 = (inp[8]) ? node60 : node57;
									assign node57 = (inp[11]) ? 3'b000 : 3'b100;
									assign node60 = (inp[11]) ? 3'b100 : 3'b010;
								assign node63 = (inp[8]) ? node71 : node64;
									assign node64 = (inp[3]) ? 3'b000 : node65;
										assign node65 = (inp[4]) ? 3'b000 : node66;
											assign node66 = (inp[11]) ? 3'b000 : 3'b100;
									assign node71 = (inp[11]) ? node79 : node72;
										assign node72 = (inp[3]) ? 3'b100 : node73;
											assign node73 = (inp[4]) ? node75 : 3'b010;
												assign node75 = (inp[5]) ? 3'b100 : 3'b010;
										assign node79 = (inp[3]) ? 3'b000 : node80;
											assign node80 = (inp[5]) ? 3'b000 : 3'b100;
						assign node84 = (inp[1]) ? 3'b000 : node85;
							assign node85 = (inp[8]) ? node87 : 3'b000;
								assign node87 = (inp[11]) ? node99 : node88;
									assign node88 = (inp[4]) ? node94 : node89;
										assign node89 = (inp[3]) ? 3'b100 : node90;
											assign node90 = (inp[2]) ? 3'b100 : 3'b010;
										assign node94 = (inp[3]) ? node96 : 3'b100;
											assign node96 = (inp[5]) ? 3'b100 : 3'b000;
									assign node99 = (inp[3]) ? 3'b000 : node100;
										assign node100 = (inp[2]) ? 3'b000 : node101;
											assign node101 = (inp[4]) ? node103 : 3'b100;
												assign node103 = (inp[5]) ? 3'b000 : 3'b100;
					assign node109 = (inp[10]) ? node189 : node110;
						assign node110 = (inp[1]) ? node152 : node111;
							assign node111 = (inp[8]) ? node133 : node112;
								assign node112 = (inp[11]) ? node122 : node113;
									assign node113 = (inp[2]) ? node117 : node114;
										assign node114 = (inp[3]) ? 3'b001 : 3'b101;
										assign node117 = (inp[3]) ? node119 : 3'b001;
											assign node119 = (inp[4]) ? 3'b110 : 3'b001;
									assign node122 = (inp[4]) ? node124 : 3'b110;
										assign node124 = (inp[3]) ? node130 : node125;
											assign node125 = (inp[5]) ? 3'b110 : node126;
												assign node126 = (inp[2]) ? 3'b110 : 3'b001;
											assign node130 = (inp[2]) ? 3'b010 : 3'b110;
								assign node133 = (inp[11]) ? node147 : node134;
									assign node134 = (inp[2]) ? node142 : node135;
										assign node135 = (inp[3]) ? 3'b101 : node136;
											assign node136 = (inp[4]) ? node138 : 3'b011;
												assign node138 = (inp[5]) ? 3'b101 : 3'b011;
										assign node142 = (inp[3]) ? node144 : 3'b101;
											assign node144 = (inp[5]) ? 3'b001 : 3'b101;
									assign node147 = (inp[3]) ? 3'b001 : node148;
										assign node148 = (inp[2]) ? 3'b001 : 3'b101;
							assign node152 = (inp[8]) ? node166 : node153;
								assign node153 = (inp[11]) ? node161 : node154;
									assign node154 = (inp[2]) ? node156 : 3'b110;
										assign node156 = (inp[3]) ? 3'b010 : node157;
											assign node157 = (inp[5]) ? 3'b010 : 3'b110;
									assign node161 = (inp[2]) ? node163 : 3'b010;
										assign node163 = (inp[3]) ? 3'b100 : 3'b010;
								assign node166 = (inp[11]) ? node178 : node167;
									assign node167 = (inp[2]) ? node175 : node168;
										assign node168 = (inp[4]) ? 3'b001 : node169;
											assign node169 = (inp[3]) ? 3'b001 : node170;
												assign node170 = (inp[5]) ? 3'b001 : 3'b101;
										assign node175 = (inp[3]) ? 3'b110 : 3'b001;
									assign node178 = (inp[5]) ? node184 : node179;
										assign node179 = (inp[4]) ? 3'b110 : node180;
											assign node180 = (inp[2]) ? 3'b110 : 3'b001;
										assign node184 = (inp[2]) ? node186 : 3'b110;
											assign node186 = (inp[3]) ? 3'b010 : 3'b110;
						assign node189 = (inp[1]) ? node223 : node190;
							assign node190 = (inp[8]) ? node212 : node191;
								assign node191 = (inp[11]) ? node201 : node192;
									assign node192 = (inp[3]) ? node196 : node193;
										assign node193 = (inp[2]) ? 3'b010 : 3'b110;
										assign node196 = (inp[4]) ? node198 : 3'b010;
											assign node198 = (inp[2]) ? 3'b100 : 3'b010;
									assign node201 = (inp[4]) ? node203 : 3'b100;
										assign node203 = (inp[2]) ? node207 : node204;
											assign node204 = (inp[3]) ? 3'b100 : 3'b010;
											assign node207 = (inp[3]) ? node209 : 3'b100;
												assign node209 = (inp[5]) ? 3'b000 : 3'b100;
								assign node212 = (inp[11]) ? node218 : node213;
									assign node213 = (inp[3]) ? 3'b110 : node214;
										assign node214 = (inp[2]) ? 3'b110 : 3'b001;
									assign node218 = (inp[3]) ? 3'b010 : node219;
										assign node219 = (inp[2]) ? 3'b010 : 3'b110;
							assign node223 = (inp[8]) ? node239 : node224;
								assign node224 = (inp[11]) ? node230 : node225;
									assign node225 = (inp[2]) ? node227 : 3'b100;
										assign node227 = (inp[3]) ? 3'b000 : 3'b100;
									assign node230 = (inp[3]) ? 3'b000 : node231;
										assign node231 = (inp[5]) ? 3'b000 : node232;
											assign node232 = (inp[4]) ? 3'b000 : node233;
												assign node233 = (inp[2]) ? 3'b000 : 3'b100;
								assign node239 = (inp[11]) ? node249 : node240;
									assign node240 = (inp[2]) ? node242 : 3'b010;
										assign node242 = (inp[3]) ? node244 : 3'b010;
											assign node244 = (inp[4]) ? 3'b100 : node245;
												assign node245 = (inp[5]) ? 3'b100 : 3'b010;
									assign node249 = (inp[3]) ? node251 : 3'b100;
										assign node251 = (inp[5]) ? node253 : 3'b100;
											assign node253 = (inp[2]) ? 3'b000 : 3'b100;
				assign node256 = (inp[7]) ? node272 : node257;
					assign node257 = (inp[2]) ? 3'b000 : node258;
						assign node258 = (inp[8]) ? node260 : 3'b000;
							assign node260 = (inp[1]) ? 3'b000 : node261;
								assign node261 = (inp[10]) ? 3'b000 : node262;
									assign node262 = (inp[11]) ? 3'b000 : node263;
										assign node263 = (inp[4]) ? node265 : 3'b100;
											assign node265 = (inp[3]) ? 3'b000 : 3'b100;
					assign node272 = (inp[10]) ? node330 : node273;
						assign node273 = (inp[1]) ? node309 : node274;
							assign node274 = (inp[8]) ? node294 : node275;
								assign node275 = (inp[11]) ? node285 : node276;
									assign node276 = (inp[2]) ? 3'b100 : node277;
										assign node277 = (inp[3]) ? node279 : 3'b010;
											assign node279 = (inp[5]) ? node281 : 3'b010;
												assign node281 = (inp[4]) ? 3'b100 : 3'b010;
									assign node285 = (inp[2]) ? node287 : 3'b100;
										assign node287 = (inp[5]) ? 3'b000 : node288;
											assign node288 = (inp[4]) ? 3'b000 : node289;
												assign node289 = (inp[3]) ? 3'b000 : 3'b100;
								assign node294 = (inp[11]) ? node302 : node295;
									assign node295 = (inp[2]) ? node297 : 3'b110;
										assign node297 = (inp[4]) ? 3'b010 : node298;
											assign node298 = (inp[3]) ? 3'b010 : 3'b110;
									assign node302 = (inp[2]) ? node304 : 3'b010;
										assign node304 = (inp[3]) ? 3'b100 : node305;
											assign node305 = (inp[4]) ? 3'b100 : 3'b010;
							assign node309 = (inp[8]) ? node317 : node310;
								assign node310 = (inp[11]) ? 3'b000 : node311;
									assign node311 = (inp[2]) ? 3'b000 : node312;
										assign node312 = (inp[3]) ? 3'b000 : 3'b100;
								assign node317 = (inp[11]) ? node325 : node318;
									assign node318 = (inp[2]) ? 3'b100 : node319;
										assign node319 = (inp[3]) ? node321 : 3'b010;
											assign node321 = (inp[5]) ? 3'b100 : 3'b010;
									assign node325 = (inp[2]) ? 3'b000 : node326;
										assign node326 = (inp[4]) ? 3'b000 : 3'b100;
						assign node330 = (inp[11]) ? 3'b000 : node331;
							assign node331 = (inp[8]) ? node333 : 3'b000;
								assign node333 = (inp[1]) ? 3'b000 : node334;
									assign node334 = (inp[2]) ? node336 : 3'b100;
										assign node336 = (inp[4]) ? 3'b000 : node337;
											assign node337 = (inp[3]) ? 3'b000 : 3'b100;
			assign node343 = (inp[0]) ? 3'b000 : node344;
				assign node344 = (inp[10]) ? 3'b000 : node345;
					assign node345 = (inp[7]) ? node347 : 3'b000;
						assign node347 = (inp[1]) ? node371 : node348;
							assign node348 = (inp[8]) ? node356 : node349;
								assign node349 = (inp[3]) ? 3'b000 : node350;
									assign node350 = (inp[2]) ? 3'b000 : node351;
										assign node351 = (inp[11]) ? 3'b000 : 3'b100;
								assign node356 = (inp[11]) ? node364 : node357;
									assign node357 = (inp[2]) ? 3'b100 : node358;
										assign node358 = (inp[3]) ? node360 : 3'b010;
											assign node360 = (inp[4]) ? 3'b100 : 3'b010;
									assign node364 = (inp[2]) ? 3'b000 : node365;
										assign node365 = (inp[3]) ? node367 : 3'b100;
											assign node367 = (inp[4]) ? 3'b000 : 3'b100;
							assign node371 = (inp[11]) ? 3'b000 : node372;
								assign node372 = (inp[3]) ? 3'b000 : node373;
									assign node373 = (inp[4]) ? 3'b000 : node374;
										assign node374 = (inp[2]) ? 3'b000 : node375;
											assign node375 = (inp[8]) ? 3'b100 : 3'b000;
		assign node384 = (inp[9]) ? node896 : node385;
			assign node385 = (inp[0]) ? node611 : node386;
				assign node386 = (inp[7]) ? node538 : node387;
					assign node387 = (inp[10]) ? node453 : node388;
						assign node388 = (inp[1]) ? node416 : node389;
							assign node389 = (inp[11]) ? node397 : node390;
								assign node390 = (inp[8]) ? 3'b111 : node391;
									assign node391 = (inp[3]) ? 3'b011 : node392;
										assign node392 = (inp[2]) ? 3'b011 : 3'b111;
								assign node397 = (inp[8]) ? node407 : node398;
									assign node398 = (inp[2]) ? 3'b101 : node399;
										assign node399 = (inp[3]) ? node401 : 3'b011;
											assign node401 = (inp[4]) ? 3'b101 : node402;
												assign node402 = (inp[5]) ? 3'b101 : 3'b011;
									assign node407 = (inp[2]) ? 3'b011 : node408;
										assign node408 = (inp[3]) ? node410 : 3'b111;
											assign node410 = (inp[4]) ? 3'b011 : node411;
												assign node411 = (inp[5]) ? 3'b011 : 3'b111;
							assign node416 = (inp[8]) ? node432 : node417;
								assign node417 = (inp[11]) ? node425 : node418;
									assign node418 = (inp[4]) ? node420 : 3'b101;
										assign node420 = (inp[3]) ? node422 : 3'b101;
											assign node422 = (inp[2]) ? 3'b001 : 3'b101;
									assign node425 = (inp[4]) ? node427 : 3'b001;
										assign node427 = (inp[3]) ? node429 : 3'b001;
											assign node429 = (inp[2]) ? 3'b110 : 3'b001;
								assign node432 = (inp[11]) ? node444 : node433;
									assign node433 = (inp[2]) ? node439 : node434;
										assign node434 = (inp[3]) ? 3'b011 : node435;
											assign node435 = (inp[5]) ? 3'b011 : 3'b111;
										assign node439 = (inp[4]) ? node441 : 3'b011;
											assign node441 = (inp[3]) ? 3'b101 : 3'b011;
									assign node444 = (inp[2]) ? node448 : node445;
										assign node445 = (inp[3]) ? 3'b101 : 3'b011;
										assign node448 = (inp[3]) ? node450 : 3'b101;
											assign node450 = (inp[4]) ? 3'b001 : 3'b101;
						assign node453 = (inp[1]) ? node487 : node454;
							assign node454 = (inp[8]) ? node474 : node455;
								assign node455 = (inp[11]) ? node465 : node456;
									assign node456 = (inp[2]) ? 3'b001 : node457;
										assign node457 = (inp[3]) ? node459 : 3'b101;
											assign node459 = (inp[5]) ? 3'b001 : node460;
												assign node460 = (inp[4]) ? 3'b001 : 3'b101;
									assign node465 = (inp[2]) ? 3'b110 : node466;
										assign node466 = (inp[3]) ? node468 : 3'b001;
											assign node468 = (inp[4]) ? 3'b110 : node469;
												assign node469 = (inp[5]) ? 3'b110 : 3'b001;
								assign node474 = (inp[11]) ? node480 : node475;
									assign node475 = (inp[2]) ? 3'b101 : node476;
										assign node476 = (inp[3]) ? 3'b101 : 3'b011;
									assign node480 = (inp[2]) ? 3'b001 : node481;
										assign node481 = (inp[3]) ? node483 : 3'b101;
											assign node483 = (inp[4]) ? 3'b001 : 3'b101;
							assign node487 = (inp[8]) ? node515 : node488;
								assign node488 = (inp[11]) ? node500 : node489;
									assign node489 = (inp[2]) ? node495 : node490;
										assign node490 = (inp[3]) ? 3'b110 : node491;
											assign node491 = (inp[5]) ? 3'b001 : 3'b110;
										assign node495 = (inp[3]) ? node497 : 3'b110;
											assign node497 = (inp[4]) ? 3'b010 : 3'b110;
									assign node500 = (inp[4]) ? node506 : node501;
										assign node501 = (inp[2]) ? 3'b010 : node502;
											assign node502 = (inp[3]) ? 3'b010 : 3'b110;
										assign node506 = (inp[3]) ? node512 : node507;
											assign node507 = (inp[2]) ? 3'b010 : node508;
												assign node508 = (inp[5]) ? 3'b010 : 3'b110;
											assign node512 = (inp[2]) ? 3'b100 : 3'b010;
								assign node515 = (inp[11]) ? node527 : node516;
									assign node516 = (inp[3]) ? node520 : node517;
										assign node517 = (inp[2]) ? 3'b001 : 3'b101;
										assign node520 = (inp[2]) ? node522 : 3'b001;
											assign node522 = (inp[4]) ? node524 : 3'b001;
												assign node524 = (inp[5]) ? 3'b110 : 3'b001;
									assign node527 = (inp[2]) ? node531 : node528;
										assign node528 = (inp[3]) ? 3'b110 : 3'b001;
										assign node531 = (inp[5]) ? node533 : 3'b110;
											assign node533 = (inp[4]) ? node535 : 3'b110;
												assign node535 = (inp[3]) ? 3'b010 : 3'b110;
					assign node538 = (inp[10]) ? node562 : node539;
						assign node539 = (inp[1]) ? node541 : 3'b111;
							assign node541 = (inp[8]) ? 3'b111 : node542;
								assign node542 = (inp[11]) ? node550 : node543;
									assign node543 = (inp[2]) ? node545 : 3'b111;
										assign node545 = (inp[3]) ? node547 : 3'b111;
											assign node547 = (inp[4]) ? 3'b011 : 3'b111;
									assign node550 = (inp[2]) ? node554 : node551;
										assign node551 = (inp[3]) ? 3'b011 : 3'b111;
										assign node554 = (inp[3]) ? node556 : 3'b011;
											assign node556 = (inp[5]) ? node558 : 3'b011;
												assign node558 = (inp[4]) ? 3'b101 : 3'b011;
						assign node562 = (inp[1]) ? node584 : node563;
							assign node563 = (inp[8]) ? node575 : node564;
								assign node564 = (inp[2]) ? node568 : node565;
									assign node565 = (inp[11]) ? 3'b011 : 3'b111;
									assign node568 = (inp[11]) ? node570 : 3'b011;
										assign node570 = (inp[4]) ? 3'b101 : node571;
											assign node571 = (inp[5]) ? 3'b101 : 3'b011;
								assign node575 = (inp[11]) ? node577 : 3'b111;
									assign node577 = (inp[2]) ? node579 : 3'b111;
										assign node579 = (inp[3]) ? 3'b011 : node580;
											assign node580 = (inp[4]) ? 3'b011 : 3'b111;
							assign node584 = (inp[8]) ? node596 : node585;
								assign node585 = (inp[11]) ? node591 : node586;
									assign node586 = (inp[2]) ? 3'b101 : node587;
										assign node587 = (inp[3]) ? 3'b101 : 3'b011;
									assign node591 = (inp[2]) ? 3'b001 : node592;
										assign node592 = (inp[3]) ? 3'b001 : 3'b101;
								assign node596 = (inp[11]) ? node604 : node597;
									assign node597 = (inp[2]) ? 3'b011 : node598;
										assign node598 = (inp[3]) ? node600 : 3'b111;
											assign node600 = (inp[4]) ? 3'b011 : 3'b111;
									assign node604 = (inp[2]) ? 3'b101 : node605;
										assign node605 = (inp[3]) ? node607 : 3'b011;
											assign node607 = (inp[4]) ? 3'b101 : 3'b011;
				assign node611 = (inp[7]) ? node745 : node612;
					assign node612 = (inp[10]) ? node684 : node613;
						assign node613 = (inp[1]) ? node647 : node614;
							assign node614 = (inp[8]) ? node632 : node615;
								assign node615 = (inp[11]) ? node623 : node616;
									assign node616 = (inp[2]) ? node618 : 3'b001;
										assign node618 = (inp[4]) ? 3'b110 : node619;
											assign node619 = (inp[3]) ? 3'b110 : 3'b001;
									assign node623 = (inp[2]) ? node625 : 3'b110;
										assign node625 = (inp[3]) ? 3'b010 : node626;
											assign node626 = (inp[4]) ? node628 : 3'b110;
												assign node628 = (inp[5]) ? 3'b010 : 3'b110;
								assign node632 = (inp[11]) ? node642 : node633;
									assign node633 = (inp[2]) ? node635 : 3'b101;
										assign node635 = (inp[3]) ? 3'b001 : node636;
											assign node636 = (inp[4]) ? node638 : 3'b101;
												assign node638 = (inp[5]) ? 3'b001 : 3'b101;
									assign node642 = (inp[3]) ? node644 : 3'b001;
										assign node644 = (inp[2]) ? 3'b110 : 3'b001;
							assign node647 = (inp[11]) ? node663 : node648;
								assign node648 = (inp[8]) ? node656 : node649;
									assign node649 = (inp[2]) ? 3'b010 : node650;
										assign node650 = (inp[3]) ? node652 : 3'b110;
											assign node652 = (inp[4]) ? 3'b010 : 3'b110;
									assign node656 = (inp[2]) ? node658 : 3'b001;
										assign node658 = (inp[3]) ? 3'b110 : node659;
											assign node659 = (inp[4]) ? 3'b110 : 3'b001;
								assign node663 = (inp[8]) ? node671 : node664;
									assign node664 = (inp[2]) ? 3'b100 : node665;
										assign node665 = (inp[5]) ? node667 : 3'b010;
											assign node667 = (inp[3]) ? 3'b100 : 3'b010;
									assign node671 = (inp[2]) ? node679 : node672;
										assign node672 = (inp[5]) ? node674 : 3'b110;
											assign node674 = (inp[4]) ? node676 : 3'b110;
												assign node676 = (inp[3]) ? 3'b010 : 3'b110;
										assign node679 = (inp[4]) ? 3'b010 : node680;
											assign node680 = (inp[5]) ? 3'b010 : 3'b110;
						assign node684 = (inp[1]) ? node716 : node685;
							assign node685 = (inp[8]) ? node701 : node686;
								assign node686 = (inp[11]) ? node696 : node687;
									assign node687 = (inp[2]) ? node689 : 3'b010;
										assign node689 = (inp[3]) ? 3'b100 : node690;
											assign node690 = (inp[5]) ? node692 : 3'b010;
												assign node692 = (inp[4]) ? 3'b100 : 3'b010;
									assign node696 = (inp[2]) ? node698 : 3'b100;
										assign node698 = (inp[3]) ? 3'b000 : 3'b100;
								assign node701 = (inp[11]) ? node707 : node702;
									assign node702 = (inp[3]) ? node704 : 3'b110;
										assign node704 = (inp[2]) ? 3'b010 : 3'b110;
									assign node707 = (inp[4]) ? 3'b010 : node708;
										assign node708 = (inp[2]) ? 3'b100 : node709;
											assign node709 = (inp[5]) ? 3'b010 : node710;
												assign node710 = (inp[3]) ? 3'b010 : 3'b110;
							assign node716 = (inp[8]) ? node728 : node717;
								assign node717 = (inp[11]) ? 3'b000 : node718;
									assign node718 = (inp[2]) ? node720 : 3'b100;
										assign node720 = (inp[5]) ? 3'b000 : node721;
											assign node721 = (inp[3]) ? 3'b000 : node722;
												assign node722 = (inp[4]) ? 3'b000 : 3'b100;
								assign node728 = (inp[11]) ? node738 : node729;
									assign node729 = (inp[2]) ? node731 : 3'b010;
										assign node731 = (inp[5]) ? 3'b100 : node732;
											assign node732 = (inp[3]) ? 3'b100 : node733;
												assign node733 = (inp[4]) ? 3'b100 : 3'b010;
									assign node738 = (inp[2]) ? node740 : 3'b100;
										assign node740 = (inp[3]) ? 3'b000 : node741;
											assign node741 = (inp[4]) ? 3'b000 : 3'b100;
					assign node745 = (inp[10]) ? node821 : node746;
						assign node746 = (inp[1]) ? node790 : node747;
							assign node747 = (inp[8]) ? node771 : node748;
								assign node748 = (inp[11]) ? node758 : node749;
									assign node749 = (inp[3]) ? node755 : node750;
										assign node750 = (inp[2]) ? 3'b011 : node751;
											assign node751 = (inp[4]) ? 3'b011 : 3'b111;
										assign node755 = (inp[2]) ? 3'b101 : 3'b011;
									assign node758 = (inp[3]) ? node764 : node759;
										assign node759 = (inp[4]) ? 3'b101 : node760;
											assign node760 = (inp[5]) ? 3'b101 : 3'b011;
										assign node764 = (inp[2]) ? node766 : 3'b101;
											assign node766 = (inp[4]) ? 3'b001 : node767;
												assign node767 = (inp[5]) ? 3'b001 : 3'b101;
								assign node771 = (inp[11]) ? node779 : node772;
									assign node772 = (inp[3]) ? node774 : 3'b111;
										assign node774 = (inp[2]) ? node776 : 3'b111;
											assign node776 = (inp[5]) ? 3'b011 : 3'b111;
									assign node779 = (inp[4]) ? node785 : node780;
										assign node780 = (inp[3]) ? 3'b011 : node781;
											assign node781 = (inp[2]) ? 3'b011 : 3'b111;
										assign node785 = (inp[2]) ? node787 : 3'b011;
											assign node787 = (inp[3]) ? 3'b101 : 3'b011;
							assign node790 = (inp[8]) ? node806 : node791;
								assign node791 = (inp[11]) ? node799 : node792;
									assign node792 = (inp[2]) ? node794 : 3'b101;
										assign node794 = (inp[3]) ? 3'b001 : node795;
											assign node795 = (inp[4]) ? 3'b001 : 3'b101;
									assign node799 = (inp[2]) ? node801 : 3'b001;
										assign node801 = (inp[4]) ? 3'b110 : node802;
											assign node802 = (inp[3]) ? 3'b110 : 3'b001;
								assign node806 = (inp[11]) ? node814 : node807;
									assign node807 = (inp[2]) ? node809 : 3'b011;
										assign node809 = (inp[3]) ? 3'b101 : node810;
											assign node810 = (inp[4]) ? 3'b101 : 3'b011;
									assign node814 = (inp[2]) ? node816 : 3'b101;
										assign node816 = (inp[3]) ? 3'b001 : node817;
											assign node817 = (inp[4]) ? 3'b001 : 3'b101;
						assign node821 = (inp[1]) ? node869 : node822;
							assign node822 = (inp[8]) ? node848 : node823;
								assign node823 = (inp[11]) ? node839 : node824;
									assign node824 = (inp[2]) ? node832 : node825;
										assign node825 = (inp[3]) ? 3'b001 : node826;
											assign node826 = (inp[5]) ? 3'b001 : node827;
												assign node827 = (inp[4]) ? 3'b001 : 3'b101;
										assign node832 = (inp[3]) ? node834 : 3'b001;
											assign node834 = (inp[5]) ? 3'b110 : node835;
												assign node835 = (inp[4]) ? 3'b110 : 3'b001;
									assign node839 = (inp[4]) ? node843 : node840;
										assign node840 = (inp[3]) ? 3'b110 : 3'b001;
										assign node843 = (inp[2]) ? node845 : 3'b110;
											assign node845 = (inp[3]) ? 3'b010 : 3'b110;
								assign node848 = (inp[11]) ? node864 : node849;
									assign node849 = (inp[5]) ? node857 : node850;
										assign node850 = (inp[2]) ? node852 : 3'b101;
											assign node852 = (inp[3]) ? node854 : 3'b101;
												assign node854 = (inp[4]) ? 3'b001 : 3'b101;
										assign node857 = (inp[3]) ? node861 : node858;
											assign node858 = (inp[4]) ? 3'b101 : 3'b011;
											assign node861 = (inp[4]) ? 3'b001 : 3'b101;
									assign node864 = (inp[2]) ? 3'b001 : node865;
										assign node865 = (inp[3]) ? 3'b001 : 3'b101;
							assign node869 = (inp[8]) ? node885 : node870;
								assign node870 = (inp[11]) ? node878 : node871;
									assign node871 = (inp[2]) ? node873 : 3'b110;
										assign node873 = (inp[4]) ? 3'b010 : node874;
											assign node874 = (inp[3]) ? 3'b010 : 3'b110;
									assign node878 = (inp[2]) ? node880 : 3'b010;
										assign node880 = (inp[3]) ? 3'b100 : node881;
											assign node881 = (inp[5]) ? 3'b100 : 3'b010;
								assign node885 = (inp[11]) ? node891 : node886;
									assign node886 = (inp[2]) ? node888 : 3'b001;
										assign node888 = (inp[3]) ? 3'b110 : 3'b001;
									assign node891 = (inp[2]) ? node893 : 3'b110;
										assign node893 = (inp[3]) ? 3'b010 : 3'b110;
			assign node896 = (inp[0]) ? node1122 : node897;
				assign node897 = (inp[7]) ? node1005 : node898;
					assign node898 = (inp[10]) ? node962 : node899;
						assign node899 = (inp[1]) ? node933 : node900;
							assign node900 = (inp[8]) ? node912 : node901;
								assign node901 = (inp[11]) ? node905 : node902;
									assign node902 = (inp[2]) ? 3'b010 : 3'b110;
									assign node905 = (inp[2]) ? 3'b100 : node906;
										assign node906 = (inp[4]) ? node908 : 3'b010;
											assign node908 = (inp[3]) ? 3'b100 : 3'b010;
								assign node912 = (inp[2]) ? node924 : node913;
									assign node913 = (inp[11]) ? node919 : node914;
										assign node914 = (inp[5]) ? node916 : 3'b001;
											assign node916 = (inp[3]) ? 3'b110 : 3'b001;
										assign node919 = (inp[3]) ? node921 : 3'b110;
											assign node921 = (inp[5]) ? 3'b010 : 3'b110;
									assign node924 = (inp[11]) ? node926 : 3'b110;
										assign node926 = (inp[5]) ? 3'b010 : node927;
											assign node927 = (inp[4]) ? 3'b010 : node928;
												assign node928 = (inp[3]) ? 3'b010 : 3'b110;
							assign node933 = (inp[11]) ? node951 : node934;
								assign node934 = (inp[8]) ? node946 : node935;
									assign node935 = (inp[3]) ? node941 : node936;
										assign node936 = (inp[4]) ? 3'b100 : node937;
											assign node937 = (inp[2]) ? 3'b100 : 3'b010;
										assign node941 = (inp[4]) ? node943 : 3'b100;
											assign node943 = (inp[2]) ? 3'b000 : 3'b100;
									assign node946 = (inp[3]) ? 3'b010 : node947;
										assign node947 = (inp[2]) ? 3'b010 : 3'b110;
								assign node951 = (inp[8]) ? node957 : node952;
									assign node952 = (inp[4]) ? 3'b000 : node953;
										assign node953 = (inp[2]) ? 3'b000 : 3'b100;
									assign node957 = (inp[3]) ? 3'b100 : node958;
										assign node958 = (inp[2]) ? 3'b100 : 3'b010;
						assign node962 = (inp[1]) ? node992 : node963;
							assign node963 = (inp[8]) ? node973 : node964;
								assign node964 = (inp[2]) ? 3'b000 : node965;
									assign node965 = (inp[11]) ? 3'b000 : node966;
										assign node966 = (inp[5]) ? node968 : 3'b100;
											assign node968 = (inp[4]) ? 3'b000 : 3'b100;
								assign node973 = (inp[11]) ? node983 : node974;
									assign node974 = (inp[2]) ? 3'b100 : node975;
										assign node975 = (inp[3]) ? node977 : 3'b010;
											assign node977 = (inp[4]) ? node979 : 3'b010;
												assign node979 = (inp[5]) ? 3'b100 : 3'b010;
									assign node983 = (inp[2]) ? node985 : 3'b100;
										assign node985 = (inp[5]) ? 3'b000 : node986;
											assign node986 = (inp[3]) ? 3'b000 : node987;
												assign node987 = (inp[4]) ? 3'b000 : 3'b100;
							assign node992 = (inp[11]) ? 3'b000 : node993;
								assign node993 = (inp[8]) ? node995 : 3'b000;
									assign node995 = (inp[2]) ? 3'b000 : node996;
										assign node996 = (inp[3]) ? node998 : 3'b100;
											assign node998 = (inp[4]) ? 3'b000 : node999;
												assign node999 = (inp[5]) ? 3'b000 : 3'b100;
					assign node1005 = (inp[10]) ? node1067 : node1006;
						assign node1006 = (inp[1]) ? node1038 : node1007;
							assign node1007 = (inp[8]) ? node1023 : node1008;
								assign node1008 = (inp[11]) ? node1016 : node1009;
									assign node1009 = (inp[2]) ? 3'b001 : node1010;
										assign node1010 = (inp[3]) ? node1012 : 3'b101;
											assign node1012 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1016 = (inp[2]) ? node1018 : 3'b001;
										assign node1018 = (inp[4]) ? 3'b110 : node1019;
											assign node1019 = (inp[3]) ? 3'b110 : 3'b001;
								assign node1023 = (inp[11]) ? node1031 : node1024;
									assign node1024 = (inp[2]) ? node1026 : 3'b011;
										assign node1026 = (inp[4]) ? 3'b101 : node1027;
											assign node1027 = (inp[3]) ? 3'b101 : 3'b011;
									assign node1031 = (inp[2]) ? node1033 : 3'b101;
										assign node1033 = (inp[3]) ? 3'b001 : node1034;
											assign node1034 = (inp[4]) ? 3'b001 : 3'b101;
							assign node1038 = (inp[8]) ? node1052 : node1039;
								assign node1039 = (inp[11]) ? node1045 : node1040;
									assign node1040 = (inp[3]) ? 3'b110 : node1041;
										assign node1041 = (inp[2]) ? 3'b110 : 3'b001;
									assign node1045 = (inp[2]) ? 3'b010 : node1046;
										assign node1046 = (inp[5]) ? node1048 : 3'b110;
											assign node1048 = (inp[3]) ? 3'b010 : 3'b110;
								assign node1052 = (inp[11]) ? node1060 : node1053;
									assign node1053 = (inp[2]) ? 3'b001 : node1054;
										assign node1054 = (inp[4]) ? node1056 : 3'b101;
											assign node1056 = (inp[3]) ? 3'b001 : 3'b101;
									assign node1060 = (inp[2]) ? 3'b110 : node1061;
										assign node1061 = (inp[4]) ? node1063 : 3'b001;
											assign node1063 = (inp[5]) ? 3'b110 : 3'b001;
						assign node1067 = (inp[1]) ? node1095 : node1068;
							assign node1068 = (inp[11]) ? node1082 : node1069;
								assign node1069 = (inp[8]) ? node1077 : node1070;
									assign node1070 = (inp[2]) ? node1072 : 3'b110;
										assign node1072 = (inp[3]) ? 3'b010 : node1073;
											assign node1073 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1077 = (inp[3]) ? node1079 : 3'b001;
										assign node1079 = (inp[2]) ? 3'b110 : 3'b001;
								assign node1082 = (inp[8]) ? node1090 : node1083;
									assign node1083 = (inp[2]) ? node1085 : 3'b010;
										assign node1085 = (inp[3]) ? 3'b100 : node1086;
											assign node1086 = (inp[4]) ? 3'b100 : 3'b010;
									assign node1090 = (inp[2]) ? node1092 : 3'b110;
										assign node1092 = (inp[3]) ? 3'b010 : 3'b110;
							assign node1095 = (inp[11]) ? node1111 : node1096;
								assign node1096 = (inp[8]) ? node1104 : node1097;
									assign node1097 = (inp[2]) ? 3'b100 : node1098;
										assign node1098 = (inp[4]) ? node1100 : 3'b010;
											assign node1100 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1104 = (inp[2]) ? 3'b010 : node1105;
										assign node1105 = (inp[3]) ? node1107 : 3'b110;
											assign node1107 = (inp[4]) ? 3'b010 : 3'b110;
								assign node1111 = (inp[8]) ? node1119 : node1112;
									assign node1112 = (inp[2]) ? 3'b000 : node1113;
										assign node1113 = (inp[4]) ? node1115 : 3'b100;
											assign node1115 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1119 = (inp[2]) ? 3'b100 : 3'b010;
				assign node1122 = (inp[7]) ? node1148 : node1123;
					assign node1123 = (inp[10]) ? 3'b000 : node1124;
						assign node1124 = (inp[8]) ? node1126 : 3'b000;
							assign node1126 = (inp[1]) ? 3'b000 : node1127;
								assign node1127 = (inp[11]) ? node1139 : node1128;
									assign node1128 = (inp[2]) ? node1136 : node1129;
										assign node1129 = (inp[5]) ? 3'b100 : node1130;
											assign node1130 = (inp[3]) ? 3'b100 : node1131;
												assign node1131 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1136 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1139 = (inp[3]) ? 3'b000 : node1140;
										assign node1140 = (inp[4]) ? 3'b000 : node1141;
											assign node1141 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1148 = (inp[10]) ? node1224 : node1149;
						assign node1149 = (inp[1]) ? node1195 : node1150;
							assign node1150 = (inp[8]) ? node1174 : node1151;
								assign node1151 = (inp[11]) ? node1163 : node1152;
									assign node1152 = (inp[2]) ? node1158 : node1153;
										assign node1153 = (inp[4]) ? 3'b010 : node1154;
											assign node1154 = (inp[3]) ? 3'b010 : 3'b110;
										assign node1158 = (inp[3]) ? node1160 : 3'b010;
											assign node1160 = (inp[4]) ? 3'b100 : 3'b010;
									assign node1163 = (inp[2]) ? node1171 : node1164;
										assign node1164 = (inp[3]) ? 3'b100 : node1165;
											assign node1165 = (inp[4]) ? node1167 : 3'b010;
												assign node1167 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1171 = (inp[3]) ? 3'b000 : 3'b100;
								assign node1174 = (inp[11]) ? node1190 : node1175;
									assign node1175 = (inp[3]) ? node1183 : node1176;
										assign node1176 = (inp[2]) ? 3'b110 : node1177;
											assign node1177 = (inp[5]) ? node1179 : 3'b001;
												assign node1179 = (inp[4]) ? 3'b110 : 3'b001;
										assign node1183 = (inp[4]) ? node1185 : 3'b110;
											assign node1185 = (inp[5]) ? node1187 : 3'b110;
												assign node1187 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1190 = (inp[2]) ? 3'b010 : node1191;
										assign node1191 = (inp[3]) ? 3'b010 : 3'b110;
							assign node1195 = (inp[8]) ? node1207 : node1196;
								assign node1196 = (inp[11]) ? 3'b000 : node1197;
									assign node1197 = (inp[2]) ? node1199 : 3'b100;
										assign node1199 = (inp[3]) ? 3'b000 : node1200;
											assign node1200 = (inp[4]) ? node1202 : 3'b100;
												assign node1202 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1207 = (inp[11]) ? node1213 : node1208;
									assign node1208 = (inp[3]) ? node1210 : 3'b010;
										assign node1210 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1213 = (inp[3]) ? node1221 : node1214;
										assign node1214 = (inp[5]) ? 3'b100 : node1215;
											assign node1215 = (inp[4]) ? 3'b100 : node1216;
												assign node1216 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1221 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1224 = (inp[1]) ? 3'b000 : node1225;
							assign node1225 = (inp[8]) ? node1235 : node1226;
								assign node1226 = (inp[2]) ? 3'b000 : node1227;
									assign node1227 = (inp[3]) ? 3'b000 : node1228;
										assign node1228 = (inp[11]) ? 3'b000 : node1229;
											assign node1229 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1235 = (inp[11]) ? node1241 : node1236;
									assign node1236 = (inp[2]) ? 3'b100 : node1237;
										assign node1237 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1241 = (inp[3]) ? 3'b000 : node1242;
										assign node1242 = (inp[2]) ? 3'b000 : 3'b100;

endmodule