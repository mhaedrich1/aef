module dtc_split66_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node15;
	wire [4-1:0] node16;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node41;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node65;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node70;
	wire [4-1:0] node73;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node97;
	wire [4-1:0] node100;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node110;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node121;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node147;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node152;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node159;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node167;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node173;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node180;
	wire [4-1:0] node183;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node196;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node205;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node211;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node227;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node234;
	wire [4-1:0] node237;
	wire [4-1:0] node240;
	wire [4-1:0] node241;
	wire [4-1:0] node244;
	wire [4-1:0] node246;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node254;
	wire [4-1:0] node257;
	wire [4-1:0] node259;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node271;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node275;
	wire [4-1:0] node280;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node285;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node300;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node307;
	wire [4-1:0] node309;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node316;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node325;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node331;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node342;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node362;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node370;
	wire [4-1:0] node373;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node393;
	wire [4-1:0] node396;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node421;
	wire [4-1:0] node423;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node506;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node513;
	wire [4-1:0] node515;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node533;
	wire [4-1:0] node536;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node544;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node551;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node573;
	wire [4-1:0] node575;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node584;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node598;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node609;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node632;
	wire [4-1:0] node634;
	wire [4-1:0] node636;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node684;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node690;
	wire [4-1:0] node692;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node713;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node727;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node766;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node775;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node793;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node806;
	wire [4-1:0] node809;
	wire [4-1:0] node811;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node822;
	wire [4-1:0] node825;
	wire [4-1:0] node826;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node848;
	wire [4-1:0] node850;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node864;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node876;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node920;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node927;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node936;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node945;
	wire [4-1:0] node948;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node954;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node969;
	wire [4-1:0] node972;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node987;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node994;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1009;
	wire [4-1:0] node1011;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1026;
	wire [4-1:0] node1028;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1042;
	wire [4-1:0] node1045;
	wire [4-1:0] node1048;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1055;
	wire [4-1:0] node1057;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1064;
	wire [4-1:0] node1067;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1090;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1137;
	wire [4-1:0] node1139;
	wire [4-1:0] node1141;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1150;
	wire [4-1:0] node1153;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1165;
	wire [4-1:0] node1167;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1203;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1270;
	wire [4-1:0] node1272;
	wire [4-1:0] node1275;
	wire [4-1:0] node1277;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1283;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1297;
	wire [4-1:0] node1299;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1314;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1330;
	wire [4-1:0] node1333;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1368;
	wire [4-1:0] node1370;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1377;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1387;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1394;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1403;
	wire [4-1:0] node1407;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1435;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1448;
	wire [4-1:0] node1449;
	wire [4-1:0] node1451;
	wire [4-1:0] node1454;
	wire [4-1:0] node1456;
	wire [4-1:0] node1459;
	wire [4-1:0] node1461;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1470;
	wire [4-1:0] node1471;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1481;
	wire [4-1:0] node1483;
	wire [4-1:0] node1486;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1499;
	wire [4-1:0] node1500;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1505;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1524;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1541;
	wire [4-1:0] node1543;
	wire [4-1:0] node1546;
	wire [4-1:0] node1548;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1554;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1564;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1570;
	wire [4-1:0] node1573;
	wire [4-1:0] node1575;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1597;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1605;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1612;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1619;
	wire [4-1:0] node1621;
	wire [4-1:0] node1624;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1630;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1652;
	wire [4-1:0] node1655;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1672;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1681;
	wire [4-1:0] node1684;
	wire [4-1:0] node1686;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1698;
	wire [4-1:0] node1700;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1706;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1731;
	wire [4-1:0] node1734;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1740;
	wire [4-1:0] node1744;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1753;
	wire [4-1:0] node1754;
	wire [4-1:0] node1757;
	wire [4-1:0] node1760;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1765;
	wire [4-1:0] node1768;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1774;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1790;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1798;
	wire [4-1:0] node1801;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1812;
	wire [4-1:0] node1814;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1826;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1831;
	wire [4-1:0] node1834;
	wire [4-1:0] node1835;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1848;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1869;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1890;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1897;
	wire [4-1:0] node1901;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1918;
	wire [4-1:0] node1920;
	wire [4-1:0] node1923;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1937;
	wire [4-1:0] node1940;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1945;
	wire [4-1:0] node1946;
	wire [4-1:0] node1949;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1957;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1964;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1996;
	wire [4-1:0] node1997;
	wire [4-1:0] node2000;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2006;
	wire [4-1:0] node2008;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2045;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2053;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2062;
	wire [4-1:0] node2065;
	wire [4-1:0] node2068;
	wire [4-1:0] node2069;
	wire [4-1:0] node2072;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2110;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2138;
	wire [4-1:0] node2141;
	wire [4-1:0] node2143;
	wire [4-1:0] node2145;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2151;
	wire [4-1:0] node2152;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2167;
	wire [4-1:0] node2168;
	wire [4-1:0] node2170;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2179;
	wire [4-1:0] node2182;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2203;
	wire [4-1:0] node2206;
	wire [4-1:0] node2207;
	wire [4-1:0] node2208;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2218;
	wire [4-1:0] node2221;
	wire [4-1:0] node2223;
	wire [4-1:0] node2225;
	wire [4-1:0] node2228;
	wire [4-1:0] node2229;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2235;
	wire [4-1:0] node2237;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2243;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2257;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2263;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2272;
	wire [4-1:0] node2273;
	wire [4-1:0] node2274;
	wire [4-1:0] node2278;
	wire [4-1:0] node2281;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2286;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2294;
	wire [4-1:0] node2295;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2309;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;
	wire [4-1:0] node2315;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2324;
	wire [4-1:0] node2326;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2339;
	wire [4-1:0] node2342;
	wire [4-1:0] node2343;
	wire [4-1:0] node2344;
	wire [4-1:0] node2345;
	wire [4-1:0] node2348;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2357;
	wire [4-1:0] node2360;
	wire [4-1:0] node2361;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2367;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2379;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2395;
	wire [4-1:0] node2397;
	wire [4-1:0] node2399;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2416;
	wire [4-1:0] node2420;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2430;
	wire [4-1:0] node2433;
	wire [4-1:0] node2435;
	wire [4-1:0] node2437;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2449;
	wire [4-1:0] node2451;
	wire [4-1:0] node2454;
	wire [4-1:0] node2455;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2467;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2472;
	wire [4-1:0] node2473;
	wire [4-1:0] node2474;
	wire [4-1:0] node2475;
	wire [4-1:0] node2479;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2498;
	wire [4-1:0] node2501;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2506;
	wire [4-1:0] node2507;
	wire [4-1:0] node2508;
	wire [4-1:0] node2511;
	wire [4-1:0] node2514;
	wire [4-1:0] node2517;
	wire [4-1:0] node2518;
	wire [4-1:0] node2521;
	wire [4-1:0] node2524;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2529;
	wire [4-1:0] node2532;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2538;
	wire [4-1:0] node2541;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2549;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2559;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2573;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2579;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2587;
	wire [4-1:0] node2588;
	wire [4-1:0] node2590;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2597;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2614;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2630;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2635;
	wire [4-1:0] node2636;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2644;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2650;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2664;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2679;
	wire [4-1:0] node2681;
	wire [4-1:0] node2684;
	wire [4-1:0] node2686;
	wire [4-1:0] node2688;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2704;
	wire [4-1:0] node2707;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2724;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2732;
	wire [4-1:0] node2736;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2753;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2760;
	wire [4-1:0] node2762;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2772;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2778;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2801;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2818;
	wire [4-1:0] node2821;
	wire [4-1:0] node2823;
	wire [4-1:0] node2825;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2835;
	wire [4-1:0] node2839;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2848;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2869;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2882;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2889;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2908;
	wire [4-1:0] node2911;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2917;
	wire [4-1:0] node2921;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2934;
	wire [4-1:0] node2937;
	wire [4-1:0] node2940;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2947;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2959;
	wire [4-1:0] node2960;
	wire [4-1:0] node2961;
	wire [4-1:0] node2962;
	wire [4-1:0] node2965;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2970;
	wire [4-1:0] node2974;
	wire [4-1:0] node2976;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2981;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2991;
	wire [4-1:0] node2993;
	wire [4-1:0] node2996;
	wire [4-1:0] node2997;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3006;
	wire [4-1:0] node3007;
	wire [4-1:0] node3010;
	wire [4-1:0] node3012;
	wire [4-1:0] node3015;
	wire [4-1:0] node3016;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3038;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3060;
	wire [4-1:0] node3061;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3071;
	wire [4-1:0] node3074;
	wire [4-1:0] node3076;
	wire [4-1:0] node3079;
	wire [4-1:0] node3080;
	wire [4-1:0] node3082;
	wire [4-1:0] node3086;
	wire [4-1:0] node3087;
	wire [4-1:0] node3088;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3096;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3106;
	wire [4-1:0] node3109;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3112;
	wire [4-1:0] node3115;
	wire [4-1:0] node3117;
	wire [4-1:0] node3120;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3125;
	wire [4-1:0] node3128;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3150;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3173;
	wire [4-1:0] node3175;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3180;
	wire [4-1:0] node3182;
	wire [4-1:0] node3185;
	wire [4-1:0] node3188;
	wire [4-1:0] node3190;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3199;
	wire [4-1:0] node3201;
	wire [4-1:0] node3204;
	wire [4-1:0] node3205;
	wire [4-1:0] node3207;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3215;
	wire [4-1:0] node3216;
	wire [4-1:0] node3219;
	wire [4-1:0] node3220;
	wire [4-1:0] node3222;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3235;
	wire [4-1:0] node3238;
	wire [4-1:0] node3239;
	wire [4-1:0] node3240;
	wire [4-1:0] node3243;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3263;
	wire [4-1:0] node3264;
	wire [4-1:0] node3267;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3278;
	wire [4-1:0] node3281;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3288;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3292;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3300;
	wire [4-1:0] node3301;
	wire [4-1:0] node3304;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3315;
	wire [4-1:0] node3316;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3323;
	wire [4-1:0] node3326;
	wire [4-1:0] node3327;
	wire [4-1:0] node3330;
	wire [4-1:0] node3331;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3341;
	wire [4-1:0] node3343;
	wire [4-1:0] node3346;
	wire [4-1:0] node3348;
	wire [4-1:0] node3350;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3364;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3379;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3386;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3396;
	wire [4-1:0] node3398;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3404;
	wire [4-1:0] node3407;
	wire [4-1:0] node3409;
	wire [4-1:0] node3412;
	wire [4-1:0] node3413;
	wire [4-1:0] node3414;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3421;
	wire [4-1:0] node3423;
	wire [4-1:0] node3426;
	wire [4-1:0] node3427;
	wire [4-1:0] node3429;
	wire [4-1:0] node3430;
	wire [4-1:0] node3434;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3444;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3449;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3453;
	wire [4-1:0] node3455;
	wire [4-1:0] node3458;
	wire [4-1:0] node3459;
	wire [4-1:0] node3460;
	wire [4-1:0] node3463;
	wire [4-1:0] node3466;
	wire [4-1:0] node3469;
	wire [4-1:0] node3470;
	wire [4-1:0] node3472;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3488;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3500;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3507;
	wire [4-1:0] node3510;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3517;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3528;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3553;
	wire [4-1:0] node3555;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3560;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3571;
	wire [4-1:0] node3573;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3579;
	wire [4-1:0] node3582;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3587;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3595;
	wire [4-1:0] node3597;
	wire [4-1:0] node3599;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3607;
	wire [4-1:0] node3608;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3615;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3622;
	wire [4-1:0] node3624;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3630;
	wire [4-1:0] node3633;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3640;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3646;
	wire [4-1:0] node3649;
	wire [4-1:0] node3650;
	wire [4-1:0] node3653;
	wire [4-1:0] node3655;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3660;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3664;
	wire [4-1:0] node3668;
	wire [4-1:0] node3669;
	wire [4-1:0] node3672;
	wire [4-1:0] node3673;
	wire [4-1:0] node3676;
	wire [4-1:0] node3679;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3684;
	wire [4-1:0] node3686;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3691;
	wire [4-1:0] node3696;
	wire [4-1:0] node3697;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3706;
	wire [4-1:0] node3709;
	wire [4-1:0] node3710;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3722;
	wire [4-1:0] node3725;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3732;
	wire [4-1:0] node3733;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3742;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3755;
	wire [4-1:0] node3756;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3763;
	wire [4-1:0] node3765;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3770;
	wire [4-1:0] node3771;
	wire [4-1:0] node3773;
	wire [4-1:0] node3776;
	wire [4-1:0] node3779;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3786;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3793;
	wire [4-1:0] node3795;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3803;
	wire [4-1:0] node3806;
	wire [4-1:0] node3807;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3823;
	wire [4-1:0] node3824;
	wire [4-1:0] node3827;
	wire [4-1:0] node3830;
	wire [4-1:0] node3831;
	wire [4-1:0] node3832;
	wire [4-1:0] node3833;
	wire [4-1:0] node3836;
	wire [4-1:0] node3839;
	wire [4-1:0] node3841;
	wire [4-1:0] node3844;
	wire [4-1:0] node3845;
	wire [4-1:0] node3846;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3860;
	wire [4-1:0] node3863;
	wire [4-1:0] node3866;
	wire [4-1:0] node3868;
	wire [4-1:0] node3870;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3876;
	wire [4-1:0] node3878;
	wire [4-1:0] node3881;
	wire [4-1:0] node3883;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3891;
	wire [4-1:0] node3892;
	wire [4-1:0] node3893;
	wire [4-1:0] node3894;
	wire [4-1:0] node3897;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3911;
	wire [4-1:0] node3912;
	wire [4-1:0] node3913;
	wire [4-1:0] node3915;
	wire [4-1:0] node3918;
	wire [4-1:0] node3921;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3928;
	wire [4-1:0] node3929;
	wire [4-1:0] node3930;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3938;
	wire [4-1:0] node3942;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3946;
	wire [4-1:0] node3949;
	wire [4-1:0] node3952;
	wire [4-1:0] node3953;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3969;
	wire [4-1:0] node3971;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3979;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3988;
	wire [4-1:0] node3991;
	wire [4-1:0] node3992;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3997;
	wire [4-1:0] node3998;
	wire [4-1:0] node4001;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4020;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4039;
	wire [4-1:0] node4040;
	wire [4-1:0] node4042;
	wire [4-1:0] node4045;
	wire [4-1:0] node4047;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4055;
	wire [4-1:0] node4058;
	wire [4-1:0] node4059;
	wire [4-1:0] node4063;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4073;
	wire [4-1:0] node4076;
	wire [4-1:0] node4078;
	wire [4-1:0] node4081;
	wire [4-1:0] node4082;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4093;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4102;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4107;
	wire [4-1:0] node4110;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4122;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4137;
	wire [4-1:0] node4138;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4145;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4151;
	wire [4-1:0] node4156;
	wire [4-1:0] node4158;
	wire [4-1:0] node4160;
	wire [4-1:0] node4163;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4168;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4176;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4184;
	wire [4-1:0] node4185;
	wire [4-1:0] node4186;
	wire [4-1:0] node4188;
	wire [4-1:0] node4191;
	wire [4-1:0] node4194;
	wire [4-1:0] node4196;
	wire [4-1:0] node4198;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4204;
	wire [4-1:0] node4205;
	wire [4-1:0] node4208;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4214;
	wire [4-1:0] node4217;
	wire [4-1:0] node4219;
	wire [4-1:0] node4222;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4227;
	wire [4-1:0] node4230;
	wire [4-1:0] node4233;
	wire [4-1:0] node4234;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4243;
	wire [4-1:0] node4246;
	wire [4-1:0] node4248;
	wire [4-1:0] node4251;
	wire [4-1:0] node4252;
	wire [4-1:0] node4253;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4260;
	wire [4-1:0] node4263;
	wire [4-1:0] node4265;
	wire [4-1:0] node4268;
	wire [4-1:0] node4269;
	wire [4-1:0] node4270;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4275;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4282;
	wire [4-1:0] node4285;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4294;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4301;
	wire [4-1:0] node4302;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4321;
	wire [4-1:0] node4324;
	wire [4-1:0] node4326;
	wire [4-1:0] node4329;
	wire [4-1:0] node4330;
	wire [4-1:0] node4331;
	wire [4-1:0] node4332;
	wire [4-1:0] node4335;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4342;
	wire [4-1:0] node4345;
	wire [4-1:0] node4346;
	wire [4-1:0] node4347;
	wire [4-1:0] node4352;
	wire [4-1:0] node4353;
	wire [4-1:0] node4354;
	wire [4-1:0] node4355;
	wire [4-1:0] node4358;
	wire [4-1:0] node4361;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4369;
	wire [4-1:0] node4372;
	wire [4-1:0] node4373;
	wire [4-1:0] node4374;
	wire [4-1:0] node4377;
	wire [4-1:0] node4380;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4391;
	wire [4-1:0] node4392;
	wire [4-1:0] node4395;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4401;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4409;
	wire [4-1:0] node4412;
	wire [4-1:0] node4414;
	wire [4-1:0] node4417;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4421;
	wire [4-1:0] node4422;
	wire [4-1:0] node4425;
	wire [4-1:0] node4429;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4439;
	wire [4-1:0] node4442;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4450;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4456;
	wire [4-1:0] node4457;
	wire [4-1:0] node4460;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4468;
	wire [4-1:0] node4470;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4477;
	wire [4-1:0] node4480;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4484;
	wire [4-1:0] node4487;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4495;
	wire [4-1:0] node4497;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4511;
	wire [4-1:0] node4512;
	wire [4-1:0] node4513;
	wire [4-1:0] node4516;
	wire [4-1:0] node4519;
	wire [4-1:0] node4520;
	wire [4-1:0] node4523;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4533;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4543;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4547;
	wire [4-1:0] node4550;
	wire [4-1:0] node4551;
	wire [4-1:0] node4552;
	wire [4-1:0] node4555;
	wire [4-1:0] node4559;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4562;
	wire [4-1:0] node4565;
	wire [4-1:0] node4569;
	wire [4-1:0] node4571;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4576;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4583;
	wire [4-1:0] node4585;
	wire [4-1:0] node4588;
	wire [4-1:0] node4590;
	wire [4-1:0] node4592;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4599;
	wire [4-1:0] node4602;
	wire [4-1:0] node4603;
	wire [4-1:0] node4606;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4611;
	wire [4-1:0] node4614;
	wire [4-1:0] node4617;
	wire [4-1:0] node4619;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4626;
	wire [4-1:0] node4628;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4635;
	wire [4-1:0] node4638;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4648;
	wire [4-1:0] node4651;
	wire [4-1:0] node4654;
	wire [4-1:0] node4656;
	wire [4-1:0] node4659;
	wire [4-1:0] node4661;
	wire [4-1:0] node4662;
	wire [4-1:0] node4666;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4673;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4683;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4690;
	wire [4-1:0] node4691;
	wire [4-1:0] node4692;
	wire [4-1:0] node4695;
	wire [4-1:0] node4698;
	wire [4-1:0] node4700;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4705;
	wire [4-1:0] node4706;
	wire [4-1:0] node4707;
	wire [4-1:0] node4708;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4713;
	wire [4-1:0] node4716;
	wire [4-1:0] node4717;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4724;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4731;
	wire [4-1:0] node4734;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4740;
	wire [4-1:0] node4743;
	wire [4-1:0] node4744;
	wire [4-1:0] node4747;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4753;
	wire [4-1:0] node4755;
	wire [4-1:0] node4759;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4769;
	wire [4-1:0] node4772;
	wire [4-1:0] node4773;
	wire [4-1:0] node4776;
	wire [4-1:0] node4777;
	wire [4-1:0] node4780;
	wire [4-1:0] node4782;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4788;
	wire [4-1:0] node4790;
	wire [4-1:0] node4793;
	wire [4-1:0] node4794;
	wire [4-1:0] node4796;
	wire [4-1:0] node4800;
	wire [4-1:0] node4802;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4810;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4819;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4830;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4839;
	wire [4-1:0] node4842;
	wire [4-1:0] node4843;
	wire [4-1:0] node4844;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4852;
	wire [4-1:0] node4853;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4861;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4875;
	wire [4-1:0] node4879;
	wire [4-1:0] node4880;
	wire [4-1:0] node4882;
	wire [4-1:0] node4884;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4894;
	wire [4-1:0] node4896;
	wire [4-1:0] node4899;
	wire [4-1:0] node4902;
	wire [4-1:0] node4904;
	wire [4-1:0] node4905;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4911;
	wire [4-1:0] node4914;
	wire [4-1:0] node4917;
	wire [4-1:0] node4918;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4928;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4935;
	wire [4-1:0] node4938;
	wire [4-1:0] node4939;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4951;
	wire [4-1:0] node4954;
	wire [4-1:0] node4955;
	wire [4-1:0] node4956;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4975;
	wire [4-1:0] node4978;
	wire [4-1:0] node4981;
	wire [4-1:0] node4982;
	wire [4-1:0] node4984;
	wire [4-1:0] node4987;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4992;
	wire [4-1:0] node4993;
	wire [4-1:0] node4997;
	wire [4-1:0] node5000;
	wire [4-1:0] node5002;
	wire [4-1:0] node5004;
	wire [4-1:0] node5007;
	wire [4-1:0] node5008;
	wire [4-1:0] node5009;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5014;
	wire [4-1:0] node5017;
	wire [4-1:0] node5018;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5029;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5038;
	wire [4-1:0] node5041;
	wire [4-1:0] node5043;
	wire [4-1:0] node5046;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5060;
	wire [4-1:0] node5061;
	wire [4-1:0] node5064;
	wire [4-1:0] node5067;
	wire [4-1:0] node5068;
	wire [4-1:0] node5069;
	wire [4-1:0] node5070;
	wire [4-1:0] node5073;
	wire [4-1:0] node5077;
	wire [4-1:0] node5079;
	wire [4-1:0] node5080;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5088;
	wire [4-1:0] node5089;
	wire [4-1:0] node5092;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5097;
	wire [4-1:0] node5100;
	wire [4-1:0] node5103;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5111;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5122;
	wire [4-1:0] node5123;
	wire [4-1:0] node5124;
	wire [4-1:0] node5125;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5134;
	wire [4-1:0] node5137;
	wire [4-1:0] node5138;
	wire [4-1:0] node5141;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5148;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5158;
	wire [4-1:0] node5161;
	wire [4-1:0] node5163;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5169;
	wire [4-1:0] node5171;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5177;
	wire [4-1:0] node5180;
	wire [4-1:0] node5183;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5191;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5200;
	wire [4-1:0] node5201;
	wire [4-1:0] node5204;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5217;
	wire [4-1:0] node5221;
	wire [4-1:0] node5222;
	wire [4-1:0] node5223;
	wire [4-1:0] node5225;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5232;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5238;
	wire [4-1:0] node5239;
	wire [4-1:0] node5242;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5260;
	wire [4-1:0] node5261;
	wire [4-1:0] node5263;
	wire [4-1:0] node5266;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5271;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5279;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5283;
	wire [4-1:0] node5287;
	wire [4-1:0] node5288;
	wire [4-1:0] node5289;
	wire [4-1:0] node5294;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5300;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5308;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5312;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5322;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5328;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5333;
	wire [4-1:0] node5334;
	wire [4-1:0] node5336;
	wire [4-1:0] node5338;
	wire [4-1:0] node5341;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5346;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5353;
	wire [4-1:0] node5355;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5360;
	wire [4-1:0] node5363;
	wire [4-1:0] node5366;
	wire [4-1:0] node5368;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5378;
	wire [4-1:0] node5380;
	wire [4-1:0] node5382;
	wire [4-1:0] node5385;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5392;
	wire [4-1:0] node5395;
	wire [4-1:0] node5397;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5407;
	wire [4-1:0] node5408;
	wire [4-1:0] node5410;
	wire [4-1:0] node5413;
	wire [4-1:0] node5416;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5420;
	wire [4-1:0] node5423;
	wire [4-1:0] node5425;
	wire [4-1:0] node5429;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5434;
	wire [4-1:0] node5437;
	wire [4-1:0] node5438;
	wire [4-1:0] node5442;
	wire [4-1:0] node5443;
	wire [4-1:0] node5445;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5455;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5463;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5471;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5478;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5484;
	wire [4-1:0] node5486;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5493;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5498;
	wire [4-1:0] node5499;
	wire [4-1:0] node5500;
	wire [4-1:0] node5505;
	wire [4-1:0] node5506;
	wire [4-1:0] node5509;
	wire [4-1:0] node5512;
	wire [4-1:0] node5513;
	wire [4-1:0] node5514;
	wire [4-1:0] node5517;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5525;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5531;
	wire [4-1:0] node5532;
	wire [4-1:0] node5533;
	wire [4-1:0] node5534;
	wire [4-1:0] node5536;
	wire [4-1:0] node5538;
	wire [4-1:0] node5541;
	wire [4-1:0] node5542;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5555;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5563;
	wire [4-1:0] node5564;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5571;
	wire [4-1:0] node5574;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5579;
	wire [4-1:0] node5582;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5588;
	wire [4-1:0] node5592;
	wire [4-1:0] node5595;
	wire [4-1:0] node5596;
	wire [4-1:0] node5599;
	wire [4-1:0] node5600;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5609;
	wire [4-1:0] node5612;
	wire [4-1:0] node5615;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5622;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5627;
	wire [4-1:0] node5629;
	wire [4-1:0] node5633;
	wire [4-1:0] node5635;
	wire [4-1:0] node5638;
	wire [4-1:0] node5639;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5645;
	wire [4-1:0] node5649;
	wire [4-1:0] node5650;
	wire [4-1:0] node5652;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5659;
	wire [4-1:0] node5661;
	wire [4-1:0] node5664;
	wire [4-1:0] node5666;
	wire [4-1:0] node5669;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5675;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5681;
	wire [4-1:0] node5684;
	wire [4-1:0] node5685;
	wire [4-1:0] node5688;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5694;
	wire [4-1:0] node5697;
	wire [4-1:0] node5698;
	wire [4-1:0] node5701;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5706;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5720;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5737;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5745;
	wire [4-1:0] node5748;
	wire [4-1:0] node5749;
	wire [4-1:0] node5750;
	wire [4-1:0] node5753;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5760;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5777;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5782;
	wire [4-1:0] node5785;
	wire [4-1:0] node5786;
	wire [4-1:0] node5789;
	wire [4-1:0] node5792;
	wire [4-1:0] node5793;
	wire [4-1:0] node5794;
	wire [4-1:0] node5795;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5800;
	wire [4-1:0] node5803;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5819;
	wire [4-1:0] node5823;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5827;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5834;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5841;
	wire [4-1:0] node5843;
	wire [4-1:0] node5844;
	wire [4-1:0] node5847;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5856;
	wire [4-1:0] node5859;
	wire [4-1:0] node5860;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5867;
	wire [4-1:0] node5871;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5878;
	wire [4-1:0] node5881;
	wire [4-1:0] node5884;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5889;
	wire [4-1:0] node5892;
	wire [4-1:0] node5893;
	wire [4-1:0] node5896;
	wire [4-1:0] node5898;
	wire [4-1:0] node5901;
	wire [4-1:0] node5902;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5905;
	wire [4-1:0] node5906;
	wire [4-1:0] node5907;
	wire [4-1:0] node5910;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5920;
	wire [4-1:0] node5921;
	wire [4-1:0] node5924;
	wire [4-1:0] node5927;
	wire [4-1:0] node5928;
	wire [4-1:0] node5930;
	wire [4-1:0] node5931;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5938;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5945;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5952;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5964;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5971;
	wire [4-1:0] node5972;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5976;
	wire [4-1:0] node5977;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5983;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5991;
	wire [4-1:0] node5994;
	wire [4-1:0] node5995;
	wire [4-1:0] node5997;
	wire [4-1:0] node6000;
	wire [4-1:0] node6001;
	wire [4-1:0] node6003;
	wire [4-1:0] node6006;
	wire [4-1:0] node6008;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6018;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6031;
	wire [4-1:0] node6033;
	wire [4-1:0] node6036;
	wire [4-1:0] node6037;
	wire [4-1:0] node6041;
	wire [4-1:0] node6043;
	wire [4-1:0] node6044;
	wire [4-1:0] node6047;
	wire [4-1:0] node6050;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6061;
	wire [4-1:0] node6064;
	wire [4-1:0] node6066;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6076;
	wire [4-1:0] node6079;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6085;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6093;
	wire [4-1:0] node6096;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6104;
	wire [4-1:0] node6108;
	wire [4-1:0] node6109;
	wire [4-1:0] node6110;
	wire [4-1:0] node6114;
	wire [4-1:0] node6115;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6124;
	wire [4-1:0] node6127;
	wire [4-1:0] node6129;
	wire [4-1:0] node6131;
	wire [4-1:0] node6134;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6138;
	wire [4-1:0] node6141;
	wire [4-1:0] node6143;
	wire [4-1:0] node6146;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6151;
	wire [4-1:0] node6154;
	wire [4-1:0] node6155;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6163;
	wire [4-1:0] node6164;
	wire [4-1:0] node6168;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6173;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6181;
	wire [4-1:0] node6182;
	wire [4-1:0] node6184;
	wire [4-1:0] node6186;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6201;
	wire [4-1:0] node6204;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6210;
	wire [4-1:0] node6213;
	wire [4-1:0] node6214;
	wire [4-1:0] node6218;
	wire [4-1:0] node6219;
	wire [4-1:0] node6220;
	wire [4-1:0] node6222;
	wire [4-1:0] node6225;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6231;
	wire [4-1:0] node6235;
	wire [4-1:0] node6236;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6242;
	wire [4-1:0] node6246;
	wire [4-1:0] node6247;
	wire [4-1:0] node6250;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6260;
	wire [4-1:0] node6262;
	wire [4-1:0] node6265;
	wire [4-1:0] node6267;
	wire [4-1:0] node6268;
	wire [4-1:0] node6271;
	wire [4-1:0] node6274;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6279;
	wire [4-1:0] node6282;
	wire [4-1:0] node6283;
	wire [4-1:0] node6286;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6293;
	wire [4-1:0] node6297;
	wire [4-1:0] node6299;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6311;
	wire [4-1:0] node6314;
	wire [4-1:0] node6315;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6322;
	wire [4-1:0] node6325;
	wire [4-1:0] node6326;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6336;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6342;
	wire [4-1:0] node6345;
	wire [4-1:0] node6346;
	wire [4-1:0] node6349;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6356;
	wire [4-1:0] node6357;
	wire [4-1:0] node6361;
	wire [4-1:0] node6363;
	wire [4-1:0] node6366;
	wire [4-1:0] node6367;
	wire [4-1:0] node6369;
	wire [4-1:0] node6371;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6378;
	wire [4-1:0] node6381;
	wire [4-1:0] node6382;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6388;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6397;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6405;
	wire [4-1:0] node6406;
	wire [4-1:0] node6407;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6412;
	wire [4-1:0] node6415;
	wire [4-1:0] node6417;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6425;
	wire [4-1:0] node6428;
	wire [4-1:0] node6430;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6435;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6443;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6449;
	wire [4-1:0] node6450;
	wire [4-1:0] node6451;
	wire [4-1:0] node6455;
	wire [4-1:0] node6457;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6463;
	wire [4-1:0] node6466;
	wire [4-1:0] node6468;
	wire [4-1:0] node6471;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6475;
	wire [4-1:0] node6476;
	wire [4-1:0] node6479;
	wire [4-1:0] node6482;
	wire [4-1:0] node6484;
	wire [4-1:0] node6485;
	wire [4-1:0] node6488;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6497;
	wire [4-1:0] node6498;
	wire [4-1:0] node6501;
	wire [4-1:0] node6503;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6511;
	wire [4-1:0] node6514;
	wire [4-1:0] node6515;
	wire [4-1:0] node6518;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6528;
	wire [4-1:0] node6531;
	wire [4-1:0] node6533;
	wire [4-1:0] node6536;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6541;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6550;
	wire [4-1:0] node6553;
	wire [4-1:0] node6554;
	wire [4-1:0] node6557;
	wire [4-1:0] node6560;
	wire [4-1:0] node6561;
	wire [4-1:0] node6563;
	wire [4-1:0] node6565;
	wire [4-1:0] node6568;
	wire [4-1:0] node6569;
	wire [4-1:0] node6572;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6579;
	wire [4-1:0] node6580;
	wire [4-1:0] node6582;
	wire [4-1:0] node6583;
	wire [4-1:0] node6586;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6593;
	wire [4-1:0] node6596;
	wire [4-1:0] node6597;
	wire [4-1:0] node6600;
	wire [4-1:0] node6602;
	wire [4-1:0] node6603;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6609;
	wire [4-1:0] node6610;
	wire [4-1:0] node6614;
	wire [4-1:0] node6615;
	wire [4-1:0] node6616;
	wire [4-1:0] node6619;
	wire [4-1:0] node6622;
	wire [4-1:0] node6623;
	wire [4-1:0] node6626;
	wire [4-1:0] node6629;
	wire [4-1:0] node6630;
	wire [4-1:0] node6631;
	wire [4-1:0] node6634;
	wire [4-1:0] node6636;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6652;
	wire [4-1:0] node6653;
	wire [4-1:0] node6654;
	wire [4-1:0] node6658;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6665;
	wire [4-1:0] node6666;
	wire [4-1:0] node6669;
	wire [4-1:0] node6671;
	wire [4-1:0] node6674;
	wire [4-1:0] node6675;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6683;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6689;
	wire [4-1:0] node6692;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6696;
	wire [4-1:0] node6700;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6717;
	wire [4-1:0] node6718;
	wire [4-1:0] node6721;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6727;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6736;
	wire [4-1:0] node6739;
	wire [4-1:0] node6740;
	wire [4-1:0] node6741;
	wire [4-1:0] node6745;
	wire [4-1:0] node6746;
	wire [4-1:0] node6750;
	wire [4-1:0] node6751;
	wire [4-1:0] node6753;
	wire [4-1:0] node6754;
	wire [4-1:0] node6757;
	wire [4-1:0] node6760;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6765;
	wire [4-1:0] node6769;
	wire [4-1:0] node6770;
	wire [4-1:0] node6771;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6781;
	wire [4-1:0] node6782;
	wire [4-1:0] node6785;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6792;
	wire [4-1:0] node6796;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6802;
	wire [4-1:0] node6805;
	wire [4-1:0] node6806;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6809;
	wire [4-1:0] node6813;
	wire [4-1:0] node6816;
	wire [4-1:0] node6818;
	wire [4-1:0] node6820;
	wire [4-1:0] node6823;
	wire [4-1:0] node6824;
	wire [4-1:0] node6825;
	wire [4-1:0] node6827;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6836;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6842;
	wire [4-1:0] node6845;
	wire [4-1:0] node6848;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6854;
	wire [4-1:0] node6858;
	wire [4-1:0] node6859;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6871;
	wire [4-1:0] node6872;
	wire [4-1:0] node6875;
	wire [4-1:0] node6878;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6888;
	wire [4-1:0] node6889;
	wire [4-1:0] node6892;
	wire [4-1:0] node6895;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6901;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6921;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6928;
	wire [4-1:0] node6931;
	wire [4-1:0] node6932;
	wire [4-1:0] node6935;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6945;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6950;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6961;
	wire [4-1:0] node6962;
	wire [4-1:0] node6966;
	wire [4-1:0] node6968;
	wire [4-1:0] node6969;
	wire [4-1:0] node6973;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6978;
	wire [4-1:0] node6982;
	wire [4-1:0] node6983;
	wire [4-1:0] node6984;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6995;
	wire [4-1:0] node6998;
	wire [4-1:0] node6999;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7003;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7009;
	wire [4-1:0] node7012;
	wire [4-1:0] node7016;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7023;
	wire [4-1:0] node7024;
	wire [4-1:0] node7025;
	wire [4-1:0] node7027;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7033;
	wire [4-1:0] node7035;
	wire [4-1:0] node7038;
	wire [4-1:0] node7039;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7049;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7054;
	wire [4-1:0] node7058;
	wire [4-1:0] node7059;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7066;
	wire [4-1:0] node7067;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7075;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7081;
	wire [4-1:0] node7082;
	wire [4-1:0] node7083;
	wire [4-1:0] node7085;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7098;
	wire [4-1:0] node7101;
	wire [4-1:0] node7103;
	wire [4-1:0] node7104;
	wire [4-1:0] node7107;
	wire [4-1:0] node7110;
	wire [4-1:0] node7111;
	wire [4-1:0] node7112;
	wire [4-1:0] node7114;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7120;
	wire [4-1:0] node7122;
	wire [4-1:0] node7125;
	wire [4-1:0] node7126;
	wire [4-1:0] node7129;
	wire [4-1:0] node7132;
	wire [4-1:0] node7134;
	wire [4-1:0] node7136;
	wire [4-1:0] node7137;
	wire [4-1:0] node7141;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7147;
	wire [4-1:0] node7149;
	wire [4-1:0] node7150;
	wire [4-1:0] node7153;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7162;
	wire [4-1:0] node7163;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7175;
	wire [4-1:0] node7179;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7185;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7196;
	wire [4-1:0] node7197;
	wire [4-1:0] node7198;
	wire [4-1:0] node7199;
	wire [4-1:0] node7200;
	wire [4-1:0] node7203;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7208;
	wire [4-1:0] node7209;
	wire [4-1:0] node7213;
	wire [4-1:0] node7214;
	wire [4-1:0] node7217;
	wire [4-1:0] node7220;
	wire [4-1:0] node7221;
	wire [4-1:0] node7222;
	wire [4-1:0] node7225;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7232;
	wire [4-1:0] node7235;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7252;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7260;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7277;
	wire [4-1:0] node7278;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7284;
	wire [4-1:0] node7287;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7293;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7299;
	wire [4-1:0] node7300;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7308;
	wire [4-1:0] node7311;
	wire [4-1:0] node7312;
	wire [4-1:0] node7315;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7320;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7329;
	wire [4-1:0] node7330;
	wire [4-1:0] node7331;
	wire [4-1:0] node7332;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7338;
	wire [4-1:0] node7339;
	wire [4-1:0] node7343;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7348;
	wire [4-1:0] node7351;
	wire [4-1:0] node7353;
	wire [4-1:0] node7356;
	wire [4-1:0] node7357;
	wire [4-1:0] node7359;
	wire [4-1:0] node7361;
	wire [4-1:0] node7364;
	wire [4-1:0] node7365;
	wire [4-1:0] node7366;
	wire [4-1:0] node7369;
	wire [4-1:0] node7372;
	wire [4-1:0] node7373;
	wire [4-1:0] node7377;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7383;
	wire [4-1:0] node7385;
	wire [4-1:0] node7388;
	wire [4-1:0] node7390;
	wire [4-1:0] node7392;
	wire [4-1:0] node7395;
	wire [4-1:0] node7396;
	wire [4-1:0] node7397;
	wire [4-1:0] node7401;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7407;
	wire [4-1:0] node7410;
	wire [4-1:0] node7411;
	wire [4-1:0] node7412;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7417;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7424;
	wire [4-1:0] node7427;
	wire [4-1:0] node7428;
	wire [4-1:0] node7429;
	wire [4-1:0] node7432;
	wire [4-1:0] node7435;
	wire [4-1:0] node7436;
	wire [4-1:0] node7438;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7446;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7452;
	wire [4-1:0] node7455;
	wire [4-1:0] node7456;
	wire [4-1:0] node7457;
	wire [4-1:0] node7461;
	wire [4-1:0] node7463;
	wire [4-1:0] node7466;
	wire [4-1:0] node7467;
	wire [4-1:0] node7468;
	wire [4-1:0] node7469;
	wire [4-1:0] node7473;
	wire [4-1:0] node7476;
	wire [4-1:0] node7477;
	wire [4-1:0] node7480;
	wire [4-1:0] node7481;
	wire [4-1:0] node7484;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7496;
	wire [4-1:0] node7497;
	wire [4-1:0] node7499;
	wire [4-1:0] node7502;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7508;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7514;
	wire [4-1:0] node7517;
	wire [4-1:0] node7519;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7528;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7541;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7553;
	wire [4-1:0] node7556;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7561;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7569;
	wire [4-1:0] node7572;
	wire [4-1:0] node7573;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7584;
	wire [4-1:0] node7585;
	wire [4-1:0] node7586;
	wire [4-1:0] node7590;
	wire [4-1:0] node7593;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7603;
	wire [4-1:0] node7604;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7612;
	wire [4-1:0] node7615;
	wire [4-1:0] node7616;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7621;
	wire [4-1:0] node7625;
	wire [4-1:0] node7627;
	wire [4-1:0] node7628;
	wire [4-1:0] node7631;
	wire [4-1:0] node7634;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7640;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7648;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7653;
	wire [4-1:0] node7654;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7663;
	wire [4-1:0] node7666;
	wire [4-1:0] node7669;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7672;
	wire [4-1:0] node7674;
	wire [4-1:0] node7677;
	wire [4-1:0] node7678;
	wire [4-1:0] node7681;
	wire [4-1:0] node7684;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7689;
	wire [4-1:0] node7692;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7703;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7711;
	wire [4-1:0] node7714;
	wire [4-1:0] node7717;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7723;
	wire [4-1:0] node7726;
	wire [4-1:0] node7727;
	wire [4-1:0] node7728;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7741;
	wire [4-1:0] node7746;
	wire [4-1:0] node7747;
	wire [4-1:0] node7750;
	wire [4-1:0] node7753;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7756;
	wire [4-1:0] node7758;
	wire [4-1:0] node7762;
	wire [4-1:0] node7763;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7772;
	wire [4-1:0] node7775;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7783;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7809;
	wire [4-1:0] node7812;
	wire [4-1:0] node7815;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7818;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7823;
	wire [4-1:0] node7826;
	wire [4-1:0] node7827;
	wire [4-1:0] node7831;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7836;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7843;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7849;
	wire [4-1:0] node7852;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7859;
	wire [4-1:0] node7862;
	wire [4-1:0] node7863;
	wire [4-1:0] node7864;
	wire [4-1:0] node7867;
	wire [4-1:0] node7868;
	wire [4-1:0] node7871;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7876;
	wire [4-1:0] node7880;
	wire [4-1:0] node7883;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7887;
	wire [4-1:0] node7891;
	wire [4-1:0] node7893;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7899;
	wire [4-1:0] node7902;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7914;
	wire [4-1:0] node7915;
	wire [4-1:0] node7916;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7924;
	wire [4-1:0] node7927;
	wire [4-1:0] node7928;
	wire [4-1:0] node7932;
	wire [4-1:0] node7933;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7937;
	wire [4-1:0] node7938;
	wire [4-1:0] node7941;
	wire [4-1:0] node7943;
	wire [4-1:0] node7946;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7950;
	wire [4-1:0] node7953;
	wire [4-1:0] node7954;
	wire [4-1:0] node7957;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7967;
	wire [4-1:0] node7968;
	wire [4-1:0] node7970;
	wire [4-1:0] node7974;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7979;
	wire [4-1:0] node7982;
	wire [4-1:0] node7983;
	wire [4-1:0] node7986;
	wire [4-1:0] node7989;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7993;
	wire [4-1:0] node7996;
	wire [4-1:0] node7997;
	wire [4-1:0] node8000;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8005;
	wire [4-1:0] node8008;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8019;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8026;
	wire [4-1:0] node8027;
	wire [4-1:0] node8030;
	wire [4-1:0] node8033;
	wire [4-1:0] node8034;
	wire [4-1:0] node8036;
	wire [4-1:0] node8039;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8056;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8061;
	wire [4-1:0] node8064;
	wire [4-1:0] node8067;
	wire [4-1:0] node8068;
	wire [4-1:0] node8072;
	wire [4-1:0] node8075;
	wire [4-1:0] node8076;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8086;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8094;
	wire [4-1:0] node8095;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8101;
	wire [4-1:0] node8104;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8110;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8115;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8122;
	wire [4-1:0] node8123;
	wire [4-1:0] node8125;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8132;
	wire [4-1:0] node8135;
	wire [4-1:0] node8138;
	wire [4-1:0] node8140;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8146;
	wire [4-1:0] node8149;
	wire [4-1:0] node8151;
	wire [4-1:0] node8154;
	wire [4-1:0] node8155;
	wire [4-1:0] node8156;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8162;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8170;
	wire [4-1:0] node8171;
	wire [4-1:0] node8172;
	wire [4-1:0] node8176;
	wire [4-1:0] node8177;
	wire [4-1:0] node8180;
	wire [4-1:0] node8183;
	wire [4-1:0] node8184;
	wire [4-1:0] node8185;
	wire [4-1:0] node8188;
	wire [4-1:0] node8191;
	wire [4-1:0] node8192;
	wire [4-1:0] node8196;
	wire [4-1:0] node8197;
	wire [4-1:0] node8198;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8209;
	wire [4-1:0] node8210;
	wire [4-1:0] node8211;
	wire [4-1:0] node8214;
	wire [4-1:0] node8218;
	wire [4-1:0] node8219;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8224;
	wire [4-1:0] node8228;
	wire [4-1:0] node8230;
	wire [4-1:0] node8231;
	wire [4-1:0] node8235;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8242;
	wire [4-1:0] node8243;
	wire [4-1:0] node8246;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8251;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8268;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8276;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8283;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8290;
	wire [4-1:0] node8293;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8304;
	wire [4-1:0] node8307;
	wire [4-1:0] node8308;
	wire [4-1:0] node8309;
	wire [4-1:0] node8312;
	wire [4-1:0] node8313;
	wire [4-1:0] node8316;
	wire [4-1:0] node8318;
	wire [4-1:0] node8321;
	wire [4-1:0] node8324;
	wire [4-1:0] node8325;
	wire [4-1:0] node8326;
	wire [4-1:0] node8327;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8335;
	wire [4-1:0] node8336;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8345;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8351;
	wire [4-1:0] node8354;
	wire [4-1:0] node8355;
	wire [4-1:0] node8356;
	wire [4-1:0] node8360;
	wire [4-1:0] node8362;
	wire [4-1:0] node8365;
	wire [4-1:0] node8366;
	wire [4-1:0] node8367;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8373;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8379;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8386;
	wire [4-1:0] node8389;
	wire [4-1:0] node8390;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8397;
	wire [4-1:0] node8399;
	wire [4-1:0] node8401;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8410;
	wire [4-1:0] node8413;
	wire [4-1:0] node8415;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8421;
	wire [4-1:0] node8424;
	wire [4-1:0] node8425;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8434;
	wire [4-1:0] node8435;
	wire [4-1:0] node8436;
	wire [4-1:0] node8439;
	wire [4-1:0] node8441;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8447;
	wire [4-1:0] node8451;
	wire [4-1:0] node8452;
	wire [4-1:0] node8453;
	wire [4-1:0] node8454;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8460;
	wire [4-1:0] node8461;
	wire [4-1:0] node8462;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8470;
	wire [4-1:0] node8473;
	wire [4-1:0] node8476;
	wire [4-1:0] node8477;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8482;
	wire [4-1:0] node8486;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8490;
	wire [4-1:0] node8494;
	wire [4-1:0] node8495;
	wire [4-1:0] node8496;
	wire [4-1:0] node8501;
	wire [4-1:0] node8502;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8507;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8515;
	wire [4-1:0] node8516;
	wire [4-1:0] node8517;
	wire [4-1:0] node8521;
	wire [4-1:0] node8523;
	wire [4-1:0] node8526;
	wire [4-1:0] node8527;
	wire [4-1:0] node8529;
	wire [4-1:0] node8532;
	wire [4-1:0] node8534;
	wire [4-1:0] node8536;
	wire [4-1:0] node8539;
	wire [4-1:0] node8540;
	wire [4-1:0] node8541;
	wire [4-1:0] node8542;
	wire [4-1:0] node8543;
	wire [4-1:0] node8546;
	wire [4-1:0] node8550;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8556;
	wire [4-1:0] node8559;
	wire [4-1:0] node8560;
	wire [4-1:0] node8564;
	wire [4-1:0] node8565;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8571;
	wire [4-1:0] node8574;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8584;
	wire [4-1:0] node8587;
	wire [4-1:0] node8588;
	wire [4-1:0] node8591;
	wire [4-1:0] node8594;
	wire [4-1:0] node8595;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8606;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8614;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8629;
	wire [4-1:0] node8631;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8639;
	wire [4-1:0] node8640;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8648;
	wire [4-1:0] node8649;
	wire [4-1:0] node8652;
	wire [4-1:0] node8654;
	wire [4-1:0] node8657;
	wire [4-1:0] node8659;
	wire [4-1:0] node8660;
	wire [4-1:0] node8661;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8670;
	wire [4-1:0] node8671;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8676;
	wire [4-1:0] node8679;
	wire [4-1:0] node8681;
	wire [4-1:0] node8683;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8690;
	wire [4-1:0] node8691;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8700;
	wire [4-1:0] node8704;
	wire [4-1:0] node8705;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8713;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8724;
	wire [4-1:0] node8725;
	wire [4-1:0] node8726;
	wire [4-1:0] node8727;
	wire [4-1:0] node8729;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8736;
	wire [4-1:0] node8740;
	wire [4-1:0] node8741;
	wire [4-1:0] node8745;
	wire [4-1:0] node8746;
	wire [4-1:0] node8748;
	wire [4-1:0] node8749;
	wire [4-1:0] node8753;
	wire [4-1:0] node8755;
	wire [4-1:0] node8756;
	wire [4-1:0] node8760;
	wire [4-1:0] node8761;
	wire [4-1:0] node8762;
	wire [4-1:0] node8764;
	wire [4-1:0] node8765;
	wire [4-1:0] node8769;
	wire [4-1:0] node8770;
	wire [4-1:0] node8774;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8778;
	wire [4-1:0] node8781;
	wire [4-1:0] node8784;
	wire [4-1:0] node8785;
	wire [4-1:0] node8789;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8795;
	wire [4-1:0] node8798;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8807;
	wire [4-1:0] node8809;
	wire [4-1:0] node8812;
	wire [4-1:0] node8813;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8816;
	wire [4-1:0] node8821;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8835;
	wire [4-1:0] node8838;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8845;
	wire [4-1:0] node8846;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8852;
	wire [4-1:0] node8855;
	wire [4-1:0] node8857;
	wire [4-1:0] node8860;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8866;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8873;
	wire [4-1:0] node8875;
	wire [4-1:0] node8879;
	wire [4-1:0] node8880;
	wire [4-1:0] node8881;
	wire [4-1:0] node8883;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8894;
	wire [4-1:0] node8896;
	wire [4-1:0] node8900;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8907;
	wire [4-1:0] node8908;
	wire [4-1:0] node8911;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8928;
	wire [4-1:0] node8932;
	wire [4-1:0] node8933;
	wire [4-1:0] node8934;
	wire [4-1:0] node8938;
	wire [4-1:0] node8940;
	wire [4-1:0] node8943;
	wire [4-1:0] node8944;
	wire [4-1:0] node8946;
	wire [4-1:0] node8949;
	wire [4-1:0] node8950;
	wire [4-1:0] node8951;
	wire [4-1:0] node8954;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8961;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8971;
	wire [4-1:0] node8974;
	wire [4-1:0] node8976;
	wire [4-1:0] node8977;
	wire [4-1:0] node8980;
	wire [4-1:0] node8983;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8987;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8994;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node9002;
	wire [4-1:0] node9003;
	wire [4-1:0] node9005;
	wire [4-1:0] node9006;
	wire [4-1:0] node9007;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9016;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9021;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9027;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9034;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9043;
	wire [4-1:0] node9044;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9059;
	wire [4-1:0] node9062;
	wire [4-1:0] node9063;
	wire [4-1:0] node9066;
	wire [4-1:0] node9069;
	wire [4-1:0] node9070;
	wire [4-1:0] node9071;
	wire [4-1:0] node9072;
	wire [4-1:0] node9075;
	wire [4-1:0] node9078;
	wire [4-1:0] node9079;
	wire [4-1:0] node9083;
	wire [4-1:0] node9084;
	wire [4-1:0] node9085;
	wire [4-1:0] node9089;
	wire [4-1:0] node9090;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9099;
	wire [4-1:0] node9102;
	wire [4-1:0] node9104;
	wire [4-1:0] node9107;
	wire [4-1:0] node9108;
	wire [4-1:0] node9110;
	wire [4-1:0] node9112;
	wire [4-1:0] node9115;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9131;
	wire [4-1:0] node9135;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9148;
	wire [4-1:0] node9152;
	wire [4-1:0] node9153;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9165;
	wire [4-1:0] node9166;
	wire [4-1:0] node9167;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9176;
	wire [4-1:0] node9179;
	wire [4-1:0] node9180;
	wire [4-1:0] node9181;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9189;
	wire [4-1:0] node9192;
	wire [4-1:0] node9193;
	wire [4-1:0] node9195;
	wire [4-1:0] node9197;
	wire [4-1:0] node9200;
	wire [4-1:0] node9201;
	wire [4-1:0] node9203;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9209;
	wire [4-1:0] node9212;
	wire [4-1:0] node9215;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9221;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9228;
	wire [4-1:0] node9231;
	wire [4-1:0] node9233;
	wire [4-1:0] node9235;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9242;
	wire [4-1:0] node9245;
	wire [4-1:0] node9246;
	wire [4-1:0] node9249;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9255;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9262;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9268;
	wire [4-1:0] node9269;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9277;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9284;
	wire [4-1:0] node9286;
	wire [4-1:0] node9289;
	wire [4-1:0] node9290;
	wire [4-1:0] node9291;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9300;
	wire [4-1:0] node9301;
	wire [4-1:0] node9302;
	wire [4-1:0] node9303;
	wire [4-1:0] node9304;
	wire [4-1:0] node9305;
	wire [4-1:0] node9306;
	wire [4-1:0] node9307;
	wire [4-1:0] node9310;
	wire [4-1:0] node9312;
	wire [4-1:0] node9315;
	wire [4-1:0] node9316;
	wire [4-1:0] node9318;
	wire [4-1:0] node9319;
	wire [4-1:0] node9323;
	wire [4-1:0] node9326;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9329;
	wire [4-1:0] node9330;
	wire [4-1:0] node9334;
	wire [4-1:0] node9336;
	wire [4-1:0] node9339;
	wire [4-1:0] node9340;
	wire [4-1:0] node9343;
	wire [4-1:0] node9345;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9351;
	wire [4-1:0] node9352;
	wire [4-1:0] node9356;
	wire [4-1:0] node9357;
	wire [4-1:0] node9361;
	wire [4-1:0] node9362;
	wire [4-1:0] node9363;
	wire [4-1:0] node9364;
	wire [4-1:0] node9367;
	wire [4-1:0] node9369;
	wire [4-1:0] node9372;
	wire [4-1:0] node9373;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9386;
	wire [4-1:0] node9389;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9397;
	wire [4-1:0] node9400;
	wire [4-1:0] node9403;
	wire [4-1:0] node9404;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9414;
	wire [4-1:0] node9415;
	wire [4-1:0] node9416;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9421;
	wire [4-1:0] node9423;
	wire [4-1:0] node9426;
	wire [4-1:0] node9427;
	wire [4-1:0] node9429;
	wire [4-1:0] node9432;
	wire [4-1:0] node9433;
	wire [4-1:0] node9436;
	wire [4-1:0] node9439;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9447;
	wire [4-1:0] node9449;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9455;
	wire [4-1:0] node9458;
	wire [4-1:0] node9461;
	wire [4-1:0] node9462;
	wire [4-1:0] node9464;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9469;
	wire [4-1:0] node9473;
	wire [4-1:0] node9474;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9480;
	wire [4-1:0] node9481;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9486;
	wire [4-1:0] node9489;
	wire [4-1:0] node9492;
	wire [4-1:0] node9493;
	wire [4-1:0] node9496;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9511;
	wire [4-1:0] node9512;
	wire [4-1:0] node9514;
	wire [4-1:0] node9518;
	wire [4-1:0] node9519;
	wire [4-1:0] node9520;
	wire [4-1:0] node9521;
	wire [4-1:0] node9522;
	wire [4-1:0] node9525;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9532;
	wire [4-1:0] node9535;
	wire [4-1:0] node9538;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9544;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9551;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9557;
	wire [4-1:0] node9558;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9567;
	wire [4-1:0] node9568;
	wire [4-1:0] node9569;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9576;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9582;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9591;
	wire [4-1:0] node9593;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9601;
	wire [4-1:0] node9602;
	wire [4-1:0] node9603;
	wire [4-1:0] node9606;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9615;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9624;
	wire [4-1:0] node9627;
	wire [4-1:0] node9628;
	wire [4-1:0] node9630;
	wire [4-1:0] node9633;
	wire [4-1:0] node9634;
	wire [4-1:0] node9635;
	wire [4-1:0] node9639;
	wire [4-1:0] node9640;
	wire [4-1:0] node9643;
	wire [4-1:0] node9646;
	wire [4-1:0] node9647;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9650;
	wire [4-1:0] node9655;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9660;
	wire [4-1:0] node9663;
	wire [4-1:0] node9664;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9671;
	wire [4-1:0] node9673;
	wire [4-1:0] node9676;
	wire [4-1:0] node9678;
	wire [4-1:0] node9679;
	wire [4-1:0] node9682;
	wire [4-1:0] node9685;
	wire [4-1:0] node9686;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9689;
	wire [4-1:0] node9690;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9711;
	wire [4-1:0] node9714;
	wire [4-1:0] node9717;
	wire [4-1:0] node9720;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9723;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9731;
	wire [4-1:0] node9734;
	wire [4-1:0] node9735;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9742;
	wire [4-1:0] node9745;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9750;
	wire [4-1:0] node9753;
	wire [4-1:0] node9754;
	wire [4-1:0] node9757;
	wire [4-1:0] node9760;
	wire [4-1:0] node9762;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9771;
	wire [4-1:0] node9774;
	wire [4-1:0] node9775;
	wire [4-1:0] node9778;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9786;
	wire [4-1:0] node9789;
	wire [4-1:0] node9790;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9801;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9805;
	wire [4-1:0] node9807;
	wire [4-1:0] node9812;
	wire [4-1:0] node9813;
	wire [4-1:0] node9814;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9820;
	wire [4-1:0] node9825;
	wire [4-1:0] node9826;
	wire [4-1:0] node9828;
	wire [4-1:0] node9829;
	wire [4-1:0] node9832;
	wire [4-1:0] node9835;
	wire [4-1:0] node9836;
	wire [4-1:0] node9837;
	wire [4-1:0] node9840;
	wire [4-1:0] node9842;
	wire [4-1:0] node9845;
	wire [4-1:0] node9848;
	wire [4-1:0] node9849;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9853;
	wire [4-1:0] node9856;
	wire [4-1:0] node9857;
	wire [4-1:0] node9858;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9867;
	wire [4-1:0] node9868;
	wire [4-1:0] node9869;
	wire [4-1:0] node9871;
	wire [4-1:0] node9874;
	wire [4-1:0] node9875;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9882;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9891;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9897;
	wire [4-1:0] node9898;
	wire [4-1:0] node9902;
	wire [4-1:0] node9903;
	wire [4-1:0] node9904;
	wire [4-1:0] node9909;
	wire [4-1:0] node9910;
	wire [4-1:0] node9911;
	wire [4-1:0] node9912;
	wire [4-1:0] node9913;
	wire [4-1:0] node9915;
	wire [4-1:0] node9918;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9924;
	wire [4-1:0] node9927;
	wire [4-1:0] node9928;
	wire [4-1:0] node9929;
	wire [4-1:0] node9933;
	wire [4-1:0] node9935;
	wire [4-1:0] node9938;
	wire [4-1:0] node9939;
	wire [4-1:0] node9940;
	wire [4-1:0] node9942;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9948;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9956;
	wire [4-1:0] node9957;
	wire [4-1:0] node9959;
	wire [4-1:0] node9960;
	wire [4-1:0] node9964;
	wire [4-1:0] node9965;
	wire [4-1:0] node9968;
	wire [4-1:0] node9971;
	wire [4-1:0] node9972;
	wire [4-1:0] node9973;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9979;
	wire [4-1:0] node9981;
	wire [4-1:0] node9984;
	wire [4-1:0] node9985;
	wire [4-1:0] node9986;
	wire [4-1:0] node9990;
	wire [4-1:0] node9991;
	wire [4-1:0] node9995;
	wire [4-1:0] node9996;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10003;
	wire [4-1:0] node10004;
	wire [4-1:0] node10005;
	wire [4-1:0] node10007;
	wire [4-1:0] node10010;
	wire [4-1:0] node10011;
	wire [4-1:0] node10014;
	wire [4-1:0] node10017;
	wire [4-1:0] node10018;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10025;
	wire [4-1:0] node10026;
	wire [4-1:0] node10027;
	wire [4-1:0] node10028;
	wire [4-1:0] node10030;
	wire [4-1:0] node10032;
	wire [4-1:0] node10034;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10045;
	wire [4-1:0] node10047;
	wire [4-1:0] node10050;
	wire [4-1:0] node10051;
	wire [4-1:0] node10053;
	wire [4-1:0] node10056;
	wire [4-1:0] node10057;
	wire [4-1:0] node10058;
	wire [4-1:0] node10060;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10069;
	wire [4-1:0] node10072;
	wire [4-1:0] node10074;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10080;
	wire [4-1:0] node10081;
	wire [4-1:0] node10084;
	wire [4-1:0] node10086;
	wire [4-1:0] node10089;
	wire [4-1:0] node10090;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10097;
	wire [4-1:0] node10100;
	wire [4-1:0] node10101;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10114;
	wire [4-1:0] node10117;
	wire [4-1:0] node10120;
	wire [4-1:0] node10121;
	wire [4-1:0] node10125;
	wire [4-1:0] node10126;
	wire [4-1:0] node10127;
	wire [4-1:0] node10129;
	wire [4-1:0] node10132;
	wire [4-1:0] node10134;
	wire [4-1:0] node10137;
	wire [4-1:0] node10138;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10145;
	wire [4-1:0] node10146;
	wire [4-1:0] node10148;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10155;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10168;
	wire [4-1:0] node10169;
	wire [4-1:0] node10172;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10179;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10191;
	wire [4-1:0] node10192;
	wire [4-1:0] node10196;
	wire [4-1:0] node10197;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10202;
	wire [4-1:0] node10205;
	wire [4-1:0] node10209;
	wire [4-1:0] node10210;
	wire [4-1:0] node10211;
	wire [4-1:0] node10214;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10220;
	wire [4-1:0] node10223;
	wire [4-1:0] node10225;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10235;
	wire [4-1:0] node10238;
	wire [4-1:0] node10239;
	wire [4-1:0] node10240;
	wire [4-1:0] node10244;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10251;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10257;
	wire [4-1:0] node10259;
	wire [4-1:0] node10262;
	wire [4-1:0] node10263;
	wire [4-1:0] node10264;
	wire [4-1:0] node10268;
	wire [4-1:0] node10271;
	wire [4-1:0] node10272;
	wire [4-1:0] node10274;
	wire [4-1:0] node10275;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10284;
	wire [4-1:0] node10285;
	wire [4-1:0] node10286;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10296;
	wire [4-1:0] node10298;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10309;
	wire [4-1:0] node10312;
	wire [4-1:0] node10315;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10324;
	wire [4-1:0] node10325;
	wire [4-1:0] node10326;
	wire [4-1:0] node10327;
	wire [4-1:0] node10331;
	wire [4-1:0] node10334;
	wire [4-1:0] node10335;
	wire [4-1:0] node10338;
	wire [4-1:0] node10341;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10357;
	wire [4-1:0] node10358;
	wire [4-1:0] node10359;
	wire [4-1:0] node10362;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10369;
	wire [4-1:0] node10370;
	wire [4-1:0] node10372;
	wire [4-1:0] node10374;
	wire [4-1:0] node10378;
	wire [4-1:0] node10379;
	wire [4-1:0] node10381;
	wire [4-1:0] node10384;
	wire [4-1:0] node10386;
	wire [4-1:0] node10389;
	wire [4-1:0] node10390;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10394;
	wire [4-1:0] node10397;
	wire [4-1:0] node10398;
	wire [4-1:0] node10401;
	wire [4-1:0] node10404;
	wire [4-1:0] node10405;
	wire [4-1:0] node10406;
	wire [4-1:0] node10411;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10416;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10422;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10431;
	wire [4-1:0] node10434;
	wire [4-1:0] node10438;
	wire [4-1:0] node10440;
	wire [4-1:0] node10442;
	wire [4-1:0] node10445;
	wire [4-1:0] node10446;
	wire [4-1:0] node10447;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10459;
	wire [4-1:0] node10461;
	wire [4-1:0] node10464;
	wire [4-1:0] node10465;
	wire [4-1:0] node10466;
	wire [4-1:0] node10468;
	wire [4-1:0] node10470;
	wire [4-1:0] node10473;
	wire [4-1:0] node10474;
	wire [4-1:0] node10477;
	wire [4-1:0] node10478;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10484;
	wire [4-1:0] node10487;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10501;
	wire [4-1:0] node10504;
	wire [4-1:0] node10505;
	wire [4-1:0] node10506;
	wire [4-1:0] node10509;
	wire [4-1:0] node10511;
	wire [4-1:0] node10514;
	wire [4-1:0] node10515;
	wire [4-1:0] node10519;
	wire [4-1:0] node10520;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10539;
	wire [4-1:0] node10540;
	wire [4-1:0] node10544;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10549;
	wire [4-1:0] node10554;
	wire [4-1:0] node10555;
	wire [4-1:0] node10556;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10563;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10570;
	wire [4-1:0] node10573;
	wire [4-1:0] node10574;
	wire [4-1:0] node10576;
	wire [4-1:0] node10579;
	wire [4-1:0] node10580;
	wire [4-1:0] node10581;
	wire [4-1:0] node10584;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10591;
	wire [4-1:0] node10594;
	wire [4-1:0] node10597;
	wire [4-1:0] node10598;
	wire [4-1:0] node10601;
	wire [4-1:0] node10602;
	wire [4-1:0] node10605;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10612;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10625;
	wire [4-1:0] node10626;
	wire [4-1:0] node10627;
	wire [4-1:0] node10629;
	wire [4-1:0] node10632;
	wire [4-1:0] node10634;
	wire [4-1:0] node10635;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10646;
	wire [4-1:0] node10647;
	wire [4-1:0] node10650;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10659;
	wire [4-1:0] node10662;
	wire [4-1:0] node10663;
	wire [4-1:0] node10664;
	wire [4-1:0] node10666;
	wire [4-1:0] node10667;
	wire [4-1:0] node10670;
	wire [4-1:0] node10673;
	wire [4-1:0] node10674;
	wire [4-1:0] node10675;
	wire [4-1:0] node10679;
	wire [4-1:0] node10680;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10686;
	wire [4-1:0] node10688;
	wire [4-1:0] node10691;
	wire [4-1:0] node10695;
	wire [4-1:0] node10696;
	wire [4-1:0] node10697;
	wire [4-1:0] node10698;
	wire [4-1:0] node10699;
	wire [4-1:0] node10702;
	wire [4-1:0] node10704;
	wire [4-1:0] node10707;
	wire [4-1:0] node10708;
	wire [4-1:0] node10712;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10724;
	wire [4-1:0] node10726;
	wire [4-1:0] node10729;
	wire [4-1:0] node10730;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10733;
	wire [4-1:0] node10736;
	wire [4-1:0] node10739;
	wire [4-1:0] node10741;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10753;
	wire [4-1:0] node10754;
	wire [4-1:0] node10756;
	wire [4-1:0] node10760;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10763;
	wire [4-1:0] node10764;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10769;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10774;
	wire [4-1:0] node10777;
	wire [4-1:0] node10780;
	wire [4-1:0] node10781;
	wire [4-1:0] node10783;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10791;
	wire [4-1:0] node10794;
	wire [4-1:0] node10797;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10804;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10808;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10818;
	wire [4-1:0] node10821;
	wire [4-1:0] node10823;
	wire [4-1:0] node10826;
	wire [4-1:0] node10827;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10832;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10840;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10846;
	wire [4-1:0] node10849;
	wire [4-1:0] node10851;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10857;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10865;
	wire [4-1:0] node10868;
	wire [4-1:0] node10869;
	wire [4-1:0] node10872;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10877;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10890;
	wire [4-1:0] node10893;
	wire [4-1:0] node10895;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10901;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10907;
	wire [4-1:0] node10909;
	wire [4-1:0] node10912;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10917;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10924;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10931;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10939;
	wire [4-1:0] node10940;
	wire [4-1:0] node10944;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10947;
	wire [4-1:0] node10948;
	wire [4-1:0] node10949;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10961;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10968;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10974;
	wire [4-1:0] node10975;
	wire [4-1:0] node10976;
	wire [4-1:0] node10980;
	wire [4-1:0] node10982;
	wire [4-1:0] node10985;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10992;
	wire [4-1:0] node10993;
	wire [4-1:0] node10994;
	wire [4-1:0] node10997;
	wire [4-1:0] node11000;
	wire [4-1:0] node11001;
	wire [4-1:0] node11004;
	wire [4-1:0] node11007;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11010;
	wire [4-1:0] node11012;
	wire [4-1:0] node11013;
	wire [4-1:0] node11016;
	wire [4-1:0] node11019;
	wire [4-1:0] node11021;
	wire [4-1:0] node11022;
	wire [4-1:0] node11026;
	wire [4-1:0] node11027;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11034;
	wire [4-1:0] node11035;
	wire [4-1:0] node11039;
	wire [4-1:0] node11040;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11044;
	wire [4-1:0] node11047;
	wire [4-1:0] node11051;
	wire [4-1:0] node11052;
	wire [4-1:0] node11053;
	wire [4-1:0] node11056;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11063;
	wire [4-1:0] node11064;
	wire [4-1:0] node11065;
	wire [4-1:0] node11067;
	wire [4-1:0] node11070;
	wire [4-1:0] node11071;
	wire [4-1:0] node11075;
	wire [4-1:0] node11076;
	wire [4-1:0] node11079;
	wire [4-1:0] node11082;
	wire [4-1:0] node11083;
	wire [4-1:0] node11085;
	wire [4-1:0] node11087;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11094;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11112;
	wire [4-1:0] node11116;
	wire [4-1:0] node11118;
	wire [4-1:0] node11121;
	wire [4-1:0] node11122;
	wire [4-1:0] node11126;
	wire [4-1:0] node11127;
	wire [4-1:0] node11128;
	wire [4-1:0] node11129;
	wire [4-1:0] node11130;
	wire [4-1:0] node11132;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11139;
	wire [4-1:0] node11142;
	wire [4-1:0] node11145;
	wire [4-1:0] node11146;
	wire [4-1:0] node11148;
	wire [4-1:0] node11149;
	wire [4-1:0] node11154;
	wire [4-1:0] node11155;
	wire [4-1:0] node11156;
	wire [4-1:0] node11158;
	wire [4-1:0] node11160;
	wire [4-1:0] node11163;
	wire [4-1:0] node11165;
	wire [4-1:0] node11168;
	wire [4-1:0] node11169;
	wire [4-1:0] node11171;
	wire [4-1:0] node11173;
	wire [4-1:0] node11176;
	wire [4-1:0] node11177;
	wire [4-1:0] node11178;
	wire [4-1:0] node11183;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11186;
	wire [4-1:0] node11187;
	wire [4-1:0] node11188;
	wire [4-1:0] node11189;
	wire [4-1:0] node11190;
	wire [4-1:0] node11193;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11200;
	wire [4-1:0] node11203;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11206;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11213;
	wire [4-1:0] node11215;
	wire [4-1:0] node11218;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11223;
	wire [4-1:0] node11226;
	wire [4-1:0] node11228;
	wire [4-1:0] node11231;
	wire [4-1:0] node11232;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11237;
	wire [4-1:0] node11242;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11245;
	wire [4-1:0] node11246;
	wire [4-1:0] node11247;
	wire [4-1:0] node11251;
	wire [4-1:0] node11252;
	wire [4-1:0] node11256;
	wire [4-1:0] node11259;
	wire [4-1:0] node11261;
	wire [4-1:0] node11263;
	wire [4-1:0] node11265;
	wire [4-1:0] node11268;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11272;
	wire [4-1:0] node11275;
	wire [4-1:0] node11276;
	wire [4-1:0] node11279;
	wire [4-1:0] node11281;
	wire [4-1:0] node11284;
	wire [4-1:0] node11285;
	wire [4-1:0] node11287;
	wire [4-1:0] node11290;
	wire [4-1:0] node11292;
	wire [4-1:0] node11295;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11299;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11307;
	wire [4-1:0] node11308;
	wire [4-1:0] node11310;
	wire [4-1:0] node11313;
	wire [4-1:0] node11315;
	wire [4-1:0] node11318;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11323;
	wire [4-1:0] node11326;
	wire [4-1:0] node11327;
	wire [4-1:0] node11328;
	wire [4-1:0] node11331;
	wire [4-1:0] node11335;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11338;
	wire [4-1:0] node11339;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11347;
	wire [4-1:0] node11348;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11356;
	wire [4-1:0] node11357;
	wire [4-1:0] node11359;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11370;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11382;
	wire [4-1:0] node11385;
	wire [4-1:0] node11386;
	wire [4-1:0] node11389;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11398;
	wire [4-1:0] node11399;
	wire [4-1:0] node11401;
	wire [4-1:0] node11404;
	wire [4-1:0] node11406;
	wire [4-1:0] node11409;
	wire [4-1:0] node11411;
	wire [4-1:0] node11413;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11419;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11425;
	wire [4-1:0] node11428;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11435;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11440;
	wire [4-1:0] node11441;
	wire [4-1:0] node11445;
	wire [4-1:0] node11446;
	wire [4-1:0] node11447;
	wire [4-1:0] node11452;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11457;
	wire [4-1:0] node11460;
	wire [4-1:0] node11462;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11471;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11480;
	wire [4-1:0] node11481;
	wire [4-1:0] node11485;
	wire [4-1:0] node11486;
	wire [4-1:0] node11488;
	wire [4-1:0] node11491;
	wire [4-1:0] node11492;
	wire [4-1:0] node11493;
	wire [4-1:0] node11497;
	wire [4-1:0] node11500;
	wire [4-1:0] node11501;
	wire [4-1:0] node11502;
	wire [4-1:0] node11503;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11506;
	wire [4-1:0] node11509;
	wire [4-1:0] node11512;
	wire [4-1:0] node11514;
	wire [4-1:0] node11517;
	wire [4-1:0] node11518;
	wire [4-1:0] node11520;
	wire [4-1:0] node11523;
	wire [4-1:0] node11524;
	wire [4-1:0] node11527;
	wire [4-1:0] node11530;
	wire [4-1:0] node11531;
	wire [4-1:0] node11532;
	wire [4-1:0] node11534;
	wire [4-1:0] node11538;
	wire [4-1:0] node11540;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11545;
	wire [4-1:0] node11547;
	wire [4-1:0] node11550;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11555;
	wire [4-1:0] node11558;
	wire [4-1:0] node11559;
	wire [4-1:0] node11562;
	wire [4-1:0] node11565;
	wire [4-1:0] node11566;
	wire [4-1:0] node11567;
	wire [4-1:0] node11568;
	wire [4-1:0] node11572;
	wire [4-1:0] node11574;
	wire [4-1:0] node11577;
	wire [4-1:0] node11578;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11585;
	wire [4-1:0] node11586;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11599;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11603;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11611;
	wire [4-1:0] node11613;
	wire [4-1:0] node11616;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11619;
	wire [4-1:0] node11621;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11628;
	wire [4-1:0] node11631;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11637;
	wire [4-1:0] node11640;
	wire [4-1:0] node11642;
	wire [4-1:0] node11644;
	wire [4-1:0] node11647;
	wire [4-1:0] node11648;
	wire [4-1:0] node11649;
	wire [4-1:0] node11650;
	wire [4-1:0] node11651;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11655;
	wire [4-1:0] node11658;
	wire [4-1:0] node11661;
	wire [4-1:0] node11662;
	wire [4-1:0] node11663;
	wire [4-1:0] node11664;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11676;
	wire [4-1:0] node11679;
	wire [4-1:0] node11680;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11686;
	wire [4-1:0] node11688;
	wire [4-1:0] node11691;
	wire [4-1:0] node11694;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11698;
	wire [4-1:0] node11701;
	wire [4-1:0] node11704;
	wire [4-1:0] node11705;
	wire [4-1:0] node11707;
	wire [4-1:0] node11710;
	wire [4-1:0] node11713;
	wire [4-1:0] node11714;
	wire [4-1:0] node11715;
	wire [4-1:0] node11716;
	wire [4-1:0] node11717;
	wire [4-1:0] node11719;
	wire [4-1:0] node11723;
	wire [4-1:0] node11724;
	wire [4-1:0] node11725;
	wire [4-1:0] node11728;
	wire [4-1:0] node11731;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11741;
	wire [4-1:0] node11744;
	wire [4-1:0] node11745;
	wire [4-1:0] node11746;
	wire [4-1:0] node11749;
	wire [4-1:0] node11752;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11779;
	wire [4-1:0] node11781;
	wire [4-1:0] node11783;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11791;
	wire [4-1:0] node11794;
	wire [4-1:0] node11796;
	wire [4-1:0] node11799;
	wire [4-1:0] node11800;
	wire [4-1:0] node11801;
	wire [4-1:0] node11806;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11811;
	wire [4-1:0] node11812;
	wire [4-1:0] node11815;
	wire [4-1:0] node11818;
	wire [4-1:0] node11819;
	wire [4-1:0] node11820;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11827;
	wire [4-1:0] node11828;
	wire [4-1:0] node11829;
	wire [4-1:0] node11834;
	wire [4-1:0] node11836;
	wire [4-1:0] node11838;
	wire [4-1:0] node11841;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11847;
	wire [4-1:0] node11848;
	wire [4-1:0] node11851;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11863;
	wire [4-1:0] node11866;
	wire [4-1:0] node11867;
	wire [4-1:0] node11870;
	wire [4-1:0] node11872;
	wire [4-1:0] node11875;
	wire [4-1:0] node11876;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11883;
	wire [4-1:0] node11884;
	wire [4-1:0] node11887;
	wire [4-1:0] node11889;
	wire [4-1:0] node11892;
	wire [4-1:0] node11893;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11896;
	wire [4-1:0] node11900;
	wire [4-1:0] node11903;
	wire [4-1:0] node11904;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11915;
	wire [4-1:0] node11916;
	wire [4-1:0] node11917;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11920;
	wire [4-1:0] node11923;
	wire [4-1:0] node11926;
	wire [4-1:0] node11927;
	wire [4-1:0] node11928;
	wire [4-1:0] node11929;
	wire [4-1:0] node11932;
	wire [4-1:0] node11935;
	wire [4-1:0] node11936;
	wire [4-1:0] node11939;
	wire [4-1:0] node11942;
	wire [4-1:0] node11943;
	wire [4-1:0] node11945;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11952;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11957;
	wire [4-1:0] node11958;
	wire [4-1:0] node11961;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11976;
	wire [4-1:0] node11978;
	wire [4-1:0] node11981;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11987;
	wire [4-1:0] node11990;
	wire [4-1:0] node11991;
	wire [4-1:0] node11992;
	wire [4-1:0] node11993;
	wire [4-1:0] node11994;
	wire [4-1:0] node11996;
	wire [4-1:0] node12000;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12013;
	wire [4-1:0] node12017;
	wire [4-1:0] node12018;
	wire [4-1:0] node12022;
	wire [4-1:0] node12023;
	wire [4-1:0] node12024;
	wire [4-1:0] node12025;
	wire [4-1:0] node12029;
	wire [4-1:0] node12031;
	wire [4-1:0] node12034;
	wire [4-1:0] node12035;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12041;
	wire [4-1:0] node12044;
	wire [4-1:0] node12045;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12052;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12058;
	wire [4-1:0] node12061;
	wire [4-1:0] node12063;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12076;
	wire [4-1:0] node12079;
	wire [4-1:0] node12080;
	wire [4-1:0] node12081;
	wire [4-1:0] node12082;
	wire [4-1:0] node12086;
	wire [4-1:0] node12087;
	wire [4-1:0] node12091;
	wire [4-1:0] node12092;
	wire [4-1:0] node12095;
	wire [4-1:0] node12096;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12103;
	wire [4-1:0] node12105;
	wire [4-1:0] node12108;
	wire [4-1:0] node12109;
	wire [4-1:0] node12112;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12119;
	wire [4-1:0] node12122;
	wire [4-1:0] node12123;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12132;
	wire [4-1:0] node12135;
	wire [4-1:0] node12136;
	wire [4-1:0] node12137;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12145;
	wire [4-1:0] node12147;
	wire [4-1:0] node12150;
	wire [4-1:0] node12152;
	wire [4-1:0] node12155;
	wire [4-1:0] node12156;
	wire [4-1:0] node12157;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12164;
	wire [4-1:0] node12165;
	wire [4-1:0] node12167;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12173;
	wire [4-1:0] node12177;
	wire [4-1:0] node12178;
	wire [4-1:0] node12179;
	wire [4-1:0] node12183;
	wire [4-1:0] node12186;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12190;
	wire [4-1:0] node12191;
	wire [4-1:0] node12192;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12196;
	wire [4-1:0] node12197;
	wire [4-1:0] node12200;
	wire [4-1:0] node12203;
	wire [4-1:0] node12205;
	wire [4-1:0] node12208;
	wire [4-1:0] node12209;
	wire [4-1:0] node12210;
	wire [4-1:0] node12212;
	wire [4-1:0] node12215;
	wire [4-1:0] node12216;
	wire [4-1:0] node12219;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12226;
	wire [4-1:0] node12229;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12232;
	wire [4-1:0] node12233;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12241;
	wire [4-1:0] node12244;
	wire [4-1:0] node12245;
	wire [4-1:0] node12246;
	wire [4-1:0] node12249;
	wire [4-1:0] node12252;
	wire [4-1:0] node12254;
	wire [4-1:0] node12257;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12261;
	wire [4-1:0] node12264;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12271;
	wire [4-1:0] node12274;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12278;
	wire [4-1:0] node12281;
	wire [4-1:0] node12284;
	wire [4-1:0] node12285;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12295;
	wire [4-1:0] node12296;
	wire [4-1:0] node12299;
	wire [4-1:0] node12300;
	wire [4-1:0] node12303;
	wire [4-1:0] node12306;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12314;
	wire [4-1:0] node12316;
	wire [4-1:0] node12319;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12324;
	wire [4-1:0] node12327;
	wire [4-1:0] node12329;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12334;
	wire [4-1:0] node12335;
	wire [4-1:0] node12337;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12348;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12355;
	wire [4-1:0] node12356;
	wire [4-1:0] node12360;
	wire [4-1:0] node12361;
	wire [4-1:0] node12362;
	wire [4-1:0] node12363;
	wire [4-1:0] node12366;
	wire [4-1:0] node12369;
	wire [4-1:0] node12370;
	wire [4-1:0] node12374;
	wire [4-1:0] node12375;
	wire [4-1:0] node12376;
	wire [4-1:0] node12379;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12386;
	wire [4-1:0] node12389;
	wire [4-1:0] node12390;
	wire [4-1:0] node12391;
	wire [4-1:0] node12392;
	wire [4-1:0] node12393;
	wire [4-1:0] node12396;
	wire [4-1:0] node12397;
	wire [4-1:0] node12399;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12409;
	wire [4-1:0] node12410;
	wire [4-1:0] node12413;
	wire [4-1:0] node12416;
	wire [4-1:0] node12417;
	wire [4-1:0] node12420;
	wire [4-1:0] node12423;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12433;
	wire [4-1:0] node12434;
	wire [4-1:0] node12438;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12445;
	wire [4-1:0] node12448;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12454;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12459;
	wire [4-1:0] node12463;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12472;
	wire [4-1:0] node12473;
	wire [4-1:0] node12476;
	wire [4-1:0] node12479;
	wire [4-1:0] node12481;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12490;
	wire [4-1:0] node12491;
	wire [4-1:0] node12492;
	wire [4-1:0] node12496;
	wire [4-1:0] node12497;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12504;
	wire [4-1:0] node12505;
	wire [4-1:0] node12507;
	wire [4-1:0] node12510;
	wire [4-1:0] node12513;
	wire [4-1:0] node12515;
	wire [4-1:0] node12517;
	wire [4-1:0] node12520;
	wire [4-1:0] node12521;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12527;
	wire [4-1:0] node12530;
	wire [4-1:0] node12531;
	wire [4-1:0] node12532;
	wire [4-1:0] node12533;
	wire [4-1:0] node12536;
	wire [4-1:0] node12539;
	wire [4-1:0] node12541;
	wire [4-1:0] node12544;
	wire [4-1:0] node12547;
	wire [4-1:0] node12548;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12551;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12559;
	wire [4-1:0] node12562;
	wire [4-1:0] node12563;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12568;
	wire [4-1:0] node12573;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12579;
	wire [4-1:0] node12582;
	wire [4-1:0] node12583;
	wire [4-1:0] node12586;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12594;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12601;
	wire [4-1:0] node12604;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12608;
	wire [4-1:0] node12609;
	wire [4-1:0] node12612;
	wire [4-1:0] node12615;
	wire [4-1:0] node12616;
	wire [4-1:0] node12617;
	wire [4-1:0] node12618;
	wire [4-1:0] node12619;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12628;
	wire [4-1:0] node12631;
	wire [4-1:0] node12632;
	wire [4-1:0] node12633;
	wire [4-1:0] node12634;
	wire [4-1:0] node12637;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12645;
	wire [4-1:0] node12647;
	wire [4-1:0] node12650;
	wire [4-1:0] node12651;
	wire [4-1:0] node12654;
	wire [4-1:0] node12657;
	wire [4-1:0] node12658;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12667;
	wire [4-1:0] node12671;
	wire [4-1:0] node12672;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12678;
	wire [4-1:0] node12682;
	wire [4-1:0] node12683;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12689;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12701;
	wire [4-1:0] node12704;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12707;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12730;
	wire [4-1:0] node12732;
	wire [4-1:0] node12733;
	wire [4-1:0] node12736;
	wire [4-1:0] node12739;
	wire [4-1:0] node12740;
	wire [4-1:0] node12744;
	wire [4-1:0] node12745;
	wire [4-1:0] node12746;
	wire [4-1:0] node12747;
	wire [4-1:0] node12750;
	wire [4-1:0] node12754;
	wire [4-1:0] node12755;
	wire [4-1:0] node12757;
	wire [4-1:0] node12760;
	wire [4-1:0] node12762;
	wire [4-1:0] node12765;
	wire [4-1:0] node12766;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12769;
	wire [4-1:0] node12772;
	wire [4-1:0] node12775;
	wire [4-1:0] node12776;
	wire [4-1:0] node12779;
	wire [4-1:0] node12782;
	wire [4-1:0] node12783;
	wire [4-1:0] node12786;
	wire [4-1:0] node12789;
	wire [4-1:0] node12790;
	wire [4-1:0] node12791;
	wire [4-1:0] node12794;
	wire [4-1:0] node12797;
	wire [4-1:0] node12798;
	wire [4-1:0] node12799;
	wire [4-1:0] node12804;
	wire [4-1:0] node12805;
	wire [4-1:0] node12806;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12811;
	wire [4-1:0] node12814;
	wire [4-1:0] node12816;
	wire [4-1:0] node12817;
	wire [4-1:0] node12820;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12827;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12832;
	wire [4-1:0] node12835;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12843;
	wire [4-1:0] node12846;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12856;
	wire [4-1:0] node12858;
	wire [4-1:0] node12861;
	wire [4-1:0] node12863;
	wire [4-1:0] node12866;
	wire [4-1:0] node12867;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12873;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12879;
	wire [4-1:0] node12883;
	wire [4-1:0] node12884;
	wire [4-1:0] node12886;
	wire [4-1:0] node12887;
	wire [4-1:0] node12889;
	wire [4-1:0] node12892;
	wire [4-1:0] node12893;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12899;
	wire [4-1:0] node12901;
	wire [4-1:0] node12905;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12910;
	wire [4-1:0] node12914;
	wire [4-1:0] node12915;
	wire [4-1:0] node12916;
	wire [4-1:0] node12917;
	wire [4-1:0] node12918;
	wire [4-1:0] node12919;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12933;
	wire [4-1:0] node12934;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12948;
	wire [4-1:0] node12952;
	wire [4-1:0] node12953;
	wire [4-1:0] node12954;
	wire [4-1:0] node12955;
	wire [4-1:0] node12957;
	wire [4-1:0] node12960;
	wire [4-1:0] node12962;
	wire [4-1:0] node12963;
	wire [4-1:0] node12967;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12972;
	wire [4-1:0] node12975;
	wire [4-1:0] node12976;
	wire [4-1:0] node12978;
	wire [4-1:0] node12981;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12986;
	wire [4-1:0] node12988;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12996;
	wire [4-1:0] node12997;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13003;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13013;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13018;
	wire [4-1:0] node13021;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13027;
	wire [4-1:0] node13030;
	wire [4-1:0] node13033;
	wire [4-1:0] node13034;
	wire [4-1:0] node13035;
	wire [4-1:0] node13038;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13045;
	wire [4-1:0] node13046;
	wire [4-1:0] node13050;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13053;
	wire [4-1:0] node13056;
	wire [4-1:0] node13059;
	wire [4-1:0] node13060;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13066;
	wire [4-1:0] node13069;
	wire [4-1:0] node13072;
	wire [4-1:0] node13073;
	wire [4-1:0] node13075;
	wire [4-1:0] node13078;
	wire [4-1:0] node13079;
	wire [4-1:0] node13080;
	wire [4-1:0] node13083;
	wire [4-1:0] node13086;
	wire [4-1:0] node13088;
	wire [4-1:0] node13091;
	wire [4-1:0] node13092;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13101;
	wire [4-1:0] node13102;
	wire [4-1:0] node13104;
	wire [4-1:0] node13107;
	wire [4-1:0] node13108;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13117;
	wire [4-1:0] node13119;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13124;
	wire [4-1:0] node13127;
	wire [4-1:0] node13130;
	wire [4-1:0] node13132;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13137;
	wire [4-1:0] node13138;
	wire [4-1:0] node13141;
	wire [4-1:0] node13143;
	wire [4-1:0] node13146;
	wire [4-1:0] node13147;
	wire [4-1:0] node13150;
	wire [4-1:0] node13151;
	wire [4-1:0] node13155;
	wire [4-1:0] node13157;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13161;
	wire [4-1:0] node13164;
	wire [4-1:0] node13165;
	wire [4-1:0] node13168;
	wire [4-1:0] node13171;
	wire [4-1:0] node13172;
	wire [4-1:0] node13175;
	wire [4-1:0] node13178;
	wire [4-1:0] node13179;
	wire [4-1:0] node13180;
	wire [4-1:0] node13181;
	wire [4-1:0] node13182;
	wire [4-1:0] node13183;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13190;
	wire [4-1:0] node13192;
	wire [4-1:0] node13193;
	wire [4-1:0] node13196;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13203;
	wire [4-1:0] node13204;
	wire [4-1:0] node13207;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13214;
	wire [4-1:0] node13217;
	wire [4-1:0] node13220;
	wire [4-1:0] node13222;
	wire [4-1:0] node13223;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13230;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13237;
	wire [4-1:0] node13238;
	wire [4-1:0] node13241;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13248;
	wire [4-1:0] node13249;
	wire [4-1:0] node13252;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13257;
	wire [4-1:0] node13260;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13266;
	wire [4-1:0] node13269;
	wire [4-1:0] node13270;
	wire [4-1:0] node13274;
	wire [4-1:0] node13275;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13279;
	wire [4-1:0] node13283;
	wire [4-1:0] node13284;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13292;
	wire [4-1:0] node13295;
	wire [4-1:0] node13296;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13307;
	wire [4-1:0] node13308;
	wire [4-1:0] node13311;
	wire [4-1:0] node13312;
	wire [4-1:0] node13315;
	wire [4-1:0] node13318;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13321;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13327;
	wire [4-1:0] node13328;
	wire [4-1:0] node13333;
	wire [4-1:0] node13334;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13341;
	wire [4-1:0] node13342;
	wire [4-1:0] node13346;
	wire [4-1:0] node13347;
	wire [4-1:0] node13348;
	wire [4-1:0] node13352;
	wire [4-1:0] node13355;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13358;
	wire [4-1:0] node13359;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13365;
	wire [4-1:0] node13368;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13373;
	wire [4-1:0] node13376;
	wire [4-1:0] node13378;
	wire [4-1:0] node13381;
	wire [4-1:0] node13382;
	wire [4-1:0] node13383;
	wire [4-1:0] node13386;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13401;
	wire [4-1:0] node13404;
	wire [4-1:0] node13405;
	wire [4-1:0] node13406;
	wire [4-1:0] node13409;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13416;
	wire [4-1:0] node13419;
	wire [4-1:0] node13420;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13424;
	wire [4-1:0] node13427;
	wire [4-1:0] node13431;
	wire [4-1:0] node13433;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13441;
	wire [4-1:0] node13444;
	wire [4-1:0] node13446;
	wire [4-1:0] node13449;
	wire [4-1:0] node13450;
	wire [4-1:0] node13451;
	wire [4-1:0] node13453;
	wire [4-1:0] node13456;
	wire [4-1:0] node13457;
	wire [4-1:0] node13460;
	wire [4-1:0] node13463;
	wire [4-1:0] node13464;
	wire [4-1:0] node13467;
	wire [4-1:0] node13468;
	wire [4-1:0] node13471;
	wire [4-1:0] node13474;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13477;
	wire [4-1:0] node13478;
	wire [4-1:0] node13480;
	wire [4-1:0] node13482;
	wire [4-1:0] node13485;
	wire [4-1:0] node13486;
	wire [4-1:0] node13487;
	wire [4-1:0] node13491;
	wire [4-1:0] node13494;
	wire [4-1:0] node13495;
	wire [4-1:0] node13497;
	wire [4-1:0] node13499;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13510;
	wire [4-1:0] node13511;
	wire [4-1:0] node13514;
	wire [4-1:0] node13517;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13524;
	wire [4-1:0] node13527;
	wire [4-1:0] node13528;
	wire [4-1:0] node13531;
	wire [4-1:0] node13533;
	wire [4-1:0] node13536;
	wire [4-1:0] node13537;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13541;
	wire [4-1:0] node13544;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13552;
	wire [4-1:0] node13553;
	wire [4-1:0] node13555;
	wire [4-1:0] node13558;
	wire [4-1:0] node13559;
	wire [4-1:0] node13562;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13567;
	wire [4-1:0] node13570;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13575;
	wire [4-1:0] node13578;
	wire [4-1:0] node13581;
	wire [4-1:0] node13584;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13598;
	wire [4-1:0] node13601;
	wire [4-1:0] node13602;
	wire [4-1:0] node13605;
	wire [4-1:0] node13608;
	wire [4-1:0] node13609;
	wire [4-1:0] node13611;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13616;
	wire [4-1:0] node13619;
	wire [4-1:0] node13622;
	wire [4-1:0] node13623;
	wire [4-1:0] node13626;
	wire [4-1:0] node13629;
	wire [4-1:0] node13630;
	wire [4-1:0] node13631;
	wire [4-1:0] node13632;
	wire [4-1:0] node13633;
	wire [4-1:0] node13634;
	wire [4-1:0] node13636;
	wire [4-1:0] node13639;
	wire [4-1:0] node13641;
	wire [4-1:0] node13644;
	wire [4-1:0] node13645;
	wire [4-1:0] node13646;
	wire [4-1:0] node13650;
	wire [4-1:0] node13651;
	wire [4-1:0] node13654;
	wire [4-1:0] node13657;
	wire [4-1:0] node13658;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13663;
	wire [4-1:0] node13666;
	wire [4-1:0] node13667;
	wire [4-1:0] node13671;
	wire [4-1:0] node13672;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13680;
	wire [4-1:0] node13681;
	wire [4-1:0] node13684;
	wire [4-1:0] node13687;
	wire [4-1:0] node13689;
	wire [4-1:0] node13692;
	wire [4-1:0] node13693;
	wire [4-1:0] node13695;
	wire [4-1:0] node13698;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13704;
	wire [4-1:0] node13708;
	wire [4-1:0] node13710;
	wire [4-1:0] node13713;
	wire [4-1:0] node13716;
	wire [4-1:0] node13717;
	wire [4-1:0] node13720;
	wire [4-1:0] node13723;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13726;
	wire [4-1:0] node13727;
	wire [4-1:0] node13730;
	wire [4-1:0] node13731;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13737;
	wire [4-1:0] node13740;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13748;
	wire [4-1:0] node13749;
	wire [4-1:0] node13752;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13758;
	wire [4-1:0] node13759;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13767;
	wire [4-1:0] node13770;
	wire [4-1:0] node13771;
	wire [4-1:0] node13772;
	wire [4-1:0] node13775;
	wire [4-1:0] node13778;
	wire [4-1:0] node13779;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13796;
	wire [4-1:0] node13799;
	wire [4-1:0] node13801;
	wire [4-1:0] node13804;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13807;
	wire [4-1:0] node13808;
	wire [4-1:0] node13809;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13813;
	wire [4-1:0] node13814;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13822;
	wire [4-1:0] node13826;
	wire [4-1:0] node13827;
	wire [4-1:0] node13828;
	wire [4-1:0] node13829;
	wire [4-1:0] node13834;
	wire [4-1:0] node13836;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13843;
	wire [4-1:0] node13844;
	wire [4-1:0] node13845;
	wire [4-1:0] node13846;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13853;
	wire [4-1:0] node13856;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13862;
	wire [4-1:0] node13864;
	wire [4-1:0] node13867;
	wire [4-1:0] node13868;
	wire [4-1:0] node13869;
	wire [4-1:0] node13874;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13879;
	wire [4-1:0] node13882;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13888;
	wire [4-1:0] node13891;
	wire [4-1:0] node13892;
	wire [4-1:0] node13893;
	wire [4-1:0] node13895;
	wire [4-1:0] node13898;
	wire [4-1:0] node13900;
	wire [4-1:0] node13903;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13915;
	wire [4-1:0] node13918;
	wire [4-1:0] node13919;
	wire [4-1:0] node13920;
	wire [4-1:0] node13922;
	wire [4-1:0] node13924;
	wire [4-1:0] node13928;
	wire [4-1:0] node13929;
	wire [4-1:0] node13930;
	wire [4-1:0] node13931;
	wire [4-1:0] node13934;
	wire [4-1:0] node13938;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13943;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13950;
	wire [4-1:0] node13953;
	wire [4-1:0] node13954;
	wire [4-1:0] node13955;
	wire [4-1:0] node13956;
	wire [4-1:0] node13957;
	wire [4-1:0] node13959;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13972;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13979;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13986;
	wire [4-1:0] node13989;
	wire [4-1:0] node13991;
	wire [4-1:0] node13992;
	wire [4-1:0] node13995;
	wire [4-1:0] node13998;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14005;
	wire [4-1:0] node14006;
	wire [4-1:0] node14009;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14015;
	wire [4-1:0] node14018;
	wire [4-1:0] node14019;
	wire [4-1:0] node14022;
	wire [4-1:0] node14025;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14029;
	wire [4-1:0] node14030;
	wire [4-1:0] node14031;
	wire [4-1:0] node14035;
	wire [4-1:0] node14038;
	wire [4-1:0] node14039;
	wire [4-1:0] node14040;
	wire [4-1:0] node14043;
	wire [4-1:0] node14045;
	wire [4-1:0] node14048;
	wire [4-1:0] node14049;
	wire [4-1:0] node14051;
	wire [4-1:0] node14054;
	wire [4-1:0] node14057;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14060;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14068;
	wire [4-1:0] node14069;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14077;
	wire [4-1:0] node14079;
	wire [4-1:0] node14082;
	wire [4-1:0] node14083;
	wire [4-1:0] node14084;
	wire [4-1:0] node14085;
	wire [4-1:0] node14086;
	wire [4-1:0] node14088;
	wire [4-1:0] node14089;
	wire [4-1:0] node14092;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14099;
	wire [4-1:0] node14102;
	wire [4-1:0] node14103;
	wire [4-1:0] node14104;
	wire [4-1:0] node14105;
	wire [4-1:0] node14107;
	wire [4-1:0] node14110;
	wire [4-1:0] node14111;
	wire [4-1:0] node14114;
	wire [4-1:0] node14117;
	wire [4-1:0] node14118;
	wire [4-1:0] node14119;
	wire [4-1:0] node14122;
	wire [4-1:0] node14126;
	wire [4-1:0] node14127;
	wire [4-1:0] node14128;
	wire [4-1:0] node14131;
	wire [4-1:0] node14134;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14144;
	wire [4-1:0] node14147;
	wire [4-1:0] node14149;
	wire [4-1:0] node14152;
	wire [4-1:0] node14153;
	wire [4-1:0] node14155;
	wire [4-1:0] node14159;
	wire [4-1:0] node14160;
	wire [4-1:0] node14161;
	wire [4-1:0] node14162;
	wire [4-1:0] node14165;
	wire [4-1:0] node14168;
	wire [4-1:0] node14169;
	wire [4-1:0] node14173;
	wire [4-1:0] node14174;
	wire [4-1:0] node14175;
	wire [4-1:0] node14179;
	wire [4-1:0] node14181;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14188;
	wire [4-1:0] node14190;
	wire [4-1:0] node14191;
	wire [4-1:0] node14194;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14201;
	wire [4-1:0] node14202;
	wire [4-1:0] node14205;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14211;
	wire [4-1:0] node14213;
	wire [4-1:0] node14214;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14224;
	wire [4-1:0] node14227;
	wire [4-1:0] node14229;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14234;
	wire [4-1:0] node14237;
	wire [4-1:0] node14239;
	wire [4-1:0] node14242;
	wire [4-1:0] node14243;
	wire [4-1:0] node14245;
	wire [4-1:0] node14248;
	wire [4-1:0] node14250;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14255;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14258;
	wire [4-1:0] node14259;
	wire [4-1:0] node14260;
	wire [4-1:0] node14263;
	wire [4-1:0] node14266;
	wire [4-1:0] node14269;
	wire [4-1:0] node14270;
	wire [4-1:0] node14271;
	wire [4-1:0] node14274;
	wire [4-1:0] node14277;
	wire [4-1:0] node14278;
	wire [4-1:0] node14282;
	wire [4-1:0] node14283;
	wire [4-1:0] node14284;
	wire [4-1:0] node14285;
	wire [4-1:0] node14288;
	wire [4-1:0] node14289;
	wire [4-1:0] node14292;
	wire [4-1:0] node14295;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14302;
	wire [4-1:0] node14303;
	wire [4-1:0] node14306;
	wire [4-1:0] node14308;
	wire [4-1:0] node14310;
	wire [4-1:0] node14313;
	wire [4-1:0] node14314;
	wire [4-1:0] node14315;
	wire [4-1:0] node14318;
	wire [4-1:0] node14319;
	wire [4-1:0] node14321;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14334;
	wire [4-1:0] node14336;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14342;
	wire [4-1:0] node14345;
	wire [4-1:0] node14347;
	wire [4-1:0] node14350;
	wire [4-1:0] node14351;
	wire [4-1:0] node14352;
	wire [4-1:0] node14353;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14359;
	wire [4-1:0] node14360;
	wire [4-1:0] node14364;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14367;
	wire [4-1:0] node14372;
	wire [4-1:0] node14374;
	wire [4-1:0] node14375;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14381;
	wire [4-1:0] node14383;
	wire [4-1:0] node14386;
	wire [4-1:0] node14388;
	wire [4-1:0] node14391;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14397;
	wire [4-1:0] node14400;
	wire [4-1:0] node14401;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14405;
	wire [4-1:0] node14408;
	wire [4-1:0] node14410;
	wire [4-1:0] node14413;
	wire [4-1:0] node14414;
	wire [4-1:0] node14416;
	wire [4-1:0] node14419;
	wire [4-1:0] node14421;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14426;
	wire [4-1:0] node14427;
	wire [4-1:0] node14430;
	wire [4-1:0] node14433;
	wire [4-1:0] node14434;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14442;
	wire [4-1:0] node14445;
	wire [4-1:0] node14446;
	wire [4-1:0] node14447;
	wire [4-1:0] node14448;
	wire [4-1:0] node14449;
	wire [4-1:0] node14451;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14463;
	wire [4-1:0] node14464;
	wire [4-1:0] node14469;
	wire [4-1:0] node14470;
	wire [4-1:0] node14472;
	wire [4-1:0] node14475;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14482;
	wire [4-1:0] node14486;
	wire [4-1:0] node14489;
	wire [4-1:0] node14490;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14496;
	wire [4-1:0] node14499;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14507;
	wire [4-1:0] node14508;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14515;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14521;
	wire [4-1:0] node14523;
	wire [4-1:0] node14526;
	wire [4-1:0] node14527;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14531;
	wire [4-1:0] node14535;
	wire [4-1:0] node14536;
	wire [4-1:0] node14539;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14548;
	wire [4-1:0] node14550;
	wire [4-1:0] node14551;
	wire [4-1:0] node14555;
	wire [4-1:0] node14556;
	wire [4-1:0] node14557;
	wire [4-1:0] node14558;
	wire [4-1:0] node14561;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14567;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14574;
	wire [4-1:0] node14577;
	wire [4-1:0] node14578;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14583;
	wire [4-1:0] node14586;
	wire [4-1:0] node14587;
	wire [4-1:0] node14590;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14595;
	wire [4-1:0] node14598;
	wire [4-1:0] node14601;
	wire [4-1:0] node14603;
	wire [4-1:0] node14606;
	wire [4-1:0] node14607;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14612;
	wire [4-1:0] node14613;
	wire [4-1:0] node14614;
	wire [4-1:0] node14618;
	wire [4-1:0] node14619;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14632;
	wire [4-1:0] node14633;
	wire [4-1:0] node14636;
	wire [4-1:0] node14640;
	wire [4-1:0] node14641;
	wire [4-1:0] node14643;
	wire [4-1:0] node14646;
	wire [4-1:0] node14648;
	wire [4-1:0] node14651;
	wire [4-1:0] node14652;
	wire [4-1:0] node14653;
	wire [4-1:0] node14654;
	wire [4-1:0] node14655;
	wire [4-1:0] node14659;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14665;
	wire [4-1:0] node14668;
	wire [4-1:0] node14670;
	wire [4-1:0] node14673;
	wire [4-1:0] node14674;
	wire [4-1:0] node14675;
	wire [4-1:0] node14676;
	wire [4-1:0] node14680;
	wire [4-1:0] node14682;
	wire [4-1:0] node14685;
	wire [4-1:0] node14686;
	wire [4-1:0] node14688;
	wire [4-1:0] node14691;
	wire [4-1:0] node14693;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14700;
	wire [4-1:0] node14702;
	wire [4-1:0] node14705;
	wire [4-1:0] node14707;
	wire [4-1:0] node14710;
	wire [4-1:0] node14711;
	wire [4-1:0] node14713;
	wire [4-1:0] node14717;
	wire [4-1:0] node14718;
	wire [4-1:0] node14719;
	wire [4-1:0] node14722;
	wire [4-1:0] node14725;
	wire [4-1:0] node14726;
	wire [4-1:0] node14727;
	wire [4-1:0] node14730;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14736;
	wire [4-1:0] node14737;
	wire [4-1:0] node14738;
	wire [4-1:0] node14741;
	wire [4-1:0] node14745;
	wire [4-1:0] node14746;
	wire [4-1:0] node14747;
	wire [4-1:0] node14748;
	wire [4-1:0] node14751;
	wire [4-1:0] node14756;
	wire [4-1:0] node14757;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14760;
	wire [4-1:0] node14763;
	wire [4-1:0] node14766;
	wire [4-1:0] node14767;
	wire [4-1:0] node14770;
	wire [4-1:0] node14774;
	wire [4-1:0] node14775;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14787;
	wire [4-1:0] node14788;
	wire [4-1:0] node14789;
	wire [4-1:0] node14790;
	wire [4-1:0] node14791;
	wire [4-1:0] node14794;
	wire [4-1:0] node14798;
	wire [4-1:0] node14799;
	wire [4-1:0] node14801;
	wire [4-1:0] node14804;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14814;
	wire [4-1:0] node14816;
	wire [4-1:0] node14819;
	wire [4-1:0] node14821;
	wire [4-1:0] node14825;
	wire [4-1:0] node14827;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14832;
	wire [4-1:0] node14833;
	wire [4-1:0] node14834;
	wire [4-1:0] node14837;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14845;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14854;
	wire [4-1:0] node14858;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14863;
	wire [4-1:0] node14866;
	wire [4-1:0] node14867;
	wire [4-1:0] node14868;
	wire [4-1:0] node14872;
	wire [4-1:0] node14873;
	wire [4-1:0] node14877;
	wire [4-1:0] node14878;
	wire [4-1:0] node14879;
	wire [4-1:0] node14880;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14890;
	wire [4-1:0] node14891;
	wire [4-1:0] node14894;
	wire [4-1:0] node14898;
	wire [4-1:0] node14899;
	wire [4-1:0] node14900;
	wire [4-1:0] node14901;
	wire [4-1:0] node14902;
	wire [4-1:0] node14905;
	wire [4-1:0] node14908;
	wire [4-1:0] node14909;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14917;
	wire [4-1:0] node14918;
	wire [4-1:0] node14920;
	wire [4-1:0] node14921;
	wire [4-1:0] node14924;
	wire [4-1:0] node14927;
	wire [4-1:0] node14928;
	wire [4-1:0] node14931;
	wire [4-1:0] node14935;
	wire [4-1:0] node14936;
	wire [4-1:0] node14937;
	wire [4-1:0] node14938;
	wire [4-1:0] node14941;
	wire [4-1:0] node14944;
	wire [4-1:0] node14945;
	wire [4-1:0] node14946;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14954;
	wire [4-1:0] node14958;
	wire [4-1:0] node14959;
	wire [4-1:0] node14960;
	wire [4-1:0] node14961;
	wire [4-1:0] node14962;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14965;
	wire [4-1:0] node14969;
	wire [4-1:0] node14970;
	wire [4-1:0] node14973;
	wire [4-1:0] node14976;
	wire [4-1:0] node14977;
	wire [4-1:0] node14980;
	wire [4-1:0] node14983;
	wire [4-1:0] node14984;
	wire [4-1:0] node14985;
	wire [4-1:0] node14987;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14994;
	wire [4-1:0] node14997;
	wire [4-1:0] node14998;
	wire [4-1:0] node14999;
	wire [4-1:0] node15000;
	wire [4-1:0] node15005;
	wire [4-1:0] node15006;
	wire [4-1:0] node15010;
	wire [4-1:0] node15011;
	wire [4-1:0] node15012;
	wire [4-1:0] node15013;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15020;
	wire [4-1:0] node15021;
	wire [4-1:0] node15024;
	wire [4-1:0] node15027;
	wire [4-1:0] node15028;
	wire [4-1:0] node15029;
	wire [4-1:0] node15032;
	wire [4-1:0] node15035;
	wire [4-1:0] node15037;
	wire [4-1:0] node15038;
	wire [4-1:0] node15042;
	wire [4-1:0] node15043;
	wire [4-1:0] node15044;
	wire [4-1:0] node15045;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15053;
	wire [4-1:0] node15056;
	wire [4-1:0] node15057;
	wire [4-1:0] node15060;
	wire [4-1:0] node15061;
	wire [4-1:0] node15065;
	wire [4-1:0] node15066;
	wire [4-1:0] node15067;
	wire [4-1:0] node15068;
	wire [4-1:0] node15069;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15076;
	wire [4-1:0] node15077;
	wire [4-1:0] node15078;
	wire [4-1:0] node15081;
	wire [4-1:0] node15085;
	wire [4-1:0] node15086;
	wire [4-1:0] node15089;
	wire [4-1:0] node15092;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15096;
	wire [4-1:0] node15099;
	wire [4-1:0] node15100;
	wire [4-1:0] node15103;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15112;
	wire [4-1:0] node15116;
	wire [4-1:0] node15118;
	wire [4-1:0] node15121;
	wire [4-1:0] node15122;
	wire [4-1:0] node15123;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15129;
	wire [4-1:0] node15132;
	wire [4-1:0] node15133;
	wire [4-1:0] node15135;
	wire [4-1:0] node15137;
	wire [4-1:0] node15140;
	wire [4-1:0] node15142;
	wire [4-1:0] node15143;
	wire [4-1:0] node15146;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15151;
	wire [4-1:0] node15152;
	wire [4-1:0] node15154;
	wire [4-1:0] node15157;
	wire [4-1:0] node15158;
	wire [4-1:0] node15161;
	wire [4-1:0] node15164;
	wire [4-1:0] node15165;
	wire [4-1:0] node15169;
	wire [4-1:0] node15170;
	wire [4-1:0] node15173;
	wire [4-1:0] node15176;
	wire [4-1:0] node15177;
	wire [4-1:0] node15178;
	wire [4-1:0] node15179;
	wire [4-1:0] node15180;
	wire [4-1:0] node15181;
	wire [4-1:0] node15182;
	wire [4-1:0] node15183;
	wire [4-1:0] node15187;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15195;
	wire [4-1:0] node15196;
	wire [4-1:0] node15198;
	wire [4-1:0] node15200;
	wire [4-1:0] node15203;
	wire [4-1:0] node15204;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15211;
	wire [4-1:0] node15214;
	wire [4-1:0] node15217;
	wire [4-1:0] node15219;
	wire [4-1:0] node15220;
	wire [4-1:0] node15224;
	wire [4-1:0] node15226;
	wire [4-1:0] node15227;
	wire [4-1:0] node15228;
	wire [4-1:0] node15231;
	wire [4-1:0] node15235;
	wire [4-1:0] node15236;
	wire [4-1:0] node15237;
	wire [4-1:0] node15238;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15246;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15252;
	wire [4-1:0] node15253;
	wire [4-1:0] node15255;
	wire [4-1:0] node15259;
	wire [4-1:0] node15260;
	wire [4-1:0] node15261;
	wire [4-1:0] node15262;
	wire [4-1:0] node15264;
	wire [4-1:0] node15267;
	wire [4-1:0] node15270;
	wire [4-1:0] node15272;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15277;
	wire [4-1:0] node15279;
	wire [4-1:0] node15282;
	wire [4-1:0] node15283;
	wire [4-1:0] node15287;
	wire [4-1:0] node15288;
	wire [4-1:0] node15292;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15295;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15301;
	wire [4-1:0] node15302;
	wire [4-1:0] node15306;
	wire [4-1:0] node15307;
	wire [4-1:0] node15310;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15315;
	wire [4-1:0] node15318;
	wire [4-1:0] node15321;
	wire [4-1:0] node15323;
	wire [4-1:0] node15324;
	wire [4-1:0] node15325;
	wire [4-1:0] node15329;
	wire [4-1:0] node15331;
	wire [4-1:0] node15334;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15341;
	wire [4-1:0] node15344;
	wire [4-1:0] node15345;
	wire [4-1:0] node15347;
	wire [4-1:0] node15350;
	wire [4-1:0] node15351;
	wire [4-1:0] node15354;
	wire [4-1:0] node15357;
	wire [4-1:0] node15359;
	wire [4-1:0] node15360;
	wire [4-1:0] node15364;
	wire [4-1:0] node15365;
	wire [4-1:0] node15366;
	wire [4-1:0] node15369;
	wire [4-1:0] node15372;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15376;
	wire [4-1:0] node15379;
	wire [4-1:0] node15380;
	wire [4-1:0] node15384;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15391;
	wire [4-1:0] node15392;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15395;
	wire [4-1:0] node15396;
	wire [4-1:0] node15397;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15400;
	wire [4-1:0] node15401;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15407;
	wire [4-1:0] node15409;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15420;
	wire [4-1:0] node15421;
	wire [4-1:0] node15422;
	wire [4-1:0] node15427;
	wire [4-1:0] node15428;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15434;
	wire [4-1:0] node15435;
	wire [4-1:0] node15436;
	wire [4-1:0] node15439;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15446;
	wire [4-1:0] node15449;
	wire [4-1:0] node15451;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15457;
	wire [4-1:0] node15458;
	wire [4-1:0] node15459;
	wire [4-1:0] node15460;
	wire [4-1:0] node15464;
	wire [4-1:0] node15467;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15472;
	wire [4-1:0] node15475;
	wire [4-1:0] node15476;
	wire [4-1:0] node15477;
	wire [4-1:0] node15482;
	wire [4-1:0] node15483;
	wire [4-1:0] node15484;
	wire [4-1:0] node15486;
	wire [4-1:0] node15488;
	wire [4-1:0] node15491;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15497;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15502;
	wire [4-1:0] node15503;
	wire [4-1:0] node15507;
	wire [4-1:0] node15510;
	wire [4-1:0] node15511;
	wire [4-1:0] node15514;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15521;
	wire [4-1:0] node15522;
	wire [4-1:0] node15525;
	wire [4-1:0] node15527;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15533;
	wire [4-1:0] node15537;
	wire [4-1:0] node15538;
	wire [4-1:0] node15539;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15550;
	wire [4-1:0] node15553;
	wire [4-1:0] node15554;
	wire [4-1:0] node15558;
	wire [4-1:0] node15559;
	wire [4-1:0] node15560;
	wire [4-1:0] node15562;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15576;
	wire [4-1:0] node15577;
	wire [4-1:0] node15578;
	wire [4-1:0] node15582;
	wire [4-1:0] node15583;
	wire [4-1:0] node15587;
	wire [4-1:0] node15588;
	wire [4-1:0] node15589;
	wire [4-1:0] node15590;
	wire [4-1:0] node15591;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15600;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15604;
	wire [4-1:0] node15607;
	wire [4-1:0] node15608;
	wire [4-1:0] node15612;
	wire [4-1:0] node15613;
	wire [4-1:0] node15616;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15622;
	wire [4-1:0] node15625;
	wire [4-1:0] node15628;
	wire [4-1:0] node15630;
	wire [4-1:0] node15631;
	wire [4-1:0] node15634;
	wire [4-1:0] node15637;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15644;
	wire [4-1:0] node15646;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15653;
	wire [4-1:0] node15655;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15661;
	wire [4-1:0] node15662;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15668;
	wire [4-1:0] node15669;
	wire [4-1:0] node15671;
	wire [4-1:0] node15675;
	wire [4-1:0] node15676;
	wire [4-1:0] node15679;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15687;
	wire [4-1:0] node15688;
	wire [4-1:0] node15690;
	wire [4-1:0] node15693;
	wire [4-1:0] node15695;
	wire [4-1:0] node15698;
	wire [4-1:0] node15699;
	wire [4-1:0] node15701;
	wire [4-1:0] node15704;
	wire [4-1:0] node15705;
	wire [4-1:0] node15709;
	wire [4-1:0] node15710;
	wire [4-1:0] node15711;
	wire [4-1:0] node15713;
	wire [4-1:0] node15714;
	wire [4-1:0] node15717;
	wire [4-1:0] node15718;
	wire [4-1:0] node15722;
	wire [4-1:0] node15723;
	wire [4-1:0] node15724;
	wire [4-1:0] node15726;
	wire [4-1:0] node15730;
	wire [4-1:0] node15731;
	wire [4-1:0] node15735;
	wire [4-1:0] node15736;
	wire [4-1:0] node15737;
	wire [4-1:0] node15739;
	wire [4-1:0] node15742;
	wire [4-1:0] node15743;
	wire [4-1:0] node15747;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15750;
	wire [4-1:0] node15755;
	wire [4-1:0] node15757;
	wire [4-1:0] node15759;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15766;
	wire [4-1:0] node15767;
	wire [4-1:0] node15770;
	wire [4-1:0] node15773;
	wire [4-1:0] node15775;
	wire [4-1:0] node15777;
	wire [4-1:0] node15780;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15784;
	wire [4-1:0] node15787;
	wire [4-1:0] node15789;
	wire [4-1:0] node15792;
	wire [4-1:0] node15794;
	wire [4-1:0] node15797;
	wire [4-1:0] node15798;
	wire [4-1:0] node15799;
	wire [4-1:0] node15801;
	wire [4-1:0] node15804;
	wire [4-1:0] node15805;
	wire [4-1:0] node15806;
	wire [4-1:0] node15811;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15815;
	wire [4-1:0] node15819;
	wire [4-1:0] node15820;
	wire [4-1:0] node15822;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15829;
	wire [4-1:0] node15830;
	wire [4-1:0] node15832;
	wire [4-1:0] node15835;
	wire [4-1:0] node15837;
	wire [4-1:0] node15840;
	wire [4-1:0] node15841;
	wire [4-1:0] node15842;
	wire [4-1:0] node15847;
	wire [4-1:0] node15849;
	wire [4-1:0] node15851;
	wire [4-1:0] node15853;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15859;
	wire [4-1:0] node15862;
	wire [4-1:0] node15865;
	wire [4-1:0] node15866;
	wire [4-1:0] node15868;
	wire [4-1:0] node15871;
	wire [4-1:0] node15873;
	wire [4-1:0] node15876;
	wire [4-1:0] node15877;
	wire [4-1:0] node15878;
	wire [4-1:0] node15879;
	wire [4-1:0] node15883;
	wire [4-1:0] node15886;
	wire [4-1:0] node15888;
	wire [4-1:0] node15889;
	wire [4-1:0] node15893;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15896;
	wire [4-1:0] node15897;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15900;
	wire [4-1:0] node15901;
	wire [4-1:0] node15904;
	wire [4-1:0] node15908;
	wire [4-1:0] node15909;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15916;
	wire [4-1:0] node15919;
	wire [4-1:0] node15920;
	wire [4-1:0] node15922;
	wire [4-1:0] node15926;
	wire [4-1:0] node15927;
	wire [4-1:0] node15928;
	wire [4-1:0] node15931;
	wire [4-1:0] node15932;
	wire [4-1:0] node15936;
	wire [4-1:0] node15937;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15944;
	wire [4-1:0] node15947;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15950;
	wire [4-1:0] node15951;
	wire [4-1:0] node15954;
	wire [4-1:0] node15956;
	wire [4-1:0] node15959;
	wire [4-1:0] node15960;
	wire [4-1:0] node15963;
	wire [4-1:0] node15964;
	wire [4-1:0] node15968;
	wire [4-1:0] node15969;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15978;
	wire [4-1:0] node15979;
	wire [4-1:0] node15983;
	wire [4-1:0] node15984;
	wire [4-1:0] node15985;
	wire [4-1:0] node15986;
	wire [4-1:0] node15990;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15997;
	wire [4-1:0] node15998;
	wire [4-1:0] node15999;
	wire [4-1:0] node16002;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16009;
	wire [4-1:0] node16012;
	wire [4-1:0] node16013;
	wire [4-1:0] node16014;
	wire [4-1:0] node16015;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16024;
	wire [4-1:0] node16027;
	wire [4-1:0] node16028;
	wire [4-1:0] node16030;
	wire [4-1:0] node16033;
	wire [4-1:0] node16036;
	wire [4-1:0] node16037;
	wire [4-1:0] node16038;
	wire [4-1:0] node16041;
	wire [4-1:0] node16042;
	wire [4-1:0] node16045;
	wire [4-1:0] node16048;
	wire [4-1:0] node16049;
	wire [4-1:0] node16050;
	wire [4-1:0] node16054;
	wire [4-1:0] node16056;
	wire [4-1:0] node16059;
	wire [4-1:0] node16060;
	wire [4-1:0] node16061;
	wire [4-1:0] node16062;
	wire [4-1:0] node16065;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16070;
	wire [4-1:0] node16074;
	wire [4-1:0] node16076;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16081;
	wire [4-1:0] node16085;
	wire [4-1:0] node16086;
	wire [4-1:0] node16087;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16094;
	wire [4-1:0] node16095;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16102;
	wire [4-1:0] node16103;
	wire [4-1:0] node16106;
	wire [4-1:0] node16109;
	wire [4-1:0] node16111;
	wire [4-1:0] node16112;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16118;
	wire [4-1:0] node16121;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16128;
	wire [4-1:0] node16129;
	wire [4-1:0] node16131;
	wire [4-1:0] node16133;
	wire [4-1:0] node16136;
	wire [4-1:0] node16137;
	wire [4-1:0] node16141;
	wire [4-1:0] node16142;
	wire [4-1:0] node16143;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16152;
	wire [4-1:0] node16153;
	wire [4-1:0] node16157;
	wire [4-1:0] node16158;
	wire [4-1:0] node16162;
	wire [4-1:0] node16163;
	wire [4-1:0] node16164;
	wire [4-1:0] node16168;
	wire [4-1:0] node16169;
	wire [4-1:0] node16170;
	wire [4-1:0] node16175;
	wire [4-1:0] node16176;
	wire [4-1:0] node16177;
	wire [4-1:0] node16178;
	wire [4-1:0] node16179;
	wire [4-1:0] node16183;
	wire [4-1:0] node16184;
	wire [4-1:0] node16187;
	wire [4-1:0] node16190;
	wire [4-1:0] node16192;
	wire [4-1:0] node16195;
	wire [4-1:0] node16197;
	wire [4-1:0] node16198;
	wire [4-1:0] node16201;
	wire [4-1:0] node16204;
	wire [4-1:0] node16205;
	wire [4-1:0] node16206;
	wire [4-1:0] node16207;
	wire [4-1:0] node16208;
	wire [4-1:0] node16211;
	wire [4-1:0] node16214;
	wire [4-1:0] node16215;
	wire [4-1:0] node16216;
	wire [4-1:0] node16219;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16225;
	wire [4-1:0] node16230;
	wire [4-1:0] node16231;
	wire [4-1:0] node16232;
	wire [4-1:0] node16233;
	wire [4-1:0] node16234;
	wire [4-1:0] node16238;
	wire [4-1:0] node16239;
	wire [4-1:0] node16243;
	wire [4-1:0] node16245;
	wire [4-1:0] node16248;
	wire [4-1:0] node16250;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16264;
	wire [4-1:0] node16268;
	wire [4-1:0] node16269;
	wire [4-1:0] node16270;
	wire [4-1:0] node16274;
	wire [4-1:0] node16276;
	wire [4-1:0] node16279;
	wire [4-1:0] node16280;
	wire [4-1:0] node16281;
	wire [4-1:0] node16283;
	wire [4-1:0] node16288;
	wire [4-1:0] node16289;
	wire [4-1:0] node16290;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16295;
	wire [4-1:0] node16299;
	wire [4-1:0] node16300;
	wire [4-1:0] node16302;
	wire [4-1:0] node16305;
	wire [4-1:0] node16308;
	wire [4-1:0] node16309;
	wire [4-1:0] node16310;
	wire [4-1:0] node16313;
	wire [4-1:0] node16316;
	wire [4-1:0] node16317;
	wire [4-1:0] node16318;
	wire [4-1:0] node16321;
	wire [4-1:0] node16324;
	wire [4-1:0] node16325;
	wire [4-1:0] node16328;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16333;
	wire [4-1:0] node16334;
	wire [4-1:0] node16335;
	wire [4-1:0] node16337;
	wire [4-1:0] node16340;
	wire [4-1:0] node16342;
	wire [4-1:0] node16346;
	wire [4-1:0] node16347;
	wire [4-1:0] node16349;
	wire [4-1:0] node16350;
	wire [4-1:0] node16354;
	wire [4-1:0] node16355;
	wire [4-1:0] node16359;
	wire [4-1:0] node16360;
	wire [4-1:0] node16361;
	wire [4-1:0] node16362;
	wire [4-1:0] node16363;
	wire [4-1:0] node16367;
	wire [4-1:0] node16370;
	wire [4-1:0] node16371;
	wire [4-1:0] node16375;
	wire [4-1:0] node16376;
	wire [4-1:0] node16378;
	wire [4-1:0] node16381;
	wire [4-1:0] node16383;
	wire [4-1:0] node16384;
	wire [4-1:0] node16387;
	wire [4-1:0] node16390;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16395;
	wire [4-1:0] node16396;
	wire [4-1:0] node16397;
	wire [4-1:0] node16398;
	wire [4-1:0] node16400;
	wire [4-1:0] node16403;
	wire [4-1:0] node16406;
	wire [4-1:0] node16408;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16413;
	wire [4-1:0] node16415;
	wire [4-1:0] node16418;
	wire [4-1:0] node16419;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16425;
	wire [4-1:0] node16429;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16436;
	wire [4-1:0] node16440;
	wire [4-1:0] node16443;
	wire [4-1:0] node16444;
	wire [4-1:0] node16447;
	wire [4-1:0] node16448;
	wire [4-1:0] node16451;
	wire [4-1:0] node16454;
	wire [4-1:0] node16455;
	wire [4-1:0] node16456;
	wire [4-1:0] node16459;
	wire [4-1:0] node16462;
	wire [4-1:0] node16464;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16470;
	wire [4-1:0] node16472;
	wire [4-1:0] node16473;
	wire [4-1:0] node16477;
	wire [4-1:0] node16479;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16484;
	wire [4-1:0] node16486;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16499;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16505;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16512;
	wire [4-1:0] node16514;
	wire [4-1:0] node16517;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16527;
	wire [4-1:0] node16528;
	wire [4-1:0] node16532;
	wire [4-1:0] node16533;
	wire [4-1:0] node16534;
	wire [4-1:0] node16535;
	wire [4-1:0] node16536;
	wire [4-1:0] node16537;
	wire [4-1:0] node16541;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16547;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16552;
	wire [4-1:0] node16554;
	wire [4-1:0] node16557;
	wire [4-1:0] node16559;
	wire [4-1:0] node16562;
	wire [4-1:0] node16563;
	wire [4-1:0] node16566;
	wire [4-1:0] node16568;
	wire [4-1:0] node16571;
	wire [4-1:0] node16572;
	wire [4-1:0] node16573;
	wire [4-1:0] node16576;
	wire [4-1:0] node16577;
	wire [4-1:0] node16578;
	wire [4-1:0] node16581;
	wire [4-1:0] node16585;
	wire [4-1:0] node16586;
	wire [4-1:0] node16588;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16593;
	wire [4-1:0] node16596;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16603;
	wire [4-1:0] node16604;
	wire [4-1:0] node16607;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16612;
	wire [4-1:0] node16617;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16625;
	wire [4-1:0] node16626;
	wire [4-1:0] node16630;
	wire [4-1:0] node16631;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16636;
	wire [4-1:0] node16639;
	wire [4-1:0] node16641;
	wire [4-1:0] node16644;
	wire [4-1:0] node16645;
	wire [4-1:0] node16646;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16656;
	wire [4-1:0] node16657;
	wire [4-1:0] node16661;
	wire [4-1:0] node16662;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16667;
	wire [4-1:0] node16669;
	wire [4-1:0] node16673;
	wire [4-1:0] node16674;
	wire [4-1:0] node16675;
	wire [4-1:0] node16680;
	wire [4-1:0] node16682;
	wire [4-1:0] node16683;
	wire [4-1:0] node16684;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16692;
	wire [4-1:0] node16695;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16701;
	wire [4-1:0] node16705;
	wire [4-1:0] node16706;
	wire [4-1:0] node16707;
	wire [4-1:0] node16709;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16716;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16722;
	wire [4-1:0] node16725;
	wire [4-1:0] node16726;
	wire [4-1:0] node16730;
	wire [4-1:0] node16731;
	wire [4-1:0] node16732;
	wire [4-1:0] node16733;
	wire [4-1:0] node16734;
	wire [4-1:0] node16737;
	wire [4-1:0] node16739;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16746;
	wire [4-1:0] node16750;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16753;
	wire [4-1:0] node16754;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16762;
	wire [4-1:0] node16765;
	wire [4-1:0] node16767;
	wire [4-1:0] node16770;
	wire [4-1:0] node16771;
	wire [4-1:0] node16773;
	wire [4-1:0] node16776;
	wire [4-1:0] node16778;
	wire [4-1:0] node16780;
	wire [4-1:0] node16783;
	wire [4-1:0] node16784;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16792;
	wire [4-1:0] node16795;
	wire [4-1:0] node16796;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16802;
	wire [4-1:0] node16804;
	wire [4-1:0] node16805;
	wire [4-1:0] node16808;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16813;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16821;
	wire [4-1:0] node16824;
	wire [4-1:0] node16827;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16830;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16835;
	wire [4-1:0] node16838;
	wire [4-1:0] node16842;
	wire [4-1:0] node16843;
	wire [4-1:0] node16844;
	wire [4-1:0] node16845;
	wire [4-1:0] node16851;
	wire [4-1:0] node16852;
	wire [4-1:0] node16853;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16859;
	wire [4-1:0] node16860;
	wire [4-1:0] node16863;
	wire [4-1:0] node16866;
	wire [4-1:0] node16867;
	wire [4-1:0] node16868;
	wire [4-1:0] node16871;
	wire [4-1:0] node16875;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16880;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16890;
	wire [4-1:0] node16891;
	wire [4-1:0] node16892;
	wire [4-1:0] node16893;
	wire [4-1:0] node16894;
	wire [4-1:0] node16895;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16903;
	wire [4-1:0] node16904;
	wire [4-1:0] node16905;
	wire [4-1:0] node16909;
	wire [4-1:0] node16912;
	wire [4-1:0] node16913;
	wire [4-1:0] node16917;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16921;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16930;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16937;
	wire [4-1:0] node16938;
	wire [4-1:0] node16939;
	wire [4-1:0] node16942;
	wire [4-1:0] node16945;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16950;
	wire [4-1:0] node16952;
	wire [4-1:0] node16953;
	wire [4-1:0] node16954;
	wire [4-1:0] node16957;
	wire [4-1:0] node16960;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16965;
	wire [4-1:0] node16966;
	wire [4-1:0] node16970;
	wire [4-1:0] node16973;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16979;
	wire [4-1:0] node16982;
	wire [4-1:0] node16983;
	wire [4-1:0] node16984;
	wire [4-1:0] node16985;
	wire [4-1:0] node16988;
	wire [4-1:0] node16989;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16995;
	wire [4-1:0] node16999;
	wire [4-1:0] node17001;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17012;
	wire [4-1:0] node17015;
	wire [4-1:0] node17016;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17019;
	wire [4-1:0] node17020;
	wire [4-1:0] node17021;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17029;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17037;
	wire [4-1:0] node17040;
	wire [4-1:0] node17041;
	wire [4-1:0] node17045;
	wire [4-1:0] node17046;
	wire [4-1:0] node17047;
	wire [4-1:0] node17048;
	wire [4-1:0] node17051;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17060;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17064;
	wire [4-1:0] node17066;
	wire [4-1:0] node17069;
	wire [4-1:0] node17071;
	wire [4-1:0] node17072;
	wire [4-1:0] node17075;
	wire [4-1:0] node17078;
	wire [4-1:0] node17079;
	wire [4-1:0] node17080;
	wire [4-1:0] node17084;
	wire [4-1:0] node17085;
	wire [4-1:0] node17088;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17095;
	wire [4-1:0] node17098;
	wire [4-1:0] node17101;
	wire [4-1:0] node17102;
	wire [4-1:0] node17105;
	wire [4-1:0] node17108;
	wire [4-1:0] node17109;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17119;
	wire [4-1:0] node17123;
	wire [4-1:0] node17124;
	wire [4-1:0] node17125;
	wire [4-1:0] node17127;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17132;
	wire [4-1:0] node17135;
	wire [4-1:0] node17138;
	wire [4-1:0] node17139;
	wire [4-1:0] node17142;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17150;
	wire [4-1:0] node17153;
	wire [4-1:0] node17155;
	wire [4-1:0] node17156;
	wire [4-1:0] node17159;
	wire [4-1:0] node17162;
	wire [4-1:0] node17163;
	wire [4-1:0] node17164;
	wire [4-1:0] node17165;
	wire [4-1:0] node17166;
	wire [4-1:0] node17167;
	wire [4-1:0] node17168;
	wire [4-1:0] node17170;
	wire [4-1:0] node17173;
	wire [4-1:0] node17176;
	wire [4-1:0] node17178;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17189;
	wire [4-1:0] node17190;
	wire [4-1:0] node17194;
	wire [4-1:0] node17195;
	wire [4-1:0] node17197;
	wire [4-1:0] node17198;
	wire [4-1:0] node17199;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17208;
	wire [4-1:0] node17209;
	wire [4-1:0] node17211;
	wire [4-1:0] node17213;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17220;
	wire [4-1:0] node17223;
	wire [4-1:0] node17224;
	wire [4-1:0] node17225;
	wire [4-1:0] node17226;
	wire [4-1:0] node17229;
	wire [4-1:0] node17231;
	wire [4-1:0] node17233;
	wire [4-1:0] node17236;
	wire [4-1:0] node17237;
	wire [4-1:0] node17238;
	wire [4-1:0] node17239;
	wire [4-1:0] node17243;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17250;
	wire [4-1:0] node17253;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17260;
	wire [4-1:0] node17262;
	wire [4-1:0] node17263;
	wire [4-1:0] node17266;
	wire [4-1:0] node17269;
	wire [4-1:0] node17270;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17277;
	wire [4-1:0] node17278;
	wire [4-1:0] node17279;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17288;
	wire [4-1:0] node17289;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17293;
	wire [4-1:0] node17294;
	wire [4-1:0] node17295;
	wire [4-1:0] node17298;
	wire [4-1:0] node17302;
	wire [4-1:0] node17303;
	wire [4-1:0] node17304;
	wire [4-1:0] node17305;
	wire [4-1:0] node17308;
	wire [4-1:0] node17311;
	wire [4-1:0] node17312;
	wire [4-1:0] node17316;
	wire [4-1:0] node17317;
	wire [4-1:0] node17320;
	wire [4-1:0] node17323;
	wire [4-1:0] node17324;
	wire [4-1:0] node17325;
	wire [4-1:0] node17326;
	wire [4-1:0] node17329;
	wire [4-1:0] node17332;
	wire [4-1:0] node17334;
	wire [4-1:0] node17335;
	wire [4-1:0] node17339;
	wire [4-1:0] node17340;
	wire [4-1:0] node17342;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17348;
	wire [4-1:0] node17352;
	wire [4-1:0] node17353;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17357;
	wire [4-1:0] node17360;
	wire [4-1:0] node17363;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17370;
	wire [4-1:0] node17373;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17380;
	wire [4-1:0] node17383;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17388;
	wire [4-1:0] node17391;
	wire [4-1:0] node17392;
	wire [4-1:0] node17393;
	wire [4-1:0] node17396;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17403;
	wire [4-1:0] node17406;
	wire [4-1:0] node17407;
	wire [4-1:0] node17408;
	wire [4-1:0] node17409;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17417;
	wire [4-1:0] node17418;
	wire [4-1:0] node17419;
	wire [4-1:0] node17423;
	wire [4-1:0] node17425;
	wire [4-1:0] node17428;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17433;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17441;
	wire [4-1:0] node17444;
	wire [4-1:0] node17447;
	wire [4-1:0] node17448;
	wire [4-1:0] node17449;
	wire [4-1:0] node17450;
	wire [4-1:0] node17451;
	wire [4-1:0] node17452;
	wire [4-1:0] node17453;
	wire [4-1:0] node17454;
	wire [4-1:0] node17455;
	wire [4-1:0] node17456;
	wire [4-1:0] node17459;
	wire [4-1:0] node17462;
	wire [4-1:0] node17463;
	wire [4-1:0] node17464;
	wire [4-1:0] node17468;
	wire [4-1:0] node17471;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17476;
	wire [4-1:0] node17479;
	wire [4-1:0] node17480;
	wire [4-1:0] node17482;
	wire [4-1:0] node17485;
	wire [4-1:0] node17488;
	wire [4-1:0] node17489;
	wire [4-1:0] node17490;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17495;
	wire [4-1:0] node17498;
	wire [4-1:0] node17501;
	wire [4-1:0] node17504;
	wire [4-1:0] node17505;
	wire [4-1:0] node17506;
	wire [4-1:0] node17507;
	wire [4-1:0] node17511;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17518;
	wire [4-1:0] node17519;
	wire [4-1:0] node17520;
	wire [4-1:0] node17523;
	wire [4-1:0] node17526;
	wire [4-1:0] node17529;
	wire [4-1:0] node17530;
	wire [4-1:0] node17531;
	wire [4-1:0] node17532;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17538;
	wire [4-1:0] node17539;
	wire [4-1:0] node17542;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17549;
	wire [4-1:0] node17550;
	wire [4-1:0] node17553;
	wire [4-1:0] node17556;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17563;
	wire [4-1:0] node17564;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17568;
	wire [4-1:0] node17572;
	wire [4-1:0] node17573;
	wire [4-1:0] node17574;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17582;
	wire [4-1:0] node17585;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17589;
	wire [4-1:0] node17594;
	wire [4-1:0] node17595;
	wire [4-1:0] node17596;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17600;
	wire [4-1:0] node17603;
	wire [4-1:0] node17604;
	wire [4-1:0] node17605;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17616;
	wire [4-1:0] node17618;
	wire [4-1:0] node17622;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17628;
	wire [4-1:0] node17629;
	wire [4-1:0] node17633;
	wire [4-1:0] node17634;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17639;
	wire [4-1:0] node17641;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17647;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17654;
	wire [4-1:0] node17657;
	wire [4-1:0] node17659;
	wire [4-1:0] node17662;
	wire [4-1:0] node17663;
	wire [4-1:0] node17664;
	wire [4-1:0] node17665;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17670;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17678;
	wire [4-1:0] node17680;
	wire [4-1:0] node17683;
	wire [4-1:0] node17684;
	wire [4-1:0] node17685;
	wire [4-1:0] node17686;
	wire [4-1:0] node17691;
	wire [4-1:0] node17693;
	wire [4-1:0] node17695;
	wire [4-1:0] node17698;
	wire [4-1:0] node17699;
	wire [4-1:0] node17700;
	wire [4-1:0] node17701;
	wire [4-1:0] node17704;
	wire [4-1:0] node17705;
	wire [4-1:0] node17708;
	wire [4-1:0] node17711;
	wire [4-1:0] node17712;
	wire [4-1:0] node17715;
	wire [4-1:0] node17717;
	wire [4-1:0] node17720;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17726;
	wire [4-1:0] node17729;
	wire [4-1:0] node17730;
	wire [4-1:0] node17731;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17737;
	wire [4-1:0] node17740;
	wire [4-1:0] node17741;
	wire [4-1:0] node17742;
	wire [4-1:0] node17743;
	wire [4-1:0] node17746;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17753;
	wire [4-1:0] node17756;
	wire [4-1:0] node17758;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17764;
	wire [4-1:0] node17769;
	wire [4-1:0] node17770;
	wire [4-1:0] node17771;
	wire [4-1:0] node17774;
	wire [4-1:0] node17777;
	wire [4-1:0] node17778;
	wire [4-1:0] node17779;
	wire [4-1:0] node17782;
	wire [4-1:0] node17786;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17789;
	wire [4-1:0] node17790;
	wire [4-1:0] node17794;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17801;
	wire [4-1:0] node17802;
	wire [4-1:0] node17803;
	wire [4-1:0] node17804;
	wire [4-1:0] node17808;
	wire [4-1:0] node17809;
	wire [4-1:0] node17813;
	wire [4-1:0] node17816;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17820;
	wire [4-1:0] node17825;
	wire [4-1:0] node17826;
	wire [4-1:0] node17828;
	wire [4-1:0] node17831;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17837;
	wire [4-1:0] node17839;
	wire [4-1:0] node17841;
	wire [4-1:0] node17844;
	wire [4-1:0] node17845;
	wire [4-1:0] node17846;
	wire [4-1:0] node17850;
	wire [4-1:0] node17852;
	wire [4-1:0] node17855;
	wire [4-1:0] node17856;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17859;
	wire [4-1:0] node17860;
	wire [4-1:0] node17863;
	wire [4-1:0] node17866;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17872;
	wire [4-1:0] node17875;
	wire [4-1:0] node17876;
	wire [4-1:0] node17877;
	wire [4-1:0] node17878;
	wire [4-1:0] node17881;
	wire [4-1:0] node17884;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17893;
	wire [4-1:0] node17894;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17900;
	wire [4-1:0] node17901;
	wire [4-1:0] node17904;
	wire [4-1:0] node17905;
	wire [4-1:0] node17908;
	wire [4-1:0] node17911;
	wire [4-1:0] node17912;
	wire [4-1:0] node17914;
	wire [4-1:0] node17917;
	wire [4-1:0] node17920;
	wire [4-1:0] node17921;
	wire [4-1:0] node17922;
	wire [4-1:0] node17925;
	wire [4-1:0] node17928;
	wire [4-1:0] node17929;
	wire [4-1:0] node17932;
	wire [4-1:0] node17935;
	wire [4-1:0] node17936;
	wire [4-1:0] node17937;
	wire [4-1:0] node17939;
	wire [4-1:0] node17941;
	wire [4-1:0] node17944;
	wire [4-1:0] node17945;
	wire [4-1:0] node17947;
	wire [4-1:0] node17949;
	wire [4-1:0] node17952;
	wire [4-1:0] node17953;
	wire [4-1:0] node17956;
	wire [4-1:0] node17958;
	wire [4-1:0] node17961;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17965;
	wire [4-1:0] node17968;
	wire [4-1:0] node17971;
	wire [4-1:0] node17974;
	wire [4-1:0] node17975;
	wire [4-1:0] node17978;
	wire [4-1:0] node17979;
	wire [4-1:0] node17982;
	wire [4-1:0] node17985;
	wire [4-1:0] node17986;
	wire [4-1:0] node17987;
	wire [4-1:0] node17988;
	wire [4-1:0] node17991;
	wire [4-1:0] node17995;
	wire [4-1:0] node17997;
	wire [4-1:0] node17998;
	wire [4-1:0] node18002;
	wire [4-1:0] node18003;
	wire [4-1:0] node18004;
	wire [4-1:0] node18005;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18008;
	wire [4-1:0] node18010;
	wire [4-1:0] node18012;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18019;
	wire [4-1:0] node18020;
	wire [4-1:0] node18024;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18029;
	wire [4-1:0] node18031;
	wire [4-1:0] node18034;
	wire [4-1:0] node18035;
	wire [4-1:0] node18036;
	wire [4-1:0] node18040;
	wire [4-1:0] node18043;
	wire [4-1:0] node18044;
	wire [4-1:0] node18045;
	wire [4-1:0] node18046;
	wire [4-1:0] node18048;
	wire [4-1:0] node18052;
	wire [4-1:0] node18053;
	wire [4-1:0] node18054;
	wire [4-1:0] node18058;
	wire [4-1:0] node18061;
	wire [4-1:0] node18062;
	wire [4-1:0] node18063;
	wire [4-1:0] node18066;
	wire [4-1:0] node18067;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18075;
	wire [4-1:0] node18077;
	wire [4-1:0] node18080;
	wire [4-1:0] node18081;
	wire [4-1:0] node18082;
	wire [4-1:0] node18083;
	wire [4-1:0] node18084;
	wire [4-1:0] node18086;
	wire [4-1:0] node18090;
	wire [4-1:0] node18091;
	wire [4-1:0] node18094;
	wire [4-1:0] node18097;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18101;
	wire [4-1:0] node18104;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18114;
	wire [4-1:0] node18115;
	wire [4-1:0] node18117;
	wire [4-1:0] node18120;
	wire [4-1:0] node18122;
	wire [4-1:0] node18125;
	wire [4-1:0] node18127;
	wire [4-1:0] node18130;
	wire [4-1:0] node18131;
	wire [4-1:0] node18133;
	wire [4-1:0] node18136;
	wire [4-1:0] node18138;
	wire [4-1:0] node18141;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18147;
	wire [4-1:0] node18150;
	wire [4-1:0] node18151;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18159;
	wire [4-1:0] node18160;
	wire [4-1:0] node18162;
	wire [4-1:0] node18165;
	wire [4-1:0] node18167;
	wire [4-1:0] node18168;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18174;
	wire [4-1:0] node18176;
	wire [4-1:0] node18178;
	wire [4-1:0] node18181;
	wire [4-1:0] node18183;
	wire [4-1:0] node18185;
	wire [4-1:0] node18188;
	wire [4-1:0] node18189;
	wire [4-1:0] node18190;
	wire [4-1:0] node18192;
	wire [4-1:0] node18196;
	wire [4-1:0] node18198;
	wire [4-1:0] node18201;
	wire [4-1:0] node18202;
	wire [4-1:0] node18203;
	wire [4-1:0] node18204;
	wire [4-1:0] node18205;
	wire [4-1:0] node18207;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18215;
	wire [4-1:0] node18217;
	wire [4-1:0] node18218;
	wire [4-1:0] node18222;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18228;
	wire [4-1:0] node18229;
	wire [4-1:0] node18231;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18238;
	wire [4-1:0] node18241;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18246;
	wire [4-1:0] node18247;
	wire [4-1:0] node18249;
	wire [4-1:0] node18253;
	wire [4-1:0] node18254;
	wire [4-1:0] node18256;
	wire [4-1:0] node18259;
	wire [4-1:0] node18260;
	wire [4-1:0] node18262;
	wire [4-1:0] node18265;
	wire [4-1:0] node18268;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18271;
	wire [4-1:0] node18272;
	wire [4-1:0] node18273;
	wire [4-1:0] node18275;
	wire [4-1:0] node18277;
	wire [4-1:0] node18280;
	wire [4-1:0] node18281;
	wire [4-1:0] node18282;
	wire [4-1:0] node18285;
	wire [4-1:0] node18289;
	wire [4-1:0] node18290;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18295;
	wire [4-1:0] node18299;
	wire [4-1:0] node18300;
	wire [4-1:0] node18303;
	wire [4-1:0] node18306;
	wire [4-1:0] node18307;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18313;
	wire [4-1:0] node18316;
	wire [4-1:0] node18318;
	wire [4-1:0] node18321;
	wire [4-1:0] node18322;
	wire [4-1:0] node18323;
	wire [4-1:0] node18327;
	wire [4-1:0] node18328;
	wire [4-1:0] node18332;
	wire [4-1:0] node18333;
	wire [4-1:0] node18335;
	wire [4-1:0] node18336;
	wire [4-1:0] node18339;
	wire [4-1:0] node18342;
	wire [4-1:0] node18343;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18349;
	wire [4-1:0] node18350;
	wire [4-1:0] node18353;
	wire [4-1:0] node18354;
	wire [4-1:0] node18356;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18364;
	wire [4-1:0] node18365;
	wire [4-1:0] node18366;
	wire [4-1:0] node18368;
	wire [4-1:0] node18371;
	wire [4-1:0] node18374;
	wire [4-1:0] node18375;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18381;
	wire [4-1:0] node18382;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18389;
	wire [4-1:0] node18392;
	wire [4-1:0] node18395;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18400;
	wire [4-1:0] node18401;
	wire [4-1:0] node18405;
	wire [4-1:0] node18406;
	wire [4-1:0] node18409;
	wire [4-1:0] node18412;
	wire [4-1:0] node18413;
	wire [4-1:0] node18414;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18420;
	wire [4-1:0] node18423;
	wire [4-1:0] node18425;
	wire [4-1:0] node18426;
	wire [4-1:0] node18430;
	wire [4-1:0] node18431;
	wire [4-1:0] node18432;
	wire [4-1:0] node18435;
	wire [4-1:0] node18436;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18451;
	wire [4-1:0] node18454;
	wire [4-1:0] node18456;
	wire [4-1:0] node18459;
	wire [4-1:0] node18460;
	wire [4-1:0] node18461;
	wire [4-1:0] node18462;
	wire [4-1:0] node18466;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18474;
	wire [4-1:0] node18475;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18482;
	wire [4-1:0] node18485;
	wire [4-1:0] node18487;
	wire [4-1:0] node18490;
	wire [4-1:0] node18491;
	wire [4-1:0] node18492;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18501;
	wire [4-1:0] node18502;
	wire [4-1:0] node18503;
	wire [4-1:0] node18506;
	wire [4-1:0] node18508;
	wire [4-1:0] node18511;
	wire [4-1:0] node18513;
	wire [4-1:0] node18516;
	wire [4-1:0] node18517;
	wire [4-1:0] node18518;
	wire [4-1:0] node18519;
	wire [4-1:0] node18521;
	wire [4-1:0] node18525;
	wire [4-1:0] node18526;
	wire [4-1:0] node18527;
	wire [4-1:0] node18530;
	wire [4-1:0] node18533;
	wire [4-1:0] node18535;
	wire [4-1:0] node18538;
	wire [4-1:0] node18539;
	wire [4-1:0] node18541;
	wire [4-1:0] node18544;
	wire [4-1:0] node18546;
	wire [4-1:0] node18547;
	wire [4-1:0] node18551;
	wire [4-1:0] node18552;
	wire [4-1:0] node18553;
	wire [4-1:0] node18554;
	wire [4-1:0] node18555;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18558;
	wire [4-1:0] node18559;
	wire [4-1:0] node18560;
	wire [4-1:0] node18563;
	wire [4-1:0] node18566;
	wire [4-1:0] node18569;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18575;
	wire [4-1:0] node18578;
	wire [4-1:0] node18579;
	wire [4-1:0] node18580;
	wire [4-1:0] node18581;
	wire [4-1:0] node18584;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18592;
	wire [4-1:0] node18593;
	wire [4-1:0] node18595;
	wire [4-1:0] node18599;
	wire [4-1:0] node18600;
	wire [4-1:0] node18601;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18607;
	wire [4-1:0] node18610;
	wire [4-1:0] node18611;
	wire [4-1:0] node18615;
	wire [4-1:0] node18616;
	wire [4-1:0] node18617;
	wire [4-1:0] node18618;
	wire [4-1:0] node18622;
	wire [4-1:0] node18625;
	wire [4-1:0] node18626;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18633;
	wire [4-1:0] node18635;
	wire [4-1:0] node18638;
	wire [4-1:0] node18639;
	wire [4-1:0] node18640;
	wire [4-1:0] node18642;
	wire [4-1:0] node18643;
	wire [4-1:0] node18646;
	wire [4-1:0] node18649;
	wire [4-1:0] node18650;
	wire [4-1:0] node18651;
	wire [4-1:0] node18653;
	wire [4-1:0] node18656;
	wire [4-1:0] node18657;
	wire [4-1:0] node18661;
	wire [4-1:0] node18664;
	wire [4-1:0] node18665;
	wire [4-1:0] node18666;
	wire [4-1:0] node18668;
	wire [4-1:0] node18671;
	wire [4-1:0] node18673;
	wire [4-1:0] node18674;
	wire [4-1:0] node18678;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18682;
	wire [4-1:0] node18685;
	wire [4-1:0] node18688;
	wire [4-1:0] node18689;
	wire [4-1:0] node18691;
	wire [4-1:0] node18694;
	wire [4-1:0] node18696;
	wire [4-1:0] node18699;
	wire [4-1:0] node18700;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18703;
	wire [4-1:0] node18704;
	wire [4-1:0] node18707;
	wire [4-1:0] node18709;
	wire [4-1:0] node18712;
	wire [4-1:0] node18713;
	wire [4-1:0] node18716;
	wire [4-1:0] node18717;
	wire [4-1:0] node18720;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18727;
	wire [4-1:0] node18731;
	wire [4-1:0] node18732;
	wire [4-1:0] node18735;
	wire [4-1:0] node18738;
	wire [4-1:0] node18739;
	wire [4-1:0] node18740;
	wire [4-1:0] node18741;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18748;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18756;
	wire [4-1:0] node18757;
	wire [4-1:0] node18758;
	wire [4-1:0] node18760;
	wire [4-1:0] node18763;
	wire [4-1:0] node18766;
	wire [4-1:0] node18768;
	wire [4-1:0] node18769;
	wire [4-1:0] node18773;
	wire [4-1:0] node18774;
	wire [4-1:0] node18775;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18780;
	wire [4-1:0] node18781;
	wire [4-1:0] node18784;
	wire [4-1:0] node18787;
	wire [4-1:0] node18789;
	wire [4-1:0] node18792;
	wire [4-1:0] node18793;
	wire [4-1:0] node18795;
	wire [4-1:0] node18796;
	wire [4-1:0] node18800;
	wire [4-1:0] node18801;
	wire [4-1:0] node18803;
	wire [4-1:0] node18806;
	wire [4-1:0] node18807;
	wire [4-1:0] node18811;
	wire [4-1:0] node18812;
	wire [4-1:0] node18813;
	wire [4-1:0] node18814;
	wire [4-1:0] node18817;
	wire [4-1:0] node18820;
	wire [4-1:0] node18821;
	wire [4-1:0] node18824;
	wire [4-1:0] node18825;
	wire [4-1:0] node18829;
	wire [4-1:0] node18830;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18836;
	wire [4-1:0] node18837;
	wire [4-1:0] node18840;
	wire [4-1:0] node18843;
	wire [4-1:0] node18844;
	wire [4-1:0] node18845;
	wire [4-1:0] node18849;
	wire [4-1:0] node18851;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18856;
	wire [4-1:0] node18857;
	wire [4-1:0] node18858;
	wire [4-1:0] node18859;
	wire [4-1:0] node18861;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18873;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18878;
	wire [4-1:0] node18882;
	wire [4-1:0] node18883;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18888;
	wire [4-1:0] node18890;
	wire [4-1:0] node18893;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18898;
	wire [4-1:0] node18901;
	wire [4-1:0] node18902;
	wire [4-1:0] node18905;
	wire [4-1:0] node18908;
	wire [4-1:0] node18909;
	wire [4-1:0] node18910;
	wire [4-1:0] node18912;
	wire [4-1:0] node18915;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18922;
	wire [4-1:0] node18925;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18930;
	wire [4-1:0] node18933;
	wire [4-1:0] node18935;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18940;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18946;
	wire [4-1:0] node18950;
	wire [4-1:0] node18951;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18958;
	wire [4-1:0] node18959;
	wire [4-1:0] node18963;
	wire [4-1:0] node18965;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18972;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18978;
	wire [4-1:0] node18981;
	wire [4-1:0] node18983;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18990;
	wire [4-1:0] node18991;
	wire [4-1:0] node18992;
	wire [4-1:0] node18996;
	wire [4-1:0] node18998;
	wire [4-1:0] node19001;
	wire [4-1:0] node19002;
	wire [4-1:0] node19005;
	wire [4-1:0] node19006;
	wire [4-1:0] node19010;
	wire [4-1:0] node19011;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19017;
	wire [4-1:0] node19020;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19027;
	wire [4-1:0] node19028;
	wire [4-1:0] node19029;
	wire [4-1:0] node19031;
	wire [4-1:0] node19034;
	wire [4-1:0] node19035;
	wire [4-1:0] node19038;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19044;
	wire [4-1:0] node19046;
	wire [4-1:0] node19049;
	wire [4-1:0] node19050;
	wire [4-1:0] node19054;
	wire [4-1:0] node19055;
	wire [4-1:0] node19056;
	wire [4-1:0] node19057;
	wire [4-1:0] node19058;
	wire [4-1:0] node19061;
	wire [4-1:0] node19065;
	wire [4-1:0] node19066;
	wire [4-1:0] node19068;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19077;
	wire [4-1:0] node19080;
	wire [4-1:0] node19081;
	wire [4-1:0] node19082;
	wire [4-1:0] node19085;
	wire [4-1:0] node19086;
	wire [4-1:0] node19087;
	wire [4-1:0] node19091;
	wire [4-1:0] node19094;
	wire [4-1:0] node19095;
	wire [4-1:0] node19096;
	wire [4-1:0] node19100;
	wire [4-1:0] node19102;
	wire [4-1:0] node19103;
	wire [4-1:0] node19107;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19113;
	wire [4-1:0] node19115;
	wire [4-1:0] node19116;
	wire [4-1:0] node19120;
	wire [4-1:0] node19121;
	wire [4-1:0] node19123;
	wire [4-1:0] node19126;
	wire [4-1:0] node19127;
	wire [4-1:0] node19130;
	wire [4-1:0] node19133;
	wire [4-1:0] node19134;
	wire [4-1:0] node19138;
	wire [4-1:0] node19139;
	wire [4-1:0] node19140;
	wire [4-1:0] node19141;
	wire [4-1:0] node19142;
	wire [4-1:0] node19145;
	wire [4-1:0] node19148;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19154;
	wire [4-1:0] node19157;
	wire [4-1:0] node19158;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19164;
	wire [4-1:0] node19168;
	wire [4-1:0] node19169;
	wire [4-1:0] node19172;
	wire [4-1:0] node19175;
	wire [4-1:0] node19176;
	wire [4-1:0] node19177;
	wire [4-1:0] node19178;
	wire [4-1:0] node19179;
	wire [4-1:0] node19182;
	wire [4-1:0] node19185;
	wire [4-1:0] node19187;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19192;
	wire [4-1:0] node19193;
	wire [4-1:0] node19198;
	wire [4-1:0] node19199;
	wire [4-1:0] node19200;
	wire [4-1:0] node19203;
	wire [4-1:0] node19206;
	wire [4-1:0] node19208;
	wire [4-1:0] node19211;
	wire [4-1:0] node19212;
	wire [4-1:0] node19213;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19220;
	wire [4-1:0] node19221;
	wire [4-1:0] node19222;
	wire [4-1:0] node19226;
	wire [4-1:0] node19229;
	wire [4-1:0] node19230;
	wire [4-1:0] node19231;
	wire [4-1:0] node19233;
	wire [4-1:0] node19236;
	wire [4-1:0] node19238;
	wire [4-1:0] node19241;
	wire [4-1:0] node19242;
	wire [4-1:0] node19243;
	wire [4-1:0] node19246;
	wire [4-1:0] node19249;
	wire [4-1:0] node19250;
	wire [4-1:0] node19253;
	wire [4-1:0] node19256;
	wire [4-1:0] node19257;
	wire [4-1:0] node19258;
	wire [4-1:0] node19259;
	wire [4-1:0] node19260;
	wire [4-1:0] node19261;
	wire [4-1:0] node19262;
	wire [4-1:0] node19265;
	wire [4-1:0] node19268;
	wire [4-1:0] node19270;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19281;
	wire [4-1:0] node19282;
	wire [4-1:0] node19285;
	wire [4-1:0] node19288;
	wire [4-1:0] node19289;
	wire [4-1:0] node19292;
	wire [4-1:0] node19295;
	wire [4-1:0] node19296;
	wire [4-1:0] node19297;
	wire [4-1:0] node19298;
	wire [4-1:0] node19300;
	wire [4-1:0] node19303;
	wire [4-1:0] node19305;
	wire [4-1:0] node19308;
	wire [4-1:0] node19309;
	wire [4-1:0] node19312;
	wire [4-1:0] node19314;
	wire [4-1:0] node19317;
	wire [4-1:0] node19318;
	wire [4-1:0] node19319;
	wire [4-1:0] node19320;
	wire [4-1:0] node19323;
	wire [4-1:0] node19326;
	wire [4-1:0] node19328;
	wire [4-1:0] node19331;
	wire [4-1:0] node19333;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19338;
	wire [4-1:0] node19339;
	wire [4-1:0] node19340;
	wire [4-1:0] node19341;
	wire [4-1:0] node19345;
	wire [4-1:0] node19346;
	wire [4-1:0] node19350;
	wire [4-1:0] node19351;
	wire [4-1:0] node19354;
	wire [4-1:0] node19355;
	wire [4-1:0] node19358;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19366;
	wire [4-1:0] node19367;
	wire [4-1:0] node19370;
	wire [4-1:0] node19373;
	wire [4-1:0] node19374;
	wire [4-1:0] node19376;
	wire [4-1:0] node19379;
	wire [4-1:0] node19382;
	wire [4-1:0] node19383;
	wire [4-1:0] node19384;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19389;
	wire [4-1:0] node19392;
	wire [4-1:0] node19393;
	wire [4-1:0] node19397;
	wire [4-1:0] node19399;
	wire [4-1:0] node19402;
	wire [4-1:0] node19403;
	wire [4-1:0] node19404;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19411;
	wire [4-1:0] node19414;
	wire [4-1:0] node19415;
	wire [4-1:0] node19416;
	wire [4-1:0] node19419;
	wire [4-1:0] node19422;
	wire [4-1:0] node19424;
	wire [4-1:0] node19427;
	wire [4-1:0] node19428;
	wire [4-1:0] node19429;
	wire [4-1:0] node19430;
	wire [4-1:0] node19431;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19437;
	wire [4-1:0] node19439;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19444;
	wire [4-1:0] node19445;
	wire [4-1:0] node19448;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19456;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19461;
	wire [4-1:0] node19463;
	wire [4-1:0] node19464;
	wire [4-1:0] node19467;
	wire [4-1:0] node19470;
	wire [4-1:0] node19471;
	wire [4-1:0] node19472;
	wire [4-1:0] node19475;
	wire [4-1:0] node19479;
	wire [4-1:0] node19480;
	wire [4-1:0] node19481;
	wire [4-1:0] node19482;
	wire [4-1:0] node19485;
	wire [4-1:0] node19489;
	wire [4-1:0] node19490;
	wire [4-1:0] node19491;
	wire [4-1:0] node19494;
	wire [4-1:0] node19497;
	wire [4-1:0] node19498;
	wire [4-1:0] node19501;
	wire [4-1:0] node19504;
	wire [4-1:0] node19505;
	wire [4-1:0] node19506;
	wire [4-1:0] node19507;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19518;
	wire [4-1:0] node19522;
	wire [4-1:0] node19525;
	wire [4-1:0] node19526;
	wire [4-1:0] node19527;
	wire [4-1:0] node19528;
	wire [4-1:0] node19529;
	wire [4-1:0] node19531;
	wire [4-1:0] node19534;
	wire [4-1:0] node19536;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19541;
	wire [4-1:0] node19544;
	wire [4-1:0] node19547;
	wire [4-1:0] node19548;
	wire [4-1:0] node19551;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19556;
	wire [4-1:0] node19557;
	wire [4-1:0] node19560;
	wire [4-1:0] node19563;
	wire [4-1:0] node19564;
	wire [4-1:0] node19565;
	wire [4-1:0] node19569;
	wire [4-1:0] node19571;
	wire [4-1:0] node19574;
	wire [4-1:0] node19575;
	wire [4-1:0] node19578;
	wire [4-1:0] node19581;
	wire [4-1:0] node19582;
	wire [4-1:0] node19583;
	wire [4-1:0] node19586;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19593;
	wire [4-1:0] node19597;
	wire [4-1:0] node19598;
	wire [4-1:0] node19599;
	wire [4-1:0] node19602;
	wire [4-1:0] node19605;
	wire [4-1:0] node19608;
	wire [4-1:0] node19609;
	wire [4-1:0] node19610;
	wire [4-1:0] node19611;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19622;
	wire [4-1:0] node19626;
	wire [4-1:0] node19629;
	wire [4-1:0] node19630;
	wire [4-1:0] node19631;
	wire [4-1:0] node19634;
	wire [4-1:0] node19635;
	wire [4-1:0] node19640;
	wire [4-1:0] node19641;
	wire [4-1:0] node19642;
	wire [4-1:0] node19644;
	wire [4-1:0] node19646;
	wire [4-1:0] node19649;
	wire [4-1:0] node19651;
	wire [4-1:0] node19652;
	wire [4-1:0] node19656;
	wire [4-1:0] node19657;
	wire [4-1:0] node19658;
	wire [4-1:0] node19662;
	wire [4-1:0] node19663;
	wire [4-1:0] node19664;
	wire [4-1:0] node19667;
	wire [4-1:0] node19670;
	wire [4-1:0] node19671;
	wire [4-1:0] node19675;
	wire [4-1:0] node19676;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19679;
	wire [4-1:0] node19680;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19689;
	wire [4-1:0] node19691;
	wire [4-1:0] node19692;
	wire [4-1:0] node19695;
	wire [4-1:0] node19698;
	wire [4-1:0] node19699;
	wire [4-1:0] node19700;
	wire [4-1:0] node19702;
	wire [4-1:0] node19705;
	wire [4-1:0] node19708;
	wire [4-1:0] node19709;
	wire [4-1:0] node19711;
	wire [4-1:0] node19714;
	wire [4-1:0] node19717;
	wire [4-1:0] node19718;
	wire [4-1:0] node19719;
	wire [4-1:0] node19721;
	wire [4-1:0] node19722;
	wire [4-1:0] node19726;
	wire [4-1:0] node19727;
	wire [4-1:0] node19728;
	wire [4-1:0] node19731;
	wire [4-1:0] node19735;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19739;
	wire [4-1:0] node19743;
	wire [4-1:0] node19746;
	wire [4-1:0] node19747;
	wire [4-1:0] node19748;
	wire [4-1:0] node19749;
	wire [4-1:0] node19750;
	wire [4-1:0] node19751;
	wire [4-1:0] node19752;
	wire [4-1:0] node19755;
	wire [4-1:0] node19759;
	wire [4-1:0] node19760;
	wire [4-1:0] node19762;
	wire [4-1:0] node19766;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19771;
	wire [4-1:0] node19774;
	wire [4-1:0] node19775;
	wire [4-1:0] node19778;
	wire [4-1:0] node19781;
	wire [4-1:0] node19782;
	wire [4-1:0] node19783;
	wire [4-1:0] node19786;
	wire [4-1:0] node19787;
	wire [4-1:0] node19788;
	wire [4-1:0] node19793;
	wire [4-1:0] node19794;
	wire [4-1:0] node19795;
	wire [4-1:0] node19796;
	wire [4-1:0] node19799;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19806;
	wire [4-1:0] node19809;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19814;
	wire [4-1:0] node19815;
	wire [4-1:0] node19817;
	wire [4-1:0] node19818;
	wire [4-1:0] node19822;
	wire [4-1:0] node19823;
	wire [4-1:0] node19827;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19837;
	wire [4-1:0] node19838;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19846;
	wire [4-1:0] node19847;
	wire [4-1:0] node19848;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19854;
	wire [4-1:0] node19855;
	wire [4-1:0] node19858;
	wire [4-1:0] node19861;
	wire [4-1:0] node19863;
	wire [4-1:0] node19864;
	wire [4-1:0] node19868;
	wire [4-1:0] node19869;
	wire [4-1:0] node19870;
	wire [4-1:0] node19874;
	wire [4-1:0] node19875;
	wire [4-1:0] node19876;
	wire [4-1:0] node19880;
	wire [4-1:0] node19881;
	wire [4-1:0] node19885;
	wire [4-1:0] node19886;
	wire [4-1:0] node19887;
	wire [4-1:0] node19888;
	wire [4-1:0] node19889;
	wire [4-1:0] node19890;
	wire [4-1:0] node19891;
	wire [4-1:0] node19894;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19899;
	wire [4-1:0] node19903;
	wire [4-1:0] node19905;
	wire [4-1:0] node19908;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19914;
	wire [4-1:0] node19915;
	wire [4-1:0] node19917;
	wire [4-1:0] node19920;
	wire [4-1:0] node19922;
	wire [4-1:0] node19925;
	wire [4-1:0] node19926;
	wire [4-1:0] node19927;
	wire [4-1:0] node19928;
	wire [4-1:0] node19931;
	wire [4-1:0] node19935;
	wire [4-1:0] node19936;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19941;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19949;
	wire [4-1:0] node19950;
	wire [4-1:0] node19953;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19958;
	wire [4-1:0] node19959;
	wire [4-1:0] node19960;
	wire [4-1:0] node19962;
	wire [4-1:0] node19966;
	wire [4-1:0] node19967;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19979;
	wire [4-1:0] node19981;
	wire [4-1:0] node19982;
	wire [4-1:0] node19985;
	wire [4-1:0] node19988;
	wire [4-1:0] node19989;
	wire [4-1:0] node19990;
	wire [4-1:0] node19991;
	wire [4-1:0] node19993;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node20001;
	wire [4-1:0] node20004;
	wire [4-1:0] node20005;
	wire [4-1:0] node20006;
	wire [4-1:0] node20008;
	wire [4-1:0] node20011;
	wire [4-1:0] node20012;
	wire [4-1:0] node20017;
	wire [4-1:0] node20018;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20024;
	wire [4-1:0] node20026;
	wire [4-1:0] node20028;
	wire [4-1:0] node20031;
	wire [4-1:0] node20032;
	wire [4-1:0] node20033;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20040;
	wire [4-1:0] node20043;
	wire [4-1:0] node20045;
	wire [4-1:0] node20047;
	wire [4-1:0] node20050;
	wire [4-1:0] node20051;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20054;
	wire [4-1:0] node20057;
	wire [4-1:0] node20061;
	wire [4-1:0] node20062;
	wire [4-1:0] node20064;
	wire [4-1:0] node20068;
	wire [4-1:0] node20069;
	wire [4-1:0] node20070;
	wire [4-1:0] node20074;
	wire [4-1:0] node20075;
	wire [4-1:0] node20076;
	wire [4-1:0] node20079;
	wire [4-1:0] node20082;
	wire [4-1:0] node20084;
	wire [4-1:0] node20087;
	wire [4-1:0] node20088;
	wire [4-1:0] node20089;
	wire [4-1:0] node20090;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20095;
	wire [4-1:0] node20099;
	wire [4-1:0] node20100;
	wire [4-1:0] node20103;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20109;
	wire [4-1:0] node20112;
	wire [4-1:0] node20113;
	wire [4-1:0] node20115;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20122;
	wire [4-1:0] node20125;
	wire [4-1:0] node20127;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20140;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20146;
	wire [4-1:0] node20147;
	wire [4-1:0] node20150;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20156;
	wire [4-1:0] node20159;
	wire [4-1:0] node20160;
	wire [4-1:0] node20164;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20167;
	wire [4-1:0] node20168;
	wire [4-1:0] node20169;
	wire [4-1:0] node20170;
	wire [4-1:0] node20173;
	wire [4-1:0] node20175;
	wire [4-1:0] node20176;
	wire [4-1:0] node20180;
	wire [4-1:0] node20181;
	wire [4-1:0] node20183;
	wire [4-1:0] node20184;
	wire [4-1:0] node20188;
	wire [4-1:0] node20189;
	wire [4-1:0] node20190;
	wire [4-1:0] node20194;
	wire [4-1:0] node20197;
	wire [4-1:0] node20198;
	wire [4-1:0] node20199;
	wire [4-1:0] node20200;
	wire [4-1:0] node20204;
	wire [4-1:0] node20205;
	wire [4-1:0] node20207;
	wire [4-1:0] node20211;
	wire [4-1:0] node20212;
	wire [4-1:0] node20213;
	wire [4-1:0] node20217;
	wire [4-1:0] node20218;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20230;
	wire [4-1:0] node20232;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20237;
	wire [4-1:0] node20238;
	wire [4-1:0] node20242;
	wire [4-1:0] node20244;
	wire [4-1:0] node20247;
	wire [4-1:0] node20249;
	wire [4-1:0] node20251;
	wire [4-1:0] node20254;
	wire [4-1:0] node20255;
	wire [4-1:0] node20256;
	wire [4-1:0] node20258;
	wire [4-1:0] node20259;
	wire [4-1:0] node20262;
	wire [4-1:0] node20265;
	wire [4-1:0] node20267;
	wire [4-1:0] node20268;
	wire [4-1:0] node20272;
	wire [4-1:0] node20273;
	wire [4-1:0] node20275;
	wire [4-1:0] node20278;
	wire [4-1:0] node20279;
	wire [4-1:0] node20282;
	wire [4-1:0] node20283;
	wire [4-1:0] node20287;
	wire [4-1:0] node20288;
	wire [4-1:0] node20289;
	wire [4-1:0] node20290;
	wire [4-1:0] node20292;
	wire [4-1:0] node20293;
	wire [4-1:0] node20294;
	wire [4-1:0] node20297;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20304;
	wire [4-1:0] node20306;
	wire [4-1:0] node20309;
	wire [4-1:0] node20311;
	wire [4-1:0] node20314;
	wire [4-1:0] node20315;
	wire [4-1:0] node20316;
	wire [4-1:0] node20317;
	wire [4-1:0] node20320;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20327;
	wire [4-1:0] node20330;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20338;
	wire [4-1:0] node20341;
	wire [4-1:0] node20342;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20346;
	wire [4-1:0] node20349;
	wire [4-1:0] node20351;
	wire [4-1:0] node20354;
	wire [4-1:0] node20355;
	wire [4-1:0] node20356;
	wire [4-1:0] node20360;
	wire [4-1:0] node20363;
	wire [4-1:0] node20364;
	wire [4-1:0] node20365;
	wire [4-1:0] node20366;
	wire [4-1:0] node20367;
	wire [4-1:0] node20372;
	wire [4-1:0] node20373;
	wire [4-1:0] node20374;
	wire [4-1:0] node20378;
	wire [4-1:0] node20379;
	wire [4-1:0] node20383;
	wire [4-1:0] node20384;
	wire [4-1:0] node20385;
	wire [4-1:0] node20386;
	wire [4-1:0] node20389;
	wire [4-1:0] node20393;
	wire [4-1:0] node20394;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20401;
	wire [4-1:0] node20402;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20407;
	wire [4-1:0] node20410;
	wire [4-1:0] node20411;
	wire [4-1:0] node20412;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20425;
	wire [4-1:0] node20428;
	wire [4-1:0] node20429;
	wire [4-1:0] node20430;
	wire [4-1:0] node20431;
	wire [4-1:0] node20434;
	wire [4-1:0] node20438;
	wire [4-1:0] node20440;
	wire [4-1:0] node20441;
	wire [4-1:0] node20444;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20449;
	wire [4-1:0] node20450;
	wire [4-1:0] node20451;
	wire [4-1:0] node20452;
	wire [4-1:0] node20455;
	wire [4-1:0] node20458;
	wire [4-1:0] node20459;
	wire [4-1:0] node20463;
	wire [4-1:0] node20465;
	wire [4-1:0] node20467;
	wire [4-1:0] node20470;
	wire [4-1:0] node20471;
	wire [4-1:0] node20473;
	wire [4-1:0] node20476;
	wire [4-1:0] node20477;
	wire [4-1:0] node20478;
	wire [4-1:0] node20482;
	wire [4-1:0] node20483;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20490;
	wire [4-1:0] node20493;
	wire [4-1:0] node20496;
	wire [4-1:0] node20498;
	wire [4-1:0] node20501;
	wire [4-1:0] node20502;
	wire [4-1:0] node20503;
	wire [4-1:0] node20506;
	wire [4-1:0] node20509;
	wire [4-1:0] node20510;
	wire [4-1:0] node20511;
	wire [4-1:0] node20514;
	wire [4-1:0] node20518;
	wire [4-1:0] node20519;
	wire [4-1:0] node20520;
	wire [4-1:0] node20521;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20530;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20542;
	wire [4-1:0] node20545;
	wire [4-1:0] node20546;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20550;
	wire [4-1:0] node20553;
	wire [4-1:0] node20556;
	wire [4-1:0] node20557;
	wire [4-1:0] node20561;
	wire [4-1:0] node20562;
	wire [4-1:0] node20563;
	wire [4-1:0] node20567;
	wire [4-1:0] node20568;
	wire [4-1:0] node20569;
	wire [4-1:0] node20573;
	wire [4-1:0] node20576;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20579;
	wire [4-1:0] node20581;
	wire [4-1:0] node20582;
	wire [4-1:0] node20585;
	wire [4-1:0] node20588;
	wire [4-1:0] node20589;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20595;
	wire [4-1:0] node20600;
	wire [4-1:0] node20601;
	wire [4-1:0] node20602;
	wire [4-1:0] node20604;
	wire [4-1:0] node20606;
	wire [4-1:0] node20609;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20615;
	wire [4-1:0] node20618;
	wire [4-1:0] node20619;
	wire [4-1:0] node20621;
	wire [4-1:0] node20624;
	wire [4-1:0] node20625;
	wire [4-1:0] node20629;
	wire [4-1:0] node20630;
	wire [4-1:0] node20631;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20634;
	wire [4-1:0] node20635;
	wire [4-1:0] node20636;
	wire [4-1:0] node20637;
	wire [4-1:0] node20640;
	wire [4-1:0] node20643;
	wire [4-1:0] node20644;
	wire [4-1:0] node20645;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20653;
	wire [4-1:0] node20656;
	wire [4-1:0] node20657;
	wire [4-1:0] node20658;
	wire [4-1:0] node20662;
	wire [4-1:0] node20664;
	wire [4-1:0] node20667;
	wire [4-1:0] node20668;
	wire [4-1:0] node20669;
	wire [4-1:0] node20670;
	wire [4-1:0] node20673;
	wire [4-1:0] node20676;
	wire [4-1:0] node20678;
	wire [4-1:0] node20681;
	wire [4-1:0] node20682;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20688;
	wire [4-1:0] node20691;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20697;
	wire [4-1:0] node20699;
	wire [4-1:0] node20702;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20705;
	wire [4-1:0] node20706;
	wire [4-1:0] node20710;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20717;
	wire [4-1:0] node20718;
	wire [4-1:0] node20720;
	wire [4-1:0] node20721;
	wire [4-1:0] node20724;
	wire [4-1:0] node20727;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20732;
	wire [4-1:0] node20736;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20743;
	wire [4-1:0] node20745;
	wire [4-1:0] node20746;
	wire [4-1:0] node20750;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20755;
	wire [4-1:0] node20758;
	wire [4-1:0] node20760;
	wire [4-1:0] node20762;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20769;
	wire [4-1:0] node20771;
	wire [4-1:0] node20772;
	wire [4-1:0] node20776;
	wire [4-1:0] node20777;
	wire [4-1:0] node20778;
	wire [4-1:0] node20782;
	wire [4-1:0] node20783;
	wire [4-1:0] node20786;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20795;
	wire [4-1:0] node20798;
	wire [4-1:0] node20799;
	wire [4-1:0] node20802;
	wire [4-1:0] node20805;
	wire [4-1:0] node20806;
	wire [4-1:0] node20808;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20814;
	wire [4-1:0] node20815;
	wire [4-1:0] node20817;
	wire [4-1:0] node20820;
	wire [4-1:0] node20822;
	wire [4-1:0] node20825;
	wire [4-1:0] node20827;
	wire [4-1:0] node20828;
	wire [4-1:0] node20831;
	wire [4-1:0] node20834;
	wire [4-1:0] node20835;
	wire [4-1:0] node20837;
	wire [4-1:0] node20839;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20844;
	wire [4-1:0] node20847;
	wire [4-1:0] node20851;
	wire [4-1:0] node20852;
	wire [4-1:0] node20853;
	wire [4-1:0] node20854;
	wire [4-1:0] node20857;
	wire [4-1:0] node20858;
	wire [4-1:0] node20862;
	wire [4-1:0] node20863;
	wire [4-1:0] node20864;
	wire [4-1:0] node20867;
	wire [4-1:0] node20870;
	wire [4-1:0] node20871;
	wire [4-1:0] node20875;
	wire [4-1:0] node20876;
	wire [4-1:0] node20877;
	wire [4-1:0] node20878;
	wire [4-1:0] node20881;
	wire [4-1:0] node20882;
	wire [4-1:0] node20885;
	wire [4-1:0] node20888;
	wire [4-1:0] node20890;
	wire [4-1:0] node20893;
	wire [4-1:0] node20894;
	wire [4-1:0] node20895;
	wire [4-1:0] node20898;
	wire [4-1:0] node20899;
	wire [4-1:0] node20902;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20907;
	wire [4-1:0] node20911;
	wire [4-1:0] node20913;
	wire [4-1:0] node20916;
	wire [4-1:0] node20917;
	wire [4-1:0] node20918;
	wire [4-1:0] node20919;
	wire [4-1:0] node20920;
	wire [4-1:0] node20921;
	wire [4-1:0] node20923;
	wire [4-1:0] node20925;
	wire [4-1:0] node20929;
	wire [4-1:0] node20930;
	wire [4-1:0] node20931;
	wire [4-1:0] node20933;
	wire [4-1:0] node20936;
	wire [4-1:0] node20937;
	wire [4-1:0] node20940;
	wire [4-1:0] node20944;
	wire [4-1:0] node20945;
	wire [4-1:0] node20946;
	wire [4-1:0] node20948;
	wire [4-1:0] node20949;
	wire [4-1:0] node20953;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20959;
	wire [4-1:0] node20962;
	wire [4-1:0] node20964;
	wire [4-1:0] node20966;
	wire [4-1:0] node20969;
	wire [4-1:0] node20970;
	wire [4-1:0] node20971;
	wire [4-1:0] node20972;
	wire [4-1:0] node20973;
	wire [4-1:0] node20975;
	wire [4-1:0] node20978;
	wire [4-1:0] node20979;
	wire [4-1:0] node20982;
	wire [4-1:0] node20985;
	wire [4-1:0] node20987;
	wire [4-1:0] node20989;
	wire [4-1:0] node20992;
	wire [4-1:0] node20993;
	wire [4-1:0] node20995;
	wire [4-1:0] node20998;
	wire [4-1:0] node21000;
	wire [4-1:0] node21003;
	wire [4-1:0] node21004;
	wire [4-1:0] node21005;
	wire [4-1:0] node21006;
	wire [4-1:0] node21009;
	wire [4-1:0] node21012;
	wire [4-1:0] node21013;
	wire [4-1:0] node21014;
	wire [4-1:0] node21018;
	wire [4-1:0] node21019;
	wire [4-1:0] node21022;
	wire [4-1:0] node21025;
	wire [4-1:0] node21026;
	wire [4-1:0] node21027;
	wire [4-1:0] node21028;
	wire [4-1:0] node21032;
	wire [4-1:0] node21034;
	wire [4-1:0] node21037;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21042;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21050;
	wire [4-1:0] node21051;
	wire [4-1:0] node21052;
	wire [4-1:0] node21053;
	wire [4-1:0] node21054;
	wire [4-1:0] node21055;
	wire [4-1:0] node21056;
	wire [4-1:0] node21059;
	wire [4-1:0] node21063;
	wire [4-1:0] node21065;
	wire [4-1:0] node21066;
	wire [4-1:0] node21069;
	wire [4-1:0] node21072;
	wire [4-1:0] node21073;
	wire [4-1:0] node21075;
	wire [4-1:0] node21076;
	wire [4-1:0] node21080;
	wire [4-1:0] node21081;
	wire [4-1:0] node21084;
	wire [4-1:0] node21087;
	wire [4-1:0] node21088;
	wire [4-1:0] node21089;
	wire [4-1:0] node21090;
	wire [4-1:0] node21094;
	wire [4-1:0] node21096;
	wire [4-1:0] node21097;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21106;
	wire [4-1:0] node21109;
	wire [4-1:0] node21110;
	wire [4-1:0] node21113;
	wire [4-1:0] node21116;
	wire [4-1:0] node21117;
	wire [4-1:0] node21118;
	wire [4-1:0] node21119;
	wire [4-1:0] node21120;
	wire [4-1:0] node21124;
	wire [4-1:0] node21125;
	wire [4-1:0] node21127;
	wire [4-1:0] node21130;
	wire [4-1:0] node21131;
	wire [4-1:0] node21134;
	wire [4-1:0] node21137;
	wire [4-1:0] node21138;
	wire [4-1:0] node21140;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21151;
	wire [4-1:0] node21152;
	wire [4-1:0] node21155;
	wire [4-1:0] node21157;
	wire [4-1:0] node21160;
	wire [4-1:0] node21161;
	wire [4-1:0] node21162;
	wire [4-1:0] node21165;
	wire [4-1:0] node21168;
	wire [4-1:0] node21169;
	wire [4-1:0] node21173;
	wire [4-1:0] node21174;
	wire [4-1:0] node21175;
	wire [4-1:0] node21176;
	wire [4-1:0] node21177;
	wire [4-1:0] node21178;
	wire [4-1:0] node21179;
	wire [4-1:0] node21181;
	wire [4-1:0] node21182;
	wire [4-1:0] node21185;
	wire [4-1:0] node21188;
	wire [4-1:0] node21190;
	wire [4-1:0] node21193;
	wire [4-1:0] node21194;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21200;
	wire [4-1:0] node21203;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21212;
	wire [4-1:0] node21215;
	wire [4-1:0] node21216;
	wire [4-1:0] node21219;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21225;
	wire [4-1:0] node21227;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21234;
	wire [4-1:0] node21236;
	wire [4-1:0] node21239;
	wire [4-1:0] node21240;
	wire [4-1:0] node21241;
	wire [4-1:0] node21242;
	wire [4-1:0] node21243;
	wire [4-1:0] node21247;
	wire [4-1:0] node21248;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21256;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21260;
	wire [4-1:0] node21264;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21271;
	wire [4-1:0] node21272;
	wire [4-1:0] node21273;
	wire [4-1:0] node21274;
	wire [4-1:0] node21277;
	wire [4-1:0] node21280;
	wire [4-1:0] node21281;
	wire [4-1:0] node21284;
	wire [4-1:0] node21287;
	wire [4-1:0] node21288;
	wire [4-1:0] node21289;
	wire [4-1:0] node21290;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21299;
	wire [4-1:0] node21300;
	wire [4-1:0] node21301;
	wire [4-1:0] node21304;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21310;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21313;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21324;
	wire [4-1:0] node21325;
	wire [4-1:0] node21326;
	wire [4-1:0] node21329;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21337;
	wire [4-1:0] node21340;
	wire [4-1:0] node21342;
	wire [4-1:0] node21345;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21348;
	wire [4-1:0] node21349;
	wire [4-1:0] node21352;
	wire [4-1:0] node21356;
	wire [4-1:0] node21358;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21369;
	wire [4-1:0] node21372;
	wire [4-1:0] node21373;
	wire [4-1:0] node21374;
	wire [4-1:0] node21375;
	wire [4-1:0] node21376;
	wire [4-1:0] node21378;
	wire [4-1:0] node21381;
	wire [4-1:0] node21382;
	wire [4-1:0] node21386;
	wire [4-1:0] node21387;
	wire [4-1:0] node21390;
	wire [4-1:0] node21393;
	wire [4-1:0] node21394;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21399;
	wire [4-1:0] node21402;
	wire [4-1:0] node21403;
	wire [4-1:0] node21407;
	wire [4-1:0] node21409;
	wire [4-1:0] node21412;
	wire [4-1:0] node21413;
	wire [4-1:0] node21414;
	wire [4-1:0] node21415;
	wire [4-1:0] node21419;
	wire [4-1:0] node21420;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21427;
	wire [4-1:0] node21432;
	wire [4-1:0] node21435;
	wire [4-1:0] node21436;
	wire [4-1:0] node21437;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21440;
	wire [4-1:0] node21441;
	wire [4-1:0] node21442;
	wire [4-1:0] node21445;
	wire [4-1:0] node21448;
	wire [4-1:0] node21449;
	wire [4-1:0] node21452;
	wire [4-1:0] node21455;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21462;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21468;
	wire [4-1:0] node21472;
	wire [4-1:0] node21473;
	wire [4-1:0] node21476;
	wire [4-1:0] node21479;
	wire [4-1:0] node21480;
	wire [4-1:0] node21481;
	wire [4-1:0] node21482;
	wire [4-1:0] node21483;
	wire [4-1:0] node21486;
	wire [4-1:0] node21490;
	wire [4-1:0] node21491;
	wire [4-1:0] node21494;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21499;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21507;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21512;
	wire [4-1:0] node21516;
	wire [4-1:0] node21517;
	wire [4-1:0] node21518;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21523;
	wire [4-1:0] node21524;
	wire [4-1:0] node21528;
	wire [4-1:0] node21529;
	wire [4-1:0] node21532;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21543;
	wire [4-1:0] node21545;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21552;
	wire [4-1:0] node21553;
	wire [4-1:0] node21557;
	wire [4-1:0] node21558;
	wire [4-1:0] node21559;
	wire [4-1:0] node21562;
	wire [4-1:0] node21566;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21571;
	wire [4-1:0] node21572;
	wire [4-1:0] node21576;
	wire [4-1:0] node21578;
	wire [4-1:0] node21579;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21589;
	wire [4-1:0] node21591;
	wire [4-1:0] node21594;
	wire [4-1:0] node21596;
	wire [4-1:0] node21597;
	wire [4-1:0] node21601;
	wire [4-1:0] node21602;
	wire [4-1:0] node21604;
	wire [4-1:0] node21605;
	wire [4-1:0] node21608;
	wire [4-1:0] node21611;
	wire [4-1:0] node21612;
	wire [4-1:0] node21616;
	wire [4-1:0] node21617;
	wire [4-1:0] node21619;
	wire [4-1:0] node21621;
	wire [4-1:0] node21622;
	wire [4-1:0] node21626;
	wire [4-1:0] node21627;
	wire [4-1:0] node21628;
	wire [4-1:0] node21631;
	wire [4-1:0] node21634;
	wire [4-1:0] node21635;
	wire [4-1:0] node21639;
	wire [4-1:0] node21640;
	wire [4-1:0] node21641;
	wire [4-1:0] node21642;
	wire [4-1:0] node21643;
	wire [4-1:0] node21646;
	wire [4-1:0] node21648;
	wire [4-1:0] node21651;
	wire [4-1:0] node21652;
	wire [4-1:0] node21653;
	wire [4-1:0] node21658;
	wire [4-1:0] node21659;
	wire [4-1:0] node21660;
	wire [4-1:0] node21661;
	wire [4-1:0] node21664;
	wire [4-1:0] node21667;
	wire [4-1:0] node21668;
	wire [4-1:0] node21672;
	wire [4-1:0] node21673;
	wire [4-1:0] node21676;
	wire [4-1:0] node21679;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21684;
	wire [4-1:0] node21687;
	wire [4-1:0] node21688;
	wire [4-1:0] node21691;
	wire [4-1:0] node21694;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21700;
	wire [4-1:0] node21703;
	wire [4-1:0] node21704;
	wire [4-1:0] node21705;
	wire [4-1:0] node21706;
	wire [4-1:0] node21709;
	wire [4-1:0] node21713;
	wire [4-1:0] node21714;
	wire [4-1:0] node21715;
	wire [4-1:0] node21718;
	wire [4-1:0] node21721;
	wire [4-1:0] node21722;
	wire [4-1:0] node21725;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21731;
	wire [4-1:0] node21732;
	wire [4-1:0] node21733;
	wire [4-1:0] node21734;
	wire [4-1:0] node21735;
	wire [4-1:0] node21736;
	wire [4-1:0] node21738;
	wire [4-1:0] node21740;
	wire [4-1:0] node21743;
	wire [4-1:0] node21745;
	wire [4-1:0] node21748;
	wire [4-1:0] node21749;
	wire [4-1:0] node21750;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21756;
	wire [4-1:0] node21759;
	wire [4-1:0] node21763;
	wire [4-1:0] node21764;
	wire [4-1:0] node21765;
	wire [4-1:0] node21766;
	wire [4-1:0] node21770;
	wire [4-1:0] node21772;
	wire [4-1:0] node21775;
	wire [4-1:0] node21776;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21782;
	wire [4-1:0] node21784;
	wire [4-1:0] node21787;
	wire [4-1:0] node21788;
	wire [4-1:0] node21789;
	wire [4-1:0] node21793;
	wire [4-1:0] node21795;
	wire [4-1:0] node21798;
	wire [4-1:0] node21799;
	wire [4-1:0] node21800;
	wire [4-1:0] node21801;
	wire [4-1:0] node21802;
	wire [4-1:0] node21804;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21810;
	wire [4-1:0] node21814;
	wire [4-1:0] node21816;
	wire [4-1:0] node21819;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21827;
	wire [4-1:0] node21830;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21833;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21841;
	wire [4-1:0] node21842;
	wire [4-1:0] node21844;
	wire [4-1:0] node21848;
	wire [4-1:0] node21849;
	wire [4-1:0] node21850;
	wire [4-1:0] node21851;
	wire [4-1:0] node21854;
	wire [4-1:0] node21857;
	wire [4-1:0] node21858;
	wire [4-1:0] node21862;
	wire [4-1:0] node21863;
	wire [4-1:0] node21865;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21875;
	wire [4-1:0] node21876;
	wire [4-1:0] node21877;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21883;
	wire [4-1:0] node21885;
	wire [4-1:0] node21888;
	wire [4-1:0] node21889;
	wire [4-1:0] node21890;
	wire [4-1:0] node21894;
	wire [4-1:0] node21897;
	wire [4-1:0] node21898;
	wire [4-1:0] node21900;
	wire [4-1:0] node21903;
	wire [4-1:0] node21904;
	wire [4-1:0] node21905;
	wire [4-1:0] node21910;
	wire [4-1:0] node21911;
	wire [4-1:0] node21912;
	wire [4-1:0] node21915;
	wire [4-1:0] node21916;
	wire [4-1:0] node21917;
	wire [4-1:0] node21921;
	wire [4-1:0] node21923;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21928;
	wire [4-1:0] node21931;
	wire [4-1:0] node21932;
	wire [4-1:0] node21936;
	wire [4-1:0] node21939;
	wire [4-1:0] node21940;
	wire [4-1:0] node21941;
	wire [4-1:0] node21942;
	wire [4-1:0] node21943;
	wire [4-1:0] node21944;
	wire [4-1:0] node21948;
	wire [4-1:0] node21949;
	wire [4-1:0] node21953;
	wire [4-1:0] node21955;
	wire [4-1:0] node21956;
	wire [4-1:0] node21959;
	wire [4-1:0] node21962;
	wire [4-1:0] node21963;
	wire [4-1:0] node21965;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21971;
	wire [4-1:0] node21974;
	wire [4-1:0] node21977;
	wire [4-1:0] node21978;
	wire [4-1:0] node21979;
	wire [4-1:0] node21980;
	wire [4-1:0] node21983;
	wire [4-1:0] node21985;
	wire [4-1:0] node21988;
	wire [4-1:0] node21989;
	wire [4-1:0] node21990;
	wire [4-1:0] node21994;
	wire [4-1:0] node21997;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22000;
	wire [4-1:0] node22004;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22009;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22017;
	wire [4-1:0] node22020;
	wire [4-1:0] node22021;
	wire [4-1:0] node22022;
	wire [4-1:0] node22023;
	wire [4-1:0] node22024;
	wire [4-1:0] node22025;
	wire [4-1:0] node22026;
	wire [4-1:0] node22030;
	wire [4-1:0] node22031;
	wire [4-1:0] node22032;
	wire [4-1:0] node22037;
	wire [4-1:0] node22038;
	wire [4-1:0] node22039;
	wire [4-1:0] node22043;
	wire [4-1:0] node22044;
	wire [4-1:0] node22047;
	wire [4-1:0] node22048;
	wire [4-1:0] node22052;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22056;
	wire [4-1:0] node22059;
	wire [4-1:0] node22060;
	wire [4-1:0] node22061;
	wire [4-1:0] node22064;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22071;
	wire [4-1:0] node22074;
	wire [4-1:0] node22075;
	wire [4-1:0] node22077;
	wire [4-1:0] node22080;
	wire [4-1:0] node22083;
	wire [4-1:0] node22084;
	wire [4-1:0] node22085;
	wire [4-1:0] node22086;
	wire [4-1:0] node22089;
	wire [4-1:0] node22090;
	wire [4-1:0] node22093;
	wire [4-1:0] node22094;
	wire [4-1:0] node22098;
	wire [4-1:0] node22099;
	wire [4-1:0] node22101;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22108;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22116;
	wire [4-1:0] node22117;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22125;
	wire [4-1:0] node22126;
	wire [4-1:0] node22127;
	wire [4-1:0] node22129;
	wire [4-1:0] node22132;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22138;
	wire [4-1:0] node22142;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22145;
	wire [4-1:0] node22146;
	wire [4-1:0] node22147;
	wire [4-1:0] node22148;
	wire [4-1:0] node22151;
	wire [4-1:0] node22155;
	wire [4-1:0] node22156;
	wire [4-1:0] node22160;
	wire [4-1:0] node22161;
	wire [4-1:0] node22162;
	wire [4-1:0] node22166;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22173;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22178;
	wire [4-1:0] node22182;
	wire [4-1:0] node22183;
	wire [4-1:0] node22184;
	wire [4-1:0] node22187;
	wire [4-1:0] node22191;
	wire [4-1:0] node22192;
	wire [4-1:0] node22193;
	wire [4-1:0] node22194;
	wire [4-1:0] node22199;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22206;
	wire [4-1:0] node22207;
	wire [4-1:0] node22208;
	wire [4-1:0] node22209;
	wire [4-1:0] node22210;
	wire [4-1:0] node22213;
	wire [4-1:0] node22215;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22220;
	wire [4-1:0] node22224;
	wire [4-1:0] node22227;
	wire [4-1:0] node22228;
	wire [4-1:0] node22229;
	wire [4-1:0] node22232;
	wire [4-1:0] node22235;
	wire [4-1:0] node22236;
	wire [4-1:0] node22237;
	wire [4-1:0] node22241;
	wire [4-1:0] node22244;
	wire [4-1:0] node22245;
	wire [4-1:0] node22246;
	wire [4-1:0] node22247;
	wire [4-1:0] node22249;
	wire [4-1:0] node22252;
	wire [4-1:0] node22256;
	wire [4-1:0] node22258;
	wire [4-1:0] node22260;
	wire [4-1:0] node22263;
	wire [4-1:0] node22264;
	wire [4-1:0] node22265;
	wire [4-1:0] node22266;
	wire [4-1:0] node22267;
	wire [4-1:0] node22268;
	wire [4-1:0] node22269;
	wire [4-1:0] node22270;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22276;
	wire [4-1:0] node22279;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22287;
	wire [4-1:0] node22288;
	wire [4-1:0] node22289;
	wire [4-1:0] node22292;
	wire [4-1:0] node22295;
	wire [4-1:0] node22298;
	wire [4-1:0] node22299;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22307;
	wire [4-1:0] node22308;
	wire [4-1:0] node22311;
	wire [4-1:0] node22314;
	wire [4-1:0] node22315;
	wire [4-1:0] node22317;
	wire [4-1:0] node22319;
	wire [4-1:0] node22322;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22327;
	wire [4-1:0] node22330;
	wire [4-1:0] node22331;
	wire [4-1:0] node22335;
	wire [4-1:0] node22336;
	wire [4-1:0] node22337;
	wire [4-1:0] node22338;
	wire [4-1:0] node22339;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22347;
	wire [4-1:0] node22348;
	wire [4-1:0] node22351;
	wire [4-1:0] node22352;
	wire [4-1:0] node22355;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22362;
	wire [4-1:0] node22363;
	wire [4-1:0] node22366;
	wire [4-1:0] node22367;
	wire [4-1:0] node22371;
	wire [4-1:0] node22372;
	wire [4-1:0] node22373;
	wire [4-1:0] node22374;
	wire [4-1:0] node22377;
	wire [4-1:0] node22380;
	wire [4-1:0] node22381;
	wire [4-1:0] node22384;
	wire [4-1:0] node22387;
	wire [4-1:0] node22388;
	wire [4-1:0] node22389;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22397;
	wire [4-1:0] node22398;
	wire [4-1:0] node22400;
	wire [4-1:0] node22403;
	wire [4-1:0] node22404;
	wire [4-1:0] node22408;
	wire [4-1:0] node22409;
	wire [4-1:0] node22410;
	wire [4-1:0] node22411;
	wire [4-1:0] node22412;
	wire [4-1:0] node22413;
	wire [4-1:0] node22414;
	wire [4-1:0] node22418;
	wire [4-1:0] node22421;
	wire [4-1:0] node22424;
	wire [4-1:0] node22425;
	wire [4-1:0] node22427;
	wire [4-1:0] node22428;
	wire [4-1:0] node22432;
	wire [4-1:0] node22433;
	wire [4-1:0] node22434;
	wire [4-1:0] node22439;
	wire [4-1:0] node22440;
	wire [4-1:0] node22441;
	wire [4-1:0] node22442;
	wire [4-1:0] node22446;
	wire [4-1:0] node22447;
	wire [4-1:0] node22449;
	wire [4-1:0] node22452;
	wire [4-1:0] node22455;
	wire [4-1:0] node22456;
	wire [4-1:0] node22457;
	wire [4-1:0] node22458;
	wire [4-1:0] node22463;
	wire [4-1:0] node22465;
	wire [4-1:0] node22467;
	wire [4-1:0] node22470;
	wire [4-1:0] node22471;
	wire [4-1:0] node22472;
	wire [4-1:0] node22473;
	wire [4-1:0] node22474;
	wire [4-1:0] node22478;
	wire [4-1:0] node22479;
	wire [4-1:0] node22482;
	wire [4-1:0] node22485;
	wire [4-1:0] node22486;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22493;
	wire [4-1:0] node22495;
	wire [4-1:0] node22498;
	wire [4-1:0] node22499;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22503;
	wire [4-1:0] node22506;
	wire [4-1:0] node22508;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22515;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22522;
	wire [4-1:0] node22523;
	wire [4-1:0] node22525;
	wire [4-1:0] node22529;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22532;
	wire [4-1:0] node22533;
	wire [4-1:0] node22534;
	wire [4-1:0] node22535;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22547;
	wire [4-1:0] node22549;
	wire [4-1:0] node22552;
	wire [4-1:0] node22553;
	wire [4-1:0] node22554;
	wire [4-1:0] node22557;
	wire [4-1:0] node22559;
	wire [4-1:0] node22562;
	wire [4-1:0] node22565;
	wire [4-1:0] node22566;
	wire [4-1:0] node22567;
	wire [4-1:0] node22568;
	wire [4-1:0] node22570;
	wire [4-1:0] node22573;
	wire [4-1:0] node22575;
	wire [4-1:0] node22578;
	wire [4-1:0] node22580;
	wire [4-1:0] node22583;
	wire [4-1:0] node22584;
	wire [4-1:0] node22586;
	wire [4-1:0] node22589;
	wire [4-1:0] node22590;
	wire [4-1:0] node22593;
	wire [4-1:0] node22595;
	wire [4-1:0] node22598;
	wire [4-1:0] node22599;
	wire [4-1:0] node22600;
	wire [4-1:0] node22603;
	wire [4-1:0] node22604;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22610;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22618;
	wire [4-1:0] node22621;
	wire [4-1:0] node22622;
	wire [4-1:0] node22625;
	wire [4-1:0] node22628;
	wire [4-1:0] node22629;
	wire [4-1:0] node22630;
	wire [4-1:0] node22632;
	wire [4-1:0] node22634;
	wire [4-1:0] node22637;
	wire [4-1:0] node22639;
	wire [4-1:0] node22640;
	wire [4-1:0] node22644;
	wire [4-1:0] node22645;
	wire [4-1:0] node22646;
	wire [4-1:0] node22648;
	wire [4-1:0] node22651;
	wire [4-1:0] node22652;
	wire [4-1:0] node22655;
	wire [4-1:0] node22658;
	wire [4-1:0] node22659;
	wire [4-1:0] node22662;
	wire [4-1:0] node22665;
	wire [4-1:0] node22666;
	wire [4-1:0] node22667;
	wire [4-1:0] node22668;
	wire [4-1:0] node22669;
	wire [4-1:0] node22671;
	wire [4-1:0] node22673;
	wire [4-1:0] node22676;
	wire [4-1:0] node22677;
	wire [4-1:0] node22680;
	wire [4-1:0] node22682;
	wire [4-1:0] node22685;
	wire [4-1:0] node22686;
	wire [4-1:0] node22687;
	wire [4-1:0] node22688;
	wire [4-1:0] node22691;
	wire [4-1:0] node22694;
	wire [4-1:0] node22697;
	wire [4-1:0] node22698;
	wire [4-1:0] node22700;
	wire [4-1:0] node22703;
	wire [4-1:0] node22705;
	wire [4-1:0] node22708;
	wire [4-1:0] node22709;
	wire [4-1:0] node22710;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22716;
	wire [4-1:0] node22717;
	wire [4-1:0] node22720;
	wire [4-1:0] node22723;
	wire [4-1:0] node22725;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22731;
	wire [4-1:0] node22734;
	wire [4-1:0] node22738;
	wire [4-1:0] node22739;
	wire [4-1:0] node22740;
	wire [4-1:0] node22743;
	wire [4-1:0] node22746;
	wire [4-1:0] node22749;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22752;
	wire [4-1:0] node22753;
	wire [4-1:0] node22754;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22763;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22769;
	wire [4-1:0] node22773;
	wire [4-1:0] node22774;
	wire [4-1:0] node22778;
	wire [4-1:0] node22779;
	wire [4-1:0] node22781;
	wire [4-1:0] node22785;
	wire [4-1:0] node22786;
	wire [4-1:0] node22787;
	wire [4-1:0] node22788;
	wire [4-1:0] node22791;
	wire [4-1:0] node22792;
	wire [4-1:0] node22795;
	wire [4-1:0] node22798;
	wire [4-1:0] node22799;
	wire [4-1:0] node22800;
	wire [4-1:0] node22804;
	wire [4-1:0] node22805;
	wire [4-1:0] node22808;
	wire [4-1:0] node22811;
	wire [4-1:0] node22812;
	wire [4-1:0] node22813;
	wire [4-1:0] node22814;
	wire [4-1:0] node22818;
	wire [4-1:0] node22819;
	wire [4-1:0] node22822;
	wire [4-1:0] node22825;
	wire [4-1:0] node22826;
	wire [4-1:0] node22827;
	wire [4-1:0] node22830;
	wire [4-1:0] node22834;
	wire [4-1:0] node22835;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22838;
	wire [4-1:0] node22839;
	wire [4-1:0] node22840;
	wire [4-1:0] node22841;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22848;
	wire [4-1:0] node22851;
	wire [4-1:0] node22854;
	wire [4-1:0] node22855;
	wire [4-1:0] node22858;
	wire [4-1:0] node22861;
	wire [4-1:0] node22862;
	wire [4-1:0] node22863;
	wire [4-1:0] node22867;
	wire [4-1:0] node22868;
	wire [4-1:0] node22871;
	wire [4-1:0] node22874;
	wire [4-1:0] node22875;
	wire [4-1:0] node22876;
	wire [4-1:0] node22877;
	wire [4-1:0] node22879;
	wire [4-1:0] node22882;
	wire [4-1:0] node22883;
	wire [4-1:0] node22886;
	wire [4-1:0] node22889;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22895;
	wire [4-1:0] node22898;
	wire [4-1:0] node22900;
	wire [4-1:0] node22901;
	wire [4-1:0] node22902;
	wire [4-1:0] node22906;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22911;
	wire [4-1:0] node22912;
	wire [4-1:0] node22913;
	wire [4-1:0] node22916;
	wire [4-1:0] node22918;
	wire [4-1:0] node22921;
	wire [4-1:0] node22922;
	wire [4-1:0] node22925;
	wire [4-1:0] node22928;
	wire [4-1:0] node22929;
	wire [4-1:0] node22930;
	wire [4-1:0] node22933;
	wire [4-1:0] node22936;
	wire [4-1:0] node22937;
	wire [4-1:0] node22938;
	wire [4-1:0] node22942;
	wire [4-1:0] node22944;
	wire [4-1:0] node22947;
	wire [4-1:0] node22948;
	wire [4-1:0] node22949;
	wire [4-1:0] node22950;
	wire [4-1:0] node22953;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22961;
	wire [4-1:0] node22962;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22968;
	wire [4-1:0] node22969;
	wire [4-1:0] node22974;
	wire [4-1:0] node22975;
	wire [4-1:0] node22976;
	wire [4-1:0] node22977;
	wire [4-1:0] node22978;
	wire [4-1:0] node22979;
	wire [4-1:0] node22982;
	wire [4-1:0] node22985;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22991;
	wire [4-1:0] node22992;
	wire [4-1:0] node22993;
	wire [4-1:0] node22997;
	wire [4-1:0] node22998;
	wire [4-1:0] node23002;
	wire [4-1:0] node23003;
	wire [4-1:0] node23004;
	wire [4-1:0] node23007;
	wire [4-1:0] node23011;
	wire [4-1:0] node23012;
	wire [4-1:0] node23013;
	wire [4-1:0] node23014;
	wire [4-1:0] node23017;
	wire [4-1:0] node23020;
	wire [4-1:0] node23021;
	wire [4-1:0] node23022;
	wire [4-1:0] node23025;
	wire [4-1:0] node23029;
	wire [4-1:0] node23030;
	wire [4-1:0] node23031;
	wire [4-1:0] node23033;
	wire [4-1:0] node23036;
	wire [4-1:0] node23039;
	wire [4-1:0] node23041;
	wire [4-1:0] node23043;
	wire [4-1:0] node23046;
	wire [4-1:0] node23047;
	wire [4-1:0] node23048;
	wire [4-1:0] node23049;
	wire [4-1:0] node23052;
	wire [4-1:0] node23054;
	wire [4-1:0] node23057;
	wire [4-1:0] node23058;
	wire [4-1:0] node23060;
	wire [4-1:0] node23063;
	wire [4-1:0] node23066;
	wire [4-1:0] node23067;
	wire [4-1:0] node23068;
	wire [4-1:0] node23070;
	wire [4-1:0] node23073;
	wire [4-1:0] node23075;
	wire [4-1:0] node23078;
	wire [4-1:0] node23079;
	wire [4-1:0] node23081;
	wire [4-1:0] node23084;
	wire [4-1:0] node23087;
	wire [4-1:0] node23088;
	wire [4-1:0] node23089;
	wire [4-1:0] node23090;
	wire [4-1:0] node23091;
	wire [4-1:0] node23092;
	wire [4-1:0] node23094;
	wire [4-1:0] node23095;
	wire [4-1:0] node23099;
	wire [4-1:0] node23100;
	wire [4-1:0] node23103;
	wire [4-1:0] node23106;
	wire [4-1:0] node23107;
	wire [4-1:0] node23108;
	wire [4-1:0] node23111;
	wire [4-1:0] node23114;
	wire [4-1:0] node23116;
	wire [4-1:0] node23119;
	wire [4-1:0] node23120;
	wire [4-1:0] node23121;
	wire [4-1:0] node23122;
	wire [4-1:0] node23125;
	wire [4-1:0] node23126;
	wire [4-1:0] node23130;
	wire [4-1:0] node23132;
	wire [4-1:0] node23135;
	wire [4-1:0] node23136;
	wire [4-1:0] node23137;
	wire [4-1:0] node23138;
	wire [4-1:0] node23143;
	wire [4-1:0] node23144;
	wire [4-1:0] node23148;
	wire [4-1:0] node23149;
	wire [4-1:0] node23150;
	wire [4-1:0] node23151;
	wire [4-1:0] node23152;
	wire [4-1:0] node23154;
	wire [4-1:0] node23157;
	wire [4-1:0] node23159;
	wire [4-1:0] node23163;
	wire [4-1:0] node23164;
	wire [4-1:0] node23165;
	wire [4-1:0] node23168;
	wire [4-1:0] node23171;
	wire [4-1:0] node23172;
	wire [4-1:0] node23173;
	wire [4-1:0] node23176;
	wire [4-1:0] node23179;
	wire [4-1:0] node23181;
	wire [4-1:0] node23184;
	wire [4-1:0] node23185;
	wire [4-1:0] node23186;
	wire [4-1:0] node23187;
	wire [4-1:0] node23188;
	wire [4-1:0] node23192;
	wire [4-1:0] node23193;
	wire [4-1:0] node23197;
	wire [4-1:0] node23198;
	wire [4-1:0] node23202;
	wire [4-1:0] node23203;
	wire [4-1:0] node23204;
	wire [4-1:0] node23205;
	wire [4-1:0] node23209;
	wire [4-1:0] node23210;
	wire [4-1:0] node23214;
	wire [4-1:0] node23215;
	wire [4-1:0] node23218;
	wire [4-1:0] node23221;
	wire [4-1:0] node23222;
	wire [4-1:0] node23223;
	wire [4-1:0] node23224;
	wire [4-1:0] node23225;
	wire [4-1:0] node23229;
	wire [4-1:0] node23230;
	wire [4-1:0] node23234;
	wire [4-1:0] node23235;
	wire [4-1:0] node23236;
	wire [4-1:0] node23240;
	wire [4-1:0] node23241;
	wire [4-1:0] node23245;
	wire [4-1:0] node23246;
	wire [4-1:0] node23247;
	wire [4-1:0] node23248;
	wire [4-1:0] node23251;
	wire [4-1:0] node23254;
	wire [4-1:0] node23256;
	wire [4-1:0] node23258;
	wire [4-1:0] node23261;
	wire [4-1:0] node23262;
	wire [4-1:0] node23263;
	wire [4-1:0] node23266;
	wire [4-1:0] node23269;
	wire [4-1:0] node23270;
	wire [4-1:0] node23271;
	wire [4-1:0] node23272;
	wire [4-1:0] node23275;
	wire [4-1:0] node23278;
	wire [4-1:0] node23280;
	wire [4-1:0] node23283;
	wire [4-1:0] node23285;
	wire [4-1:0] node23288;
	wire [4-1:0] node23289;
	wire [4-1:0] node23290;
	wire [4-1:0] node23291;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23294;
	wire [4-1:0] node23295;
	wire [4-1:0] node23296;
	wire [4-1:0] node23300;
	wire [4-1:0] node23301;
	wire [4-1:0] node23305;
	wire [4-1:0] node23306;
	wire [4-1:0] node23307;
	wire [4-1:0] node23310;
	wire [4-1:0] node23313;
	wire [4-1:0] node23314;
	wire [4-1:0] node23318;
	wire [4-1:0] node23319;
	wire [4-1:0] node23320;
	wire [4-1:0] node23321;
	wire [4-1:0] node23325;
	wire [4-1:0] node23328;
	wire [4-1:0] node23330;
	wire [4-1:0] node23333;
	wire [4-1:0] node23334;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23338;
	wire [4-1:0] node23342;
	wire [4-1:0] node23344;
	wire [4-1:0] node23345;
	wire [4-1:0] node23348;
	wire [4-1:0] node23351;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23354;
	wire [4-1:0] node23357;
	wire [4-1:0] node23360;
	wire [4-1:0] node23361;
	wire [4-1:0] node23364;
	wire [4-1:0] node23367;
	wire [4-1:0] node23368;
	wire [4-1:0] node23369;
	wire [4-1:0] node23372;
	wire [4-1:0] node23375;
	wire [4-1:0] node23378;
	wire [4-1:0] node23379;
	wire [4-1:0] node23380;
	wire [4-1:0] node23381;
	wire [4-1:0] node23383;
	wire [4-1:0] node23386;
	wire [4-1:0] node23388;
	wire [4-1:0] node23390;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23395;
	wire [4-1:0] node23398;
	wire [4-1:0] node23402;
	wire [4-1:0] node23403;
	wire [4-1:0] node23404;
	wire [4-1:0] node23407;
	wire [4-1:0] node23408;
	wire [4-1:0] node23409;
	wire [4-1:0] node23413;
	wire [4-1:0] node23416;
	wire [4-1:0] node23417;
	wire [4-1:0] node23418;
	wire [4-1:0] node23419;
	wire [4-1:0] node23424;
	wire [4-1:0] node23425;
	wire [4-1:0] node23426;
	wire [4-1:0] node23430;
	wire [4-1:0] node23431;
	wire [4-1:0] node23435;
	wire [4-1:0] node23436;
	wire [4-1:0] node23437;
	wire [4-1:0] node23438;
	wire [4-1:0] node23439;
	wire [4-1:0] node23440;
	wire [4-1:0] node23441;
	wire [4-1:0] node23445;
	wire [4-1:0] node23448;
	wire [4-1:0] node23449;
	wire [4-1:0] node23453;
	wire [4-1:0] node23454;
	wire [4-1:0] node23455;
	wire [4-1:0] node23456;
	wire [4-1:0] node23461;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23468;
	wire [4-1:0] node23469;
	wire [4-1:0] node23470;
	wire [4-1:0] node23471;
	wire [4-1:0] node23474;
	wire [4-1:0] node23478;
	wire [4-1:0] node23479;
	wire [4-1:0] node23480;
	wire [4-1:0] node23484;
	wire [4-1:0] node23485;
	wire [4-1:0] node23489;
	wire [4-1:0] node23490;
	wire [4-1:0] node23491;
	wire [4-1:0] node23492;
	wire [4-1:0] node23493;
	wire [4-1:0] node23494;
	wire [4-1:0] node23497;
	wire [4-1:0] node23501;
	wire [4-1:0] node23503;
	wire [4-1:0] node23504;
	wire [4-1:0] node23508;
	wire [4-1:0] node23509;
	wire [4-1:0] node23510;
	wire [4-1:0] node23513;
	wire [4-1:0] node23514;
	wire [4-1:0] node23519;
	wire [4-1:0] node23520;
	wire [4-1:0] node23521;
	wire [4-1:0] node23523;
	wire [4-1:0] node23524;
	wire [4-1:0] node23528;
	wire [4-1:0] node23530;
	wire [4-1:0] node23531;
	wire [4-1:0] node23535;
	wire [4-1:0] node23536;
	wire [4-1:0] node23538;
	wire [4-1:0] node23541;
	wire [4-1:0] node23543;
	wire [4-1:0] node23544;
	wire [4-1:0] node23548;
	wire [4-1:0] node23549;
	wire [4-1:0] node23550;
	wire [4-1:0] node23551;
	wire [4-1:0] node23552;
	wire [4-1:0] node23553;
	wire [4-1:0] node23554;
	wire [4-1:0] node23558;
	wire [4-1:0] node23559;
	wire [4-1:0] node23561;
	wire [4-1:0] node23565;
	wire [4-1:0] node23566;
	wire [4-1:0] node23567;
	wire [4-1:0] node23568;
	wire [4-1:0] node23573;
	wire [4-1:0] node23575;
	wire [4-1:0] node23577;
	wire [4-1:0] node23580;
	wire [4-1:0] node23581;
	wire [4-1:0] node23582;
	wire [4-1:0] node23583;
	wire [4-1:0] node23586;
	wire [4-1:0] node23589;
	wire [4-1:0] node23591;
	wire [4-1:0] node23593;
	wire [4-1:0] node23596;
	wire [4-1:0] node23597;
	wire [4-1:0] node23598;
	wire [4-1:0] node23601;
	wire [4-1:0] node23604;
	wire [4-1:0] node23607;
	wire [4-1:0] node23608;
	wire [4-1:0] node23609;
	wire [4-1:0] node23610;
	wire [4-1:0] node23611;
	wire [4-1:0] node23612;
	wire [4-1:0] node23616;
	wire [4-1:0] node23617;
	wire [4-1:0] node23621;
	wire [4-1:0] node23622;
	wire [4-1:0] node23624;
	wire [4-1:0] node23627;
	wire [4-1:0] node23628;
	wire [4-1:0] node23632;
	wire [4-1:0] node23633;
	wire [4-1:0] node23634;
	wire [4-1:0] node23636;
	wire [4-1:0] node23640;
	wire [4-1:0] node23642;
	wire [4-1:0] node23643;
	wire [4-1:0] node23647;
	wire [4-1:0] node23648;
	wire [4-1:0] node23649;
	wire [4-1:0] node23650;
	wire [4-1:0] node23651;
	wire [4-1:0] node23654;
	wire [4-1:0] node23657;
	wire [4-1:0] node23658;
	wire [4-1:0] node23661;
	wire [4-1:0] node23664;
	wire [4-1:0] node23665;
	wire [4-1:0] node23669;
	wire [4-1:0] node23670;
	wire [4-1:0] node23671;
	wire [4-1:0] node23672;
	wire [4-1:0] node23676;
	wire [4-1:0] node23677;
	wire [4-1:0] node23682;
	wire [4-1:0] node23683;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23686;
	wire [4-1:0] node23690;
	wire [4-1:0] node23691;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23697;
	wire [4-1:0] node23701;
	wire [4-1:0] node23702;
	wire [4-1:0] node23706;
	wire [4-1:0] node23707;
	wire [4-1:0] node23708;
	wire [4-1:0] node23709;
	wire [4-1:0] node23711;
	wire [4-1:0] node23714;
	wire [4-1:0] node23715;
	wire [4-1:0] node23716;
	wire [4-1:0] node23719;
	wire [4-1:0] node23722;
	wire [4-1:0] node23723;
	wire [4-1:0] node23726;
	wire [4-1:0] node23729;
	wire [4-1:0] node23730;
	wire [4-1:0] node23731;
	wire [4-1:0] node23734;
	wire [4-1:0] node23737;
	wire [4-1:0] node23738;
	wire [4-1:0] node23741;
	wire [4-1:0] node23744;
	wire [4-1:0] node23745;
	wire [4-1:0] node23746;
	wire [4-1:0] node23747;
	wire [4-1:0] node23751;
	wire [4-1:0] node23752;
	wire [4-1:0] node23756;
	wire [4-1:0] node23758;
	wire [4-1:0] node23760;
	wire [4-1:0] node23763;
	wire [4-1:0] node23764;
	wire [4-1:0] node23765;
	wire [4-1:0] node23766;
	wire [4-1:0] node23767;
	wire [4-1:0] node23768;
	wire [4-1:0] node23769;
	wire [4-1:0] node23770;
	wire [4-1:0] node23771;
	wire [4-1:0] node23774;
	wire [4-1:0] node23775;
	wire [4-1:0] node23776;
	wire [4-1:0] node23779;
	wire [4-1:0] node23782;
	wire [4-1:0] node23784;
	wire [4-1:0] node23787;
	wire [4-1:0] node23788;
	wire [4-1:0] node23790;
	wire [4-1:0] node23793;
	wire [4-1:0] node23794;
	wire [4-1:0] node23795;
	wire [4-1:0] node23798;
	wire [4-1:0] node23801;
	wire [4-1:0] node23802;
	wire [4-1:0] node23806;
	wire [4-1:0] node23807;
	wire [4-1:0] node23808;
	wire [4-1:0] node23809;
	wire [4-1:0] node23811;
	wire [4-1:0] node23814;
	wire [4-1:0] node23816;
	wire [4-1:0] node23819;
	wire [4-1:0] node23820;
	wire [4-1:0] node23822;
	wire [4-1:0] node23825;
	wire [4-1:0] node23826;
	wire [4-1:0] node23829;
	wire [4-1:0] node23832;
	wire [4-1:0] node23833;
	wire [4-1:0] node23834;
	wire [4-1:0] node23836;
	wire [4-1:0] node23839;
	wire [4-1:0] node23841;
	wire [4-1:0] node23844;
	wire [4-1:0] node23845;
	wire [4-1:0] node23847;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23854;
	wire [4-1:0] node23857;
	wire [4-1:0] node23858;
	wire [4-1:0] node23859;
	wire [4-1:0] node23860;
	wire [4-1:0] node23862;
	wire [4-1:0] node23864;
	wire [4-1:0] node23867;
	wire [4-1:0] node23869;
	wire [4-1:0] node23872;
	wire [4-1:0] node23873;
	wire [4-1:0] node23875;
	wire [4-1:0] node23878;
	wire [4-1:0] node23879;
	wire [4-1:0] node23880;
	wire [4-1:0] node23883;
	wire [4-1:0] node23886;
	wire [4-1:0] node23887;
	wire [4-1:0] node23890;
	wire [4-1:0] node23893;
	wire [4-1:0] node23894;
	wire [4-1:0] node23895;
	wire [4-1:0] node23896;
	wire [4-1:0] node23899;
	wire [4-1:0] node23900;
	wire [4-1:0] node23903;
	wire [4-1:0] node23906;
	wire [4-1:0] node23907;
	wire [4-1:0] node23908;
	wire [4-1:0] node23911;
	wire [4-1:0] node23914;
	wire [4-1:0] node23915;
	wire [4-1:0] node23916;
	wire [4-1:0] node23919;
	wire [4-1:0] node23923;
	wire [4-1:0] node23924;
	wire [4-1:0] node23925;
	wire [4-1:0] node23927;
	wire [4-1:0] node23930;
	wire [4-1:0] node23932;
	wire [4-1:0] node23935;
	wire [4-1:0] node23936;
	wire [4-1:0] node23938;
	wire [4-1:0] node23941;
	wire [4-1:0] node23942;
	wire [4-1:0] node23945;
	wire [4-1:0] node23948;
	wire [4-1:0] node23949;
	wire [4-1:0] node23950;
	wire [4-1:0] node23951;
	wire [4-1:0] node23952;
	wire [4-1:0] node23954;
	wire [4-1:0] node23956;
	wire [4-1:0] node23959;
	wire [4-1:0] node23961;
	wire [4-1:0] node23964;
	wire [4-1:0] node23965;
	wire [4-1:0] node23967;
	wire [4-1:0] node23968;
	wire [4-1:0] node23971;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23976;
	wire [4-1:0] node23979;
	wire [4-1:0] node23982;
	wire [4-1:0] node23983;
	wire [4-1:0] node23986;
	wire [4-1:0] node23989;
	wire [4-1:0] node23990;
	wire [4-1:0] node23991;
	wire [4-1:0] node23992;
	wire [4-1:0] node23995;
	wire [4-1:0] node23996;
	wire [4-1:0] node23999;
	wire [4-1:0] node24002;
	wire [4-1:0] node24003;
	wire [4-1:0] node24004;
	wire [4-1:0] node24007;
	wire [4-1:0] node24010;
	wire [4-1:0] node24011;
	wire [4-1:0] node24014;
	wire [4-1:0] node24017;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24021;
	wire [4-1:0] node24024;
	wire [4-1:0] node24025;
	wire [4-1:0] node24028;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24033;
	wire [4-1:0] node24036;
	wire [4-1:0] node24039;
	wire [4-1:0] node24040;
	wire [4-1:0] node24043;
	wire [4-1:0] node24046;
	wire [4-1:0] node24047;
	wire [4-1:0] node24048;
	wire [4-1:0] node24049;
	wire [4-1:0] node24051;
	wire [4-1:0] node24053;
	wire [4-1:0] node24056;
	wire [4-1:0] node24058;
	wire [4-1:0] node24061;
	wire [4-1:0] node24062;
	wire [4-1:0] node24063;
	wire [4-1:0] node24066;
	wire [4-1:0] node24069;
	wire [4-1:0] node24070;
	wire [4-1:0] node24071;
	wire [4-1:0] node24074;
	wire [4-1:0] node24077;
	wire [4-1:0] node24078;
	wire [4-1:0] node24082;
	wire [4-1:0] node24083;
	wire [4-1:0] node24084;
	wire [4-1:0] node24085;
	wire [4-1:0] node24088;
	wire [4-1:0] node24089;
	wire [4-1:0] node24092;
	wire [4-1:0] node24095;
	wire [4-1:0] node24096;
	wire [4-1:0] node24097;
	wire [4-1:0] node24100;
	wire [4-1:0] node24103;
	wire [4-1:0] node24104;
	wire [4-1:0] node24105;
	wire [4-1:0] node24108;
	wire [4-1:0] node24111;
	wire [4-1:0] node24112;
	wire [4-1:0] node24113;
	wire [4-1:0] node24116;
	wire [4-1:0] node24120;
	wire [4-1:0] node24121;
	wire [4-1:0] node24122;
	wire [4-1:0] node24124;
	wire [4-1:0] node24127;
	wire [4-1:0] node24128;
	wire [4-1:0] node24131;
	wire [4-1:0] node24134;
	wire [4-1:0] node24135;
	wire [4-1:0] node24136;
	wire [4-1:0] node24140;
	wire [4-1:0] node24141;
	wire [4-1:0] node24144;
	wire [4-1:0] node24147;
	wire [4-1:0] node24148;
	wire [4-1:0] node24149;
	wire [4-1:0] node24150;
	wire [4-1:0] node24151;
	wire [4-1:0] node24152;
	wire [4-1:0] node24153;
	wire [4-1:0] node24156;
	wire [4-1:0] node24158;
	wire [4-1:0] node24161;
	wire [4-1:0] node24162;
	wire [4-1:0] node24165;
	wire [4-1:0] node24167;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24172;
	wire [4-1:0] node24173;
	wire [4-1:0] node24176;
	wire [4-1:0] node24179;
	wire [4-1:0] node24180;
	wire [4-1:0] node24182;
	wire [4-1:0] node24183;
	wire [4-1:0] node24187;
	wire [4-1:0] node24189;
	wire [4-1:0] node24192;
	wire [4-1:0] node24193;
	wire [4-1:0] node24196;
	wire [4-1:0] node24198;
	wire [4-1:0] node24201;
	wire [4-1:0] node24202;
	wire [4-1:0] node24203;
	wire [4-1:0] node24204;
	wire [4-1:0] node24205;
	wire [4-1:0] node24206;
	wire [4-1:0] node24210;
	wire [4-1:0] node24213;
	wire [4-1:0] node24214;
	wire [4-1:0] node24215;
	wire [4-1:0] node24219;
	wire [4-1:0] node24222;
	wire [4-1:0] node24223;
	wire [4-1:0] node24225;
	wire [4-1:0] node24226;
	wire [4-1:0] node24227;
	wire [4-1:0] node24231;
	wire [4-1:0] node24234;
	wire [4-1:0] node24235;
	wire [4-1:0] node24236;
	wire [4-1:0] node24240;
	wire [4-1:0] node24243;
	wire [4-1:0] node24244;
	wire [4-1:0] node24245;
	wire [4-1:0] node24246;
	wire [4-1:0] node24250;
	wire [4-1:0] node24253;
	wire [4-1:0] node24254;
	wire [4-1:0] node24255;
	wire [4-1:0] node24256;
	wire [4-1:0] node24259;
	wire [4-1:0] node24262;
	wire [4-1:0] node24264;
	wire [4-1:0] node24266;
	wire [4-1:0] node24269;
	wire [4-1:0] node24270;
	wire [4-1:0] node24273;
	wire [4-1:0] node24276;
	wire [4-1:0] node24277;
	wire [4-1:0] node24278;
	wire [4-1:0] node24279;
	wire [4-1:0] node24280;
	wire [4-1:0] node24282;
	wire [4-1:0] node24283;
	wire [4-1:0] node24286;
	wire [4-1:0] node24289;
	wire [4-1:0] node24290;
	wire [4-1:0] node24291;
	wire [4-1:0] node24295;
	wire [4-1:0] node24296;
	wire [4-1:0] node24298;
	wire [4-1:0] node24302;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24306;
	wire [4-1:0] node24309;
	wire [4-1:0] node24312;
	wire [4-1:0] node24314;
	wire [4-1:0] node24317;
	wire [4-1:0] node24318;
	wire [4-1:0] node24321;
	wire [4-1:0] node24324;
	wire [4-1:0] node24326;
	wire [4-1:0] node24327;
	wire [4-1:0] node24330;
	wire [4-1:0] node24333;
	wire [4-1:0] node24334;
	wire [4-1:0] node24337;
	wire [4-1:0] node24340;
	wire [4-1:0] node24341;
	wire [4-1:0] node24342;
	wire [4-1:0] node24343;
	wire [4-1:0] node24345;
	wire [4-1:0] node24346;
	wire [4-1:0] node24349;
	wire [4-1:0] node24352;
	wire [4-1:0] node24353;
	wire [4-1:0] node24355;
	wire [4-1:0] node24356;
	wire [4-1:0] node24359;
	wire [4-1:0] node24362;
	wire [4-1:0] node24363;
	wire [4-1:0] node24367;
	wire [4-1:0] node24368;
	wire [4-1:0] node24369;
	wire [4-1:0] node24370;
	wire [4-1:0] node24373;
	wire [4-1:0] node24376;
	wire [4-1:0] node24377;
	wire [4-1:0] node24381;
	wire [4-1:0] node24382;
	wire [4-1:0] node24383;
	wire [4-1:0] node24384;
	wire [4-1:0] node24387;
	wire [4-1:0] node24390;
	wire [4-1:0] node24391;
	wire [4-1:0] node24394;
	wire [4-1:0] node24397;
	wire [4-1:0] node24398;
	wire [4-1:0] node24401;
	wire [4-1:0] node24404;
	wire [4-1:0] node24405;
	wire [4-1:0] node24406;
	wire [4-1:0] node24407;
	wire [4-1:0] node24408;
	wire [4-1:0] node24409;
	wire [4-1:0] node24415;
	wire [4-1:0] node24416;
	wire [4-1:0] node24418;
	wire [4-1:0] node24421;
	wire [4-1:0] node24422;
	wire [4-1:0] node24423;
	wire [4-1:0] node24426;
	wire [4-1:0] node24429;
	wire [4-1:0] node24430;
	wire [4-1:0] node24434;
	wire [4-1:0] node24435;
	wire [4-1:0] node24438;
	wire [4-1:0] node24441;
	wire [4-1:0] node24442;
	wire [4-1:0] node24443;
	wire [4-1:0] node24444;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24447;
	wire [4-1:0] node24450;
	wire [4-1:0] node24453;
	wire [4-1:0] node24454;
	wire [4-1:0] node24457;
	wire [4-1:0] node24460;
	wire [4-1:0] node24461;
	wire [4-1:0] node24462;
	wire [4-1:0] node24464;
	wire [4-1:0] node24465;
	wire [4-1:0] node24468;
	wire [4-1:0] node24471;
	wire [4-1:0] node24473;
	wire [4-1:0] node24476;
	wire [4-1:0] node24477;
	wire [4-1:0] node24478;
	wire [4-1:0] node24479;
	wire [4-1:0] node24484;
	wire [4-1:0] node24486;
	wire [4-1:0] node24489;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24492;
	wire [4-1:0] node24493;
	wire [4-1:0] node24494;
	wire [4-1:0] node24498;
	wire [4-1:0] node24499;
	wire [4-1:0] node24502;
	wire [4-1:0] node24505;
	wire [4-1:0] node24506;
	wire [4-1:0] node24509;
	wire [4-1:0] node24512;
	wire [4-1:0] node24513;
	wire [4-1:0] node24514;
	wire [4-1:0] node24515;
	wire [4-1:0] node24518;
	wire [4-1:0] node24522;
	wire [4-1:0] node24523;
	wire [4-1:0] node24526;
	wire [4-1:0] node24529;
	wire [4-1:0] node24530;
	wire [4-1:0] node24531;
	wire [4-1:0] node24532;
	wire [4-1:0] node24535;
	wire [4-1:0] node24538;
	wire [4-1:0] node24539;
	wire [4-1:0] node24543;
	wire [4-1:0] node24544;
	wire [4-1:0] node24546;
	wire [4-1:0] node24547;
	wire [4-1:0] node24551;
	wire [4-1:0] node24554;
	wire [4-1:0] node24555;
	wire [4-1:0] node24556;
	wire [4-1:0] node24557;
	wire [4-1:0] node24558;
	wire [4-1:0] node24561;
	wire [4-1:0] node24564;
	wire [4-1:0] node24565;
	wire [4-1:0] node24566;
	wire [4-1:0] node24568;
	wire [4-1:0] node24572;
	wire [4-1:0] node24573;
	wire [4-1:0] node24574;
	wire [4-1:0] node24578;
	wire [4-1:0] node24579;
	wire [4-1:0] node24582;
	wire [4-1:0] node24585;
	wire [4-1:0] node24586;
	wire [4-1:0] node24587;
	wire [4-1:0] node24588;
	wire [4-1:0] node24591;
	wire [4-1:0] node24594;
	wire [4-1:0] node24595;
	wire [4-1:0] node24598;
	wire [4-1:0] node24601;
	wire [4-1:0] node24602;
	wire [4-1:0] node24605;
	wire [4-1:0] node24608;
	wire [4-1:0] node24609;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24614;
	wire [4-1:0] node24617;
	wire [4-1:0] node24619;
	wire [4-1:0] node24620;
	wire [4-1:0] node24621;
	wire [4-1:0] node24624;
	wire [4-1:0] node24627;
	wire [4-1:0] node24629;
	wire [4-1:0] node24632;
	wire [4-1:0] node24633;
	wire [4-1:0] node24634;
	wire [4-1:0] node24637;
	wire [4-1:0] node24640;
	wire [4-1:0] node24641;
	wire [4-1:0] node24644;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24649;
	wire [4-1:0] node24650;
	wire [4-1:0] node24651;
	wire [4-1:0] node24654;
	wire [4-1:0] node24657;
	wire [4-1:0] node24658;
	wire [4-1:0] node24661;
	wire [4-1:0] node24664;
	wire [4-1:0] node24665;
	wire [4-1:0] node24666;
	wire [4-1:0] node24668;
	wire [4-1:0] node24669;
	wire [4-1:0] node24672;
	wire [4-1:0] node24675;
	wire [4-1:0] node24676;
	wire [4-1:0] node24679;
	wire [4-1:0] node24682;
	wire [4-1:0] node24683;
	wire [4-1:0] node24686;
	wire [4-1:0] node24689;
	wire [4-1:0] node24690;
	wire [4-1:0] node24691;
	wire [4-1:0] node24692;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24698;
	wire [4-1:0] node24699;
	wire [4-1:0] node24700;
	wire [4-1:0] node24704;
	wire [4-1:0] node24705;
	wire [4-1:0] node24709;
	wire [4-1:0] node24710;
	wire [4-1:0] node24711;
	wire [4-1:0] node24712;
	wire [4-1:0] node24715;
	wire [4-1:0] node24718;
	wire [4-1:0] node24719;
	wire [4-1:0] node24722;
	wire [4-1:0] node24725;
	wire [4-1:0] node24726;
	wire [4-1:0] node24728;
	wire [4-1:0] node24731;
	wire [4-1:0] node24732;
	wire [4-1:0] node24736;
	wire [4-1:0] node24737;
	wire [4-1:0] node24738;
	wire [4-1:0] node24739;
	wire [4-1:0] node24744;
	wire [4-1:0] node24745;
	wire [4-1:0] node24748;
	wire [4-1:0] node24751;
	wire [4-1:0] node24752;
	wire [4-1:0] node24753;
	wire [4-1:0] node24754;
	wire [4-1:0] node24755;
	wire [4-1:0] node24756;
	wire [4-1:0] node24760;
	wire [4-1:0] node24761;
	wire [4-1:0] node24765;
	wire [4-1:0] node24766;
	wire [4-1:0] node24767;
	wire [4-1:0] node24772;
	wire [4-1:0] node24773;
	wire [4-1:0] node24774;
	wire [4-1:0] node24775;
	wire [4-1:0] node24779;
	wire [4-1:0] node24780;
	wire [4-1:0] node24783;
	wire [4-1:0] node24787;
	wire [4-1:0] node24788;
	wire [4-1:0] node24789;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24794;
	wire [4-1:0] node24798;
	wire [4-1:0] node24800;
	wire [4-1:0] node24801;
	wire [4-1:0] node24805;
	wire [4-1:0] node24806;
	wire [4-1:0] node24807;
	wire [4-1:0] node24809;
	wire [4-1:0] node24812;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24819;
	wire [4-1:0] node24822;
	wire [4-1:0] node24823;
	wire [4-1:0] node24824;
	wire [4-1:0] node24825;
	wire [4-1:0] node24826;
	wire [4-1:0] node24827;
	wire [4-1:0] node24830;
	wire [4-1:0] node24833;
	wire [4-1:0] node24834;
	wire [4-1:0] node24835;
	wire [4-1:0] node24836;
	wire [4-1:0] node24837;
	wire [4-1:0] node24838;
	wire [4-1:0] node24841;
	wire [4-1:0] node24844;
	wire [4-1:0] node24846;
	wire [4-1:0] node24847;
	wire [4-1:0] node24850;
	wire [4-1:0] node24853;
	wire [4-1:0] node24854;
	wire [4-1:0] node24857;
	wire [4-1:0] node24860;
	wire [4-1:0] node24861;
	wire [4-1:0] node24862;
	wire [4-1:0] node24865;
	wire [4-1:0] node24868;
	wire [4-1:0] node24869;
	wire [4-1:0] node24870;
	wire [4-1:0] node24871;
	wire [4-1:0] node24875;
	wire [4-1:0] node24877;
	wire [4-1:0] node24880;
	wire [4-1:0] node24881;
	wire [4-1:0] node24884;
	wire [4-1:0] node24887;
	wire [4-1:0] node24888;
	wire [4-1:0] node24889;
	wire [4-1:0] node24890;
	wire [4-1:0] node24893;
	wire [4-1:0] node24896;
	wire [4-1:0] node24897;
	wire [4-1:0] node24898;
	wire [4-1:0] node24901;
	wire [4-1:0] node24905;
	wire [4-1:0] node24906;
	wire [4-1:0] node24907;
	wire [4-1:0] node24908;
	wire [4-1:0] node24909;
	wire [4-1:0] node24912;
	wire [4-1:0] node24916;
	wire [4-1:0] node24917;
	wire [4-1:0] node24920;
	wire [4-1:0] node24923;
	wire [4-1:0] node24924;
	wire [4-1:0] node24928;
	wire [4-1:0] node24929;
	wire [4-1:0] node24930;
	wire [4-1:0] node24931;
	wire [4-1:0] node24932;
	wire [4-1:0] node24934;
	wire [4-1:0] node24937;
	wire [4-1:0] node24938;
	wire [4-1:0] node24940;
	wire [4-1:0] node24942;
	wire [4-1:0] node24945;
	wire [4-1:0] node24946;
	wire [4-1:0] node24950;
	wire [4-1:0] node24951;
	wire [4-1:0] node24953;
	wire [4-1:0] node24956;
	wire [4-1:0] node24957;
	wire [4-1:0] node24960;
	wire [4-1:0] node24963;
	wire [4-1:0] node24964;
	wire [4-1:0] node24965;
	wire [4-1:0] node24967;
	wire [4-1:0] node24970;
	wire [4-1:0] node24971;
	wire [4-1:0] node24972;
	wire [4-1:0] node24975;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24982;
	wire [4-1:0] node24985;
	wire [4-1:0] node24986;
	wire [4-1:0] node24988;
	wire [4-1:0] node24991;
	wire [4-1:0] node24992;
	wire [4-1:0] node24995;
	wire [4-1:0] node24996;
	wire [4-1:0] node25000;
	wire [4-1:0] node25001;
	wire [4-1:0] node25002;
	wire [4-1:0] node25003;
	wire [4-1:0] node25005;
	wire [4-1:0] node25008;
	wire [4-1:0] node25010;
	wire [4-1:0] node25013;
	wire [4-1:0] node25014;
	wire [4-1:0] node25015;
	wire [4-1:0] node25016;
	wire [4-1:0] node25019;
	wire [4-1:0] node25022;
	wire [4-1:0] node25023;
	wire [4-1:0] node25027;
	wire [4-1:0] node25029;
	wire [4-1:0] node25031;
	wire [4-1:0] node25032;
	wire [4-1:0] node25035;
	wire [4-1:0] node25038;
	wire [4-1:0] node25039;
	wire [4-1:0] node25040;
	wire [4-1:0] node25042;
	wire [4-1:0] node25045;
	wire [4-1:0] node25046;
	wire [4-1:0] node25047;
	wire [4-1:0] node25049;
	wire [4-1:0] node25052;
	wire [4-1:0] node25054;
	wire [4-1:0] node25057;
	wire [4-1:0] node25058;
	wire [4-1:0] node25061;
	wire [4-1:0] node25064;
	wire [4-1:0] node25065;
	wire [4-1:0] node25067;
	wire [4-1:0] node25070;
	wire [4-1:0] node25071;
	wire [4-1:0] node25075;
	wire [4-1:0] node25076;
	wire [4-1:0] node25077;
	wire [4-1:0] node25078;
	wire [4-1:0] node25081;
	wire [4-1:0] node25084;
	wire [4-1:0] node25085;
	wire [4-1:0] node25086;
	wire [4-1:0] node25087;
	wire [4-1:0] node25088;
	wire [4-1:0] node25090;
	wire [4-1:0] node25093;
	wire [4-1:0] node25095;
	wire [4-1:0] node25098;
	wire [4-1:0] node25099;
	wire [4-1:0] node25100;
	wire [4-1:0] node25101;
	wire [4-1:0] node25104;
	wire [4-1:0] node25109;
	wire [4-1:0] node25110;
	wire [4-1:0] node25113;
	wire [4-1:0] node25116;
	wire [4-1:0] node25117;
	wire [4-1:0] node25118;
	wire [4-1:0] node25119;
	wire [4-1:0] node25120;
	wire [4-1:0] node25121;
	wire [4-1:0] node25126;
	wire [4-1:0] node25128;
	wire [4-1:0] node25131;
	wire [4-1:0] node25132;
	wire [4-1:0] node25133;
	wire [4-1:0] node25137;
	wire [4-1:0] node25138;
	wire [4-1:0] node25142;
	wire [4-1:0] node25143;
	wire [4-1:0] node25144;
	wire [4-1:0] node25145;
	wire [4-1:0] node25149;
	wire [4-1:0] node25150;
	wire [4-1:0] node25152;
	wire [4-1:0] node25155;
	wire [4-1:0] node25156;
	wire [4-1:0] node25160;
	wire [4-1:0] node25161;
	wire [4-1:0] node25162;
	wire [4-1:0] node25165;
	wire [4-1:0] node25168;
	wire [4-1:0] node25169;
	wire [4-1:0] node25170;
	wire [4-1:0] node25173;
	wire [4-1:0] node25176;
	wire [4-1:0] node25178;
	wire [4-1:0] node25181;
	wire [4-1:0] node25182;
	wire [4-1:0] node25183;
	wire [4-1:0] node25184;
	wire [4-1:0] node25185;
	wire [4-1:0] node25187;
	wire [4-1:0] node25189;
	wire [4-1:0] node25190;
	wire [4-1:0] node25193;
	wire [4-1:0] node25196;
	wire [4-1:0] node25197;
	wire [4-1:0] node25198;
	wire [4-1:0] node25202;
	wire [4-1:0] node25203;
	wire [4-1:0] node25204;
	wire [4-1:0] node25207;
	wire [4-1:0] node25210;
	wire [4-1:0] node25211;
	wire [4-1:0] node25215;
	wire [4-1:0] node25216;
	wire [4-1:0] node25217;
	wire [4-1:0] node25219;
	wire [4-1:0] node25222;
	wire [4-1:0] node25225;
	wire [4-1:0] node25226;
	wire [4-1:0] node25229;
	wire [4-1:0] node25231;
	wire [4-1:0] node25232;
	wire [4-1:0] node25236;
	wire [4-1:0] node25237;
	wire [4-1:0] node25238;
	wire [4-1:0] node25239;
	wire [4-1:0] node25240;
	wire [4-1:0] node25242;
	wire [4-1:0] node25245;
	wire [4-1:0] node25246;
	wire [4-1:0] node25249;
	wire [4-1:0] node25252;
	wire [4-1:0] node25253;
	wire [4-1:0] node25257;
	wire [4-1:0] node25258;
	wire [4-1:0] node25261;
	wire [4-1:0] node25262;
	wire [4-1:0] node25263;
	wire [4-1:0] node25267;
	wire [4-1:0] node25269;
	wire [4-1:0] node25272;
	wire [4-1:0] node25273;
	wire [4-1:0] node25274;
	wire [4-1:0] node25275;
	wire [4-1:0] node25277;
	wire [4-1:0] node25280;
	wire [4-1:0] node25281;
	wire [4-1:0] node25285;
	wire [4-1:0] node25286;
	wire [4-1:0] node25287;
	wire [4-1:0] node25292;
	wire [4-1:0] node25294;
	wire [4-1:0] node25296;
	wire [4-1:0] node25299;
	wire [4-1:0] node25300;
	wire [4-1:0] node25301;
	wire [4-1:0] node25302;
	wire [4-1:0] node25303;
	wire [4-1:0] node25304;
	wire [4-1:0] node25305;
	wire [4-1:0] node25309;
	wire [4-1:0] node25312;
	wire [4-1:0] node25313;
	wire [4-1:0] node25316;
	wire [4-1:0] node25319;
	wire [4-1:0] node25320;
	wire [4-1:0] node25323;
	wire [4-1:0] node25324;
	wire [4-1:0] node25328;
	wire [4-1:0] node25329;
	wire [4-1:0] node25330;
	wire [4-1:0] node25332;
	wire [4-1:0] node25333;
	wire [4-1:0] node25337;
	wire [4-1:0] node25339;
	wire [4-1:0] node25342;
	wire [4-1:0] node25343;
	wire [4-1:0] node25344;
	wire [4-1:0] node25347;
	wire [4-1:0] node25350;
	wire [4-1:0] node25351;
	wire [4-1:0] node25354;
	wire [4-1:0] node25357;
	wire [4-1:0] node25358;
	wire [4-1:0] node25359;
	wire [4-1:0] node25360;
	wire [4-1:0] node25362;
	wire [4-1:0] node25364;
	wire [4-1:0] node25367;
	wire [4-1:0] node25368;
	wire [4-1:0] node25369;
	wire [4-1:0] node25372;
	wire [4-1:0] node25376;
	wire [4-1:0] node25377;
	wire [4-1:0] node25378;
	wire [4-1:0] node25379;
	wire [4-1:0] node25382;
	wire [4-1:0] node25385;
	wire [4-1:0] node25386;
	wire [4-1:0] node25389;
	wire [4-1:0] node25392;
	wire [4-1:0] node25393;
	wire [4-1:0] node25396;
	wire [4-1:0] node25399;
	wire [4-1:0] node25400;
	wire [4-1:0] node25401;
	wire [4-1:0] node25404;
	wire [4-1:0] node25407;
	wire [4-1:0] node25408;
	wire [4-1:0] node25409;
	wire [4-1:0] node25412;
	wire [4-1:0] node25415;
	wire [4-1:0] node25416;
	wire [4-1:0] node25419;
	wire [4-1:0] node25421;
	wire [4-1:0] node25424;
	wire [4-1:0] node25425;
	wire [4-1:0] node25426;
	wire [4-1:0] node25427;
	wire [4-1:0] node25428;
	wire [4-1:0] node25429;
	wire [4-1:0] node25430;
	wire [4-1:0] node25431;
	wire [4-1:0] node25435;
	wire [4-1:0] node25436;
	wire [4-1:0] node25440;
	wire [4-1:0] node25441;
	wire [4-1:0] node25443;
	wire [4-1:0] node25446;
	wire [4-1:0] node25448;
	wire [4-1:0] node25451;
	wire [4-1:0] node25452;
	wire [4-1:0] node25453;
	wire [4-1:0] node25454;
	wire [4-1:0] node25456;
	wire [4-1:0] node25457;
	wire [4-1:0] node25460;
	wire [4-1:0] node25463;
	wire [4-1:0] node25465;
	wire [4-1:0] node25466;
	wire [4-1:0] node25470;
	wire [4-1:0] node25472;
	wire [4-1:0] node25473;
	wire [4-1:0] node25474;
	wire [4-1:0] node25478;
	wire [4-1:0] node25480;
	wire [4-1:0] node25483;
	wire [4-1:0] node25484;
	wire [4-1:0] node25485;
	wire [4-1:0] node25486;
	wire [4-1:0] node25489;
	wire [4-1:0] node25492;
	wire [4-1:0] node25493;
	wire [4-1:0] node25494;
	wire [4-1:0] node25498;
	wire [4-1:0] node25500;
	wire [4-1:0] node25503;
	wire [4-1:0] node25504;
	wire [4-1:0] node25505;
	wire [4-1:0] node25508;
	wire [4-1:0] node25512;
	wire [4-1:0] node25513;
	wire [4-1:0] node25514;
	wire [4-1:0] node25515;
	wire [4-1:0] node25516;
	wire [4-1:0] node25518;
	wire [4-1:0] node25521;
	wire [4-1:0] node25522;
	wire [4-1:0] node25524;
	wire [4-1:0] node25527;
	wire [4-1:0] node25528;
	wire [4-1:0] node25532;
	wire [4-1:0] node25533;
	wire [4-1:0] node25536;
	wire [4-1:0] node25539;
	wire [4-1:0] node25540;
	wire [4-1:0] node25541;
	wire [4-1:0] node25542;
	wire [4-1:0] node25545;
	wire [4-1:0] node25548;
	wire [4-1:0] node25549;
	wire [4-1:0] node25550;
	wire [4-1:0] node25554;
	wire [4-1:0] node25557;
	wire [4-1:0] node25558;
	wire [4-1:0] node25559;
	wire [4-1:0] node25562;
	wire [4-1:0] node25565;
	wire [4-1:0] node25566;
	wire [4-1:0] node25568;
	wire [4-1:0] node25571;
	wire [4-1:0] node25572;
	wire [4-1:0] node25576;
	wire [4-1:0] node25577;
	wire [4-1:0] node25578;
	wire [4-1:0] node25579;
	wire [4-1:0] node25580;
	wire [4-1:0] node25583;
	wire [4-1:0] node25586;
	wire [4-1:0] node25587;
	wire [4-1:0] node25590;
	wire [4-1:0] node25593;
	wire [4-1:0] node25594;
	wire [4-1:0] node25595;
	wire [4-1:0] node25598;
	wire [4-1:0] node25602;
	wire [4-1:0] node25603;
	wire [4-1:0] node25606;
	wire [4-1:0] node25609;
	wire [4-1:0] node25610;
	wire [4-1:0] node25611;
	wire [4-1:0] node25612;
	wire [4-1:0] node25613;
	wire [4-1:0] node25614;
	wire [4-1:0] node25615;
	wire [4-1:0] node25618;
	wire [4-1:0] node25622;
	wire [4-1:0] node25623;
	wire [4-1:0] node25624;
	wire [4-1:0] node25627;
	wire [4-1:0] node25631;
	wire [4-1:0] node25633;
	wire [4-1:0] node25634;
	wire [4-1:0] node25635;
	wire [4-1:0] node25639;
	wire [4-1:0] node25640;
	wire [4-1:0] node25644;
	wire [4-1:0] node25645;
	wire [4-1:0] node25646;
	wire [4-1:0] node25647;
	wire [4-1:0] node25648;
	wire [4-1:0] node25649;
	wire [4-1:0] node25652;
	wire [4-1:0] node25656;
	wire [4-1:0] node25657;
	wire [4-1:0] node25658;
	wire [4-1:0] node25661;
	wire [4-1:0] node25664;
	wire [4-1:0] node25665;
	wire [4-1:0] node25668;
	wire [4-1:0] node25671;
	wire [4-1:0] node25672;
	wire [4-1:0] node25676;
	wire [4-1:0] node25677;
	wire [4-1:0] node25678;
	wire [4-1:0] node25679;
	wire [4-1:0] node25682;
	wire [4-1:0] node25685;
	wire [4-1:0] node25686;
	wire [4-1:0] node25687;
	wire [4-1:0] node25690;
	wire [4-1:0] node25694;
	wire [4-1:0] node25695;
	wire [4-1:0] node25699;
	wire [4-1:0] node25700;
	wire [4-1:0] node25701;
	wire [4-1:0] node25703;
	wire [4-1:0] node25704;
	wire [4-1:0] node25708;
	wire [4-1:0] node25710;
	wire [4-1:0] node25711;
	wire [4-1:0] node25715;
	wire [4-1:0] node25716;
	wire [4-1:0] node25718;
	wire [4-1:0] node25719;
	wire [4-1:0] node25723;
	wire [4-1:0] node25724;
	wire [4-1:0] node25726;
	wire [4-1:0] node25730;
	wire [4-1:0] node25731;
	wire [4-1:0] node25732;
	wire [4-1:0] node25733;
	wire [4-1:0] node25734;
	wire [4-1:0] node25735;
	wire [4-1:0] node25736;
	wire [4-1:0] node25740;
	wire [4-1:0] node25741;
	wire [4-1:0] node25744;
	wire [4-1:0] node25747;
	wire [4-1:0] node25748;
	wire [4-1:0] node25749;
	wire [4-1:0] node25752;
	wire [4-1:0] node25755;
	wire [4-1:0] node25756;
	wire [4-1:0] node25760;
	wire [4-1:0] node25761;
	wire [4-1:0] node25763;
	wire [4-1:0] node25764;
	wire [4-1:0] node25768;
	wire [4-1:0] node25770;
	wire [4-1:0] node25772;
	wire [4-1:0] node25775;
	wire [4-1:0] node25776;
	wire [4-1:0] node25777;
	wire [4-1:0] node25778;
	wire [4-1:0] node25779;
	wire [4-1:0] node25783;
	wire [4-1:0] node25784;
	wire [4-1:0] node25787;
	wire [4-1:0] node25790;
	wire [4-1:0] node25791;
	wire [4-1:0] node25792;
	wire [4-1:0] node25794;
	wire [4-1:0] node25798;
	wire [4-1:0] node25799;
	wire [4-1:0] node25800;
	wire [4-1:0] node25804;
	wire [4-1:0] node25805;
	wire [4-1:0] node25809;
	wire [4-1:0] node25810;
	wire [4-1:0] node25812;
	wire [4-1:0] node25813;
	wire [4-1:0] node25817;
	wire [4-1:0] node25818;
	wire [4-1:0] node25820;
	wire [4-1:0] node25824;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25828;
	wire [4-1:0] node25829;
	wire [4-1:0] node25833;
	wire [4-1:0] node25834;
	wire [4-1:0] node25837;
	wire [4-1:0] node25840;
	wire [4-1:0] node25841;
	wire [4-1:0] node25842;
	wire [4-1:0] node25843;
	wire [4-1:0] node25846;
	wire [4-1:0] node25849;
	wire [4-1:0] node25850;
	wire [4-1:0] node25853;
	wire [4-1:0] node25856;
	wire [4-1:0] node25857;
	wire [4-1:0] node25861;
	wire [4-1:0] node25862;
	wire [4-1:0] node25864;
	wire [4-1:0] node25865;
	wire [4-1:0] node25869;
	wire [4-1:0] node25870;
	wire [4-1:0] node25872;
	wire [4-1:0] node25876;
	wire [4-1:0] node25877;
	wire [4-1:0] node25878;
	wire [4-1:0] node25879;
	wire [4-1:0] node25880;
	wire [4-1:0] node25883;
	wire [4-1:0] node25886;
	wire [4-1:0] node25887;
	wire [4-1:0] node25888;
	wire [4-1:0] node25889;
	wire [4-1:0] node25893;
	wire [4-1:0] node25895;
	wire [4-1:0] node25898;
	wire [4-1:0] node25900;
	wire [4-1:0] node25903;
	wire [4-1:0] node25904;
	wire [4-1:0] node25906;
	wire [4-1:0] node25909;
	wire [4-1:0] node25911;
	wire [4-1:0] node25914;
	wire [4-1:0] node25915;
	wire [4-1:0] node25916;
	wire [4-1:0] node25918;
	wire [4-1:0] node25921;
	wire [4-1:0] node25922;
	wire [4-1:0] node25926;
	wire [4-1:0] node25929;
	wire [4-1:0] node25930;
	wire [4-1:0] node25931;
	wire [4-1:0] node25932;
	wire [4-1:0] node25933;
	wire [4-1:0] node25934;
	wire [4-1:0] node25935;
	wire [4-1:0] node25936;
	wire [4-1:0] node25937;
	wire [4-1:0] node25938;
	wire [4-1:0] node25942;
	wire [4-1:0] node25944;
	wire [4-1:0] node25947;
	wire [4-1:0] node25948;
	wire [4-1:0] node25950;
	wire [4-1:0] node25953;
	wire [4-1:0] node25954;
	wire [4-1:0] node25958;
	wire [4-1:0] node25959;
	wire [4-1:0] node25960;
	wire [4-1:0] node25961;
	wire [4-1:0] node25963;
	wire [4-1:0] node25966;
	wire [4-1:0] node25967;
	wire [4-1:0] node25971;
	wire [4-1:0] node25972;
	wire [4-1:0] node25973;
	wire [4-1:0] node25977;
	wire [4-1:0] node25978;
	wire [4-1:0] node25982;
	wire [4-1:0] node25983;
	wire [4-1:0] node25984;
	wire [4-1:0] node25985;
	wire [4-1:0] node25988;
	wire [4-1:0] node25991;
	wire [4-1:0] node25992;
	wire [4-1:0] node25995;
	wire [4-1:0] node25998;
	wire [4-1:0] node25999;
	wire [4-1:0] node26000;
	wire [4-1:0] node26003;
	wire [4-1:0] node26006;
	wire [4-1:0] node26007;
	wire [4-1:0] node26010;
	wire [4-1:0] node26012;
	wire [4-1:0] node26015;
	wire [4-1:0] node26016;
	wire [4-1:0] node26017;
	wire [4-1:0] node26018;
	wire [4-1:0] node26019;
	wire [4-1:0] node26023;
	wire [4-1:0] node26025;
	wire [4-1:0] node26028;
	wire [4-1:0] node26029;
	wire [4-1:0] node26030;
	wire [4-1:0] node26034;
	wire [4-1:0] node26035;
	wire [4-1:0] node26039;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26042;
	wire [4-1:0] node26045;
	wire [4-1:0] node26048;
	wire [4-1:0] node26049;
	wire [4-1:0] node26052;
	wire [4-1:0] node26055;
	wire [4-1:0] node26056;
	wire [4-1:0] node26057;
	wire [4-1:0] node26058;
	wire [4-1:0] node26059;
	wire [4-1:0] node26062;
	wire [4-1:0] node26066;
	wire [4-1:0] node26068;
	wire [4-1:0] node26069;
	wire [4-1:0] node26073;
	wire [4-1:0] node26074;
	wire [4-1:0] node26077;
	wire [4-1:0] node26080;
	wire [4-1:0] node26081;
	wire [4-1:0] node26082;
	wire [4-1:0] node26083;
	wire [4-1:0] node26084;
	wire [4-1:0] node26085;
	wire [4-1:0] node26086;
	wire [4-1:0] node26090;
	wire [4-1:0] node26091;
	wire [4-1:0] node26095;
	wire [4-1:0] node26096;
	wire [4-1:0] node26098;
	wire [4-1:0] node26099;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26106;
	wire [4-1:0] node26109;
	wire [4-1:0] node26112;
	wire [4-1:0] node26113;
	wire [4-1:0] node26115;
	wire [4-1:0] node26116;
	wire [4-1:0] node26120;
	wire [4-1:0] node26121;
	wire [4-1:0] node26123;
	wire [4-1:0] node26127;
	wire [4-1:0] node26128;
	wire [4-1:0] node26129;
	wire [4-1:0] node26131;
	wire [4-1:0] node26134;
	wire [4-1:0] node26136;
	wire [4-1:0] node26139;
	wire [4-1:0] node26140;
	wire [4-1:0] node26142;
	wire [4-1:0] node26145;
	wire [4-1:0] node26147;
	wire [4-1:0] node26150;
	wire [4-1:0] node26151;
	wire [4-1:0] node26152;
	wire [4-1:0] node26153;
	wire [4-1:0] node26154;
	wire [4-1:0] node26158;
	wire [4-1:0] node26159;
	wire [4-1:0] node26163;
	wire [4-1:0] node26164;
	wire [4-1:0] node26166;
	wire [4-1:0] node26169;
	wire [4-1:0] node26171;
	wire [4-1:0] node26174;
	wire [4-1:0] node26175;
	wire [4-1:0] node26176;
	wire [4-1:0] node26178;
	wire [4-1:0] node26181;
	wire [4-1:0] node26183;
	wire [4-1:0] node26186;
	wire [4-1:0] node26187;
	wire [4-1:0] node26189;
	wire [4-1:0] node26192;
	wire [4-1:0] node26194;
	wire [4-1:0] node26197;
	wire [4-1:0] node26198;
	wire [4-1:0] node26199;
	wire [4-1:0] node26200;
	wire [4-1:0] node26201;
	wire [4-1:0] node26202;
	wire [4-1:0] node26203;
	wire [4-1:0] node26207;
	wire [4-1:0] node26208;
	wire [4-1:0] node26212;
	wire [4-1:0] node26213;
	wire [4-1:0] node26215;
	wire [4-1:0] node26218;
	wire [4-1:0] node26219;
	wire [4-1:0] node26223;
	wire [4-1:0] node26224;
	wire [4-1:0] node26225;
	wire [4-1:0] node26227;
	wire [4-1:0] node26230;
	wire [4-1:0] node26231;
	wire [4-1:0] node26235;
	wire [4-1:0] node26236;
	wire [4-1:0] node26238;
	wire [4-1:0] node26241;
	wire [4-1:0] node26242;
	wire [4-1:0] node26246;
	wire [4-1:0] node26247;
	wire [4-1:0] node26248;
	wire [4-1:0] node26249;
	wire [4-1:0] node26251;
	wire [4-1:0] node26254;
	wire [4-1:0] node26255;
	wire [4-1:0] node26259;
	wire [4-1:0] node26260;
	wire [4-1:0] node26262;
	wire [4-1:0] node26265;
	wire [4-1:0] node26266;
	wire [4-1:0] node26270;
	wire [4-1:0] node26271;
	wire [4-1:0] node26272;
	wire [4-1:0] node26273;
	wire [4-1:0] node26274;
	wire [4-1:0] node26277;
	wire [4-1:0] node26280;
	wire [4-1:0] node26282;
	wire [4-1:0] node26285;
	wire [4-1:0] node26286;
	wire [4-1:0] node26289;
	wire [4-1:0] node26292;
	wire [4-1:0] node26293;
	wire [4-1:0] node26294;
	wire [4-1:0] node26295;
	wire [4-1:0] node26296;
	wire [4-1:0] node26299;
	wire [4-1:0] node26302;
	wire [4-1:0] node26303;
	wire [4-1:0] node26306;
	wire [4-1:0] node26309;
	wire [4-1:0] node26310;
	wire [4-1:0] node26313;
	wire [4-1:0] node26316;
	wire [4-1:0] node26318;
	wire [4-1:0] node26320;
	wire [4-1:0] node26323;
	wire [4-1:0] node26324;
	wire [4-1:0] node26325;
	wire [4-1:0] node26326;
	wire [4-1:0] node26327;
	wire [4-1:0] node26329;
	wire [4-1:0] node26332;
	wire [4-1:0] node26334;
	wire [4-1:0] node26337;
	wire [4-1:0] node26338;
	wire [4-1:0] node26340;
	wire [4-1:0] node26343;
	wire [4-1:0] node26344;
	wire [4-1:0] node26348;
	wire [4-1:0] node26349;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26352;
	wire [4-1:0] node26355;
	wire [4-1:0] node26359;
	wire [4-1:0] node26360;
	wire [4-1:0] node26363;
	wire [4-1:0] node26366;
	wire [4-1:0] node26367;
	wire [4-1:0] node26368;
	wire [4-1:0] node26372;
	wire [4-1:0] node26373;
	wire [4-1:0] node26376;
	wire [4-1:0] node26379;
	wire [4-1:0] node26380;
	wire [4-1:0] node26381;
	wire [4-1:0] node26382;
	wire [4-1:0] node26385;
	wire [4-1:0] node26388;
	wire [4-1:0] node26389;
	wire [4-1:0] node26390;
	wire [4-1:0] node26393;
	wire [4-1:0] node26396;
	wire [4-1:0] node26397;
	wire [4-1:0] node26400;
	wire [4-1:0] node26403;
	wire [4-1:0] node26404;
	wire [4-1:0] node26405;
	wire [4-1:0] node26406;
	wire [4-1:0] node26408;
	wire [4-1:0] node26409;
	wire [4-1:0] node26412;
	wire [4-1:0] node26415;
	wire [4-1:0] node26416;
	wire [4-1:0] node26419;
	wire [4-1:0] node26422;
	wire [4-1:0] node26423;
	wire [4-1:0] node26424;
	wire [4-1:0] node26427;
	wire [4-1:0] node26430;
	wire [4-1:0] node26431;
	wire [4-1:0] node26432;
	wire [4-1:0] node26435;
	wire [4-1:0] node26438;
	wire [4-1:0] node26439;
	wire [4-1:0] node26442;
	wire [4-1:0] node26445;
	wire [4-1:0] node26446;
	wire [4-1:0] node26448;
	wire [4-1:0] node26451;
	wire [4-1:0] node26452;
	wire [4-1:0] node26453;
	wire [4-1:0] node26457;
	wire [4-1:0] node26458;
	wire [4-1:0] node26462;
	wire [4-1:0] node26463;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26466;
	wire [4-1:0] node26467;
	wire [4-1:0] node26468;
	wire [4-1:0] node26469;
	wire [4-1:0] node26472;
	wire [4-1:0] node26475;
	wire [4-1:0] node26476;
	wire [4-1:0] node26479;
	wire [4-1:0] node26482;
	wire [4-1:0] node26483;
	wire [4-1:0] node26484;
	wire [4-1:0] node26488;
	wire [4-1:0] node26489;
	wire [4-1:0] node26493;
	wire [4-1:0] node26494;
	wire [4-1:0] node26495;
	wire [4-1:0] node26496;
	wire [4-1:0] node26499;
	wire [4-1:0] node26502;
	wire [4-1:0] node26503;
	wire [4-1:0] node26507;
	wire [4-1:0] node26508;
	wire [4-1:0] node26509;
	wire [4-1:0] node26513;
	wire [4-1:0] node26514;
	wire [4-1:0] node26518;
	wire [4-1:0] node26519;
	wire [4-1:0] node26520;
	wire [4-1:0] node26521;
	wire [4-1:0] node26523;
	wire [4-1:0] node26526;
	wire [4-1:0] node26527;
	wire [4-1:0] node26530;
	wire [4-1:0] node26533;
	wire [4-1:0] node26534;
	wire [4-1:0] node26538;
	wire [4-1:0] node26539;
	wire [4-1:0] node26540;
	wire [4-1:0] node26544;
	wire [4-1:0] node26545;
	wire [4-1:0] node26546;
	wire [4-1:0] node26551;
	wire [4-1:0] node26552;
	wire [4-1:0] node26553;
	wire [4-1:0] node26554;
	wire [4-1:0] node26555;
	wire [4-1:0] node26556;
	wire [4-1:0] node26559;
	wire [4-1:0] node26562;
	wire [4-1:0] node26563;
	wire [4-1:0] node26567;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26573;
	wire [4-1:0] node26574;
	wire [4-1:0] node26578;
	wire [4-1:0] node26579;
	wire [4-1:0] node26580;
	wire [4-1:0] node26581;
	wire [4-1:0] node26584;
	wire [4-1:0] node26587;
	wire [4-1:0] node26588;
	wire [4-1:0] node26591;
	wire [4-1:0] node26594;
	wire [4-1:0] node26595;
	wire [4-1:0] node26596;
	wire [4-1:0] node26599;
	wire [4-1:0] node26602;
	wire [4-1:0] node26605;
	wire [4-1:0] node26606;
	wire [4-1:0] node26607;
	wire [4-1:0] node26608;
	wire [4-1:0] node26610;
	wire [4-1:0] node26613;
	wire [4-1:0] node26614;
	wire [4-1:0] node26615;
	wire [4-1:0] node26616;
	wire [4-1:0] node26619;
	wire [4-1:0] node26623;
	wire [4-1:0] node26624;
	wire [4-1:0] node26625;
	wire [4-1:0] node26628;
	wire [4-1:0] node26631;
	wire [4-1:0] node26632;
	wire [4-1:0] node26636;
	wire [4-1:0] node26637;
	wire [4-1:0] node26641;
	wire [4-1:0] node26642;
	wire [4-1:0] node26643;
	wire [4-1:0] node26644;
	wire [4-1:0] node26647;
	wire [4-1:0] node26650;
	wire [4-1:0] node26651;
	wire [4-1:0] node26654;
	wire [4-1:0] node26657;
	wire [4-1:0] node26660;
	wire [4-1:0] node26661;
	wire [4-1:0] node26662;
	wire [4-1:0] node26663;
	wire [4-1:0] node26664;
	wire [4-1:0] node26665;
	wire [4-1:0] node26666;
	wire [4-1:0] node26669;
	wire [4-1:0] node26672;
	wire [4-1:0] node26673;
	wire [4-1:0] node26676;
	wire [4-1:0] node26679;
	wire [4-1:0] node26680;
	wire [4-1:0] node26681;
	wire [4-1:0] node26684;
	wire [4-1:0] node26687;
	wire [4-1:0] node26688;
	wire [4-1:0] node26692;
	wire [4-1:0] node26693;
	wire [4-1:0] node26694;
	wire [4-1:0] node26695;
	wire [4-1:0] node26696;
	wire [4-1:0] node26700;
	wire [4-1:0] node26702;
	wire [4-1:0] node26705;
	wire [4-1:0] node26706;
	wire [4-1:0] node26709;
	wire [4-1:0] node26712;
	wire [4-1:0] node26713;
	wire [4-1:0] node26714;
	wire [4-1:0] node26717;
	wire [4-1:0] node26720;
	wire [4-1:0] node26723;
	wire [4-1:0] node26724;
	wire [4-1:0] node26725;
	wire [4-1:0] node26726;
	wire [4-1:0] node26728;
	wire [4-1:0] node26731;
	wire [4-1:0] node26732;
	wire [4-1:0] node26735;
	wire [4-1:0] node26738;
	wire [4-1:0] node26739;
	wire [4-1:0] node26743;
	wire [4-1:0] node26744;
	wire [4-1:0] node26745;
	wire [4-1:0] node26747;
	wire [4-1:0] node26750;
	wire [4-1:0] node26753;
	wire [4-1:0] node26756;
	wire [4-1:0] node26757;
	wire [4-1:0] node26758;
	wire [4-1:0] node26759;
	wire [4-1:0] node26760;
	wire [4-1:0] node26761;
	wire [4-1:0] node26764;
	wire [4-1:0] node26767;
	wire [4-1:0] node26768;
	wire [4-1:0] node26771;
	wire [4-1:0] node26774;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26780;
	wire [4-1:0] node26781;
	wire [4-1:0] node26785;
	wire [4-1:0] node26786;
	wire [4-1:0] node26787;
	wire [4-1:0] node26788;
	wire [4-1:0] node26791;
	wire [4-1:0] node26794;
	wire [4-1:0] node26795;
	wire [4-1:0] node26799;
	wire [4-1:0] node26800;
	wire [4-1:0] node26801;
	wire [4-1:0] node26804;
	wire [4-1:0] node26807;
	wire [4-1:0] node26808;
	wire [4-1:0] node26812;
	wire [4-1:0] node26813;
	wire [4-1:0] node26814;
	wire [4-1:0] node26815;
	wire [4-1:0] node26817;
	wire [4-1:0] node26820;
	wire [4-1:0] node26821;
	wire [4-1:0] node26822;
	wire [4-1:0] node26826;
	wire [4-1:0] node26827;
	wire [4-1:0] node26830;
	wire [4-1:0] node26833;
	wire [4-1:0] node26834;
	wire [4-1:0] node26838;
	wire [4-1:0] node26839;
	wire [4-1:0] node26840;
	wire [4-1:0] node26844;
	wire [4-1:0] node26845;
	wire [4-1:0] node26846;
	wire [4-1:0] node26851;
	wire [4-1:0] node26852;
	wire [4-1:0] node26853;
	wire [4-1:0] node26854;
	wire [4-1:0] node26855;
	wire [4-1:0] node26856;
	wire [4-1:0] node26857;
	wire [4-1:0] node26858;
	wire [4-1:0] node26861;
	wire [4-1:0] node26864;
	wire [4-1:0] node26865;
	wire [4-1:0] node26868;
	wire [4-1:0] node26871;
	wire [4-1:0] node26872;
	wire [4-1:0] node26875;
	wire [4-1:0] node26878;
	wire [4-1:0] node26879;
	wire [4-1:0] node26880;
	wire [4-1:0] node26881;
	wire [4-1:0] node26883;
	wire [4-1:0] node26886;
	wire [4-1:0] node26887;
	wire [4-1:0] node26890;
	wire [4-1:0] node26893;
	wire [4-1:0] node26894;
	wire [4-1:0] node26895;
	wire [4-1:0] node26897;
	wire [4-1:0] node26898;
	wire [4-1:0] node26902;
	wire [4-1:0] node26903;
	wire [4-1:0] node26905;
	wire [4-1:0] node26909;
	wire [4-1:0] node26910;
	wire [4-1:0] node26911;
	wire [4-1:0] node26913;
	wire [4-1:0] node26916;
	wire [4-1:0] node26917;
	wire [4-1:0] node26921;
	wire [4-1:0] node26922;
	wire [4-1:0] node26923;
	wire [4-1:0] node26926;
	wire [4-1:0] node26930;
	wire [4-1:0] node26931;
	wire [4-1:0] node26932;
	wire [4-1:0] node26935;
	wire [4-1:0] node26938;
	wire [4-1:0] node26939;
	wire [4-1:0] node26942;
	wire [4-1:0] node26945;
	wire [4-1:0] node26946;
	wire [4-1:0] node26947;
	wire [4-1:0] node26948;
	wire [4-1:0] node26949;
	wire [4-1:0] node26951;
	wire [4-1:0] node26954;
	wire [4-1:0] node26955;
	wire [4-1:0] node26959;
	wire [4-1:0] node26960;
	wire [4-1:0] node26961;
	wire [4-1:0] node26965;
	wire [4-1:0] node26966;
	wire [4-1:0] node26970;
	wire [4-1:0] node26971;
	wire [4-1:0] node26972;
	wire [4-1:0] node26975;
	wire [4-1:0] node26978;
	wire [4-1:0] node26979;
	wire [4-1:0] node26981;
	wire [4-1:0] node26984;
	wire [4-1:0] node26985;
	wire [4-1:0] node26988;
	wire [4-1:0] node26991;
	wire [4-1:0] node26992;
	wire [4-1:0] node26993;
	wire [4-1:0] node26996;
	wire [4-1:0] node26999;
	wire [4-1:0] node27000;
	wire [4-1:0] node27001;
	wire [4-1:0] node27002;
	wire [4-1:0] node27006;
	wire [4-1:0] node27007;
	wire [4-1:0] node27008;
	wire [4-1:0] node27011;
	wire [4-1:0] node27013;
	wire [4-1:0] node27016;
	wire [4-1:0] node27018;
	wire [4-1:0] node27021;
	wire [4-1:0] node27022;
	wire [4-1:0] node27023;
	wire [4-1:0] node27025;
	wire [4-1:0] node27028;
	wire [4-1:0] node27029;
	wire [4-1:0] node27032;
	wire [4-1:0] node27035;
	wire [4-1:0] node27036;
	wire [4-1:0] node27037;
	wire [4-1:0] node27040;
	wire [4-1:0] node27043;
	wire [4-1:0] node27044;
	wire [4-1:0] node27046;
	wire [4-1:0] node27049;
	wire [4-1:0] node27050;
	wire [4-1:0] node27053;
	wire [4-1:0] node27056;
	wire [4-1:0] node27057;
	wire [4-1:0] node27058;
	wire [4-1:0] node27059;
	wire [4-1:0] node27060;
	wire [4-1:0] node27061;
	wire [4-1:0] node27062;
	wire [4-1:0] node27065;
	wire [4-1:0] node27068;
	wire [4-1:0] node27069;
	wire [4-1:0] node27072;
	wire [4-1:0] node27075;
	wire [4-1:0] node27076;
	wire [4-1:0] node27077;
	wire [4-1:0] node27078;
	wire [4-1:0] node27082;
	wire [4-1:0] node27083;
	wire [4-1:0] node27086;
	wire [4-1:0] node27089;
	wire [4-1:0] node27090;
	wire [4-1:0] node27093;
	wire [4-1:0] node27096;
	wire [4-1:0] node27097;
	wire [4-1:0] node27098;
	wire [4-1:0] node27101;
	wire [4-1:0] node27104;
	wire [4-1:0] node27105;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27112;
	wire [4-1:0] node27113;
	wire [4-1:0] node27114;
	wire [4-1:0] node27115;
	wire [4-1:0] node27118;
	wire [4-1:0] node27121;
	wire [4-1:0] node27122;
	wire [4-1:0] node27123;
	wire [4-1:0] node27124;
	wire [4-1:0] node27127;
	wire [4-1:0] node27131;
	wire [4-1:0] node27133;
	wire [4-1:0] node27134;
	wire [4-1:0] node27137;
	wire [4-1:0] node27140;
	wire [4-1:0] node27141;
	wire [4-1:0] node27144;
	wire [4-1:0] node27147;
	wire [4-1:0] node27148;
	wire [4-1:0] node27149;
	wire [4-1:0] node27150;
	wire [4-1:0] node27153;
	wire [4-1:0] node27156;
	wire [4-1:0] node27157;
	wire [4-1:0] node27160;
	wire [4-1:0] node27163;
	wire [4-1:0] node27164;
	wire [4-1:0] node27167;
	wire [4-1:0] node27170;
	wire [4-1:0] node27171;
	wire [4-1:0] node27172;
	wire [4-1:0] node27175;
	wire [4-1:0] node27178;
	wire [4-1:0] node27179;
	wire [4-1:0] node27180;
	wire [4-1:0] node27181;
	wire [4-1:0] node27182;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27187;
	wire [4-1:0] node27191;
	wire [4-1:0] node27192;
	wire [4-1:0] node27196;
	wire [4-1:0] node27197;
	wire [4-1:0] node27200;
	wire [4-1:0] node27203;
	wire [4-1:0] node27204;
	wire [4-1:0] node27205;
	wire [4-1:0] node27206;
	wire [4-1:0] node27210;
	wire [4-1:0] node27211;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27217;
	wire [4-1:0] node27221;
	wire [4-1:0] node27223;
	wire [4-1:0] node27225;
	wire [4-1:0] node27228;
	wire [4-1:0] node27229;
	wire [4-1:0] node27232;
	wire [4-1:0] node27235;
	wire [4-1:0] node27236;
	wire [4-1:0] node27237;
	wire [4-1:0] node27238;
	wire [4-1:0] node27239;
	wire [4-1:0] node27242;
	wire [4-1:0] node27245;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27248;
	wire [4-1:0] node27249;
	wire [4-1:0] node27252;
	wire [4-1:0] node27255;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27260;
	wire [4-1:0] node27263;
	wire [4-1:0] node27265;
	wire [4-1:0] node27266;
	wire [4-1:0] node27269;
	wire [4-1:0] node27272;
	wire [4-1:0] node27273;
	wire [4-1:0] node27276;
	wire [4-1:0] node27279;
	wire [4-1:0] node27280;
	wire [4-1:0] node27281;
	wire [4-1:0] node27284;
	wire [4-1:0] node27287;
	wire [4-1:0] node27288;
	wire [4-1:0] node27289;
	wire [4-1:0] node27290;
	wire [4-1:0] node27293;
	wire [4-1:0] node27297;
	wire [4-1:0] node27298;
	wire [4-1:0] node27300;
	wire [4-1:0] node27303;
	wire [4-1:0] node27304;
	wire [4-1:0] node27305;
	wire [4-1:0] node27309;
	wire [4-1:0] node27310;
	wire [4-1:0] node27313;
	wire [4-1:0] node27316;
	wire [4-1:0] node27317;
	wire [4-1:0] node27318;
	wire [4-1:0] node27319;
	wire [4-1:0] node27320;
	wire [4-1:0] node27324;
	wire [4-1:0] node27325;
	wire [4-1:0] node27329;
	wire [4-1:0] node27330;
	wire [4-1:0] node27331;
	wire [4-1:0] node27335;
	wire [4-1:0] node27336;
	wire [4-1:0] node27340;
	wire [4-1:0] node27341;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27344;
	wire [4-1:0] node27347;
	wire [4-1:0] node27350;
	wire [4-1:0] node27351;
	wire [4-1:0] node27352;
	wire [4-1:0] node27355;
	wire [4-1:0] node27358;
	wire [4-1:0] node27359;
	wire [4-1:0] node27363;
	wire [4-1:0] node27364;
	wire [4-1:0] node27365;
	wire [4-1:0] node27366;
	wire [4-1:0] node27370;
	wire [4-1:0] node27371;
	wire [4-1:0] node27374;
	wire [4-1:0] node27377;
	wire [4-1:0] node27379;
	wire [4-1:0] node27381;
	wire [4-1:0] node27384;
	wire [4-1:0] node27385;
	wire [4-1:0] node27386;
	wire [4-1:0] node27387;
	wire [4-1:0] node27391;
	wire [4-1:0] node27392;
	wire [4-1:0] node27396;
	wire [4-1:0] node27397;
	wire [4-1:0] node27398;
	wire [4-1:0] node27402;
	wire [4-1:0] node27403;
	wire [4-1:0] node27407;
	wire [4-1:0] node27408;
	wire [4-1:0] node27409;
	wire [4-1:0] node27413;
	wire [4-1:0] node27414;
	wire [4-1:0] node27418;
	wire [4-1:0] node27419;
	wire [4-1:0] node27420;
	wire [4-1:0] node27421;
	wire [4-1:0] node27422;
	wire [4-1:0] node27423;
	wire [4-1:0] node27424;
	wire [4-1:0] node27425;
	wire [4-1:0] node27426;
	wire [4-1:0] node27427;
	wire [4-1:0] node27428;
	wire [4-1:0] node27429;
	wire [4-1:0] node27430;
	wire [4-1:0] node27433;
	wire [4-1:0] node27436;
	wire [4-1:0] node27437;
	wire [4-1:0] node27439;
	wire [4-1:0] node27440;
	wire [4-1:0] node27444;
	wire [4-1:0] node27446;
	wire [4-1:0] node27449;
	wire [4-1:0] node27450;
	wire [4-1:0] node27451;
	wire [4-1:0] node27452;
	wire [4-1:0] node27456;
	wire [4-1:0] node27458;
	wire [4-1:0] node27461;
	wire [4-1:0] node27462;
	wire [4-1:0] node27464;
	wire [4-1:0] node27467;
	wire [4-1:0] node27469;
	wire [4-1:0] node27472;
	wire [4-1:0] node27473;
	wire [4-1:0] node27474;
	wire [4-1:0] node27476;
	wire [4-1:0] node27477;
	wire [4-1:0] node27480;
	wire [4-1:0] node27483;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27490;
	wire [4-1:0] node27491;
	wire [4-1:0] node27493;
	wire [4-1:0] node27495;
	wire [4-1:0] node27498;
	wire [4-1:0] node27500;
	wire [4-1:0] node27501;
	wire [4-1:0] node27504;
	wire [4-1:0] node27507;
	wire [4-1:0] node27508;
	wire [4-1:0] node27509;
	wire [4-1:0] node27510;
	wire [4-1:0] node27511;
	wire [4-1:0] node27515;
	wire [4-1:0] node27517;
	wire [4-1:0] node27520;
	wire [4-1:0] node27521;
	wire [4-1:0] node27523;
	wire [4-1:0] node27526;
	wire [4-1:0] node27528;
	wire [4-1:0] node27531;
	wire [4-1:0] node27532;
	wire [4-1:0] node27533;
	wire [4-1:0] node27534;
	wire [4-1:0] node27538;
	wire [4-1:0] node27539;
	wire [4-1:0] node27543;
	wire [4-1:0] node27544;
	wire [4-1:0] node27546;
	wire [4-1:0] node27549;
	wire [4-1:0] node27550;
	wire [4-1:0] node27554;
	wire [4-1:0] node27555;
	wire [4-1:0] node27556;
	wire [4-1:0] node27557;
	wire [4-1:0] node27558;
	wire [4-1:0] node27560;
	wire [4-1:0] node27562;
	wire [4-1:0] node27565;
	wire [4-1:0] node27566;
	wire [4-1:0] node27568;
	wire [4-1:0] node27571;
	wire [4-1:0] node27572;
	wire [4-1:0] node27575;
	wire [4-1:0] node27578;
	wire [4-1:0] node27579;
	wire [4-1:0] node27580;
	wire [4-1:0] node27581;
	wire [4-1:0] node27582;
	wire [4-1:0] node27586;
	wire [4-1:0] node27590;
	wire [4-1:0] node27591;
	wire [4-1:0] node27592;
	wire [4-1:0] node27596;
	wire [4-1:0] node27597;
	wire [4-1:0] node27601;
	wire [4-1:0] node27602;
	wire [4-1:0] node27603;
	wire [4-1:0] node27604;
	wire [4-1:0] node27606;
	wire [4-1:0] node27607;
	wire [4-1:0] node27611;
	wire [4-1:0] node27613;
	wire [4-1:0] node27616;
	wire [4-1:0] node27617;
	wire [4-1:0] node27619;
	wire [4-1:0] node27622;
	wire [4-1:0] node27624;
	wire [4-1:0] node27627;
	wire [4-1:0] node27628;
	wire [4-1:0] node27630;
	wire [4-1:0] node27633;
	wire [4-1:0] node27634;
	wire [4-1:0] node27635;
	wire [4-1:0] node27636;
	wire [4-1:0] node27639;
	wire [4-1:0] node27643;
	wire [4-1:0] node27644;
	wire [4-1:0] node27647;
	wire [4-1:0] node27650;
	wire [4-1:0] node27651;
	wire [4-1:0] node27652;
	wire [4-1:0] node27653;
	wire [4-1:0] node27654;
	wire [4-1:0] node27656;
	wire [4-1:0] node27659;
	wire [4-1:0] node27661;
	wire [4-1:0] node27664;
	wire [4-1:0] node27665;
	wire [4-1:0] node27667;
	wire [4-1:0] node27670;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27677;
	wire [4-1:0] node27678;
	wire [4-1:0] node27680;
	wire [4-1:0] node27683;
	wire [4-1:0] node27686;
	wire [4-1:0] node27687;
	wire [4-1:0] node27688;
	wire [4-1:0] node27689;
	wire [4-1:0] node27690;
	wire [4-1:0] node27693;
	wire [4-1:0] node27696;
	wire [4-1:0] node27698;
	wire [4-1:0] node27701;
	wire [4-1:0] node27702;
	wire [4-1:0] node27706;
	wire [4-1:0] node27707;
	wire [4-1:0] node27708;
	wire [4-1:0] node27711;
	wire [4-1:0] node27714;
	wire [4-1:0] node27715;
	wire [4-1:0] node27716;
	wire [4-1:0] node27717;
	wire [4-1:0] node27720;
	wire [4-1:0] node27723;
	wire [4-1:0] node27724;
	wire [4-1:0] node27728;
	wire [4-1:0] node27729;
	wire [4-1:0] node27731;
	wire [4-1:0] node27734;
	wire [4-1:0] node27735;
	wire [4-1:0] node27738;
	wire [4-1:0] node27741;
	wire [4-1:0] node27742;
	wire [4-1:0] node27743;
	wire [4-1:0] node27744;
	wire [4-1:0] node27745;
	wire [4-1:0] node27746;
	wire [4-1:0] node27747;
	wire [4-1:0] node27748;
	wire [4-1:0] node27750;
	wire [4-1:0] node27754;
	wire [4-1:0] node27757;
	wire [4-1:0] node27758;
	wire [4-1:0] node27760;
	wire [4-1:0] node27762;
	wire [4-1:0] node27766;
	wire [4-1:0] node27767;
	wire [4-1:0] node27768;
	wire [4-1:0] node27770;
	wire [4-1:0] node27772;
	wire [4-1:0] node27775;
	wire [4-1:0] node27776;
	wire [4-1:0] node27780;
	wire [4-1:0] node27781;
	wire [4-1:0] node27782;
	wire [4-1:0] node27786;
	wire [4-1:0] node27787;
	wire [4-1:0] node27790;
	wire [4-1:0] node27793;
	wire [4-1:0] node27794;
	wire [4-1:0] node27795;
	wire [4-1:0] node27796;
	wire [4-1:0] node27797;
	wire [4-1:0] node27801;
	wire [4-1:0] node27802;
	wire [4-1:0] node27803;
	wire [4-1:0] node27806;
	wire [4-1:0] node27809;
	wire [4-1:0] node27810;
	wire [4-1:0] node27813;
	wire [4-1:0] node27816;
	wire [4-1:0] node27818;
	wire [4-1:0] node27820;
	wire [4-1:0] node27821;
	wire [4-1:0] node27824;
	wire [4-1:0] node27827;
	wire [4-1:0] node27828;
	wire [4-1:0] node27829;
	wire [4-1:0] node27831;
	wire [4-1:0] node27832;
	wire [4-1:0] node27836;
	wire [4-1:0] node27838;
	wire [4-1:0] node27841;
	wire [4-1:0] node27842;
	wire [4-1:0] node27843;
	wire [4-1:0] node27844;
	wire [4-1:0] node27848;
	wire [4-1:0] node27851;
	wire [4-1:0] node27852;
	wire [4-1:0] node27856;
	wire [4-1:0] node27857;
	wire [4-1:0] node27858;
	wire [4-1:0] node27859;
	wire [4-1:0] node27860;
	wire [4-1:0] node27863;
	wire [4-1:0] node27866;
	wire [4-1:0] node27867;
	wire [4-1:0] node27868;
	wire [4-1:0] node27872;
	wire [4-1:0] node27874;
	wire [4-1:0] node27877;
	wire [4-1:0] node27878;
	wire [4-1:0] node27879;
	wire [4-1:0] node27880;
	wire [4-1:0] node27884;
	wire [4-1:0] node27885;
	wire [4-1:0] node27889;
	wire [4-1:0] node27890;
	wire [4-1:0] node27893;
	wire [4-1:0] node27894;
	wire [4-1:0] node27898;
	wire [4-1:0] node27899;
	wire [4-1:0] node27900;
	wire [4-1:0] node27901;
	wire [4-1:0] node27902;
	wire [4-1:0] node27906;
	wire [4-1:0] node27909;
	wire [4-1:0] node27910;
	wire [4-1:0] node27911;
	wire [4-1:0] node27915;
	wire [4-1:0] node27916;
	wire [4-1:0] node27918;
	wire [4-1:0] node27921;
	wire [4-1:0] node27924;
	wire [4-1:0] node27925;
	wire [4-1:0] node27926;
	wire [4-1:0] node27927;
	wire [4-1:0] node27930;
	wire [4-1:0] node27933;
	wire [4-1:0] node27935;
	wire [4-1:0] node27938;
	wire [4-1:0] node27939;
	wire [4-1:0] node27940;
	wire [4-1:0] node27943;
	wire [4-1:0] node27947;
	wire [4-1:0] node27948;
	wire [4-1:0] node27949;
	wire [4-1:0] node27950;
	wire [4-1:0] node27951;
	wire [4-1:0] node27952;
	wire [4-1:0] node27953;
	wire [4-1:0] node27956;
	wire [4-1:0] node27957;
	wire [4-1:0] node27960;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27966;
	wire [4-1:0] node27969;
	wire [4-1:0] node27970;
	wire [4-1:0] node27973;
	wire [4-1:0] node27976;
	wire [4-1:0] node27977;
	wire [4-1:0] node27980;
	wire [4-1:0] node27982;
	wire [4-1:0] node27983;
	wire [4-1:0] node27987;
	wire [4-1:0] node27988;
	wire [4-1:0] node27989;
	wire [4-1:0] node27990;
	wire [4-1:0] node27994;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node27999;
	wire [4-1:0] node28000;
	wire [4-1:0] node28004;
	wire [4-1:0] node28008;
	wire [4-1:0] node28009;
	wire [4-1:0] node28010;
	wire [4-1:0] node28011;
	wire [4-1:0] node28012;
	wire [4-1:0] node28013;
	wire [4-1:0] node28016;
	wire [4-1:0] node28019;
	wire [4-1:0] node28021;
	wire [4-1:0] node28024;
	wire [4-1:0] node28025;
	wire [4-1:0] node28028;
	wire [4-1:0] node28031;
	wire [4-1:0] node28032;
	wire [4-1:0] node28033;
	wire [4-1:0] node28035;
	wire [4-1:0] node28038;
	wire [4-1:0] node28039;
	wire [4-1:0] node28043;
	wire [4-1:0] node28044;
	wire [4-1:0] node28045;
	wire [4-1:0] node28048;
	wire [4-1:0] node28052;
	wire [4-1:0] node28053;
	wire [4-1:0] node28054;
	wire [4-1:0] node28055;
	wire [4-1:0] node28056;
	wire [4-1:0] node28061;
	wire [4-1:0] node28062;
	wire [4-1:0] node28065;
	wire [4-1:0] node28068;
	wire [4-1:0] node28069;
	wire [4-1:0] node28070;
	wire [4-1:0] node28073;
	wire [4-1:0] node28076;
	wire [4-1:0] node28077;
	wire [4-1:0] node28078;
	wire [4-1:0] node28082;
	wire [4-1:0] node28084;
	wire [4-1:0] node28087;
	wire [4-1:0] node28088;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28091;
	wire [4-1:0] node28092;
	wire [4-1:0] node28094;
	wire [4-1:0] node28097;
	wire [4-1:0] node28099;
	wire [4-1:0] node28103;
	wire [4-1:0] node28104;
	wire [4-1:0] node28106;
	wire [4-1:0] node28108;
	wire [4-1:0] node28111;
	wire [4-1:0] node28112;
	wire [4-1:0] node28113;
	wire [4-1:0] node28117;
	wire [4-1:0] node28120;
	wire [4-1:0] node28121;
	wire [4-1:0] node28122;
	wire [4-1:0] node28123;
	wire [4-1:0] node28125;
	wire [4-1:0] node28128;
	wire [4-1:0] node28130;
	wire [4-1:0] node28133;
	wire [4-1:0] node28135;
	wire [4-1:0] node28138;
	wire [4-1:0] node28139;
	wire [4-1:0] node28140;
	wire [4-1:0] node28144;
	wire [4-1:0] node28145;
	wire [4-1:0] node28148;
	wire [4-1:0] node28151;
	wire [4-1:0] node28152;
	wire [4-1:0] node28153;
	wire [4-1:0] node28154;
	wire [4-1:0] node28156;
	wire [4-1:0] node28159;
	wire [4-1:0] node28160;
	wire [4-1:0] node28164;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28170;
	wire [4-1:0] node28173;
	wire [4-1:0] node28174;
	wire [4-1:0] node28176;
	wire [4-1:0] node28177;
	wire [4-1:0] node28180;
	wire [4-1:0] node28183;
	wire [4-1:0] node28184;
	wire [4-1:0] node28188;
	wire [4-1:0] node28189;
	wire [4-1:0] node28190;
	wire [4-1:0] node28191;
	wire [4-1:0] node28192;
	wire [4-1:0] node28193;
	wire [4-1:0] node28194;
	wire [4-1:0] node28195;
	wire [4-1:0] node28198;
	wire [4-1:0] node28201;
	wire [4-1:0] node28203;
	wire [4-1:0] node28205;
	wire [4-1:0] node28208;
	wire [4-1:0] node28209;
	wire [4-1:0] node28210;
	wire [4-1:0] node28211;
	wire [4-1:0] node28212;
	wire [4-1:0] node28216;
	wire [4-1:0] node28217;
	wire [4-1:0] node28220;
	wire [4-1:0] node28223;
	wire [4-1:0] node28224;
	wire [4-1:0] node28228;
	wire [4-1:0] node28229;
	wire [4-1:0] node28230;
	wire [4-1:0] node28235;
	wire [4-1:0] node28236;
	wire [4-1:0] node28237;
	wire [4-1:0] node28238;
	wire [4-1:0] node28240;
	wire [4-1:0] node28241;
	wire [4-1:0] node28244;
	wire [4-1:0] node28247;
	wire [4-1:0] node28248;
	wire [4-1:0] node28251;
	wire [4-1:0] node28254;
	wire [4-1:0] node28255;
	wire [4-1:0] node28256;
	wire [4-1:0] node28258;
	wire [4-1:0] node28262;
	wire [4-1:0] node28263;
	wire [4-1:0] node28266;
	wire [4-1:0] node28267;
	wire [4-1:0] node28271;
	wire [4-1:0] node28272;
	wire [4-1:0] node28273;
	wire [4-1:0] node28275;
	wire [4-1:0] node28278;
	wire [4-1:0] node28279;
	wire [4-1:0] node28282;
	wire [4-1:0] node28283;
	wire [4-1:0] node28287;
	wire [4-1:0] node28288;
	wire [4-1:0] node28289;
	wire [4-1:0] node28291;
	wire [4-1:0] node28295;
	wire [4-1:0] node28296;
	wire [4-1:0] node28297;
	wire [4-1:0] node28300;
	wire [4-1:0] node28303;
	wire [4-1:0] node28304;
	wire [4-1:0] node28308;
	wire [4-1:0] node28309;
	wire [4-1:0] node28310;
	wire [4-1:0] node28311;
	wire [4-1:0] node28312;
	wire [4-1:0] node28315;
	wire [4-1:0] node28316;
	wire [4-1:0] node28320;
	wire [4-1:0] node28321;
	wire [4-1:0] node28324;
	wire [4-1:0] node28327;
	wire [4-1:0] node28328;
	wire [4-1:0] node28329;
	wire [4-1:0] node28331;
	wire [4-1:0] node28334;
	wire [4-1:0] node28337;
	wire [4-1:0] node28338;
	wire [4-1:0] node28339;
	wire [4-1:0] node28340;
	wire [4-1:0] node28345;
	wire [4-1:0] node28346;
	wire [4-1:0] node28350;
	wire [4-1:0] node28351;
	wire [4-1:0] node28352;
	wire [4-1:0] node28353;
	wire [4-1:0] node28354;
	wire [4-1:0] node28357;
	wire [4-1:0] node28360;
	wire [4-1:0] node28361;
	wire [4-1:0] node28364;
	wire [4-1:0] node28367;
	wire [4-1:0] node28369;
	wire [4-1:0] node28372;
	wire [4-1:0] node28373;
	wire [4-1:0] node28374;
	wire [4-1:0] node28377;
	wire [4-1:0] node28378;
	wire [4-1:0] node28382;
	wire [4-1:0] node28383;
	wire [4-1:0] node28385;
	wire [4-1:0] node28388;
	wire [4-1:0] node28390;
	wire [4-1:0] node28393;
	wire [4-1:0] node28394;
	wire [4-1:0] node28395;
	wire [4-1:0] node28396;
	wire [4-1:0] node28397;
	wire [4-1:0] node28398;
	wire [4-1:0] node28399;
	wire [4-1:0] node28402;
	wire [4-1:0] node28405;
	wire [4-1:0] node28406;
	wire [4-1:0] node28410;
	wire [4-1:0] node28411;
	wire [4-1:0] node28412;
	wire [4-1:0] node28413;
	wire [4-1:0] node28416;
	wire [4-1:0] node28421;
	wire [4-1:0] node28422;
	wire [4-1:0] node28424;
	wire [4-1:0] node28425;
	wire [4-1:0] node28429;
	wire [4-1:0] node28430;
	wire [4-1:0] node28431;
	wire [4-1:0] node28435;
	wire [4-1:0] node28436;
	wire [4-1:0] node28440;
	wire [4-1:0] node28441;
	wire [4-1:0] node28442;
	wire [4-1:0] node28443;
	wire [4-1:0] node28444;
	wire [4-1:0] node28447;
	wire [4-1:0] node28450;
	wire [4-1:0] node28451;
	wire [4-1:0] node28455;
	wire [4-1:0] node28456;
	wire [4-1:0] node28457;
	wire [4-1:0] node28458;
	wire [4-1:0] node28461;
	wire [4-1:0] node28465;
	wire [4-1:0] node28466;
	wire [4-1:0] node28467;
	wire [4-1:0] node28470;
	wire [4-1:0] node28474;
	wire [4-1:0] node28475;
	wire [4-1:0] node28476;
	wire [4-1:0] node28478;
	wire [4-1:0] node28481;
	wire [4-1:0] node28482;
	wire [4-1:0] node28486;
	wire [4-1:0] node28487;
	wire [4-1:0] node28488;
	wire [4-1:0] node28490;
	wire [4-1:0] node28493;
	wire [4-1:0] node28494;
	wire [4-1:0] node28498;
	wire [4-1:0] node28499;
	wire [4-1:0] node28500;
	wire [4-1:0] node28505;
	wire [4-1:0] node28506;
	wire [4-1:0] node28507;
	wire [4-1:0] node28508;
	wire [4-1:0] node28509;
	wire [4-1:0] node28511;
	wire [4-1:0] node28514;
	wire [4-1:0] node28517;
	wire [4-1:0] node28519;
	wire [4-1:0] node28520;
	wire [4-1:0] node28522;
	wire [4-1:0] node28525;
	wire [4-1:0] node28528;
	wire [4-1:0] node28530;
	wire [4-1:0] node28531;
	wire [4-1:0] node28532;
	wire [4-1:0] node28534;
	wire [4-1:0] node28537;
	wire [4-1:0] node28541;
	wire [4-1:0] node28542;
	wire [4-1:0] node28543;
	wire [4-1:0] node28544;
	wire [4-1:0] node28547;
	wire [4-1:0] node28550;
	wire [4-1:0] node28551;
	wire [4-1:0] node28552;
	wire [4-1:0] node28554;
	wire [4-1:0] node28557;
	wire [4-1:0] node28558;
	wire [4-1:0] node28562;
	wire [4-1:0] node28563;
	wire [4-1:0] node28566;
	wire [4-1:0] node28569;
	wire [4-1:0] node28570;
	wire [4-1:0] node28571;
	wire [4-1:0] node28574;
	wire [4-1:0] node28577;
	wire [4-1:0] node28579;
	wire [4-1:0] node28580;
	wire [4-1:0] node28583;
	wire [4-1:0] node28586;
	wire [4-1:0] node28587;
	wire [4-1:0] node28588;
	wire [4-1:0] node28589;
	wire [4-1:0] node28590;
	wire [4-1:0] node28591;
	wire [4-1:0] node28592;
	wire [4-1:0] node28595;
	wire [4-1:0] node28596;
	wire [4-1:0] node28600;
	wire [4-1:0] node28601;
	wire [4-1:0] node28602;
	wire [4-1:0] node28604;
	wire [4-1:0] node28608;
	wire [4-1:0] node28609;
	wire [4-1:0] node28610;
	wire [4-1:0] node28613;
	wire [4-1:0] node28617;
	wire [4-1:0] node28618;
	wire [4-1:0] node28619;
	wire [4-1:0] node28621;
	wire [4-1:0] node28622;
	wire [4-1:0] node28625;
	wire [4-1:0] node28629;
	wire [4-1:0] node28630;
	wire [4-1:0] node28631;
	wire [4-1:0] node28632;
	wire [4-1:0] node28635;
	wire [4-1:0] node28638;
	wire [4-1:0] node28640;
	wire [4-1:0] node28643;
	wire [4-1:0] node28644;
	wire [4-1:0] node28646;
	wire [4-1:0] node28649;
	wire [4-1:0] node28650;
	wire [4-1:0] node28653;
	wire [4-1:0] node28656;
	wire [4-1:0] node28657;
	wire [4-1:0] node28658;
	wire [4-1:0] node28659;
	wire [4-1:0] node28661;
	wire [4-1:0] node28664;
	wire [4-1:0] node28667;
	wire [4-1:0] node28668;
	wire [4-1:0] node28669;
	wire [4-1:0] node28672;
	wire [4-1:0] node28675;
	wire [4-1:0] node28676;
	wire [4-1:0] node28680;
	wire [4-1:0] node28681;
	wire [4-1:0] node28682;
	wire [4-1:0] node28683;
	wire [4-1:0] node28687;
	wire [4-1:0] node28689;
	wire [4-1:0] node28690;
	wire [4-1:0] node28693;
	wire [4-1:0] node28696;
	wire [4-1:0] node28698;
	wire [4-1:0] node28699;
	wire [4-1:0] node28700;
	wire [4-1:0] node28703;
	wire [4-1:0] node28707;
	wire [4-1:0] node28708;
	wire [4-1:0] node28709;
	wire [4-1:0] node28710;
	wire [4-1:0] node28711;
	wire [4-1:0] node28712;
	wire [4-1:0] node28716;
	wire [4-1:0] node28717;
	wire [4-1:0] node28720;
	wire [4-1:0] node28723;
	wire [4-1:0] node28724;
	wire [4-1:0] node28725;
	wire [4-1:0] node28726;
	wire [4-1:0] node28730;
	wire [4-1:0] node28732;
	wire [4-1:0] node28735;
	wire [4-1:0] node28736;
	wire [4-1:0] node28737;
	wire [4-1:0] node28742;
	wire [4-1:0] node28743;
	wire [4-1:0] node28744;
	wire [4-1:0] node28746;
	wire [4-1:0] node28748;
	wire [4-1:0] node28751;
	wire [4-1:0] node28752;
	wire [4-1:0] node28753;
	wire [4-1:0] node28756;
	wire [4-1:0] node28760;
	wire [4-1:0] node28761;
	wire [4-1:0] node28764;
	wire [4-1:0] node28767;
	wire [4-1:0] node28768;
	wire [4-1:0] node28770;
	wire [4-1:0] node28771;
	wire [4-1:0] node28772;
	wire [4-1:0] node28773;
	wire [4-1:0] node28777;
	wire [4-1:0] node28779;
	wire [4-1:0] node28783;
	wire [4-1:0] node28784;
	wire [4-1:0] node28785;
	wire [4-1:0] node28786;
	wire [4-1:0] node28789;
	wire [4-1:0] node28792;
	wire [4-1:0] node28794;
	wire [4-1:0] node28796;
	wire [4-1:0] node28799;
	wire [4-1:0] node28800;
	wire [4-1:0] node28801;
	wire [4-1:0] node28805;
	wire [4-1:0] node28807;
	wire [4-1:0] node28810;
	wire [4-1:0] node28811;
	wire [4-1:0] node28812;
	wire [4-1:0] node28813;
	wire [4-1:0] node28814;
	wire [4-1:0] node28816;
	wire [4-1:0] node28817;
	wire [4-1:0] node28821;
	wire [4-1:0] node28823;
	wire [4-1:0] node28824;
	wire [4-1:0] node28825;
	wire [4-1:0] node28829;
	wire [4-1:0] node28831;
	wire [4-1:0] node28834;
	wire [4-1:0] node28835;
	wire [4-1:0] node28837;
	wire [4-1:0] node28839;
	wire [4-1:0] node28842;
	wire [4-1:0] node28844;
	wire [4-1:0] node28846;
	wire [4-1:0] node28849;
	wire [4-1:0] node28850;
	wire [4-1:0] node28851;
	wire [4-1:0] node28852;
	wire [4-1:0] node28853;
	wire [4-1:0] node28857;
	wire [4-1:0] node28858;
	wire [4-1:0] node28861;
	wire [4-1:0] node28864;
	wire [4-1:0] node28865;
	wire [4-1:0] node28866;
	wire [4-1:0] node28867;
	wire [4-1:0] node28870;
	wire [4-1:0] node28873;
	wire [4-1:0] node28874;
	wire [4-1:0] node28877;
	wire [4-1:0] node28880;
	wire [4-1:0] node28882;
	wire [4-1:0] node28884;
	wire [4-1:0] node28887;
	wire [4-1:0] node28888;
	wire [4-1:0] node28889;
	wire [4-1:0] node28892;
	wire [4-1:0] node28895;
	wire [4-1:0] node28897;
	wire [4-1:0] node28898;
	wire [4-1:0] node28899;
	wire [4-1:0] node28902;
	wire [4-1:0] node28905;
	wire [4-1:0] node28906;
	wire [4-1:0] node28909;
	wire [4-1:0] node28912;
	wire [4-1:0] node28913;
	wire [4-1:0] node28914;
	wire [4-1:0] node28915;
	wire [4-1:0] node28916;
	wire [4-1:0] node28917;
	wire [4-1:0] node28919;
	wire [4-1:0] node28922;
	wire [4-1:0] node28925;
	wire [4-1:0] node28926;
	wire [4-1:0] node28930;
	wire [4-1:0] node28932;
	wire [4-1:0] node28934;
	wire [4-1:0] node28935;
	wire [4-1:0] node28938;
	wire [4-1:0] node28941;
	wire [4-1:0] node28942;
	wire [4-1:0] node28943;
	wire [4-1:0] node28944;
	wire [4-1:0] node28948;
	wire [4-1:0] node28949;
	wire [4-1:0] node28953;
	wire [4-1:0] node28956;
	wire [4-1:0] node28957;
	wire [4-1:0] node28958;
	wire [4-1:0] node28960;
	wire [4-1:0] node28962;
	wire [4-1:0] node28963;
	wire [4-1:0] node28966;
	wire [4-1:0] node28969;
	wire [4-1:0] node28970;
	wire [4-1:0] node28972;
	wire [4-1:0] node28975;
	wire [4-1:0] node28977;
	wire [4-1:0] node28980;
	wire [4-1:0] node28981;
	wire [4-1:0] node28982;
	wire [4-1:0] node28984;
	wire [4-1:0] node28987;
	wire [4-1:0] node28989;
	wire [4-1:0] node28992;
	wire [4-1:0] node28993;
	wire [4-1:0] node28996;
	wire [4-1:0] node28999;
	wire [4-1:0] node29000;
	wire [4-1:0] node29001;
	wire [4-1:0] node29002;
	wire [4-1:0] node29003;
	wire [4-1:0] node29004;
	wire [4-1:0] node29005;
	wire [4-1:0] node29007;
	wire [4-1:0] node29008;
	wire [4-1:0] node29009;
	wire [4-1:0] node29012;
	wire [4-1:0] node29015;
	wire [4-1:0] node29016;
	wire [4-1:0] node29017;
	wire [4-1:0] node29020;
	wire [4-1:0] node29024;
	wire [4-1:0] node29026;
	wire [4-1:0] node29027;
	wire [4-1:0] node29030;
	wire [4-1:0] node29033;
	wire [4-1:0] node29034;
	wire [4-1:0] node29036;
	wire [4-1:0] node29037;
	wire [4-1:0] node29040;
	wire [4-1:0] node29043;
	wire [4-1:0] node29045;
	wire [4-1:0] node29046;
	wire [4-1:0] node29049;
	wire [4-1:0] node29052;
	wire [4-1:0] node29053;
	wire [4-1:0] node29054;
	wire [4-1:0] node29056;
	wire [4-1:0] node29057;
	wire [4-1:0] node29059;
	wire [4-1:0] node29062;
	wire [4-1:0] node29063;
	wire [4-1:0] node29066;
	wire [4-1:0] node29069;
	wire [4-1:0] node29071;
	wire [4-1:0] node29072;
	wire [4-1:0] node29073;
	wire [4-1:0] node29075;
	wire [4-1:0] node29079;
	wire [4-1:0] node29081;
	wire [4-1:0] node29084;
	wire [4-1:0] node29085;
	wire [4-1:0] node29087;
	wire [4-1:0] node29088;
	wire [4-1:0] node29092;
	wire [4-1:0] node29094;
	wire [4-1:0] node29095;
	wire [4-1:0] node29096;
	wire [4-1:0] node29099;
	wire [4-1:0] node29102;
	wire [4-1:0] node29105;
	wire [4-1:0] node29106;
	wire [4-1:0] node29107;
	wire [4-1:0] node29108;
	wire [4-1:0] node29109;
	wire [4-1:0] node29111;
	wire [4-1:0] node29112;
	wire [4-1:0] node29116;
	wire [4-1:0] node29118;
	wire [4-1:0] node29121;
	wire [4-1:0] node29122;
	wire [4-1:0] node29123;
	wire [4-1:0] node29125;
	wire [4-1:0] node29126;
	wire [4-1:0] node29129;
	wire [4-1:0] node29132;
	wire [4-1:0] node29133;
	wire [4-1:0] node29134;
	wire [4-1:0] node29138;
	wire [4-1:0] node29139;
	wire [4-1:0] node29143;
	wire [4-1:0] node29144;
	wire [4-1:0] node29145;
	wire [4-1:0] node29149;
	wire [4-1:0] node29150;
	wire [4-1:0] node29152;
	wire [4-1:0] node29156;
	wire [4-1:0] node29157;
	wire [4-1:0] node29158;
	wire [4-1:0] node29159;
	wire [4-1:0] node29160;
	wire [4-1:0] node29164;
	wire [4-1:0] node29166;
	wire [4-1:0] node29169;
	wire [4-1:0] node29170;
	wire [4-1:0] node29172;
	wire [4-1:0] node29175;
	wire [4-1:0] node29177;
	wire [4-1:0] node29180;
	wire [4-1:0] node29181;
	wire [4-1:0] node29182;
	wire [4-1:0] node29186;
	wire [4-1:0] node29187;
	wire [4-1:0] node29189;
	wire [4-1:0] node29192;
	wire [4-1:0] node29194;
	wire [4-1:0] node29197;
	wire [4-1:0] node29198;
	wire [4-1:0] node29199;
	wire [4-1:0] node29200;
	wire [4-1:0] node29201;
	wire [4-1:0] node29202;
	wire [4-1:0] node29203;
	wire [4-1:0] node29207;
	wire [4-1:0] node29208;
	wire [4-1:0] node29212;
	wire [4-1:0] node29213;
	wire [4-1:0] node29216;
	wire [4-1:0] node29219;
	wire [4-1:0] node29220;
	wire [4-1:0] node29222;
	wire [4-1:0] node29225;
	wire [4-1:0] node29226;
	wire [4-1:0] node29227;
	wire [4-1:0] node29231;
	wire [4-1:0] node29232;
	wire [4-1:0] node29236;
	wire [4-1:0] node29237;
	wire [4-1:0] node29238;
	wire [4-1:0] node29239;
	wire [4-1:0] node29242;
	wire [4-1:0] node29245;
	wire [4-1:0] node29246;
	wire [4-1:0] node29249;
	wire [4-1:0] node29252;
	wire [4-1:0] node29254;
	wire [4-1:0] node29255;
	wire [4-1:0] node29256;
	wire [4-1:0] node29260;
	wire [4-1:0] node29262;
	wire [4-1:0] node29265;
	wire [4-1:0] node29266;
	wire [4-1:0] node29267;
	wire [4-1:0] node29268;
	wire [4-1:0] node29269;
	wire [4-1:0] node29270;
	wire [4-1:0] node29273;
	wire [4-1:0] node29276;
	wire [4-1:0] node29277;
	wire [4-1:0] node29282;
	wire [4-1:0] node29283;
	wire [4-1:0] node29286;
	wire [4-1:0] node29287;
	wire [4-1:0] node29290;
	wire [4-1:0] node29293;
	wire [4-1:0] node29294;
	wire [4-1:0] node29295;
	wire [4-1:0] node29298;
	wire [4-1:0] node29300;
	wire [4-1:0] node29303;
	wire [4-1:0] node29304;
	wire [4-1:0] node29306;
	wire [4-1:0] node29309;
	wire [4-1:0] node29310;
	wire [4-1:0] node29314;
	wire [4-1:0] node29315;
	wire [4-1:0] node29316;
	wire [4-1:0] node29317;
	wire [4-1:0] node29318;
	wire [4-1:0] node29319;
	wire [4-1:0] node29320;
	wire [4-1:0] node29322;
	wire [4-1:0] node29325;
	wire [4-1:0] node29327;
	wire [4-1:0] node29330;
	wire [4-1:0] node29331;
	wire [4-1:0] node29332;
	wire [4-1:0] node29337;
	wire [4-1:0] node29338;
	wire [4-1:0] node29339;
	wire [4-1:0] node29341;
	wire [4-1:0] node29344;
	wire [4-1:0] node29346;
	wire [4-1:0] node29349;
	wire [4-1:0] node29350;
	wire [4-1:0] node29351;
	wire [4-1:0] node29355;
	wire [4-1:0] node29357;
	wire [4-1:0] node29360;
	wire [4-1:0] node29361;
	wire [4-1:0] node29362;
	wire [4-1:0] node29363;
	wire [4-1:0] node29365;
	wire [4-1:0] node29368;
	wire [4-1:0] node29369;
	wire [4-1:0] node29373;
	wire [4-1:0] node29374;
	wire [4-1:0] node29376;
	wire [4-1:0] node29379;
	wire [4-1:0] node29381;
	wire [4-1:0] node29384;
	wire [4-1:0] node29385;
	wire [4-1:0] node29386;
	wire [4-1:0] node29388;
	wire [4-1:0] node29391;
	wire [4-1:0] node29392;
	wire [4-1:0] node29396;
	wire [4-1:0] node29397;
	wire [4-1:0] node29400;
	wire [4-1:0] node29402;
	wire [4-1:0] node29405;
	wire [4-1:0] node29406;
	wire [4-1:0] node29407;
	wire [4-1:0] node29408;
	wire [4-1:0] node29409;
	wire [4-1:0] node29410;
	wire [4-1:0] node29414;
	wire [4-1:0] node29415;
	wire [4-1:0] node29419;
	wire [4-1:0] node29420;
	wire [4-1:0] node29422;
	wire [4-1:0] node29425;
	wire [4-1:0] node29426;
	wire [4-1:0] node29430;
	wire [4-1:0] node29431;
	wire [4-1:0] node29434;
	wire [4-1:0] node29435;
	wire [4-1:0] node29437;
	wire [4-1:0] node29440;
	wire [4-1:0] node29443;
	wire [4-1:0] node29444;
	wire [4-1:0] node29445;
	wire [4-1:0] node29446;
	wire [4-1:0] node29447;
	wire [4-1:0] node29450;
	wire [4-1:0] node29453;
	wire [4-1:0] node29456;
	wire [4-1:0] node29458;
	wire [4-1:0] node29459;
	wire [4-1:0] node29462;
	wire [4-1:0] node29464;
	wire [4-1:0] node29467;
	wire [4-1:0] node29468;
	wire [4-1:0] node29469;
	wire [4-1:0] node29472;
	wire [4-1:0] node29475;
	wire [4-1:0] node29477;
	wire [4-1:0] node29480;
	wire [4-1:0] node29481;
	wire [4-1:0] node29482;
	wire [4-1:0] node29483;
	wire [4-1:0] node29484;
	wire [4-1:0] node29485;
	wire [4-1:0] node29487;
	wire [4-1:0] node29491;
	wire [4-1:0] node29493;
	wire [4-1:0] node29494;
	wire [4-1:0] node29495;
	wire [4-1:0] node29500;
	wire [4-1:0] node29501;
	wire [4-1:0] node29503;
	wire [4-1:0] node29505;
	wire [4-1:0] node29508;
	wire [4-1:0] node29510;
	wire [4-1:0] node29511;
	wire [4-1:0] node29514;
	wire [4-1:0] node29517;
	wire [4-1:0] node29518;
	wire [4-1:0] node29519;
	wire [4-1:0] node29521;
	wire [4-1:0] node29524;
	wire [4-1:0] node29525;
	wire [4-1:0] node29526;
	wire [4-1:0] node29527;
	wire [4-1:0] node29530;
	wire [4-1:0] node29534;
	wire [4-1:0] node29535;
	wire [4-1:0] node29537;
	wire [4-1:0] node29540;
	wire [4-1:0] node29541;
	wire [4-1:0] node29545;
	wire [4-1:0] node29546;
	wire [4-1:0] node29547;
	wire [4-1:0] node29549;
	wire [4-1:0] node29552;
	wire [4-1:0] node29553;
	wire [4-1:0] node29554;
	wire [4-1:0] node29557;
	wire [4-1:0] node29560;
	wire [4-1:0] node29561;
	wire [4-1:0] node29564;
	wire [4-1:0] node29567;
	wire [4-1:0] node29568;
	wire [4-1:0] node29571;
	wire [4-1:0] node29574;
	wire [4-1:0] node29575;
	wire [4-1:0] node29576;
	wire [4-1:0] node29577;
	wire [4-1:0] node29578;
	wire [4-1:0] node29579;
	wire [4-1:0] node29582;
	wire [4-1:0] node29586;
	wire [4-1:0] node29587;
	wire [4-1:0] node29588;
	wire [4-1:0] node29591;
	wire [4-1:0] node29594;
	wire [4-1:0] node29595;
	wire [4-1:0] node29597;
	wire [4-1:0] node29601;
	wire [4-1:0] node29602;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29608;
	wire [4-1:0] node29610;
	wire [4-1:0] node29611;
	wire [4-1:0] node29615;
	wire [4-1:0] node29617;
	wire [4-1:0] node29620;
	wire [4-1:0] node29621;
	wire [4-1:0] node29622;
	wire [4-1:0] node29623;
	wire [4-1:0] node29624;
	wire [4-1:0] node29625;
	wire [4-1:0] node29630;
	wire [4-1:0] node29632;
	wire [4-1:0] node29635;
	wire [4-1:0] node29636;
	wire [4-1:0] node29639;
	wire [4-1:0] node29640;
	wire [4-1:0] node29641;
	wire [4-1:0] node29645;
	wire [4-1:0] node29646;
	wire [4-1:0] node29650;
	wire [4-1:0] node29651;
	wire [4-1:0] node29652;
	wire [4-1:0] node29655;
	wire [4-1:0] node29657;
	wire [4-1:0] node29660;
	wire [4-1:0] node29661;
	wire [4-1:0] node29662;
	wire [4-1:0] node29663;
	wire [4-1:0] node29667;
	wire [4-1:0] node29668;
	wire [4-1:0] node29671;
	wire [4-1:0] node29674;
	wire [4-1:0] node29675;
	wire [4-1:0] node29676;
	wire [4-1:0] node29679;
	wire [4-1:0] node29682;
	wire [4-1:0] node29684;
	wire [4-1:0] node29687;
	wire [4-1:0] node29688;
	wire [4-1:0] node29689;
	wire [4-1:0] node29690;
	wire [4-1:0] node29691;
	wire [4-1:0] node29692;
	wire [4-1:0] node29693;
	wire [4-1:0] node29694;
	wire [4-1:0] node29695;
	wire [4-1:0] node29696;
	wire [4-1:0] node29700;
	wire [4-1:0] node29701;
	wire [4-1:0] node29705;
	wire [4-1:0] node29706;
	wire [4-1:0] node29707;
	wire [4-1:0] node29710;
	wire [4-1:0] node29713;
	wire [4-1:0] node29714;
	wire [4-1:0] node29717;
	wire [4-1:0] node29720;
	wire [4-1:0] node29721;
	wire [4-1:0] node29723;
	wire [4-1:0] node29724;
	wire [4-1:0] node29728;
	wire [4-1:0] node29729;
	wire [4-1:0] node29730;
	wire [4-1:0] node29734;
	wire [4-1:0] node29735;
	wire [4-1:0] node29739;
	wire [4-1:0] node29740;
	wire [4-1:0] node29741;
	wire [4-1:0] node29742;
	wire [4-1:0] node29746;
	wire [4-1:0] node29747;
	wire [4-1:0] node29748;
	wire [4-1:0] node29752;
	wire [4-1:0] node29755;
	wire [4-1:0] node29756;
	wire [4-1:0] node29758;
	wire [4-1:0] node29761;
	wire [4-1:0] node29762;
	wire [4-1:0] node29763;
	wire [4-1:0] node29766;
	wire [4-1:0] node29770;
	wire [4-1:0] node29771;
	wire [4-1:0] node29772;
	wire [4-1:0] node29773;
	wire [4-1:0] node29774;
	wire [4-1:0] node29778;
	wire [4-1:0] node29781;
	wire [4-1:0] node29782;
	wire [4-1:0] node29783;
	wire [4-1:0] node29786;
	wire [4-1:0] node29789;
	wire [4-1:0] node29792;
	wire [4-1:0] node29793;
	wire [4-1:0] node29794;
	wire [4-1:0] node29795;
	wire [4-1:0] node29799;
	wire [4-1:0] node29802;
	wire [4-1:0] node29803;
	wire [4-1:0] node29804;
	wire [4-1:0] node29809;
	wire [4-1:0] node29810;
	wire [4-1:0] node29811;
	wire [4-1:0] node29812;
	wire [4-1:0] node29813;
	wire [4-1:0] node29814;
	wire [4-1:0] node29815;
	wire [4-1:0] node29818;
	wire [4-1:0] node29821;
	wire [4-1:0] node29823;
	wire [4-1:0] node29826;
	wire [4-1:0] node29828;
	wire [4-1:0] node29831;
	wire [4-1:0] node29833;
	wire [4-1:0] node29834;
	wire [4-1:0] node29836;
	wire [4-1:0] node29839;
	wire [4-1:0] node29842;
	wire [4-1:0] node29843;
	wire [4-1:0] node29845;
	wire [4-1:0] node29846;
	wire [4-1:0] node29848;
	wire [4-1:0] node29851;
	wire [4-1:0] node29853;
	wire [4-1:0] node29856;
	wire [4-1:0] node29857;
	wire [4-1:0] node29858;
	wire [4-1:0] node29859;
	wire [4-1:0] node29864;
	wire [4-1:0] node29865;
	wire [4-1:0] node29866;
	wire [4-1:0] node29870;
	wire [4-1:0] node29872;
	wire [4-1:0] node29875;
	wire [4-1:0] node29876;
	wire [4-1:0] node29877;
	wire [4-1:0] node29879;
	wire [4-1:0] node29880;
	wire [4-1:0] node29884;
	wire [4-1:0] node29885;
	wire [4-1:0] node29886;
	wire [4-1:0] node29890;
	wire [4-1:0] node29891;
	wire [4-1:0] node29895;
	wire [4-1:0] node29896;
	wire [4-1:0] node29897;
	wire [4-1:0] node29898;
	wire [4-1:0] node29902;
	wire [4-1:0] node29904;
	wire [4-1:0] node29905;
	wire [4-1:0] node29908;
	wire [4-1:0] node29911;
	wire [4-1:0] node29912;
	wire [4-1:0] node29913;
	wire [4-1:0] node29914;
	wire [4-1:0] node29918;
	wire [4-1:0] node29920;
	wire [4-1:0] node29924;
	wire [4-1:0] node29925;
	wire [4-1:0] node29926;
	wire [4-1:0] node29927;
	wire [4-1:0] node29928;
	wire [4-1:0] node29929;
	wire [4-1:0] node29930;
	wire [4-1:0] node29934;
	wire [4-1:0] node29937;
	wire [4-1:0] node29938;
	wire [4-1:0] node29939;
	wire [4-1:0] node29942;
	wire [4-1:0] node29945;
	wire [4-1:0] node29946;
	wire [4-1:0] node29950;
	wire [4-1:0] node29951;
	wire [4-1:0] node29952;
	wire [4-1:0] node29955;
	wire [4-1:0] node29956;
	wire [4-1:0] node29959;
	wire [4-1:0] node29960;
	wire [4-1:0] node29964;
	wire [4-1:0] node29965;
	wire [4-1:0] node29966;
	wire [4-1:0] node29969;
	wire [4-1:0] node29972;
	wire [4-1:0] node29975;
	wire [4-1:0] node29976;
	wire [4-1:0] node29977;
	wire [4-1:0] node29978;
	wire [4-1:0] node29981;
	wire [4-1:0] node29984;
	wire [4-1:0] node29985;
	wire [4-1:0] node29988;
	wire [4-1:0] node29989;
	wire [4-1:0] node29992;
	wire [4-1:0] node29995;
	wire [4-1:0] node29996;
	wire [4-1:0] node29997;
	wire [4-1:0] node30000;
	wire [4-1:0] node30003;
	wire [4-1:0] node30004;
	wire [4-1:0] node30007;
	wire [4-1:0] node30008;
	wire [4-1:0] node30012;
	wire [4-1:0] node30013;
	wire [4-1:0] node30014;
	wire [4-1:0] node30015;
	wire [4-1:0] node30016;
	wire [4-1:0] node30018;
	wire [4-1:0] node30021;
	wire [4-1:0] node30023;
	wire [4-1:0] node30026;
	wire [4-1:0] node30027;
	wire [4-1:0] node30028;
	wire [4-1:0] node30031;
	wire [4-1:0] node30034;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30040;
	wire [4-1:0] node30042;
	wire [4-1:0] node30045;
	wire [4-1:0] node30046;
	wire [4-1:0] node30047;
	wire [4-1:0] node30050;
	wire [4-1:0] node30053;
	wire [4-1:0] node30054;
	wire [4-1:0] node30058;
	wire [4-1:0] node30059;
	wire [4-1:0] node30060;
	wire [4-1:0] node30062;
	wire [4-1:0] node30063;
	wire [4-1:0] node30064;
	wire [4-1:0] node30067;
	wire [4-1:0] node30070;
	wire [4-1:0] node30071;
	wire [4-1:0] node30074;
	wire [4-1:0] node30077;
	wire [4-1:0] node30078;
	wire [4-1:0] node30079;
	wire [4-1:0] node30080;
	wire [4-1:0] node30083;
	wire [4-1:0] node30087;
	wire [4-1:0] node30088;
	wire [4-1:0] node30092;
	wire [4-1:0] node30093;
	wire [4-1:0] node30094;
	wire [4-1:0] node30096;
	wire [4-1:0] node30099;
	wire [4-1:0] node30101;
	wire [4-1:0] node30103;
	wire [4-1:0] node30106;
	wire [4-1:0] node30107;
	wire [4-1:0] node30110;
	wire [4-1:0] node30113;
	wire [4-1:0] node30114;
	wire [4-1:0] node30115;
	wire [4-1:0] node30116;
	wire [4-1:0] node30117;
	wire [4-1:0] node30118;
	wire [4-1:0] node30120;
	wire [4-1:0] node30121;
	wire [4-1:0] node30125;
	wire [4-1:0] node30126;
	wire [4-1:0] node30128;
	wire [4-1:0] node30129;
	wire [4-1:0] node30134;
	wire [4-1:0] node30135;
	wire [4-1:0] node30136;
	wire [4-1:0] node30138;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30146;
	wire [4-1:0] node30148;
	wire [4-1:0] node30151;
	wire [4-1:0] node30152;
	wire [4-1:0] node30153;
	wire [4-1:0] node30154;
	wire [4-1:0] node30155;
	wire [4-1:0] node30159;
	wire [4-1:0] node30162;
	wire [4-1:0] node30163;
	wire [4-1:0] node30165;
	wire [4-1:0] node30166;
	wire [4-1:0] node30169;
	wire [4-1:0] node30173;
	wire [4-1:0] node30174;
	wire [4-1:0] node30175;
	wire [4-1:0] node30177;
	wire [4-1:0] node30180;
	wire [4-1:0] node30182;
	wire [4-1:0] node30185;
	wire [4-1:0] node30186;
	wire [4-1:0] node30188;
	wire [4-1:0] node30192;
	wire [4-1:0] node30193;
	wire [4-1:0] node30194;
	wire [4-1:0] node30195;
	wire [4-1:0] node30196;
	wire [4-1:0] node30197;
	wire [4-1:0] node30199;
	wire [4-1:0] node30202;
	wire [4-1:0] node30204;
	wire [4-1:0] node30207;
	wire [4-1:0] node30208;
	wire [4-1:0] node30212;
	wire [4-1:0] node30213;
	wire [4-1:0] node30214;
	wire [4-1:0] node30216;
	wire [4-1:0] node30219;
	wire [4-1:0] node30221;
	wire [4-1:0] node30224;
	wire [4-1:0] node30227;
	wire [4-1:0] node30228;
	wire [4-1:0] node30229;
	wire [4-1:0] node30232;
	wire [4-1:0] node30235;
	wire [4-1:0] node30236;
	wire [4-1:0] node30237;
	wire [4-1:0] node30239;
	wire [4-1:0] node30242;
	wire [4-1:0] node30243;
	wire [4-1:0] node30246;
	wire [4-1:0] node30249;
	wire [4-1:0] node30250;
	wire [4-1:0] node30252;
	wire [4-1:0] node30256;
	wire [4-1:0] node30257;
	wire [4-1:0] node30258;
	wire [4-1:0] node30259;
	wire [4-1:0] node30260;
	wire [4-1:0] node30264;
	wire [4-1:0] node30267;
	wire [4-1:0] node30268;
	wire [4-1:0] node30270;
	wire [4-1:0] node30273;
	wire [4-1:0] node30274;
	wire [4-1:0] node30277;
	wire [4-1:0] node30278;
	wire [4-1:0] node30282;
	wire [4-1:0] node30283;
	wire [4-1:0] node30284;
	wire [4-1:0] node30285;
	wire [4-1:0] node30289;
	wire [4-1:0] node30290;
	wire [4-1:0] node30293;
	wire [4-1:0] node30295;
	wire [4-1:0] node30298;
	wire [4-1:0] node30300;
	wire [4-1:0] node30301;
	wire [4-1:0] node30304;
	wire [4-1:0] node30305;
	wire [4-1:0] node30309;
	wire [4-1:0] node30310;
	wire [4-1:0] node30311;
	wire [4-1:0] node30312;
	wire [4-1:0] node30313;
	wire [4-1:0] node30314;
	wire [4-1:0] node30315;
	wire [4-1:0] node30318;
	wire [4-1:0] node30321;
	wire [4-1:0] node30322;
	wire [4-1:0] node30326;
	wire [4-1:0] node30327;
	wire [4-1:0] node30328;
	wire [4-1:0] node30329;
	wire [4-1:0] node30333;
	wire [4-1:0] node30336;
	wire [4-1:0] node30337;
	wire [4-1:0] node30338;
	wire [4-1:0] node30341;
	wire [4-1:0] node30344;
	wire [4-1:0] node30345;
	wire [4-1:0] node30348;
	wire [4-1:0] node30351;
	wire [4-1:0] node30352;
	wire [4-1:0] node30353;
	wire [4-1:0] node30356;
	wire [4-1:0] node30359;
	wire [4-1:0] node30361;
	wire [4-1:0] node30362;
	wire [4-1:0] node30363;
	wire [4-1:0] node30366;
	wire [4-1:0] node30370;
	wire [4-1:0] node30371;
	wire [4-1:0] node30372;
	wire [4-1:0] node30373;
	wire [4-1:0] node30374;
	wire [4-1:0] node30377;
	wire [4-1:0] node30381;
	wire [4-1:0] node30382;
	wire [4-1:0] node30383;
	wire [4-1:0] node30384;
	wire [4-1:0] node30387;
	wire [4-1:0] node30390;
	wire [4-1:0] node30391;
	wire [4-1:0] node30394;
	wire [4-1:0] node30398;
	wire [4-1:0] node30399;
	wire [4-1:0] node30400;
	wire [4-1:0] node30401;
	wire [4-1:0] node30404;
	wire [4-1:0] node30408;
	wire [4-1:0] node30409;
	wire [4-1:0] node30410;
	wire [4-1:0] node30413;
	wire [4-1:0] node30417;
	wire [4-1:0] node30418;
	wire [4-1:0] node30419;
	wire [4-1:0] node30421;
	wire [4-1:0] node30422;
	wire [4-1:0] node30424;
	wire [4-1:0] node30427;
	wire [4-1:0] node30428;
	wire [4-1:0] node30430;
	wire [4-1:0] node30433;
	wire [4-1:0] node30434;
	wire [4-1:0] node30437;
	wire [4-1:0] node30440;
	wire [4-1:0] node30441;
	wire [4-1:0] node30442;
	wire [4-1:0] node30443;
	wire [4-1:0] node30444;
	wire [4-1:0] node30448;
	wire [4-1:0] node30450;
	wire [4-1:0] node30453;
	wire [4-1:0] node30454;
	wire [4-1:0] node30455;
	wire [4-1:0] node30459;
	wire [4-1:0] node30460;
	wire [4-1:0] node30463;
	wire [4-1:0] node30466;
	wire [4-1:0] node30467;
	wire [4-1:0] node30469;
	wire [4-1:0] node30472;
	wire [4-1:0] node30473;
	wire [4-1:0] node30477;
	wire [4-1:0] node30478;
	wire [4-1:0] node30479;
	wire [4-1:0] node30480;
	wire [4-1:0] node30484;
	wire [4-1:0] node30485;
	wire [4-1:0] node30489;
	wire [4-1:0] node30490;
	wire [4-1:0] node30491;
	wire [4-1:0] node30495;
	wire [4-1:0] node30496;
	wire [4-1:0] node30500;
	wire [4-1:0] node30501;
	wire [4-1:0] node30502;
	wire [4-1:0] node30503;
	wire [4-1:0] node30504;
	wire [4-1:0] node30505;
	wire [4-1:0] node30506;
	wire [4-1:0] node30507;
	wire [4-1:0] node30508;
	wire [4-1:0] node30509;
	wire [4-1:0] node30512;
	wire [4-1:0] node30515;
	wire [4-1:0] node30516;
	wire [4-1:0] node30518;
	wire [4-1:0] node30521;
	wire [4-1:0] node30522;
	wire [4-1:0] node30525;
	wire [4-1:0] node30528;
	wire [4-1:0] node30529;
	wire [4-1:0] node30531;
	wire [4-1:0] node30532;
	wire [4-1:0] node30535;
	wire [4-1:0] node30538;
	wire [4-1:0] node30539;
	wire [4-1:0] node30540;
	wire [4-1:0] node30543;
	wire [4-1:0] node30546;
	wire [4-1:0] node30547;
	wire [4-1:0] node30550;
	wire [4-1:0] node30553;
	wire [4-1:0] node30554;
	wire [4-1:0] node30555;
	wire [4-1:0] node30556;
	wire [4-1:0] node30557;
	wire [4-1:0] node30559;
	wire [4-1:0] node30562;
	wire [4-1:0] node30564;
	wire [4-1:0] node30568;
	wire [4-1:0] node30569;
	wire [4-1:0] node30570;
	wire [4-1:0] node30573;
	wire [4-1:0] node30576;
	wire [4-1:0] node30577;
	wire [4-1:0] node30581;
	wire [4-1:0] node30582;
	wire [4-1:0] node30583;
	wire [4-1:0] node30584;
	wire [4-1:0] node30588;
	wire [4-1:0] node30590;
	wire [4-1:0] node30593;
	wire [4-1:0] node30594;
	wire [4-1:0] node30596;
	wire [4-1:0] node30599;
	wire [4-1:0] node30601;
	wire [4-1:0] node30602;
	wire [4-1:0] node30606;
	wire [4-1:0] node30607;
	wire [4-1:0] node30608;
	wire [4-1:0] node30609;
	wire [4-1:0] node30611;
	wire [4-1:0] node30612;
	wire [4-1:0] node30615;
	wire [4-1:0] node30618;
	wire [4-1:0] node30620;
	wire [4-1:0] node30621;
	wire [4-1:0] node30624;
	wire [4-1:0] node30627;
	wire [4-1:0] node30628;
	wire [4-1:0] node30630;
	wire [4-1:0] node30631;
	wire [4-1:0] node30634;
	wire [4-1:0] node30637;
	wire [4-1:0] node30639;
	wire [4-1:0] node30641;
	wire [4-1:0] node30644;
	wire [4-1:0] node30645;
	wire [4-1:0] node30646;
	wire [4-1:0] node30648;
	wire [4-1:0] node30649;
	wire [4-1:0] node30651;
	wire [4-1:0] node30655;
	wire [4-1:0] node30657;
	wire [4-1:0] node30658;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30665;
	wire [4-1:0] node30668;
	wire [4-1:0] node30670;
	wire [4-1:0] node30671;
	wire [4-1:0] node30674;
	wire [4-1:0] node30677;
	wire [4-1:0] node30678;
	wire [4-1:0] node30679;
	wire [4-1:0] node30680;
	wire [4-1:0] node30681;
	wire [4-1:0] node30682;
	wire [4-1:0] node30683;
	wire [4-1:0] node30686;
	wire [4-1:0] node30688;
	wire [4-1:0] node30692;
	wire [4-1:0] node30693;
	wire [4-1:0] node30694;
	wire [4-1:0] node30698;
	wire [4-1:0] node30699;
	wire [4-1:0] node30703;
	wire [4-1:0] node30704;
	wire [4-1:0] node30705;
	wire [4-1:0] node30707;
	wire [4-1:0] node30710;
	wire [4-1:0] node30712;
	wire [4-1:0] node30715;
	wire [4-1:0] node30716;
	wire [4-1:0] node30717;
	wire [4-1:0] node30722;
	wire [4-1:0] node30723;
	wire [4-1:0] node30724;
	wire [4-1:0] node30725;
	wire [4-1:0] node30726;
	wire [4-1:0] node30730;
	wire [4-1:0] node30733;
	wire [4-1:0] node30734;
	wire [4-1:0] node30736;
	wire [4-1:0] node30739;
	wire [4-1:0] node30741;
	wire [4-1:0] node30744;
	wire [4-1:0] node30745;
	wire [4-1:0] node30746;
	wire [4-1:0] node30747;
	wire [4-1:0] node30749;
	wire [4-1:0] node30752;
	wire [4-1:0] node30754;
	wire [4-1:0] node30758;
	wire [4-1:0] node30759;
	wire [4-1:0] node30760;
	wire [4-1:0] node30764;
	wire [4-1:0] node30766;
	wire [4-1:0] node30769;
	wire [4-1:0] node30770;
	wire [4-1:0] node30771;
	wire [4-1:0] node30772;
	wire [4-1:0] node30773;
	wire [4-1:0] node30774;
	wire [4-1:0] node30777;
	wire [4-1:0] node30781;
	wire [4-1:0] node30782;
	wire [4-1:0] node30783;
	wire [4-1:0] node30786;
	wire [4-1:0] node30787;
	wire [4-1:0] node30791;
	wire [4-1:0] node30792;
	wire [4-1:0] node30793;
	wire [4-1:0] node30797;
	wire [4-1:0] node30800;
	wire [4-1:0] node30801;
	wire [4-1:0] node30802;
	wire [4-1:0] node30805;
	wire [4-1:0] node30808;
	wire [4-1:0] node30809;
	wire [4-1:0] node30810;
	wire [4-1:0] node30813;
	wire [4-1:0] node30816;
	wire [4-1:0] node30817;
	wire [4-1:0] node30820;
	wire [4-1:0] node30823;
	wire [4-1:0] node30824;
	wire [4-1:0] node30825;
	wire [4-1:0] node30826;
	wire [4-1:0] node30827;
	wire [4-1:0] node30830;
	wire [4-1:0] node30833;
	wire [4-1:0] node30835;
	wire [4-1:0] node30836;
	wire [4-1:0] node30839;
	wire [4-1:0] node30842;
	wire [4-1:0] node30843;
	wire [4-1:0] node30844;
	wire [4-1:0] node30847;
	wire [4-1:0] node30851;
	wire [4-1:0] node30852;
	wire [4-1:0] node30853;
	wire [4-1:0] node30855;
	wire [4-1:0] node30856;
	wire [4-1:0] node30859;
	wire [4-1:0] node30862;
	wire [4-1:0] node30863;
	wire [4-1:0] node30864;
	wire [4-1:0] node30867;
	wire [4-1:0] node30871;
	wire [4-1:0] node30872;
	wire [4-1:0] node30874;
	wire [4-1:0] node30875;
	wire [4-1:0] node30878;
	wire [4-1:0] node30881;
	wire [4-1:0] node30882;
	wire [4-1:0] node30883;
	wire [4-1:0] node30886;
	wire [4-1:0] node30889;
	wire [4-1:0] node30890;
	wire [4-1:0] node30893;
	wire [4-1:0] node30896;
	wire [4-1:0] node30897;
	wire [4-1:0] node30898;
	wire [4-1:0] node30899;
	wire [4-1:0] node30900;
	wire [4-1:0] node30901;
	wire [4-1:0] node30902;
	wire [4-1:0] node30904;
	wire [4-1:0] node30907;
	wire [4-1:0] node30908;
	wire [4-1:0] node30910;
	wire [4-1:0] node30913;
	wire [4-1:0] node30916;
	wire [4-1:0] node30917;
	wire [4-1:0] node30918;
	wire [4-1:0] node30922;
	wire [4-1:0] node30924;
	wire [4-1:0] node30925;
	wire [4-1:0] node30928;
	wire [4-1:0] node30931;
	wire [4-1:0] node30932;
	wire [4-1:0] node30933;
	wire [4-1:0] node30935;
	wire [4-1:0] node30938;
	wire [4-1:0] node30941;
	wire [4-1:0] node30942;
	wire [4-1:0] node30944;
	wire [4-1:0] node30945;
	wire [4-1:0] node30949;
	wire [4-1:0] node30951;
	wire [4-1:0] node30952;
	wire [4-1:0] node30956;
	wire [4-1:0] node30957;
	wire [4-1:0] node30958;
	wire [4-1:0] node30959;
	wire [4-1:0] node30961;
	wire [4-1:0] node30964;
	wire [4-1:0] node30966;
	wire [4-1:0] node30969;
	wire [4-1:0] node30970;
	wire [4-1:0] node30971;
	wire [4-1:0] node30975;
	wire [4-1:0] node30976;
	wire [4-1:0] node30980;
	wire [4-1:0] node30981;
	wire [4-1:0] node30983;
	wire [4-1:0] node30986;
	wire [4-1:0] node30987;
	wire [4-1:0] node30988;
	wire [4-1:0] node30991;
	wire [4-1:0] node30994;
	wire [4-1:0] node30997;
	wire [4-1:0] node30998;
	wire [4-1:0] node30999;
	wire [4-1:0] node31000;
	wire [4-1:0] node31001;
	wire [4-1:0] node31002;
	wire [4-1:0] node31006;
	wire [4-1:0] node31007;
	wire [4-1:0] node31011;
	wire [4-1:0] node31012;
	wire [4-1:0] node31015;
	wire [4-1:0] node31016;
	wire [4-1:0] node31020;
	wire [4-1:0] node31021;
	wire [4-1:0] node31022;
	wire [4-1:0] node31024;
	wire [4-1:0] node31027;
	wire [4-1:0] node31029;
	wire [4-1:0] node31032;
	wire [4-1:0] node31034;
	wire [4-1:0] node31037;
	wire [4-1:0] node31038;
	wire [4-1:0] node31039;
	wire [4-1:0] node31040;
	wire [4-1:0] node31041;
	wire [4-1:0] node31042;
	wire [4-1:0] node31045;
	wire [4-1:0] node31048;
	wire [4-1:0] node31050;
	wire [4-1:0] node31054;
	wire [4-1:0] node31055;
	wire [4-1:0] node31056;
	wire [4-1:0] node31060;
	wire [4-1:0] node31061;
	wire [4-1:0] node31064;
	wire [4-1:0] node31067;
	wire [4-1:0] node31068;
	wire [4-1:0] node31069;
	wire [4-1:0] node31070;
	wire [4-1:0] node31073;
	wire [4-1:0] node31077;
	wire [4-1:0] node31078;
	wire [4-1:0] node31081;
	wire [4-1:0] node31084;
	wire [4-1:0] node31085;
	wire [4-1:0] node31086;
	wire [4-1:0] node31087;
	wire [4-1:0] node31088;
	wire [4-1:0] node31089;
	wire [4-1:0] node31092;
	wire [4-1:0] node31095;
	wire [4-1:0] node31097;
	wire [4-1:0] node31099;
	wire [4-1:0] node31100;
	wire [4-1:0] node31104;
	wire [4-1:0] node31105;
	wire [4-1:0] node31106;
	wire [4-1:0] node31107;
	wire [4-1:0] node31108;
	wire [4-1:0] node31112;
	wire [4-1:0] node31113;
	wire [4-1:0] node31116;
	wire [4-1:0] node31119;
	wire [4-1:0] node31120;
	wire [4-1:0] node31121;
	wire [4-1:0] node31124;
	wire [4-1:0] node31127;
	wire [4-1:0] node31129;
	wire [4-1:0] node31132;
	wire [4-1:0] node31133;
	wire [4-1:0] node31134;
	wire [4-1:0] node31138;
	wire [4-1:0] node31139;
	wire [4-1:0] node31140;
	wire [4-1:0] node31143;
	wire [4-1:0] node31147;
	wire [4-1:0] node31148;
	wire [4-1:0] node31149;
	wire [4-1:0] node31150;
	wire [4-1:0] node31152;
	wire [4-1:0] node31155;
	wire [4-1:0] node31156;
	wire [4-1:0] node31160;
	wire [4-1:0] node31161;
	wire [4-1:0] node31163;
	wire [4-1:0] node31166;
	wire [4-1:0] node31167;
	wire [4-1:0] node31171;
	wire [4-1:0] node31172;
	wire [4-1:0] node31174;
	wire [4-1:0] node31177;
	wire [4-1:0] node31179;
	wire [4-1:0] node31180;
	wire [4-1:0] node31182;
	wire [4-1:0] node31185;
	wire [4-1:0] node31187;
	wire [4-1:0] node31190;
	wire [4-1:0] node31191;
	wire [4-1:0] node31192;
	wire [4-1:0] node31193;
	wire [4-1:0] node31194;
	wire [4-1:0] node31197;
	wire [4-1:0] node31199;
	wire [4-1:0] node31202;
	wire [4-1:0] node31203;
	wire [4-1:0] node31205;
	wire [4-1:0] node31208;
	wire [4-1:0] node31210;
	wire [4-1:0] node31213;
	wire [4-1:0] node31214;
	wire [4-1:0] node31215;
	wire [4-1:0] node31218;
	wire [4-1:0] node31219;
	wire [4-1:0] node31223;
	wire [4-1:0] node31224;
	wire [4-1:0] node31226;
	wire [4-1:0] node31229;
	wire [4-1:0] node31231;
	wire [4-1:0] node31234;
	wire [4-1:0] node31235;
	wire [4-1:0] node31236;
	wire [4-1:0] node31237;
	wire [4-1:0] node31238;
	wire [4-1:0] node31243;
	wire [4-1:0] node31244;
	wire [4-1:0] node31245;
	wire [4-1:0] node31248;
	wire [4-1:0] node31252;
	wire [4-1:0] node31253;
	wire [4-1:0] node31254;
	wire [4-1:0] node31255;
	wire [4-1:0] node31260;
	wire [4-1:0] node31261;
	wire [4-1:0] node31262;
	wire [4-1:0] node31265;
	wire [4-1:0] node31269;
	wire [4-1:0] node31270;
	wire [4-1:0] node31271;
	wire [4-1:0] node31272;
	wire [4-1:0] node31273;
	wire [4-1:0] node31274;
	wire [4-1:0] node31275;
	wire [4-1:0] node31276;
	wire [4-1:0] node31278;
	wire [4-1:0] node31281;
	wire [4-1:0] node31282;
	wire [4-1:0] node31286;
	wire [4-1:0] node31287;
	wire [4-1:0] node31289;
	wire [4-1:0] node31292;
	wire [4-1:0] node31294;
	wire [4-1:0] node31297;
	wire [4-1:0] node31298;
	wire [4-1:0] node31299;
	wire [4-1:0] node31301;
	wire [4-1:0] node31303;
	wire [4-1:0] node31306;
	wire [4-1:0] node31307;
	wire [4-1:0] node31309;
	wire [4-1:0] node31312;
	wire [4-1:0] node31315;
	wire [4-1:0] node31316;
	wire [4-1:0] node31317;
	wire [4-1:0] node31321;
	wire [4-1:0] node31323;
	wire [4-1:0] node31325;
	wire [4-1:0] node31328;
	wire [4-1:0] node31329;
	wire [4-1:0] node31330;
	wire [4-1:0] node31331;
	wire [4-1:0] node31332;
	wire [4-1:0] node31335;
	wire [4-1:0] node31338;
	wire [4-1:0] node31339;
	wire [4-1:0] node31342;
	wire [4-1:0] node31345;
	wire [4-1:0] node31346;
	wire [4-1:0] node31347;
	wire [4-1:0] node31350;
	wire [4-1:0] node31354;
	wire [4-1:0] node31355;
	wire [4-1:0] node31356;
	wire [4-1:0] node31358;
	wire [4-1:0] node31361;
	wire [4-1:0] node31362;
	wire [4-1:0] node31364;
	wire [4-1:0] node31367;
	wire [4-1:0] node31370;
	wire [4-1:0] node31372;
	wire [4-1:0] node31375;
	wire [4-1:0] node31376;
	wire [4-1:0] node31377;
	wire [4-1:0] node31378;
	wire [4-1:0] node31379;
	wire [4-1:0] node31381;
	wire [4-1:0] node31384;
	wire [4-1:0] node31386;
	wire [4-1:0] node31389;
	wire [4-1:0] node31390;
	wire [4-1:0] node31394;
	wire [4-1:0] node31395;
	wire [4-1:0] node31396;
	wire [4-1:0] node31398;
	wire [4-1:0] node31399;
	wire [4-1:0] node31402;
	wire [4-1:0] node31405;
	wire [4-1:0] node31406;
	wire [4-1:0] node31407;
	wire [4-1:0] node31412;
	wire [4-1:0] node31413;
	wire [4-1:0] node31414;
	wire [4-1:0] node31417;
	wire [4-1:0] node31418;
	wire [4-1:0] node31422;
	wire [4-1:0] node31425;
	wire [4-1:0] node31426;
	wire [4-1:0] node31427;
	wire [4-1:0] node31429;
	wire [4-1:0] node31432;
	wire [4-1:0] node31434;
	wire [4-1:0] node31435;
	wire [4-1:0] node31439;
	wire [4-1:0] node31440;
	wire [4-1:0] node31441;
	wire [4-1:0] node31442;
	wire [4-1:0] node31446;
	wire [4-1:0] node31447;
	wire [4-1:0] node31448;
	wire [4-1:0] node31451;
	wire [4-1:0] node31455;
	wire [4-1:0] node31456;
	wire [4-1:0] node31459;
	wire [4-1:0] node31462;
	wire [4-1:0] node31463;
	wire [4-1:0] node31464;
	wire [4-1:0] node31465;
	wire [4-1:0] node31466;
	wire [4-1:0] node31467;
	wire [4-1:0] node31469;
	wire [4-1:0] node31472;
	wire [4-1:0] node31473;
	wire [4-1:0] node31477;
	wire [4-1:0] node31478;
	wire [4-1:0] node31480;
	wire [4-1:0] node31484;
	wire [4-1:0] node31485;
	wire [4-1:0] node31486;
	wire [4-1:0] node31487;
	wire [4-1:0] node31491;
	wire [4-1:0] node31492;
	wire [4-1:0] node31496;
	wire [4-1:0] node31497;
	wire [4-1:0] node31499;
	wire [4-1:0] node31502;
	wire [4-1:0] node31504;
	wire [4-1:0] node31507;
	wire [4-1:0] node31508;
	wire [4-1:0] node31509;
	wire [4-1:0] node31510;
	wire [4-1:0] node31512;
	wire [4-1:0] node31515;
	wire [4-1:0] node31516;
	wire [4-1:0] node31518;
	wire [4-1:0] node31521;
	wire [4-1:0] node31522;
	wire [4-1:0] node31526;
	wire [4-1:0] node31527;
	wire [4-1:0] node31528;
	wire [4-1:0] node31531;
	wire [4-1:0] node31535;
	wire [4-1:0] node31536;
	wire [4-1:0] node31537;
	wire [4-1:0] node31540;
	wire [4-1:0] node31542;
	wire [4-1:0] node31545;
	wire [4-1:0] node31546;
	wire [4-1:0] node31549;
	wire [4-1:0] node31551;
	wire [4-1:0] node31554;
	wire [4-1:0] node31555;
	wire [4-1:0] node31556;
	wire [4-1:0] node31557;
	wire [4-1:0] node31558;
	wire [4-1:0] node31559;
	wire [4-1:0] node31560;
	wire [4-1:0] node31564;
	wire [4-1:0] node31565;
	wire [4-1:0] node31568;
	wire [4-1:0] node31571;
	wire [4-1:0] node31572;
	wire [4-1:0] node31576;
	wire [4-1:0] node31577;
	wire [4-1:0] node31579;
	wire [4-1:0] node31582;
	wire [4-1:0] node31583;
	wire [4-1:0] node31586;
	wire [4-1:0] node31587;
	wire [4-1:0] node31591;
	wire [4-1:0] node31592;
	wire [4-1:0] node31593;
	wire [4-1:0] node31594;
	wire [4-1:0] node31596;
	wire [4-1:0] node31599;
	wire [4-1:0] node31601;
	wire [4-1:0] node31604;
	wire [4-1:0] node31605;
	wire [4-1:0] node31606;
	wire [4-1:0] node31609;
	wire [4-1:0] node31612;
	wire [4-1:0] node31615;
	wire [4-1:0] node31616;
	wire [4-1:0] node31617;
	wire [4-1:0] node31618;
	wire [4-1:0] node31622;
	wire [4-1:0] node31623;
	wire [4-1:0] node31627;
	wire [4-1:0] node31628;
	wire [4-1:0] node31631;
	wire [4-1:0] node31634;
	wire [4-1:0] node31635;
	wire [4-1:0] node31636;
	wire [4-1:0] node31637;
	wire [4-1:0] node31638;
	wire [4-1:0] node31640;
	wire [4-1:0] node31643;
	wire [4-1:0] node31644;
	wire [4-1:0] node31648;
	wire [4-1:0] node31649;
	wire [4-1:0] node31650;
	wire [4-1:0] node31653;
	wire [4-1:0] node31656;
	wire [4-1:0] node31657;
	wire [4-1:0] node31660;
	wire [4-1:0] node31663;
	wire [4-1:0] node31665;
	wire [4-1:0] node31666;
	wire [4-1:0] node31667;
	wire [4-1:0] node31670;
	wire [4-1:0] node31673;
	wire [4-1:0] node31675;
	wire [4-1:0] node31678;
	wire [4-1:0] node31679;
	wire [4-1:0] node31680;
	wire [4-1:0] node31681;
	wire [4-1:0] node31684;
	wire [4-1:0] node31687;
	wire [4-1:0] node31690;
	wire [4-1:0] node31691;
	wire [4-1:0] node31693;
	wire [4-1:0] node31696;
	wire [4-1:0] node31697;
	wire [4-1:0] node31698;
	wire [4-1:0] node31701;
	wire [4-1:0] node31705;
	wire [4-1:0] node31706;
	wire [4-1:0] node31707;
	wire [4-1:0] node31708;
	wire [4-1:0] node31709;
	wire [4-1:0] node31710;
	wire [4-1:0] node31711;
	wire [4-1:0] node31712;
	wire [4-1:0] node31713;
	wire [4-1:0] node31716;
	wire [4-1:0] node31721;
	wire [4-1:0] node31722;
	wire [4-1:0] node31723;
	wire [4-1:0] node31724;
	wire [4-1:0] node31727;
	wire [4-1:0] node31730;
	wire [4-1:0] node31731;
	wire [4-1:0] node31734;
	wire [4-1:0] node31738;
	wire [4-1:0] node31739;
	wire [4-1:0] node31740;
	wire [4-1:0] node31741;
	wire [4-1:0] node31744;
	wire [4-1:0] node31748;
	wire [4-1:0] node31749;
	wire [4-1:0] node31751;
	wire [4-1:0] node31755;
	wire [4-1:0] node31756;
	wire [4-1:0] node31757;
	wire [4-1:0] node31758;
	wire [4-1:0] node31759;
	wire [4-1:0] node31760;
	wire [4-1:0] node31763;
	wire [4-1:0] node31767;
	wire [4-1:0] node31768;
	wire [4-1:0] node31771;
	wire [4-1:0] node31774;
	wire [4-1:0] node31775;
	wire [4-1:0] node31776;
	wire [4-1:0] node31779;
	wire [4-1:0] node31782;
	wire [4-1:0] node31783;
	wire [4-1:0] node31787;
	wire [4-1:0] node31788;
	wire [4-1:0] node31789;
	wire [4-1:0] node31791;
	wire [4-1:0] node31792;
	wire [4-1:0] node31796;
	wire [4-1:0] node31797;
	wire [4-1:0] node31799;
	wire [4-1:0] node31802;
	wire [4-1:0] node31804;
	wire [4-1:0] node31807;
	wire [4-1:0] node31808;
	wire [4-1:0] node31809;
	wire [4-1:0] node31812;
	wire [4-1:0] node31815;
	wire [4-1:0] node31818;
	wire [4-1:0] node31819;
	wire [4-1:0] node31820;
	wire [4-1:0] node31821;
	wire [4-1:0] node31823;
	wire [4-1:0] node31825;
	wire [4-1:0] node31828;
	wire [4-1:0] node31829;
	wire [4-1:0] node31830;
	wire [4-1:0] node31834;
	wire [4-1:0] node31837;
	wire [4-1:0] node31838;
	wire [4-1:0] node31839;
	wire [4-1:0] node31840;
	wire [4-1:0] node31844;
	wire [4-1:0] node31845;
	wire [4-1:0] node31848;
	wire [4-1:0] node31851;
	wire [4-1:0] node31852;
	wire [4-1:0] node31854;
	wire [4-1:0] node31855;
	wire [4-1:0] node31860;
	wire [4-1:0] node31861;
	wire [4-1:0] node31862;
	wire [4-1:0] node31863;
	wire [4-1:0] node31866;
	wire [4-1:0] node31869;
	wire [4-1:0] node31870;
	wire [4-1:0] node31872;
	wire [4-1:0] node31875;
	wire [4-1:0] node31876;
	wire [4-1:0] node31877;
	wire [4-1:0] node31880;
	wire [4-1:0] node31883;
	wire [4-1:0] node31885;
	wire [4-1:0] node31888;
	wire [4-1:0] node31889;
	wire [4-1:0] node31890;
	wire [4-1:0] node31891;
	wire [4-1:0] node31895;
	wire [4-1:0] node31896;
	wire [4-1:0] node31900;
	wire [4-1:0] node31901;
	wire [4-1:0] node31905;
	wire [4-1:0] node31906;
	wire [4-1:0] node31907;
	wire [4-1:0] node31908;
	wire [4-1:0] node31909;
	wire [4-1:0] node31910;
	wire [4-1:0] node31911;
	wire [4-1:0] node31913;
	wire [4-1:0] node31918;
	wire [4-1:0] node31919;
	wire [4-1:0] node31921;
	wire [4-1:0] node31922;
	wire [4-1:0] node31926;
	wire [4-1:0] node31928;
	wire [4-1:0] node31931;
	wire [4-1:0] node31932;
	wire [4-1:0] node31933;
	wire [4-1:0] node31934;
	wire [4-1:0] node31937;
	wire [4-1:0] node31940;
	wire [4-1:0] node31941;
	wire [4-1:0] node31943;
	wire [4-1:0] node31947;
	wire [4-1:0] node31948;
	wire [4-1:0] node31949;
	wire [4-1:0] node31953;
	wire [4-1:0] node31954;
	wire [4-1:0] node31955;
	wire [4-1:0] node31959;
	wire [4-1:0] node31962;
	wire [4-1:0] node31963;
	wire [4-1:0] node31964;
	wire [4-1:0] node31965;
	wire [4-1:0] node31966;
	wire [4-1:0] node31969;
	wire [4-1:0] node31972;
	wire [4-1:0] node31973;
	wire [4-1:0] node31976;
	wire [4-1:0] node31979;
	wire [4-1:0] node31980;
	wire [4-1:0] node31981;
	wire [4-1:0] node31984;
	wire [4-1:0] node31987;
	wire [4-1:0] node31988;
	wire [4-1:0] node31991;
	wire [4-1:0] node31994;
	wire [4-1:0] node31995;
	wire [4-1:0] node31996;
	wire [4-1:0] node31999;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32006;
	wire [4-1:0] node32009;
	wire [4-1:0] node32010;
	wire [4-1:0] node32011;
	wire [4-1:0] node32012;
	wire [4-1:0] node32013;
	wire [4-1:0] node32014;
	wire [4-1:0] node32015;
	wire [4-1:0] node32018;
	wire [4-1:0] node32021;
	wire [4-1:0] node32022;
	wire [4-1:0] node32026;
	wire [4-1:0] node32028;
	wire [4-1:0] node32032;
	wire [4-1:0] node32033;
	wire [4-1:0] node32034;
	wire [4-1:0] node32037;
	wire [4-1:0] node32041;
	wire [4-1:0] node32042;
	wire [4-1:0] node32043;
	wire [4-1:0] node32044;
	wire [4-1:0] node32045;
	wire [4-1:0] node32049;
	wire [4-1:0] node32051;
	wire [4-1:0] node32055;
	wire [4-1:0] node32056;
	wire [4-1:0] node32057;
	wire [4-1:0] node32060;
	wire [4-1:0] node32064;
	wire [4-1:0] node32065;
	wire [4-1:0] node32066;
	wire [4-1:0] node32067;
	wire [4-1:0] node32068;
	wire [4-1:0] node32069;
	wire [4-1:0] node32070;
	wire [4-1:0] node32071;
	wire [4-1:0] node32072;
	wire [4-1:0] node32073;
	wire [4-1:0] node32074;
	wire [4-1:0] node32078;
	wire [4-1:0] node32080;
	wire [4-1:0] node32084;
	wire [4-1:0] node32086;
	wire [4-1:0] node32087;
	wire [4-1:0] node32090;
	wire [4-1:0] node32092;
	wire [4-1:0] node32095;
	wire [4-1:0] node32096;
	wire [4-1:0] node32097;
	wire [4-1:0] node32098;
	wire [4-1:0] node32103;
	wire [4-1:0] node32105;
	wire [4-1:0] node32106;
	wire [4-1:0] node32107;
	wire [4-1:0] node32110;
	wire [4-1:0] node32113;
	wire [4-1:0] node32114;
	wire [4-1:0] node32117;
	wire [4-1:0] node32120;
	wire [4-1:0] node32121;
	wire [4-1:0] node32122;
	wire [4-1:0] node32123;
	wire [4-1:0] node32125;
	wire [4-1:0] node32126;
	wire [4-1:0] node32131;
	wire [4-1:0] node32133;
	wire [4-1:0] node32135;
	wire [4-1:0] node32138;
	wire [4-1:0] node32139;
	wire [4-1:0] node32140;
	wire [4-1:0] node32141;
	wire [4-1:0] node32144;
	wire [4-1:0] node32148;
	wire [4-1:0] node32150;
	wire [4-1:0] node32151;
	wire [4-1:0] node32155;
	wire [4-1:0] node32156;
	wire [4-1:0] node32157;
	wire [4-1:0] node32158;
	wire [4-1:0] node32160;
	wire [4-1:0] node32162;
	wire [4-1:0] node32165;
	wire [4-1:0] node32166;
	wire [4-1:0] node32167;
	wire [4-1:0] node32170;
	wire [4-1:0] node32174;
	wire [4-1:0] node32175;
	wire [4-1:0] node32176;
	wire [4-1:0] node32177;
	wire [4-1:0] node32178;
	wire [4-1:0] node32181;
	wire [4-1:0] node32184;
	wire [4-1:0] node32185;
	wire [4-1:0] node32188;
	wire [4-1:0] node32192;
	wire [4-1:0] node32193;
	wire [4-1:0] node32195;
	wire [4-1:0] node32199;
	wire [4-1:0] node32200;
	wire [4-1:0] node32201;
	wire [4-1:0] node32202;
	wire [4-1:0] node32204;
	wire [4-1:0] node32205;
	wire [4-1:0] node32210;
	wire [4-1:0] node32211;
	wire [4-1:0] node32212;
	wire [4-1:0] node32213;
	wire [4-1:0] node32216;
	wire [4-1:0] node32220;
	wire [4-1:0] node32221;
	wire [4-1:0] node32225;
	wire [4-1:0] node32226;
	wire [4-1:0] node32227;
	wire [4-1:0] node32228;
	wire [4-1:0] node32229;
	wire [4-1:0] node32235;
	wire [4-1:0] node32236;
	wire [4-1:0] node32237;
	wire [4-1:0] node32241;
	wire [4-1:0] node32242;
	wire [4-1:0] node32245;
	wire [4-1:0] node32248;
	wire [4-1:0] node32249;
	wire [4-1:0] node32250;
	wire [4-1:0] node32251;
	wire [4-1:0] node32252;
	wire [4-1:0] node32253;
	wire [4-1:0] node32254;
	wire [4-1:0] node32255;
	wire [4-1:0] node32258;
	wire [4-1:0] node32262;
	wire [4-1:0] node32263;
	wire [4-1:0] node32264;
	wire [4-1:0] node32268;
	wire [4-1:0] node32269;
	wire [4-1:0] node32272;
	wire [4-1:0] node32275;
	wire [4-1:0] node32276;
	wire [4-1:0] node32277;
	wire [4-1:0] node32278;
	wire [4-1:0] node32281;
	wire [4-1:0] node32284;
	wire [4-1:0] node32285;
	wire [4-1:0] node32288;
	wire [4-1:0] node32291;
	wire [4-1:0] node32293;
	wire [4-1:0] node32294;
	wire [4-1:0] node32297;
	wire [4-1:0] node32300;
	wire [4-1:0] node32301;
	wire [4-1:0] node32304;
	wire [4-1:0] node32307;
	wire [4-1:0] node32308;
	wire [4-1:0] node32309;
	wire [4-1:0] node32310;
	wire [4-1:0] node32314;
	wire [4-1:0] node32315;
	wire [4-1:0] node32316;
	wire [4-1:0] node32320;
	wire [4-1:0] node32321;
	wire [4-1:0] node32325;
	wire [4-1:0] node32326;
	wire [4-1:0] node32327;
	wire [4-1:0] node32328;
	wire [4-1:0] node32332;
	wire [4-1:0] node32333;
	wire [4-1:0] node32334;
	wire [4-1:0] node32337;
	wire [4-1:0] node32340;
	wire [4-1:0] node32342;
	wire [4-1:0] node32345;
	wire [4-1:0] node32346;
	wire [4-1:0] node32347;
	wire [4-1:0] node32350;
	wire [4-1:0] node32353;
	wire [4-1:0] node32355;
	wire [4-1:0] node32358;
	wire [4-1:0] node32359;
	wire [4-1:0] node32360;
	wire [4-1:0] node32361;
	wire [4-1:0] node32362;
	wire [4-1:0] node32363;
	wire [4-1:0] node32366;
	wire [4-1:0] node32369;
	wire [4-1:0] node32371;
	wire [4-1:0] node32374;
	wire [4-1:0] node32375;
	wire [4-1:0] node32376;
	wire [4-1:0] node32379;
	wire [4-1:0] node32382;
	wire [4-1:0] node32384;
	wire [4-1:0] node32387;
	wire [4-1:0] node32388;
	wire [4-1:0] node32389;
	wire [4-1:0] node32390;
	wire [4-1:0] node32393;
	wire [4-1:0] node32396;
	wire [4-1:0] node32398;
	wire [4-1:0] node32401;
	wire [4-1:0] node32402;
	wire [4-1:0] node32404;
	wire [4-1:0] node32407;
	wire [4-1:0] node32409;
	wire [4-1:0] node32412;
	wire [4-1:0] node32413;
	wire [4-1:0] node32414;
	wire [4-1:0] node32415;
	wire [4-1:0] node32416;
	wire [4-1:0] node32417;
	wire [4-1:0] node32421;
	wire [4-1:0] node32423;
	wire [4-1:0] node32427;
	wire [4-1:0] node32428;
	wire [4-1:0] node32430;
	wire [4-1:0] node32431;
	wire [4-1:0] node32434;
	wire [4-1:0] node32437;
	wire [4-1:0] node32439;
	wire [4-1:0] node32440;
	wire [4-1:0] node32443;
	wire [4-1:0] node32446;
	wire [4-1:0] node32447;
	wire [4-1:0] node32448;
	wire [4-1:0] node32449;
	wire [4-1:0] node32452;
	wire [4-1:0] node32456;
	wire [4-1:0] node32457;
	wire [4-1:0] node32460;
	wire [4-1:0] node32463;
	wire [4-1:0] node32464;
	wire [4-1:0] node32465;
	wire [4-1:0] node32466;
	wire [4-1:0] node32467;
	wire [4-1:0] node32468;
	wire [4-1:0] node32469;
	wire [4-1:0] node32472;
	wire [4-1:0] node32475;
	wire [4-1:0] node32476;
	wire [4-1:0] node32478;
	wire [4-1:0] node32479;
	wire [4-1:0] node32482;
	wire [4-1:0] node32485;
	wire [4-1:0] node32486;
	wire [4-1:0] node32488;
	wire [4-1:0] node32491;
	wire [4-1:0] node32492;
	wire [4-1:0] node32495;
	wire [4-1:0] node32498;
	wire [4-1:0] node32499;
	wire [4-1:0] node32500;
	wire [4-1:0] node32501;
	wire [4-1:0] node32505;
	wire [4-1:0] node32506;
	wire [4-1:0] node32509;
	wire [4-1:0] node32513;
	wire [4-1:0] node32514;
	wire [4-1:0] node32515;
	wire [4-1:0] node32516;
	wire [4-1:0] node32519;
	wire [4-1:0] node32522;
	wire [4-1:0] node32523;
	wire [4-1:0] node32524;
	wire [4-1:0] node32528;
	wire [4-1:0] node32529;
	wire [4-1:0] node32532;
	wire [4-1:0] node32535;
	wire [4-1:0] node32536;
	wire [4-1:0] node32539;
	wire [4-1:0] node32542;
	wire [4-1:0] node32543;
	wire [4-1:0] node32544;
	wire [4-1:0] node32545;
	wire [4-1:0] node32546;
	wire [4-1:0] node32549;
	wire [4-1:0] node32552;
	wire [4-1:0] node32553;
	wire [4-1:0] node32555;
	wire [4-1:0] node32558;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32563;
	wire [4-1:0] node32567;
	wire [4-1:0] node32568;
	wire [4-1:0] node32569;
	wire [4-1:0] node32570;
	wire [4-1:0] node32575;
	wire [4-1:0] node32576;
	wire [4-1:0] node32577;
	wire [4-1:0] node32581;
	wire [4-1:0] node32583;
	wire [4-1:0] node32586;
	wire [4-1:0] node32587;
	wire [4-1:0] node32588;
	wire [4-1:0] node32589;
	wire [4-1:0] node32591;
	wire [4-1:0] node32594;
	wire [4-1:0] node32596;
	wire [4-1:0] node32599;
	wire [4-1:0] node32600;
	wire [4-1:0] node32602;
	wire [4-1:0] node32605;
	wire [4-1:0] node32608;
	wire [4-1:0] node32609;
	wire [4-1:0] node32610;
	wire [4-1:0] node32611;
	wire [4-1:0] node32613;
	wire [4-1:0] node32617;
	wire [4-1:0] node32619;
	wire [4-1:0] node32622;
	wire [4-1:0] node32623;
	wire [4-1:0] node32624;
	wire [4-1:0] node32625;
	wire [4-1:0] node32629;
	wire [4-1:0] node32630;
	wire [4-1:0] node32634;
	wire [4-1:0] node32636;
	wire [4-1:0] node32639;
	wire [4-1:0] node32640;
	wire [4-1:0] node32641;
	wire [4-1:0] node32642;
	wire [4-1:0] node32643;
	wire [4-1:0] node32644;
	wire [4-1:0] node32646;
	wire [4-1:0] node32649;
	wire [4-1:0] node32651;
	wire [4-1:0] node32654;
	wire [4-1:0] node32655;
	wire [4-1:0] node32657;
	wire [4-1:0] node32660;
	wire [4-1:0] node32662;
	wire [4-1:0] node32665;
	wire [4-1:0] node32666;
	wire [4-1:0] node32667;
	wire [4-1:0] node32668;
	wire [4-1:0] node32672;
	wire [4-1:0] node32673;
	wire [4-1:0] node32674;
	wire [4-1:0] node32677;
	wire [4-1:0] node32680;
	wire [4-1:0] node32681;
	wire [4-1:0] node32684;
	wire [4-1:0] node32687;
	wire [4-1:0] node32688;
	wire [4-1:0] node32691;
	wire [4-1:0] node32694;
	wire [4-1:0] node32695;
	wire [4-1:0] node32696;
	wire [4-1:0] node32697;
	wire [4-1:0] node32699;
	wire [4-1:0] node32702;
	wire [4-1:0] node32703;
	wire [4-1:0] node32707;
	wire [4-1:0] node32708;
	wire [4-1:0] node32709;
	wire [4-1:0] node32712;
	wire [4-1:0] node32715;
	wire [4-1:0] node32716;
	wire [4-1:0] node32717;
	wire [4-1:0] node32720;
	wire [4-1:0] node32724;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32727;
	wire [4-1:0] node32729;
	wire [4-1:0] node32732;
	wire [4-1:0] node32735;
	wire [4-1:0] node32736;
	wire [4-1:0] node32740;
	wire [4-1:0] node32741;
	wire [4-1:0] node32742;
	wire [4-1:0] node32744;
	wire [4-1:0] node32748;
	wire [4-1:0] node32749;
	wire [4-1:0] node32751;
	wire [4-1:0] node32755;
	wire [4-1:0] node32756;
	wire [4-1:0] node32757;
	wire [4-1:0] node32758;
	wire [4-1:0] node32759;
	wire [4-1:0] node32760;
	wire [4-1:0] node32763;
	wire [4-1:0] node32766;
	wire [4-1:0] node32767;
	wire [4-1:0] node32771;
	wire [4-1:0] node32772;
	wire [4-1:0] node32775;
	wire [4-1:0] node32778;
	wire [4-1:0] node32779;
	wire [4-1:0] node32780;
	wire [4-1:0] node32783;
	wire [4-1:0] node32786;
	wire [4-1:0] node32787;
	wire [4-1:0] node32788;
	wire [4-1:0] node32791;
	wire [4-1:0] node32794;
	wire [4-1:0] node32795;
	wire [4-1:0] node32799;
	wire [4-1:0] node32800;
	wire [4-1:0] node32801;
	wire [4-1:0] node32802;
	wire [4-1:0] node32804;
	wire [4-1:0] node32807;
	wire [4-1:0] node32809;
	wire [4-1:0] node32812;
	wire [4-1:0] node32813;
	wire [4-1:0] node32814;
	wire [4-1:0] node32818;
	wire [4-1:0] node32819;
	wire [4-1:0] node32823;
	wire [4-1:0] node32824;
	wire [4-1:0] node32825;
	wire [4-1:0] node32827;
	wire [4-1:0] node32830;
	wire [4-1:0] node32831;
	wire [4-1:0] node32834;
	wire [4-1:0] node32837;
	wire [4-1:0] node32838;
	wire [4-1:0] node32841;
	wire [4-1:0] node32843;
	wire [4-1:0] node32844;
	wire [4-1:0] node32848;
	wire [4-1:0] node32849;
	wire [4-1:0] node32850;
	wire [4-1:0] node32851;
	wire [4-1:0] node32852;
	wire [4-1:0] node32853;
	wire [4-1:0] node32854;
	wire [4-1:0] node32855;
	wire [4-1:0] node32857;
	wire [4-1:0] node32861;
	wire [4-1:0] node32862;
	wire [4-1:0] node32863;
	wire [4-1:0] node32864;
	wire [4-1:0] node32868;
	wire [4-1:0] node32869;
	wire [4-1:0] node32872;
	wire [4-1:0] node32876;
	wire [4-1:0] node32877;
	wire [4-1:0] node32878;
	wire [4-1:0] node32880;
	wire [4-1:0] node32884;
	wire [4-1:0] node32885;
	wire [4-1:0] node32886;
	wire [4-1:0] node32891;
	wire [4-1:0] node32892;
	wire [4-1:0] node32893;
	wire [4-1:0] node32894;
	wire [4-1:0] node32895;
	wire [4-1:0] node32896;
	wire [4-1:0] node32899;
	wire [4-1:0] node32903;
	wire [4-1:0] node32904;
	wire [4-1:0] node32907;
	wire [4-1:0] node32909;
	wire [4-1:0] node32912;
	wire [4-1:0] node32913;
	wire [4-1:0] node32915;
	wire [4-1:0] node32917;
	wire [4-1:0] node32920;
	wire [4-1:0] node32921;
	wire [4-1:0] node32924;
	wire [4-1:0] node32927;
	wire [4-1:0] node32928;
	wire [4-1:0] node32929;
	wire [4-1:0] node32932;
	wire [4-1:0] node32934;
	wire [4-1:0] node32936;
	wire [4-1:0] node32939;
	wire [4-1:0] node32940;
	wire [4-1:0] node32942;
	wire [4-1:0] node32945;
	wire [4-1:0] node32947;
	wire [4-1:0] node32950;
	wire [4-1:0] node32951;
	wire [4-1:0] node32952;
	wire [4-1:0] node32953;
	wire [4-1:0] node32954;
	wire [4-1:0] node32956;
	wire [4-1:0] node32959;
	wire [4-1:0] node32961;
	wire [4-1:0] node32964;
	wire [4-1:0] node32965;
	wire [4-1:0] node32966;
	wire [4-1:0] node32970;
	wire [4-1:0] node32973;
	wire [4-1:0] node32974;
	wire [4-1:0] node32975;
	wire [4-1:0] node32977;
	wire [4-1:0] node32980;
	wire [4-1:0] node32981;
	wire [4-1:0] node32985;
	wire [4-1:0] node32986;
	wire [4-1:0] node32990;
	wire [4-1:0] node32991;
	wire [4-1:0] node32992;
	wire [4-1:0] node32993;
	wire [4-1:0] node32995;
	wire [4-1:0] node32998;
	wire [4-1:0] node33000;
	wire [4-1:0] node33003;
	wire [4-1:0] node33004;
	wire [4-1:0] node33006;
	wire [4-1:0] node33009;
	wire [4-1:0] node33012;
	wire [4-1:0] node33013;
	wire [4-1:0] node33014;
	wire [4-1:0] node33016;
	wire [4-1:0] node33019;
	wire [4-1:0] node33020;
	wire [4-1:0] node33024;
	wire [4-1:0] node33025;
	wire [4-1:0] node33027;
	wire [4-1:0] node33031;
	wire [4-1:0] node33032;
	wire [4-1:0] node33033;
	wire [4-1:0] node33034;
	wire [4-1:0] node33035;
	wire [4-1:0] node33036;
	wire [4-1:0] node33037;
	wire [4-1:0] node33041;
	wire [4-1:0] node33042;
	wire [4-1:0] node33045;
	wire [4-1:0] node33048;
	wire [4-1:0] node33050;
	wire [4-1:0] node33051;
	wire [4-1:0] node33055;
	wire [4-1:0] node33056;
	wire [4-1:0] node33057;
	wire [4-1:0] node33058;
	wire [4-1:0] node33061;
	wire [4-1:0] node33064;
	wire [4-1:0] node33065;
	wire [4-1:0] node33066;
	wire [4-1:0] node33069;
	wire [4-1:0] node33073;
	wire [4-1:0] node33074;
	wire [4-1:0] node33075;
	wire [4-1:0] node33076;
	wire [4-1:0] node33079;
	wire [4-1:0] node33082;
	wire [4-1:0] node33083;
	wire [4-1:0] node33086;
	wire [4-1:0] node33089;
	wire [4-1:0] node33090;
	wire [4-1:0] node33092;
	wire [4-1:0] node33095;
	wire [4-1:0] node33096;
	wire [4-1:0] node33099;
	wire [4-1:0] node33102;
	wire [4-1:0] node33103;
	wire [4-1:0] node33106;
	wire [4-1:0] node33109;
	wire [4-1:0] node33110;
	wire [4-1:0] node33111;
	wire [4-1:0] node33112;
	wire [4-1:0] node33114;
	wire [4-1:0] node33117;
	wire [4-1:0] node33118;
	wire [4-1:0] node33119;
	wire [4-1:0] node33123;
	wire [4-1:0] node33125;
	wire [4-1:0] node33128;
	wire [4-1:0] node33129;
	wire [4-1:0] node33130;
	wire [4-1:0] node33133;
	wire [4-1:0] node33136;
	wire [4-1:0] node33137;
	wire [4-1:0] node33138;
	wire [4-1:0] node33142;
	wire [4-1:0] node33144;
	wire [4-1:0] node33147;
	wire [4-1:0] node33148;
	wire [4-1:0] node33149;
	wire [4-1:0] node33150;
	wire [4-1:0] node33151;
	wire [4-1:0] node33153;
	wire [4-1:0] node33156;
	wire [4-1:0] node33157;
	wire [4-1:0] node33162;
	wire [4-1:0] node33163;
	wire [4-1:0] node33164;
	wire [4-1:0] node33169;
	wire [4-1:0] node33170;
	wire [4-1:0] node33171;
	wire [4-1:0] node33173;
	wire [4-1:0] node33177;
	wire [4-1:0] node33178;
	wire [4-1:0] node33179;
	wire [4-1:0] node33182;
	wire [4-1:0] node33186;
	wire [4-1:0] node33187;
	wire [4-1:0] node33188;
	wire [4-1:0] node33189;
	wire [4-1:0] node33190;
	wire [4-1:0] node33191;
	wire [4-1:0] node33192;
	wire [4-1:0] node33193;
	wire [4-1:0] node33196;
	wire [4-1:0] node33199;
	wire [4-1:0] node33201;
	wire [4-1:0] node33204;
	wire [4-1:0] node33205;
	wire [4-1:0] node33206;
	wire [4-1:0] node33210;
	wire [4-1:0] node33211;
	wire [4-1:0] node33214;
	wire [4-1:0] node33217;
	wire [4-1:0] node33218;
	wire [4-1:0] node33219;
	wire [4-1:0] node33220;
	wire [4-1:0] node33221;
	wire [4-1:0] node33224;
	wire [4-1:0] node33229;
	wire [4-1:0] node33230;
	wire [4-1:0] node33231;
	wire [4-1:0] node33236;
	wire [4-1:0] node33237;
	wire [4-1:0] node33238;
	wire [4-1:0] node33239;
	wire [4-1:0] node33240;
	wire [4-1:0] node33244;
	wire [4-1:0] node33245;
	wire [4-1:0] node33249;
	wire [4-1:0] node33250;
	wire [4-1:0] node33252;
	wire [4-1:0] node33256;
	wire [4-1:0] node33257;
	wire [4-1:0] node33258;
	wire [4-1:0] node33260;
	wire [4-1:0] node33263;
	wire [4-1:0] node33266;
	wire [4-1:0] node33267;
	wire [4-1:0] node33268;
	wire [4-1:0] node33272;
	wire [4-1:0] node33275;
	wire [4-1:0] node33276;
	wire [4-1:0] node33277;
	wire [4-1:0] node33278;
	wire [4-1:0] node33279;
	wire [4-1:0] node33280;
	wire [4-1:0] node33281;
	wire [4-1:0] node33284;
	wire [4-1:0] node33287;
	wire [4-1:0] node33288;
	wire [4-1:0] node33292;
	wire [4-1:0] node33293;
	wire [4-1:0] node33294;
	wire [4-1:0] node33297;
	wire [4-1:0] node33301;
	wire [4-1:0] node33302;
	wire [4-1:0] node33305;
	wire [4-1:0] node33308;
	wire [4-1:0] node33309;
	wire [4-1:0] node33310;
	wire [4-1:0] node33311;
	wire [4-1:0] node33313;
	wire [4-1:0] node33316;
	wire [4-1:0] node33318;
	wire [4-1:0] node33322;
	wire [4-1:0] node33323;
	wire [4-1:0] node33324;
	wire [4-1:0] node33328;
	wire [4-1:0] node33329;
	wire [4-1:0] node33330;
	wire [4-1:0] node33333;
	wire [4-1:0] node33337;
	wire [4-1:0] node33338;
	wire [4-1:0] node33339;
	wire [4-1:0] node33340;
	wire [4-1:0] node33341;
	wire [4-1:0] node33345;
	wire [4-1:0] node33346;
	wire [4-1:0] node33350;
	wire [4-1:0] node33351;
	wire [4-1:0] node33353;
	wire [4-1:0] node33356;
	wire [4-1:0] node33357;
	wire [4-1:0] node33361;
	wire [4-1:0] node33362;
	wire [4-1:0] node33363;
	wire [4-1:0] node33364;
	wire [4-1:0] node33367;
	wire [4-1:0] node33370;
	wire [4-1:0] node33371;
	wire [4-1:0] node33374;
	wire [4-1:0] node33377;
	wire [4-1:0] node33378;
	wire [4-1:0] node33380;
	wire [4-1:0] node33383;
	wire [4-1:0] node33384;
	wire [4-1:0] node33388;
	wire [4-1:0] node33389;
	wire [4-1:0] node33390;
	wire [4-1:0] node33391;
	wire [4-1:0] node33392;
	wire [4-1:0] node33393;
	wire [4-1:0] node33396;
	wire [4-1:0] node33397;
	wire [4-1:0] node33401;
	wire [4-1:0] node33402;
	wire [4-1:0] node33403;
	wire [4-1:0] node33407;
	wire [4-1:0] node33408;
	wire [4-1:0] node33412;
	wire [4-1:0] node33413;
	wire [4-1:0] node33414;
	wire [4-1:0] node33417;
	wire [4-1:0] node33420;
	wire [4-1:0] node33421;
	wire [4-1:0] node33423;
	wire [4-1:0] node33427;
	wire [4-1:0] node33428;
	wire [4-1:0] node33429;
	wire [4-1:0] node33431;
	wire [4-1:0] node33432;
	wire [4-1:0] node33436;
	wire [4-1:0] node33437;
	wire [4-1:0] node33439;
	wire [4-1:0] node33441;
	wire [4-1:0] node33445;
	wire [4-1:0] node33446;
	wire [4-1:0] node33447;
	wire [4-1:0] node33450;
	wire [4-1:0] node33453;
	wire [4-1:0] node33454;
	wire [4-1:0] node33457;
	wire [4-1:0] node33458;
	wire [4-1:0] node33462;
	wire [4-1:0] node33463;
	wire [4-1:0] node33464;
	wire [4-1:0] node33465;
	wire [4-1:0] node33466;
	wire [4-1:0] node33467;
	wire [4-1:0] node33470;
	wire [4-1:0] node33471;
	wire [4-1:0] node33475;
	wire [4-1:0] node33476;
	wire [4-1:0] node33477;
	wire [4-1:0] node33480;
	wire [4-1:0] node33483;
	wire [4-1:0] node33484;
	wire [4-1:0] node33487;
	wire [4-1:0] node33490;
	wire [4-1:0] node33491;
	wire [4-1:0] node33492;
	wire [4-1:0] node33496;
	wire [4-1:0] node33497;
	wire [4-1:0] node33501;
	wire [4-1:0] node33502;
	wire [4-1:0] node33503;
	wire [4-1:0] node33506;
	wire [4-1:0] node33509;
	wire [4-1:0] node33510;
	wire [4-1:0] node33513;
	wire [4-1:0] node33516;
	wire [4-1:0] node33517;
	wire [4-1:0] node33520;
	wire [4-1:0] node33523;
	wire [4-1:0] node33524;
	wire [4-1:0] node33525;
	wire [4-1:0] node33526;
	wire [4-1:0] node33527;
	wire [4-1:0] node33528;
	wire [4-1:0] node33529;
	wire [4-1:0] node33530;
	wire [4-1:0] node33531;
	wire [4-1:0] node33534;
	wire [4-1:0] node33535;
	wire [4-1:0] node33538;
	wire [4-1:0] node33539;
	wire [4-1:0] node33542;
	wire [4-1:0] node33545;
	wire [4-1:0] node33546;
	wire [4-1:0] node33549;
	wire [4-1:0] node33550;
	wire [4-1:0] node33553;
	wire [4-1:0] node33554;
	wire [4-1:0] node33557;
	wire [4-1:0] node33560;
	wire [4-1:0] node33561;
	wire [4-1:0] node33562;
	wire [4-1:0] node33565;
	wire [4-1:0] node33566;
	wire [4-1:0] node33569;
	wire [4-1:0] node33570;
	wire [4-1:0] node33574;
	wire [4-1:0] node33575;
	wire [4-1:0] node33578;
	wire [4-1:0] node33579;
	wire [4-1:0] node33582;
	wire [4-1:0] node33583;
	wire [4-1:0] node33586;
	wire [4-1:0] node33589;
	wire [4-1:0] node33590;
	wire [4-1:0] node33591;
	wire [4-1:0] node33592;
	wire [4-1:0] node33593;
	wire [4-1:0] node33595;
	wire [4-1:0] node33598;
	wire [4-1:0] node33599;
	wire [4-1:0] node33600;
	wire [4-1:0] node33601;
	wire [4-1:0] node33604;
	wire [4-1:0] node33607;
	wire [4-1:0] node33608;
	wire [4-1:0] node33611;
	wire [4-1:0] node33614;
	wire [4-1:0] node33616;
	wire [4-1:0] node33619;
	wire [4-1:0] node33620;
	wire [4-1:0] node33621;
	wire [4-1:0] node33622;
	wire [4-1:0] node33623;
	wire [4-1:0] node33628;
	wire [4-1:0] node33629;
	wire [4-1:0] node33632;
	wire [4-1:0] node33635;
	wire [4-1:0] node33636;
	wire [4-1:0] node33637;
	wire [4-1:0] node33640;
	wire [4-1:0] node33643;
	wire [4-1:0] node33645;
	wire [4-1:0] node33648;
	wire [4-1:0] node33649;
	wire [4-1:0] node33650;
	wire [4-1:0] node33651;
	wire [4-1:0] node33653;
	wire [4-1:0] node33656;
	wire [4-1:0] node33658;
	wire [4-1:0] node33661;
	wire [4-1:0] node33662;
	wire [4-1:0] node33663;
	wire [4-1:0] node33664;
	wire [4-1:0] node33667;
	wire [4-1:0] node33671;
	wire [4-1:0] node33673;
	wire [4-1:0] node33674;
	wire [4-1:0] node33677;
	wire [4-1:0] node33680;
	wire [4-1:0] node33681;
	wire [4-1:0] node33682;
	wire [4-1:0] node33683;
	wire [4-1:0] node33685;
	wire [4-1:0] node33688;
	wire [4-1:0] node33690;
	wire [4-1:0] node33693;
	wire [4-1:0] node33695;
	wire [4-1:0] node33696;
	wire [4-1:0] node33699;
	wire [4-1:0] node33702;
	wire [4-1:0] node33703;
	wire [4-1:0] node33704;
	wire [4-1:0] node33707;
	wire [4-1:0] node33710;
	wire [4-1:0] node33712;
	wire [4-1:0] node33714;
	wire [4-1:0] node33717;
	wire [4-1:0] node33718;
	wire [4-1:0] node33719;
	wire [4-1:0] node33720;
	wire [4-1:0] node33721;
	wire [4-1:0] node33722;
	wire [4-1:0] node33723;
	wire [4-1:0] node33726;
	wire [4-1:0] node33729;
	wire [4-1:0] node33730;
	wire [4-1:0] node33733;
	wire [4-1:0] node33736;
	wire [4-1:0] node33737;
	wire [4-1:0] node33740;
	wire [4-1:0] node33743;
	wire [4-1:0] node33744;
	wire [4-1:0] node33747;
	wire [4-1:0] node33750;
	wire [4-1:0] node33751;
	wire [4-1:0] node33752;
	wire [4-1:0] node33755;
	wire [4-1:0] node33758;
	wire [4-1:0] node33759;
	wire [4-1:0] node33762;
	wire [4-1:0] node33765;
	wire [4-1:0] node33766;
	wire [4-1:0] node33767;
	wire [4-1:0] node33768;
	wire [4-1:0] node33769;
	wire [4-1:0] node33771;
	wire [4-1:0] node33774;
	wire [4-1:0] node33775;
	wire [4-1:0] node33778;
	wire [4-1:0] node33782;
	wire [4-1:0] node33783;
	wire [4-1:0] node33785;
	wire [4-1:0] node33787;
	wire [4-1:0] node33790;
	wire [4-1:0] node33791;
	wire [4-1:0] node33795;
	wire [4-1:0] node33796;
	wire [4-1:0] node33797;
	wire [4-1:0] node33798;
	wire [4-1:0] node33799;
	wire [4-1:0] node33802;
	wire [4-1:0] node33805;
	wire [4-1:0] node33806;
	wire [4-1:0] node33809;
	wire [4-1:0] node33812;
	wire [4-1:0] node33813;
	wire [4-1:0] node33817;
	wire [4-1:0] node33818;
	wire [4-1:0] node33819;
	wire [4-1:0] node33822;
	wire [4-1:0] node33825;
	wire [4-1:0] node33826;
	wire [4-1:0] node33830;
	wire [4-1:0] node33831;
	wire [4-1:0] node33832;
	wire [4-1:0] node33833;
	wire [4-1:0] node33834;
	wire [4-1:0] node33835;
	wire [4-1:0] node33838;
	wire [4-1:0] node33839;
	wire [4-1:0] node33843;
	wire [4-1:0] node33844;
	wire [4-1:0] node33847;
	wire [4-1:0] node33848;
	wire [4-1:0] node33852;
	wire [4-1:0] node33853;
	wire [4-1:0] node33854;
	wire [4-1:0] node33857;
	wire [4-1:0] node33858;
	wire [4-1:0] node33862;
	wire [4-1:0] node33863;
	wire [4-1:0] node33864;
	wire [4-1:0] node33867;
	wire [4-1:0] node33870;
	wire [4-1:0] node33871;
	wire [4-1:0] node33874;
	wire [4-1:0] node33877;
	wire [4-1:0] node33878;
	wire [4-1:0] node33879;
	wire [4-1:0] node33880;
	wire [4-1:0] node33882;
	wire [4-1:0] node33885;
	wire [4-1:0] node33888;
	wire [4-1:0] node33889;
	wire [4-1:0] node33891;
	wire [4-1:0] node33894;
	wire [4-1:0] node33897;
	wire [4-1:0] node33898;
	wire [4-1:0] node33899;
	wire [4-1:0] node33901;
	wire [4-1:0] node33904;
	wire [4-1:0] node33907;
	wire [4-1:0] node33908;
	wire [4-1:0] node33910;
	wire [4-1:0] node33913;
	wire [4-1:0] node33916;
	wire [4-1:0] node33917;
	wire [4-1:0] node33918;
	wire [4-1:0] node33919;
	wire [4-1:0] node33920;
	wire [4-1:0] node33921;
	wire [4-1:0] node33922;
	wire [4-1:0] node33926;
	wire [4-1:0] node33927;
	wire [4-1:0] node33930;
	wire [4-1:0] node33933;
	wire [4-1:0] node33934;
	wire [4-1:0] node33937;
	wire [4-1:0] node33940;
	wire [4-1:0] node33941;
	wire [4-1:0] node33942;
	wire [4-1:0] node33945;
	wire [4-1:0] node33948;
	wire [4-1:0] node33949;
	wire [4-1:0] node33952;
	wire [4-1:0] node33955;
	wire [4-1:0] node33956;
	wire [4-1:0] node33957;
	wire [4-1:0] node33958;
	wire [4-1:0] node33959;
	wire [4-1:0] node33962;
	wire [4-1:0] node33965;
	wire [4-1:0] node33966;
	wire [4-1:0] node33969;
	wire [4-1:0] node33972;
	wire [4-1:0] node33973;
	wire [4-1:0] node33974;
	wire [4-1:0] node33977;
	wire [4-1:0] node33981;
	wire [4-1:0] node33982;
	wire [4-1:0] node33983;
	wire [4-1:0] node33986;
	wire [4-1:0] node33989;
	wire [4-1:0] node33990;
	wire [4-1:0] node33993;
	wire [4-1:0] node33996;
	wire [4-1:0] node33997;
	wire [4-1:0] node33998;
	wire [4-1:0] node33999;
	wire [4-1:0] node34000;
	wire [4-1:0] node34003;
	wire [4-1:0] node34006;
	wire [4-1:0] node34007;
	wire [4-1:0] node34010;
	wire [4-1:0] node34013;
	wire [4-1:0] node34014;
	wire [4-1:0] node34016;
	wire [4-1:0] node34019;
	wire [4-1:0] node34020;
	wire [4-1:0] node34023;
	wire [4-1:0] node34026;
	wire [4-1:0] node34027;
	wire [4-1:0] node34028;
	wire [4-1:0] node34029;
	wire [4-1:0] node34030;
	wire [4-1:0] node34033;
	wire [4-1:0] node34036;
	wire [4-1:0] node34037;
	wire [4-1:0] node34041;
	wire [4-1:0] node34042;
	wire [4-1:0] node34043;
	wire [4-1:0] node34046;
	wire [4-1:0] node34049;
	wire [4-1:0] node34050;
	wire [4-1:0] node34053;
	wire [4-1:0] node34056;
	wire [4-1:0] node34057;
	wire [4-1:0] node34059;
	wire [4-1:0] node34060;
	wire [4-1:0] node34063;
	wire [4-1:0] node34066;
	wire [4-1:0] node34067;
	wire [4-1:0] node34068;
	wire [4-1:0] node34071;
	wire [4-1:0] node34074;
	wire [4-1:0] node34075;
	wire [4-1:0] node34078;
	wire [4-1:0] node34081;
	wire [4-1:0] node34082;
	wire [4-1:0] node34083;
	wire [4-1:0] node34084;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34090;
	wire [4-1:0] node34092;
	wire [4-1:0] node34095;
	wire [4-1:0] node34096;
	wire [4-1:0] node34097;
	wire [4-1:0] node34098;
	wire [4-1:0] node34099;
	wire [4-1:0] node34105;
	wire [4-1:0] node34106;
	wire [4-1:0] node34107;
	wire [4-1:0] node34108;
	wire [4-1:0] node34111;
	wire [4-1:0] node34114;
	wire [4-1:0] node34116;
	wire [4-1:0] node34119;
	wire [4-1:0] node34120;
	wire [4-1:0] node34123;
	wire [4-1:0] node34126;
	wire [4-1:0] node34127;
	wire [4-1:0] node34128;
	wire [4-1:0] node34130;
	wire [4-1:0] node34133;
	wire [4-1:0] node34135;
	wire [4-1:0] node34138;
	wire [4-1:0] node34139;
	wire [4-1:0] node34140;
	wire [4-1:0] node34143;
	wire [4-1:0] node34146;
	wire [4-1:0] node34147;
	wire [4-1:0] node34151;
	wire [4-1:0] node34152;
	wire [4-1:0] node34153;
	wire [4-1:0] node34155;
	wire [4-1:0] node34158;
	wire [4-1:0] node34159;
	wire [4-1:0] node34161;
	wire [4-1:0] node34165;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34169;
	wire [4-1:0] node34172;
	wire [4-1:0] node34173;
	wire [4-1:0] node34177;
	wire [4-1:0] node34178;
	wire [4-1:0] node34182;
	wire [4-1:0] node34183;
	wire [4-1:0] node34184;
	wire [4-1:0] node34185;
	wire [4-1:0] node34186;
	wire [4-1:0] node34189;
	wire [4-1:0] node34190;
	wire [4-1:0] node34193;
	wire [4-1:0] node34196;
	wire [4-1:0] node34197;
	wire [4-1:0] node34198;
	wire [4-1:0] node34202;
	wire [4-1:0] node34203;
	wire [4-1:0] node34206;
	wire [4-1:0] node34209;
	wire [4-1:0] node34210;
	wire [4-1:0] node34211;
	wire [4-1:0] node34212;
	wire [4-1:0] node34215;
	wire [4-1:0] node34218;
	wire [4-1:0] node34219;
	wire [4-1:0] node34222;
	wire [4-1:0] node34225;
	wire [4-1:0] node34226;
	wire [4-1:0] node34227;
	wire [4-1:0] node34231;
	wire [4-1:0] node34232;
	wire [4-1:0] node34235;
	wire [4-1:0] node34238;
	wire [4-1:0] node34239;
	wire [4-1:0] node34240;
	wire [4-1:0] node34242;
	wire [4-1:0] node34245;
	wire [4-1:0] node34247;
	wire [4-1:0] node34248;
	wire [4-1:0] node34252;
	wire [4-1:0] node34253;
	wire [4-1:0] node34254;
	wire [4-1:0] node34255;
	wire [4-1:0] node34259;
	wire [4-1:0] node34260;
	wire [4-1:0] node34261;
	wire [4-1:0] node34264;
	wire [4-1:0] node34267;
	wire [4-1:0] node34270;
	wire [4-1:0] node34271;
	wire [4-1:0] node34274;
	wire [4-1:0] node34277;
	wire [4-1:0] node34278;
	wire [4-1:0] node34279;
	wire [4-1:0] node34280;
	wire [4-1:0] node34281;
	wire [4-1:0] node34282;
	wire [4-1:0] node34284;
	wire [4-1:0] node34287;
	wire [4-1:0] node34288;
	wire [4-1:0] node34292;
	wire [4-1:0] node34293;
	wire [4-1:0] node34294;
	wire [4-1:0] node34297;
	wire [4-1:0] node34300;
	wire [4-1:0] node34301;
	wire [4-1:0] node34304;
	wire [4-1:0] node34307;
	wire [4-1:0] node34308;
	wire [4-1:0] node34309;
	wire [4-1:0] node34310;
	wire [4-1:0] node34313;
	wire [4-1:0] node34316;
	wire [4-1:0] node34317;
	wire [4-1:0] node34320;
	wire [4-1:0] node34323;
	wire [4-1:0] node34324;
	wire [4-1:0] node34326;
	wire [4-1:0] node34329;
	wire [4-1:0] node34330;
	wire [4-1:0] node34334;
	wire [4-1:0] node34335;
	wire [4-1:0] node34336;
	wire [4-1:0] node34338;
	wire [4-1:0] node34341;
	wire [4-1:0] node34342;
	wire [4-1:0] node34343;
	wire [4-1:0] node34347;
	wire [4-1:0] node34348;
	wire [4-1:0] node34350;
	wire [4-1:0] node34353;
	wire [4-1:0] node34354;
	wire [4-1:0] node34355;
	wire [4-1:0] node34358;
	wire [4-1:0] node34361;
	wire [4-1:0] node34362;
	wire [4-1:0] node34365;
	wire [4-1:0] node34368;
	wire [4-1:0] node34369;
	wire [4-1:0] node34370;
	wire [4-1:0] node34372;
	wire [4-1:0] node34376;
	wire [4-1:0] node34377;
	wire [4-1:0] node34381;
	wire [4-1:0] node34382;
	wire [4-1:0] node34383;
	wire [4-1:0] node34384;
	wire [4-1:0] node34385;
	wire [4-1:0] node34388;
	wire [4-1:0] node34389;
	wire [4-1:0] node34390;
	wire [4-1:0] node34393;
	wire [4-1:0] node34394;
	wire [4-1:0] node34398;
	wire [4-1:0] node34399;
	wire [4-1:0] node34400;
	wire [4-1:0] node34405;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34410;
	wire [4-1:0] node34413;
	wire [4-1:0] node34414;
	wire [4-1:0] node34417;
	wire [4-1:0] node34420;
	wire [4-1:0] node34421;
	wire [4-1:0] node34422;
	wire [4-1:0] node34423;
	wire [4-1:0] node34426;
	wire [4-1:0] node34429;
	wire [4-1:0] node34430;
	wire [4-1:0] node34434;
	wire [4-1:0] node34435;
	wire [4-1:0] node34437;
	wire [4-1:0] node34440;
	wire [4-1:0] node34441;
	wire [4-1:0] node34445;
	wire [4-1:0] node34446;
	wire [4-1:0] node34447;
	wire [4-1:0] node34450;
	wire [4-1:0] node34451;
	wire [4-1:0] node34452;
	wire [4-1:0] node34455;
	wire [4-1:0] node34458;
	wire [4-1:0] node34459;
	wire [4-1:0] node34463;
	wire [4-1:0] node34464;
	wire [4-1:0] node34465;
	wire [4-1:0] node34466;
	wire [4-1:0] node34469;
	wire [4-1:0] node34472;
	wire [4-1:0] node34473;
	wire [4-1:0] node34474;
	wire [4-1:0] node34477;
	wire [4-1:0] node34479;
	wire [4-1:0] node34483;
	wire [4-1:0] node34484;
	wire [4-1:0] node34487;
	wire [4-1:0] node34490;
	wire [4-1:0] node34491;
	wire [4-1:0] node34492;
	wire [4-1:0] node34493;
	wire [4-1:0] node34494;
	wire [4-1:0] node34495;
	wire [4-1:0] node34496;
	wire [4-1:0] node34497;
	wire [4-1:0] node34498;
	wire [4-1:0] node34501;
	wire [4-1:0] node34503;
	wire [4-1:0] node34506;
	wire [4-1:0] node34508;
	wire [4-1:0] node34509;
	wire [4-1:0] node34512;
	wire [4-1:0] node34515;
	wire [4-1:0] node34516;
	wire [4-1:0] node34517;
	wire [4-1:0] node34518;
	wire [4-1:0] node34522;
	wire [4-1:0] node34523;
	wire [4-1:0] node34526;
	wire [4-1:0] node34529;
	wire [4-1:0] node34530;
	wire [4-1:0] node34531;
	wire [4-1:0] node34534;
	wire [4-1:0] node34537;
	wire [4-1:0] node34538;
	wire [4-1:0] node34542;
	wire [4-1:0] node34543;
	wire [4-1:0] node34544;
	wire [4-1:0] node34545;
	wire [4-1:0] node34546;
	wire [4-1:0] node34547;
	wire [4-1:0] node34552;
	wire [4-1:0] node34553;
	wire [4-1:0] node34554;
	wire [4-1:0] node34557;
	wire [4-1:0] node34560;
	wire [4-1:0] node34561;
	wire [4-1:0] node34565;
	wire [4-1:0] node34566;
	wire [4-1:0] node34567;
	wire [4-1:0] node34570;
	wire [4-1:0] node34573;
	wire [4-1:0] node34574;
	wire [4-1:0] node34577;
	wire [4-1:0] node34580;
	wire [4-1:0] node34581;
	wire [4-1:0] node34582;
	wire [4-1:0] node34583;
	wire [4-1:0] node34586;
	wire [4-1:0] node34589;
	wire [4-1:0] node34590;
	wire [4-1:0] node34593;
	wire [4-1:0] node34595;
	wire [4-1:0] node34598;
	wire [4-1:0] node34599;
	wire [4-1:0] node34600;
	wire [4-1:0] node34602;
	wire [4-1:0] node34606;
	wire [4-1:0] node34608;
	wire [4-1:0] node34609;
	wire [4-1:0] node34612;
	wire [4-1:0] node34615;
	wire [4-1:0] node34616;
	wire [4-1:0] node34617;
	wire [4-1:0] node34618;
	wire [4-1:0] node34619;
	wire [4-1:0] node34620;
	wire [4-1:0] node34621;
	wire [4-1:0] node34624;
	wire [4-1:0] node34627;
	wire [4-1:0] node34628;
	wire [4-1:0] node34632;
	wire [4-1:0] node34635;
	wire [4-1:0] node34636;
	wire [4-1:0] node34637;
	wire [4-1:0] node34640;
	wire [4-1:0] node34641;
	wire [4-1:0] node34645;
	wire [4-1:0] node34646;
	wire [4-1:0] node34649;
	wire [4-1:0] node34652;
	wire [4-1:0] node34653;
	wire [4-1:0] node34654;
	wire [4-1:0] node34655;
	wire [4-1:0] node34658;
	wire [4-1:0] node34661;
	wire [4-1:0] node34662;
	wire [4-1:0] node34665;
	wire [4-1:0] node34668;
	wire [4-1:0] node34669;
	wire [4-1:0] node34672;
	wire [4-1:0] node34673;
	wire [4-1:0] node34674;
	wire [4-1:0] node34677;
	wire [4-1:0] node34680;
	wire [4-1:0] node34682;
	wire [4-1:0] node34685;
	wire [4-1:0] node34686;
	wire [4-1:0] node34687;
	wire [4-1:0] node34688;
	wire [4-1:0] node34689;
	wire [4-1:0] node34693;
	wire [4-1:0] node34694;
	wire [4-1:0] node34696;
	wire [4-1:0] node34699;
	wire [4-1:0] node34700;
	wire [4-1:0] node34703;
	wire [4-1:0] node34706;
	wire [4-1:0] node34708;
	wire [4-1:0] node34709;
	wire [4-1:0] node34712;
	wire [4-1:0] node34715;
	wire [4-1:0] node34716;
	wire [4-1:0] node34717;
	wire [4-1:0] node34718;
	wire [4-1:0] node34719;
	wire [4-1:0] node34722;
	wire [4-1:0] node34726;
	wire [4-1:0] node34727;
	wire [4-1:0] node34730;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34736;
	wire [4-1:0] node34737;
	wire [4-1:0] node34740;
	wire [4-1:0] node34743;
	wire [4-1:0] node34744;
	wire [4-1:0] node34746;
	wire [4-1:0] node34749;
	wire [4-1:0] node34752;
	wire [4-1:0] node34753;
	wire [4-1:0] node34754;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34757;
	wire [4-1:0] node34758;
	wire [4-1:0] node34761;
	wire [4-1:0] node34763;
	wire [4-1:0] node34767;
	wire [4-1:0] node34768;
	wire [4-1:0] node34771;
	wire [4-1:0] node34774;
	wire [4-1:0] node34775;
	wire [4-1:0] node34776;
	wire [4-1:0] node34777;
	wire [4-1:0] node34781;
	wire [4-1:0] node34782;
	wire [4-1:0] node34783;
	wire [4-1:0] node34787;
	wire [4-1:0] node34790;
	wire [4-1:0] node34791;
	wire [4-1:0] node34794;
	wire [4-1:0] node34795;
	wire [4-1:0] node34799;
	wire [4-1:0] node34800;
	wire [4-1:0] node34801;
	wire [4-1:0] node34804;
	wire [4-1:0] node34805;
	wire [4-1:0] node34807;
	wire [4-1:0] node34810;
	wire [4-1:0] node34811;
	wire [4-1:0] node34815;
	wire [4-1:0] node34816;
	wire [4-1:0] node34817;
	wire [4-1:0] node34818;
	wire [4-1:0] node34821;
	wire [4-1:0] node34824;
	wire [4-1:0] node34827;
	wire [4-1:0] node34828;
	wire [4-1:0] node34830;
	wire [4-1:0] node34833;
	wire [4-1:0] node34835;
	wire [4-1:0] node34838;
	wire [4-1:0] node34839;
	wire [4-1:0] node34840;
	wire [4-1:0] node34841;
	wire [4-1:0] node34842;
	wire [4-1:0] node34845;
	wire [4-1:0] node34847;
	wire [4-1:0] node34850;
	wire [4-1:0] node34852;
	wire [4-1:0] node34853;
	wire [4-1:0] node34856;
	wire [4-1:0] node34859;
	wire [4-1:0] node34860;
	wire [4-1:0] node34861;
	wire [4-1:0] node34862;
	wire [4-1:0] node34866;
	wire [4-1:0] node34867;
	wire [4-1:0] node34870;
	wire [4-1:0] node34873;
	wire [4-1:0] node34874;
	wire [4-1:0] node34875;
	wire [4-1:0] node34879;
	wire [4-1:0] node34881;
	wire [4-1:0] node34882;
	wire [4-1:0] node34885;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34890;
	wire [4-1:0] node34893;
	wire [4-1:0] node34895;
	wire [4-1:0] node34896;
	wire [4-1:0] node34900;
	wire [4-1:0] node34901;
	wire [4-1:0] node34902;
	wire [4-1:0] node34903;
	wire [4-1:0] node34906;
	wire [4-1:0] node34909;
	wire [4-1:0] node34910;
	wire [4-1:0] node34913;
	wire [4-1:0] node34916;
	wire [4-1:0] node34917;
	wire [4-1:0] node34919;
	wire [4-1:0] node34922;
	wire [4-1:0] node34924;
	wire [4-1:0] node34927;
	wire [4-1:0] node34928;
	wire [4-1:0] node34929;
	wire [4-1:0] node34930;
	wire [4-1:0] node34931;
	wire [4-1:0] node34934;
	wire [4-1:0] node34935;
	wire [4-1:0] node34937;
	wire [4-1:0] node34940;
	wire [4-1:0] node34941;
	wire [4-1:0] node34945;
	wire [4-1:0] node34946;
	wire [4-1:0] node34947;
	wire [4-1:0] node34948;
	wire [4-1:0] node34949;
	wire [4-1:0] node34952;
	wire [4-1:0] node34956;
	wire [4-1:0] node34957;
	wire [4-1:0] node34958;
	wire [4-1:0] node34961;
	wire [4-1:0] node34964;
	wire [4-1:0] node34965;
	wire [4-1:0] node34968;
	wire [4-1:0] node34971;
	wire [4-1:0] node34972;
	wire [4-1:0] node34973;
	wire [4-1:0] node34977;
	wire [4-1:0] node34979;
	wire [4-1:0] node34982;
	wire [4-1:0] node34983;
	wire [4-1:0] node34984;
	wire [4-1:0] node34987;
	wire [4-1:0] node34988;
	wire [4-1:0] node34990;
	wire [4-1:0] node34993;
	wire [4-1:0] node34994;
	wire [4-1:0] node34998;
	wire [4-1:0] node34999;
	wire [4-1:0] node35000;
	wire [4-1:0] node35001;
	wire [4-1:0] node35004;
	wire [4-1:0] node35007;
	wire [4-1:0] node35008;
	wire [4-1:0] node35010;
	wire [4-1:0] node35013;
	wire [4-1:0] node35015;
	wire [4-1:0] node35016;
	wire [4-1:0] node35020;
	wire [4-1:0] node35021;
	wire [4-1:0] node35022;
	wire [4-1:0] node35026;
	wire [4-1:0] node35027;
	wire [4-1:0] node35031;
	wire [4-1:0] node35032;
	wire [4-1:0] node35033;
	wire [4-1:0] node35034;
	wire [4-1:0] node35037;
	wire [4-1:0] node35038;
	wire [4-1:0] node35040;
	wire [4-1:0] node35043;
	wire [4-1:0] node35044;
	wire [4-1:0] node35048;
	wire [4-1:0] node35049;
	wire [4-1:0] node35050;
	wire [4-1:0] node35052;
	wire [4-1:0] node35054;
	wire [4-1:0] node35055;
	wire [4-1:0] node35058;
	wire [4-1:0] node35061;
	wire [4-1:0] node35062;
	wire [4-1:0] node35065;
	wire [4-1:0] node35068;
	wire [4-1:0] node35069;
	wire [4-1:0] node35070;
	wire [4-1:0] node35074;
	wire [4-1:0] node35075;
	wire [4-1:0] node35079;
	wire [4-1:0] node35080;
	wire [4-1:0] node35081;
	wire [4-1:0] node35084;
	wire [4-1:0] node35085;
	wire [4-1:0] node35087;
	wire [4-1:0] node35090;
	wire [4-1:0] node35091;
	wire [4-1:0] node35095;
	wire [4-1:0] node35096;
	wire [4-1:0] node35097;
	wire [4-1:0] node35098;
	wire [4-1:0] node35099;
	wire [4-1:0] node35102;
	wire [4-1:0] node35105;
	wire [4-1:0] node35107;
	wire [4-1:0] node35110;
	wire [4-1:0] node35111;
	wire [4-1:0] node35114;
	wire [4-1:0] node35117;
	wire [4-1:0] node35118;
	wire [4-1:0] node35120;
	wire [4-1:0] node35123;
	wire [4-1:0] node35124;
	wire [4-1:0] node35128;
	wire [4-1:0] node35129;
	wire [4-1:0] node35130;
	wire [4-1:0] node35131;
	wire [4-1:0] node35132;
	wire [4-1:0] node35133;
	wire [4-1:0] node35134;
	wire [4-1:0] node35136;
	wire [4-1:0] node35137;
	wire [4-1:0] node35140;
	wire [4-1:0] node35143;
	wire [4-1:0] node35144;
	wire [4-1:0] node35147;
	wire [4-1:0] node35150;
	wire [4-1:0] node35151;
	wire [4-1:0] node35152;
	wire [4-1:0] node35154;
	wire [4-1:0] node35156;
	wire [4-1:0] node35159;
	wire [4-1:0] node35161;
	wire [4-1:0] node35164;
	wire [4-1:0] node35165;
	wire [4-1:0] node35166;
	wire [4-1:0] node35169;
	wire [4-1:0] node35172;
	wire [4-1:0] node35173;
	wire [4-1:0] node35177;
	wire [4-1:0] node35178;
	wire [4-1:0] node35179;
	wire [4-1:0] node35182;
	wire [4-1:0] node35183;
	wire [4-1:0] node35184;
	wire [4-1:0] node35188;
	wire [4-1:0] node35189;
	wire [4-1:0] node35193;
	wire [4-1:0] node35194;
	wire [4-1:0] node35195;
	wire [4-1:0] node35196;
	wire [4-1:0] node35200;
	wire [4-1:0] node35201;
	wire [4-1:0] node35204;
	wire [4-1:0] node35207;
	wire [4-1:0] node35208;
	wire [4-1:0] node35211;
	wire [4-1:0] node35212;
	wire [4-1:0] node35215;
	wire [4-1:0] node35218;
	wire [4-1:0] node35219;
	wire [4-1:0] node35220;
	wire [4-1:0] node35221;
	wire [4-1:0] node35222;
	wire [4-1:0] node35225;
	wire [4-1:0] node35228;
	wire [4-1:0] node35229;
	wire [4-1:0] node35232;
	wire [4-1:0] node35235;
	wire [4-1:0] node35236;
	wire [4-1:0] node35237;
	wire [4-1:0] node35239;
	wire [4-1:0] node35241;
	wire [4-1:0] node35245;
	wire [4-1:0] node35246;
	wire [4-1:0] node35247;
	wire [4-1:0] node35249;
	wire [4-1:0] node35252;
	wire [4-1:0] node35253;
	wire [4-1:0] node35256;
	wire [4-1:0] node35259;
	wire [4-1:0] node35260;
	wire [4-1:0] node35264;
	wire [4-1:0] node35265;
	wire [4-1:0] node35266;
	wire [4-1:0] node35267;
	wire [4-1:0] node35269;
	wire [4-1:0] node35272;
	wire [4-1:0] node35274;
	wire [4-1:0] node35275;
	wire [4-1:0] node35278;
	wire [4-1:0] node35281;
	wire [4-1:0] node35282;
	wire [4-1:0] node35286;
	wire [4-1:0] node35287;
	wire [4-1:0] node35288;
	wire [4-1:0] node35290;
	wire [4-1:0] node35293;
	wire [4-1:0] node35294;
	wire [4-1:0] node35298;
	wire [4-1:0] node35299;
	wire [4-1:0] node35301;
	wire [4-1:0] node35304;
	wire [4-1:0] node35305;
	wire [4-1:0] node35309;
	wire [4-1:0] node35310;
	wire [4-1:0] node35311;
	wire [4-1:0] node35312;
	wire [4-1:0] node35313;
	wire [4-1:0] node35314;
	wire [4-1:0] node35315;
	wire [4-1:0] node35318;
	wire [4-1:0] node35321;
	wire [4-1:0] node35322;
	wire [4-1:0] node35325;
	wire [4-1:0] node35328;
	wire [4-1:0] node35329;
	wire [4-1:0] node35330;
	wire [4-1:0] node35333;
	wire [4-1:0] node35337;
	wire [4-1:0] node35338;
	wire [4-1:0] node35339;
	wire [4-1:0] node35340;
	wire [4-1:0] node35344;
	wire [4-1:0] node35347;
	wire [4-1:0] node35348;
	wire [4-1:0] node35349;
	wire [4-1:0] node35352;
	wire [4-1:0] node35355;
	wire [4-1:0] node35356;
	wire [4-1:0] node35358;
	wire [4-1:0] node35361;
	wire [4-1:0] node35362;
	wire [4-1:0] node35365;
	wire [4-1:0] node35368;
	wire [4-1:0] node35369;
	wire [4-1:0] node35370;
	wire [4-1:0] node35371;
	wire [4-1:0] node35373;
	wire [4-1:0] node35374;
	wire [4-1:0] node35377;
	wire [4-1:0] node35380;
	wire [4-1:0] node35382;
	wire [4-1:0] node35383;
	wire [4-1:0] node35386;
	wire [4-1:0] node35389;
	wire [4-1:0] node35390;
	wire [4-1:0] node35391;
	wire [4-1:0] node35394;
	wire [4-1:0] node35397;
	wire [4-1:0] node35398;
	wire [4-1:0] node35401;
	wire [4-1:0] node35404;
	wire [4-1:0] node35405;
	wire [4-1:0] node35406;
	wire [4-1:0] node35407;
	wire [4-1:0] node35411;
	wire [4-1:0] node35413;
	wire [4-1:0] node35416;
	wire [4-1:0] node35417;
	wire [4-1:0] node35418;
	wire [4-1:0] node35421;
	wire [4-1:0] node35424;
	wire [4-1:0] node35425;
	wire [4-1:0] node35428;
	wire [4-1:0] node35431;
	wire [4-1:0] node35432;
	wire [4-1:0] node35433;
	wire [4-1:0] node35434;
	wire [4-1:0] node35435;
	wire [4-1:0] node35438;
	wire [4-1:0] node35441;
	wire [4-1:0] node35442;
	wire [4-1:0] node35445;
	wire [4-1:0] node35448;
	wire [4-1:0] node35449;
	wire [4-1:0] node35450;
	wire [4-1:0] node35454;
	wire [4-1:0] node35457;
	wire [4-1:0] node35458;
	wire [4-1:0] node35459;
	wire [4-1:0] node35460;
	wire [4-1:0] node35464;
	wire [4-1:0] node35467;
	wire [4-1:0] node35468;
	wire [4-1:0] node35469;
	wire [4-1:0] node35473;
	wire [4-1:0] node35476;
	wire [4-1:0] node35477;
	wire [4-1:0] node35478;
	wire [4-1:0] node35479;
	wire [4-1:0] node35480;
	wire [4-1:0] node35481;
	wire [4-1:0] node35483;
	wire [4-1:0] node35484;
	wire [4-1:0] node35487;
	wire [4-1:0] node35490;
	wire [4-1:0] node35491;
	wire [4-1:0] node35492;
	wire [4-1:0] node35495;
	wire [4-1:0] node35498;
	wire [4-1:0] node35499;
	wire [4-1:0] node35503;
	wire [4-1:0] node35504;
	wire [4-1:0] node35505;
	wire [4-1:0] node35506;
	wire [4-1:0] node35509;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35514;
	wire [4-1:0] node35517;
	wire [4-1:0] node35520;
	wire [4-1:0] node35521;
	wire [4-1:0] node35525;
	wire [4-1:0] node35526;
	wire [4-1:0] node35527;
	wire [4-1:0] node35530;
	wire [4-1:0] node35533;
	wire [4-1:0] node35535;
	wire [4-1:0] node35538;
	wire [4-1:0] node35539;
	wire [4-1:0] node35540;
	wire [4-1:0] node35541;
	wire [4-1:0] node35544;
	wire [4-1:0] node35547;
	wire [4-1:0] node35548;
	wire [4-1:0] node35549;
	wire [4-1:0] node35551;
	wire [4-1:0] node35555;
	wire [4-1:0] node35556;
	wire [4-1:0] node35558;
	wire [4-1:0] node35562;
	wire [4-1:0] node35563;
	wire [4-1:0] node35564;
	wire [4-1:0] node35565;
	wire [4-1:0] node35567;
	wire [4-1:0] node35570;
	wire [4-1:0] node35573;
	wire [4-1:0] node35574;
	wire [4-1:0] node35578;
	wire [4-1:0] node35579;
	wire [4-1:0] node35580;
	wire [4-1:0] node35584;
	wire [4-1:0] node35585;
	wire [4-1:0] node35588;
	wire [4-1:0] node35590;
	wire [4-1:0] node35593;
	wire [4-1:0] node35594;
	wire [4-1:0] node35595;
	wire [4-1:0] node35596;
	wire [4-1:0] node35597;
	wire [4-1:0] node35598;
	wire [4-1:0] node35601;
	wire [4-1:0] node35604;
	wire [4-1:0] node35605;
	wire [4-1:0] node35609;
	wire [4-1:0] node35610;
	wire [4-1:0] node35612;
	wire [4-1:0] node35615;
	wire [4-1:0] node35616;
	wire [4-1:0] node35617;
	wire [4-1:0] node35622;
	wire [4-1:0] node35623;
	wire [4-1:0] node35625;
	wire [4-1:0] node35628;
	wire [4-1:0] node35629;
	wire [4-1:0] node35630;
	wire [4-1:0] node35634;
	wire [4-1:0] node35635;
	wire [4-1:0] node35638;
	wire [4-1:0] node35641;
	wire [4-1:0] node35642;
	wire [4-1:0] node35643;
	wire [4-1:0] node35646;
	wire [4-1:0] node35649;
	wire [4-1:0] node35650;
	wire [4-1:0] node35653;
	wire [4-1:0] node35656;
	wire [4-1:0] node35657;
	wire [4-1:0] node35658;
	wire [4-1:0] node35659;
	wire [4-1:0] node35660;
	wire [4-1:0] node35662;
	wire [4-1:0] node35663;
	wire [4-1:0] node35666;
	wire [4-1:0] node35670;
	wire [4-1:0] node35671;
	wire [4-1:0] node35672;
	wire [4-1:0] node35673;
	wire [4-1:0] node35674;
	wire [4-1:0] node35677;
	wire [4-1:0] node35680;
	wire [4-1:0] node35681;
	wire [4-1:0] node35684;
	wire [4-1:0] node35687;
	wire [4-1:0] node35688;
	wire [4-1:0] node35690;
	wire [4-1:0] node35693;
	wire [4-1:0] node35694;
	wire [4-1:0] node35697;
	wire [4-1:0] node35701;
	wire [4-1:0] node35702;
	wire [4-1:0] node35703;
	wire [4-1:0] node35704;
	wire [4-1:0] node35707;
	wire [4-1:0] node35711;
	wire [4-1:0] node35712;
	wire [4-1:0] node35713;
	wire [4-1:0] node35716;
	wire [4-1:0] node35720;
	wire [4-1:0] node35721;
	wire [4-1:0] node35722;
	wire [4-1:0] node35723;
	wire [4-1:0] node35725;
	wire [4-1:0] node35727;
	wire [4-1:0] node35729;
	wire [4-1:0] node35732;
	wire [4-1:0] node35733;
	wire [4-1:0] node35736;
	wire [4-1:0] node35739;
	wire [4-1:0] node35740;
	wire [4-1:0] node35741;
	wire [4-1:0] node35743;
	wire [4-1:0] node35744;
	wire [4-1:0] node35748;
	wire [4-1:0] node35749;
	wire [4-1:0] node35751;
	wire [4-1:0] node35755;
	wire [4-1:0] node35756;
	wire [4-1:0] node35757;
	wire [4-1:0] node35759;
	wire [4-1:0] node35763;
	wire [4-1:0] node35765;
	wire [4-1:0] node35766;
	wire [4-1:0] node35770;
	wire [4-1:0] node35771;
	wire [4-1:0] node35772;
	wire [4-1:0] node35773;
	wire [4-1:0] node35775;
	wire [4-1:0] node35778;
	wire [4-1:0] node35780;
	wire [4-1:0] node35782;
	wire [4-1:0] node35785;
	wire [4-1:0] node35786;
	wire [4-1:0] node35788;
	wire [4-1:0] node35791;
	wire [4-1:0] node35793;
	wire [4-1:0] node35794;
	wire [4-1:0] node35797;
	wire [4-1:0] node35800;
	wire [4-1:0] node35801;
	wire [4-1:0] node35802;
	wire [4-1:0] node35803;
	wire [4-1:0] node35807;
	wire [4-1:0] node35808;
	wire [4-1:0] node35812;
	wire [4-1:0] node35813;
	wire [4-1:0] node35816;
	wire [4-1:0] node35817;
	wire [4-1:0] node35821;
	wire [4-1:0] node35822;
	wire [4-1:0] node35823;
	wire [4-1:0] node35824;
	wire [4-1:0] node35825;
	wire [4-1:0] node35826;
	wire [4-1:0] node35827;
	wire [4-1:0] node35828;
	wire [4-1:0] node35829;
	wire [4-1:0] node35832;
	wire [4-1:0] node35833;
	wire [4-1:0] node35834;
	wire [4-1:0] node35837;
	wire [4-1:0] node35840;
	wire [4-1:0] node35841;
	wire [4-1:0] node35842;
	wire [4-1:0] node35845;
	wire [4-1:0] node35848;
	wire [4-1:0] node35849;
	wire [4-1:0] node35853;
	wire [4-1:0] node35854;
	wire [4-1:0] node35855;
	wire [4-1:0] node35858;
	wire [4-1:0] node35861;
	wire [4-1:0] node35862;
	wire [4-1:0] node35865;
	wire [4-1:0] node35868;
	wire [4-1:0] node35869;
	wire [4-1:0] node35870;
	wire [4-1:0] node35872;
	wire [4-1:0] node35875;
	wire [4-1:0] node35877;
	wire [4-1:0] node35880;
	wire [4-1:0] node35881;
	wire [4-1:0] node35882;
	wire [4-1:0] node35885;
	wire [4-1:0] node35888;
	wire [4-1:0] node35889;
	wire [4-1:0] node35893;
	wire [4-1:0] node35894;
	wire [4-1:0] node35895;
	wire [4-1:0] node35896;
	wire [4-1:0] node35899;
	wire [4-1:0] node35902;
	wire [4-1:0] node35903;
	wire [4-1:0] node35904;
	wire [4-1:0] node35907;
	wire [4-1:0] node35910;
	wire [4-1:0] node35912;
	wire [4-1:0] node35915;
	wire [4-1:0] node35916;
	wire [4-1:0] node35917;
	wire [4-1:0] node35919;
	wire [4-1:0] node35923;
	wire [4-1:0] node35924;
	wire [4-1:0] node35928;
	wire [4-1:0] node35929;
	wire [4-1:0] node35930;
	wire [4-1:0] node35931;
	wire [4-1:0] node35932;
	wire [4-1:0] node35933;
	wire [4-1:0] node35936;
	wire [4-1:0] node35939;
	wire [4-1:0] node35940;
	wire [4-1:0] node35944;
	wire [4-1:0] node35945;
	wire [4-1:0] node35946;
	wire [4-1:0] node35949;
	wire [4-1:0] node35952;
	wire [4-1:0] node35953;
	wire [4-1:0] node35957;
	wire [4-1:0] node35958;
	wire [4-1:0] node35959;
	wire [4-1:0] node35961;
	wire [4-1:0] node35964;
	wire [4-1:0] node35965;
	wire [4-1:0] node35969;
	wire [4-1:0] node35970;
	wire [4-1:0] node35971;
	wire [4-1:0] node35974;
	wire [4-1:0] node35977;
	wire [4-1:0] node35978;
	wire [4-1:0] node35982;
	wire [4-1:0] node35983;
	wire [4-1:0] node35984;
	wire [4-1:0] node35986;
	wire [4-1:0] node35987;
	wire [4-1:0] node35991;
	wire [4-1:0] node35992;
	wire [4-1:0] node35993;
	wire [4-1:0] node35996;
	wire [4-1:0] node35999;
	wire [4-1:0] node36001;
	wire [4-1:0] node36002;
	wire [4-1:0] node36005;
	wire [4-1:0] node36008;
	wire [4-1:0] node36009;
	wire [4-1:0] node36010;
	wire [4-1:0] node36012;
	wire [4-1:0] node36016;
	wire [4-1:0] node36017;
	wire [4-1:0] node36020;
	wire [4-1:0] node36023;
	wire [4-1:0] node36024;
	wire [4-1:0] node36025;
	wire [4-1:0] node36026;
	wire [4-1:0] node36027;
	wire [4-1:0] node36028;
	wire [4-1:0] node36029;
	wire [4-1:0] node36033;
	wire [4-1:0] node36034;
	wire [4-1:0] node36036;
	wire [4-1:0] node36037;
	wire [4-1:0] node36040;
	wire [4-1:0] node36043;
	wire [4-1:0] node36044;
	wire [4-1:0] node36045;
	wire [4-1:0] node36048;
	wire [4-1:0] node36052;
	wire [4-1:0] node36053;
	wire [4-1:0] node36054;
	wire [4-1:0] node36057;
	wire [4-1:0] node36060;
	wire [4-1:0] node36063;
	wire [4-1:0] node36064;
	wire [4-1:0] node36065;
	wire [4-1:0] node36066;
	wire [4-1:0] node36070;
	wire [4-1:0] node36071;
	wire [4-1:0] node36074;
	wire [4-1:0] node36077;
	wire [4-1:0] node36078;
	wire [4-1:0] node36079;
	wire [4-1:0] node36083;
	wire [4-1:0] node36084;
	wire [4-1:0] node36088;
	wire [4-1:0] node36089;
	wire [4-1:0] node36090;
	wire [4-1:0] node36092;
	wire [4-1:0] node36095;
	wire [4-1:0] node36097;
	wire [4-1:0] node36098;
	wire [4-1:0] node36102;
	wire [4-1:0] node36103;
	wire [4-1:0] node36104;
	wire [4-1:0] node36105;
	wire [4-1:0] node36109;
	wire [4-1:0] node36110;
	wire [4-1:0] node36112;
	wire [4-1:0] node36113;
	wire [4-1:0] node36116;
	wire [4-1:0] node36119;
	wire [4-1:0] node36120;
	wire [4-1:0] node36123;
	wire [4-1:0] node36126;
	wire [4-1:0] node36127;
	wire [4-1:0] node36131;
	wire [4-1:0] node36132;
	wire [4-1:0] node36133;
	wire [4-1:0] node36134;
	wire [4-1:0] node36135;
	wire [4-1:0] node36138;
	wire [4-1:0] node36139;
	wire [4-1:0] node36142;
	wire [4-1:0] node36145;
	wire [4-1:0] node36146;
	wire [4-1:0] node36147;
	wire [4-1:0] node36148;
	wire [4-1:0] node36152;
	wire [4-1:0] node36153;
	wire [4-1:0] node36156;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36163;
	wire [4-1:0] node36166;
	wire [4-1:0] node36167;
	wire [4-1:0] node36168;
	wire [4-1:0] node36169;
	wire [4-1:0] node36172;
	wire [4-1:0] node36175;
	wire [4-1:0] node36176;
	wire [4-1:0] node36179;
	wire [4-1:0] node36182;
	wire [4-1:0] node36183;
	wire [4-1:0] node36185;
	wire [4-1:0] node36188;
	wire [4-1:0] node36189;
	wire [4-1:0] node36192;
	wire [4-1:0] node36195;
	wire [4-1:0] node36196;
	wire [4-1:0] node36197;
	wire [4-1:0] node36199;
	wire [4-1:0] node36202;
	wire [4-1:0] node36203;
	wire [4-1:0] node36204;
	wire [4-1:0] node36208;
	wire [4-1:0] node36209;
	wire [4-1:0] node36212;
	wire [4-1:0] node36215;
	wire [4-1:0] node36216;
	wire [4-1:0] node36218;
	wire [4-1:0] node36219;
	wire [4-1:0] node36223;
	wire [4-1:0] node36224;
	wire [4-1:0] node36228;
	wire [4-1:0] node36229;
	wire [4-1:0] node36230;
	wire [4-1:0] node36231;
	wire [4-1:0] node36232;
	wire [4-1:0] node36233;
	wire [4-1:0] node36234;
	wire [4-1:0] node36236;
	wire [4-1:0] node36237;
	wire [4-1:0] node36241;
	wire [4-1:0] node36242;
	wire [4-1:0] node36246;
	wire [4-1:0] node36247;
	wire [4-1:0] node36248;
	wire [4-1:0] node36252;
	wire [4-1:0] node36253;
	wire [4-1:0] node36257;
	wire [4-1:0] node36258;
	wire [4-1:0] node36259;
	wire [4-1:0] node36262;
	wire [4-1:0] node36265;
	wire [4-1:0] node36266;
	wire [4-1:0] node36267;
	wire [4-1:0] node36268;
	wire [4-1:0] node36272;
	wire [4-1:0] node36273;
	wire [4-1:0] node36274;
	wire [4-1:0] node36278;
	wire [4-1:0] node36279;
	wire [4-1:0] node36283;
	wire [4-1:0] node36284;
	wire [4-1:0] node36285;
	wire [4-1:0] node36288;
	wire [4-1:0] node36291;
	wire [4-1:0] node36293;
	wire [4-1:0] node36294;
	wire [4-1:0] node36297;
	wire [4-1:0] node36300;
	wire [4-1:0] node36301;
	wire [4-1:0] node36302;
	wire [4-1:0] node36303;
	wire [4-1:0] node36304;
	wire [4-1:0] node36305;
	wire [4-1:0] node36307;
	wire [4-1:0] node36310;
	wire [4-1:0] node36313;
	wire [4-1:0] node36314;
	wire [4-1:0] node36316;
	wire [4-1:0] node36319;
	wire [4-1:0] node36322;
	wire [4-1:0] node36324;
	wire [4-1:0] node36325;
	wire [4-1:0] node36328;
	wire [4-1:0] node36329;
	wire [4-1:0] node36333;
	wire [4-1:0] node36334;
	wire [4-1:0] node36335;
	wire [4-1:0] node36336;
	wire [4-1:0] node36337;
	wire [4-1:0] node36340;
	wire [4-1:0] node36343;
	wire [4-1:0] node36345;
	wire [4-1:0] node36348;
	wire [4-1:0] node36349;
	wire [4-1:0] node36353;
	wire [4-1:0] node36354;
	wire [4-1:0] node36355;
	wire [4-1:0] node36358;
	wire [4-1:0] node36361;
	wire [4-1:0] node36362;
	wire [4-1:0] node36365;
	wire [4-1:0] node36368;
	wire [4-1:0] node36369;
	wire [4-1:0] node36370;
	wire [4-1:0] node36371;
	wire [4-1:0] node36372;
	wire [4-1:0] node36373;
	wire [4-1:0] node36377;
	wire [4-1:0] node36378;
	wire [4-1:0] node36381;
	wire [4-1:0] node36384;
	wire [4-1:0] node36385;
	wire [4-1:0] node36386;
	wire [4-1:0] node36391;
	wire [4-1:0] node36393;
	wire [4-1:0] node36394;
	wire [4-1:0] node36395;
	wire [4-1:0] node36399;
	wire [4-1:0] node36400;
	wire [4-1:0] node36403;
	wire [4-1:0] node36406;
	wire [4-1:0] node36407;
	wire [4-1:0] node36408;
	wire [4-1:0] node36410;
	wire [4-1:0] node36414;
	wire [4-1:0] node36415;
	wire [4-1:0] node36416;
	wire [4-1:0] node36418;
	wire [4-1:0] node36421;
	wire [4-1:0] node36422;
	wire [4-1:0] node36425;
	wire [4-1:0] node36428;
	wire [4-1:0] node36429;
	wire [4-1:0] node36433;
	wire [4-1:0] node36434;
	wire [4-1:0] node36435;
	wire [4-1:0] node36436;
	wire [4-1:0] node36437;
	wire [4-1:0] node36438;
	wire [4-1:0] node36439;
	wire [4-1:0] node36441;
	wire [4-1:0] node36444;
	wire [4-1:0] node36445;
	wire [4-1:0] node36448;
	wire [4-1:0] node36451;
	wire [4-1:0] node36452;
	wire [4-1:0] node36454;
	wire [4-1:0] node36457;
	wire [4-1:0] node36459;
	wire [4-1:0] node36462;
	wire [4-1:0] node36463;
	wire [4-1:0] node36464;
	wire [4-1:0] node36466;
	wire [4-1:0] node36470;
	wire [4-1:0] node36471;
	wire [4-1:0] node36475;
	wire [4-1:0] node36476;
	wire [4-1:0] node36477;
	wire [4-1:0] node36479;
	wire [4-1:0] node36480;
	wire [4-1:0] node36484;
	wire [4-1:0] node36485;
	wire [4-1:0] node36488;
	wire [4-1:0] node36492;
	wire [4-1:0] node36493;
	wire [4-1:0] node36494;
	wire [4-1:0] node36495;
	wire [4-1:0] node36496;
	wire [4-1:0] node36498;
	wire [4-1:0] node36501;
	wire [4-1:0] node36505;
	wire [4-1:0] node36506;
	wire [4-1:0] node36507;
	wire [4-1:0] node36511;
	wire [4-1:0] node36513;
	wire [4-1:0] node36516;
	wire [4-1:0] node36517;
	wire [4-1:0] node36518;
	wire [4-1:0] node36520;
	wire [4-1:0] node36521;
	wire [4-1:0] node36524;
	wire [4-1:0] node36528;
	wire [4-1:0] node36529;
	wire [4-1:0] node36530;
	wire [4-1:0] node36535;
	wire [4-1:0] node36536;
	wire [4-1:0] node36537;
	wire [4-1:0] node36538;
	wire [4-1:0] node36539;
	wire [4-1:0] node36540;
	wire [4-1:0] node36542;
	wire [4-1:0] node36545;
	wire [4-1:0] node36546;
	wire [4-1:0] node36549;
	wire [4-1:0] node36552;
	wire [4-1:0] node36554;
	wire [4-1:0] node36555;
	wire [4-1:0] node36558;
	wire [4-1:0] node36561;
	wire [4-1:0] node36562;
	wire [4-1:0] node36565;
	wire [4-1:0] node36568;
	wire [4-1:0] node36569;
	wire [4-1:0] node36570;
	wire [4-1:0] node36571;
	wire [4-1:0] node36573;
	wire [4-1:0] node36576;
	wire [4-1:0] node36577;
	wire [4-1:0] node36580;
	wire [4-1:0] node36583;
	wire [4-1:0] node36584;
	wire [4-1:0] node36585;
	wire [4-1:0] node36588;
	wire [4-1:0] node36591;
	wire [4-1:0] node36593;
	wire [4-1:0] node36596;
	wire [4-1:0] node36597;
	wire [4-1:0] node36598;
	wire [4-1:0] node36601;
	wire [4-1:0] node36604;
	wire [4-1:0] node36605;
	wire [4-1:0] node36608;
	wire [4-1:0] node36611;
	wire [4-1:0] node36612;
	wire [4-1:0] node36613;
	wire [4-1:0] node36614;
	wire [4-1:0] node36615;
	wire [4-1:0] node36616;
	wire [4-1:0] node36621;
	wire [4-1:0] node36622;
	wire [4-1:0] node36623;
	wire [4-1:0] node36626;
	wire [4-1:0] node36630;
	wire [4-1:0] node36632;
	wire [4-1:0] node36635;
	wire [4-1:0] node36636;
	wire [4-1:0] node36637;
	wire [4-1:0] node36638;
	wire [4-1:0] node36642;
	wire [4-1:0] node36643;
	wire [4-1:0] node36647;
	wire [4-1:0] node36648;
	wire [4-1:0] node36649;
	wire [4-1:0] node36654;
	wire [4-1:0] node36655;
	wire [4-1:0] node36656;
	wire [4-1:0] node36657;
	wire [4-1:0] node36658;
	wire [4-1:0] node36659;
	wire [4-1:0] node36660;
	wire [4-1:0] node36662;
	wire [4-1:0] node36665;
	wire [4-1:0] node36667;
	wire [4-1:0] node36670;
	wire [4-1:0] node36671;
	wire [4-1:0] node36672;
	wire [4-1:0] node36676;
	wire [4-1:0] node36677;
	wire [4-1:0] node36679;
	wire [4-1:0] node36682;
	wire [4-1:0] node36683;
	wire [4-1:0] node36687;
	wire [4-1:0] node36688;
	wire [4-1:0] node36689;
	wire [4-1:0] node36692;
	wire [4-1:0] node36695;
	wire [4-1:0] node36696;
	wire [4-1:0] node36700;
	wire [4-1:0] node36701;
	wire [4-1:0] node36702;
	wire [4-1:0] node36703;
	wire [4-1:0] node36704;
	wire [4-1:0] node36709;
	wire [4-1:0] node36710;
	wire [4-1:0] node36712;
	wire [4-1:0] node36714;
	wire [4-1:0] node36717;
	wire [4-1:0] node36718;
	wire [4-1:0] node36719;
	wire [4-1:0] node36723;
	wire [4-1:0] node36724;
	wire [4-1:0] node36727;
	wire [4-1:0] node36730;
	wire [4-1:0] node36731;
	wire [4-1:0] node36734;
	wire [4-1:0] node36737;
	wire [4-1:0] node36738;
	wire [4-1:0] node36739;
	wire [4-1:0] node36740;
	wire [4-1:0] node36741;
	wire [4-1:0] node36742;
	wire [4-1:0] node36745;
	wire [4-1:0] node36748;
	wire [4-1:0] node36749;
	wire [4-1:0] node36753;
	wire [4-1:0] node36754;
	wire [4-1:0] node36757;
	wire [4-1:0] node36760;
	wire [4-1:0] node36761;
	wire [4-1:0] node36764;
	wire [4-1:0] node36767;
	wire [4-1:0] node36768;
	wire [4-1:0] node36769;
	wire [4-1:0] node36770;
	wire [4-1:0] node36774;
	wire [4-1:0] node36775;
	wire [4-1:0] node36779;
	wire [4-1:0] node36780;
	wire [4-1:0] node36781;
	wire [4-1:0] node36785;
	wire [4-1:0] node36786;
	wire [4-1:0] node36790;
	wire [4-1:0] node36791;
	wire [4-1:0] node36792;
	wire [4-1:0] node36793;
	wire [4-1:0] node36794;
	wire [4-1:0] node36797;
	wire [4-1:0] node36800;
	wire [4-1:0] node36801;
	wire [4-1:0] node36802;
	wire [4-1:0] node36805;
	wire [4-1:0] node36808;
	wire [4-1:0] node36809;
	wire [4-1:0] node36812;
	wire [4-1:0] node36815;
	wire [4-1:0] node36816;
	wire [4-1:0] node36817;
	wire [4-1:0] node36818;
	wire [4-1:0] node36822;
	wire [4-1:0] node36823;
	wire [4-1:0] node36827;
	wire [4-1:0] node36828;
	wire [4-1:0] node36829;
	wire [4-1:0] node36833;
	wire [4-1:0] node36834;
	wire [4-1:0] node36838;
	wire [4-1:0] node36839;
	wire [4-1:0] node36840;
	wire [4-1:0] node36841;
	wire [4-1:0] node36842;
	wire [4-1:0] node36844;
	wire [4-1:0] node36845;
	wire [4-1:0] node36848;
	wire [4-1:0] node36851;
	wire [4-1:0] node36852;
	wire [4-1:0] node36853;
	wire [4-1:0] node36857;
	wire [4-1:0] node36858;
	wire [4-1:0] node36862;
	wire [4-1:0] node36863;
	wire [4-1:0] node36864;
	wire [4-1:0] node36867;
	wire [4-1:0] node36870;
	wire [4-1:0] node36871;
	wire [4-1:0] node36875;
	wire [4-1:0] node36876;
	wire [4-1:0] node36877;
	wire [4-1:0] node36878;
	wire [4-1:0] node36879;
	wire [4-1:0] node36882;
	wire [4-1:0] node36885;
	wire [4-1:0] node36887;
	wire [4-1:0] node36890;
	wire [4-1:0] node36891;
	wire [4-1:0] node36892;
	wire [4-1:0] node36896;
	wire [4-1:0] node36897;
	wire [4-1:0] node36900;
	wire [4-1:0] node36903;
	wire [4-1:0] node36904;
	wire [4-1:0] node36907;
	wire [4-1:0] node36910;
	wire [4-1:0] node36911;
	wire [4-1:0] node36912;
	wire [4-1:0] node36913;
	wire [4-1:0] node36914;
	wire [4-1:0] node36917;
	wire [4-1:0] node36920;
	wire [4-1:0] node36922;
	wire [4-1:0] node36925;
	wire [4-1:0] node36926;
	wire [4-1:0] node36929;
	wire [4-1:0] node36932;
	wire [4-1:0] node36933;
	wire [4-1:0] node36934;
	wire [4-1:0] node36935;
	wire [4-1:0] node36940;
	wire [4-1:0] node36941;
	wire [4-1:0] node36942;
	wire [4-1:0] node36946;
	wire [4-1:0] node36947;
	wire [4-1:0] node36951;
	wire [4-1:0] node36952;
	wire [4-1:0] node36953;
	wire [4-1:0] node36954;
	wire [4-1:0] node36955;
	wire [4-1:0] node36956;
	wire [4-1:0] node36957;
	wire [4-1:0] node36958;
	wire [4-1:0] node36959;
	wire [4-1:0] node36962;
	wire [4-1:0] node36965;
	wire [4-1:0] node36966;
	wire [4-1:0] node36967;
	wire [4-1:0] node36970;
	wire [4-1:0] node36973;
	wire [4-1:0] node36975;
	wire [4-1:0] node36978;
	wire [4-1:0] node36979;
	wire [4-1:0] node36980;
	wire [4-1:0] node36982;
	wire [4-1:0] node36985;
	wire [4-1:0] node36988;
	wire [4-1:0] node36990;
	wire [4-1:0] node36992;
	wire [4-1:0] node36995;
	wire [4-1:0] node36996;
	wire [4-1:0] node36997;
	wire [4-1:0] node36998;
	wire [4-1:0] node37000;
	wire [4-1:0] node37003;
	wire [4-1:0] node37005;
	wire [4-1:0] node37008;
	wire [4-1:0] node37010;
	wire [4-1:0] node37011;
	wire [4-1:0] node37014;
	wire [4-1:0] node37017;
	wire [4-1:0] node37018;
	wire [4-1:0] node37019;
	wire [4-1:0] node37022;
	wire [4-1:0] node37024;
	wire [4-1:0] node37027;
	wire [4-1:0] node37028;
	wire [4-1:0] node37030;
	wire [4-1:0] node37033;
	wire [4-1:0] node37035;
	wire [4-1:0] node37038;
	wire [4-1:0] node37039;
	wire [4-1:0] node37040;
	wire [4-1:0] node37041;
	wire [4-1:0] node37042;
	wire [4-1:0] node37045;
	wire [4-1:0] node37048;
	wire [4-1:0] node37049;
	wire [4-1:0] node37052;
	wire [4-1:0] node37055;
	wire [4-1:0] node37056;
	wire [4-1:0] node37059;
	wire [4-1:0] node37062;
	wire [4-1:0] node37063;
	wire [4-1:0] node37064;
	wire [4-1:0] node37065;
	wire [4-1:0] node37067;
	wire [4-1:0] node37068;
	wire [4-1:0] node37071;
	wire [4-1:0] node37074;
	wire [4-1:0] node37075;
	wire [4-1:0] node37077;
	wire [4-1:0] node37080;
	wire [4-1:0] node37081;
	wire [4-1:0] node37085;
	wire [4-1:0] node37086;
	wire [4-1:0] node37087;
	wire [4-1:0] node37091;
	wire [4-1:0] node37092;
	wire [4-1:0] node37093;
	wire [4-1:0] node37096;
	wire [4-1:0] node37099;
	wire [4-1:0] node37100;
	wire [4-1:0] node37104;
	wire [4-1:0] node37105;
	wire [4-1:0] node37106;
	wire [4-1:0] node37107;
	wire [4-1:0] node37110;
	wire [4-1:0] node37114;
	wire [4-1:0] node37115;
	wire [4-1:0] node37118;
	wire [4-1:0] node37121;
	wire [4-1:0] node37122;
	wire [4-1:0] node37123;
	wire [4-1:0] node37124;
	wire [4-1:0] node37125;
	wire [4-1:0] node37128;
	wire [4-1:0] node37131;
	wire [4-1:0] node37132;
	wire [4-1:0] node37133;
	wire [4-1:0] node37136;
	wire [4-1:0] node37139;
	wire [4-1:0] node37140;
	wire [4-1:0] node37142;
	wire [4-1:0] node37143;
	wire [4-1:0] node37146;
	wire [4-1:0] node37149;
	wire [4-1:0] node37151;
	wire [4-1:0] node37152;
	wire [4-1:0] node37155;
	wire [4-1:0] node37158;
	wire [4-1:0] node37159;
	wire [4-1:0] node37162;
	wire [4-1:0] node37165;
	wire [4-1:0] node37166;
	wire [4-1:0] node37167;
	wire [4-1:0] node37170;
	wire [4-1:0] node37173;
	wire [4-1:0] node37174;
	wire [4-1:0] node37175;
	wire [4-1:0] node37176;
	wire [4-1:0] node37179;
	wire [4-1:0] node37182;
	wire [4-1:0] node37183;
	wire [4-1:0] node37186;
	wire [4-1:0] node37189;
	wire [4-1:0] node37190;
	wire [4-1:0] node37193;
	wire [4-1:0] node37196;
	wire [4-1:0] node37197;
	wire [4-1:0] node37198;
	wire [4-1:0] node37199;
	wire [4-1:0] node37200;
	wire [4-1:0] node37201;
	wire [4-1:0] node37202;
	wire [4-1:0] node37206;
	wire [4-1:0] node37208;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37213;
	wire [4-1:0] node37217;
	wire [4-1:0] node37219;
	wire [4-1:0] node37222;
	wire [4-1:0] node37223;
	wire [4-1:0] node37224;
	wire [4-1:0] node37225;
	wire [4-1:0] node37229;
	wire [4-1:0] node37230;
	wire [4-1:0] node37234;
	wire [4-1:0] node37235;
	wire [4-1:0] node37236;
	wire [4-1:0] node37240;
	wire [4-1:0] node37242;
	wire [4-1:0] node37245;
	wire [4-1:0] node37246;
	wire [4-1:0] node37247;
	wire [4-1:0] node37248;
	wire [4-1:0] node37249;
	wire [4-1:0] node37250;
	wire [4-1:0] node37251;
	wire [4-1:0] node37255;
	wire [4-1:0] node37256;
	wire [4-1:0] node37259;
	wire [4-1:0] node37262;
	wire [4-1:0] node37263;
	wire [4-1:0] node37266;
	wire [4-1:0] node37269;
	wire [4-1:0] node37270;
	wire [4-1:0] node37271;
	wire [4-1:0] node37274;
	wire [4-1:0] node37277;
	wire [4-1:0] node37279;
	wire [4-1:0] node37282;
	wire [4-1:0] node37283;
	wire [4-1:0] node37284;
	wire [4-1:0] node37286;
	wire [4-1:0] node37289;
	wire [4-1:0] node37292;
	wire [4-1:0] node37293;
	wire [4-1:0] node37294;
	wire [4-1:0] node37297;
	wire [4-1:0] node37301;
	wire [4-1:0] node37302;
	wire [4-1:0] node37303;
	wire [4-1:0] node37304;
	wire [4-1:0] node37305;
	wire [4-1:0] node37308;
	wire [4-1:0] node37311;
	wire [4-1:0] node37312;
	wire [4-1:0] node37316;
	wire [4-1:0] node37317;
	wire [4-1:0] node37318;
	wire [4-1:0] node37321;
	wire [4-1:0] node37324;
	wire [4-1:0] node37325;
	wire [4-1:0] node37328;
	wire [4-1:0] node37331;
	wire [4-1:0] node37332;
	wire [4-1:0] node37335;
	wire [4-1:0] node37338;
	wire [4-1:0] node37339;
	wire [4-1:0] node37340;
	wire [4-1:0] node37341;
	wire [4-1:0] node37342;
	wire [4-1:0] node37343;
	wire [4-1:0] node37346;
	wire [4-1:0] node37349;
	wire [4-1:0] node37350;
	wire [4-1:0] node37352;
	wire [4-1:0] node37355;
	wire [4-1:0] node37356;
	wire [4-1:0] node37359;
	wire [4-1:0] node37362;
	wire [4-1:0] node37363;
	wire [4-1:0] node37364;
	wire [4-1:0] node37365;
	wire [4-1:0] node37366;
	wire [4-1:0] node37369;
	wire [4-1:0] node37372;
	wire [4-1:0] node37373;
	wire [4-1:0] node37377;
	wire [4-1:0] node37378;
	wire [4-1:0] node37379;
	wire [4-1:0] node37382;
	wire [4-1:0] node37385;
	wire [4-1:0] node37386;
	wire [4-1:0] node37390;
	wire [4-1:0] node37391;
	wire [4-1:0] node37394;
	wire [4-1:0] node37397;
	wire [4-1:0] node37398;
	wire [4-1:0] node37401;
	wire [4-1:0] node37404;
	wire [4-1:0] node37405;
	wire [4-1:0] node37406;
	wire [4-1:0] node37407;
	wire [4-1:0] node37410;
	wire [4-1:0] node37413;
	wire [4-1:0] node37414;
	wire [4-1:0] node37415;
	wire [4-1:0] node37417;
	wire [4-1:0] node37418;
	wire [4-1:0] node37421;
	wire [4-1:0] node37424;
	wire [4-1:0] node37425;
	wire [4-1:0] node37428;
	wire [4-1:0] node37431;
	wire [4-1:0] node37432;
	wire [4-1:0] node37433;
	wire [4-1:0] node37436;
	wire [4-1:0] node37440;
	wire [4-1:0] node37441;
	wire [4-1:0] node37442;
	wire [4-1:0] node37444;
	wire [4-1:0] node37445;
	wire [4-1:0] node37448;
	wire [4-1:0] node37449;
	wire [4-1:0] node37453;
	wire [4-1:0] node37454;
	wire [4-1:0] node37457;
	wire [4-1:0] node37460;
	wire [4-1:0] node37461;
	wire [4-1:0] node37462;
	wire [4-1:0] node37463;
	wire [4-1:0] node37464;
	wire [4-1:0] node37467;
	wire [4-1:0] node37470;
	wire [4-1:0] node37471;
	wire [4-1:0] node37474;
	wire [4-1:0] node37477;
	wire [4-1:0] node37478;
	wire [4-1:0] node37481;
	wire [4-1:0] node37484;
	wire [4-1:0] node37485;
	wire [4-1:0] node37486;
	wire [4-1:0] node37489;
	wire [4-1:0] node37492;
	wire [4-1:0] node37494;
	wire [4-1:0] node37497;
	wire [4-1:0] node37498;
	wire [4-1:0] node37499;
	wire [4-1:0] node37500;
	wire [4-1:0] node37501;
	wire [4-1:0] node37502;
	wire [4-1:0] node37505;
	wire [4-1:0] node37508;
	wire [4-1:0] node37509;
	wire [4-1:0] node37512;
	wire [4-1:0] node37515;
	wire [4-1:0] node37516;
	wire [4-1:0] node37517;
	wire [4-1:0] node37518;
	wire [4-1:0] node37519;
	wire [4-1:0] node37523;
	wire [4-1:0] node37524;
	wire [4-1:0] node37525;
	wire [4-1:0] node37528;
	wire [4-1:0] node37531;
	wire [4-1:0] node37532;
	wire [4-1:0] node37533;
	wire [4-1:0] node37537;
	wire [4-1:0] node37539;
	wire [4-1:0] node37542;
	wire [4-1:0] node37543;
	wire [4-1:0] node37544;
	wire [4-1:0] node37547;
	wire [4-1:0] node37550;
	wire [4-1:0] node37551;
	wire [4-1:0] node37552;
	wire [4-1:0] node37553;
	wire [4-1:0] node37556;
	wire [4-1:0] node37559;
	wire [4-1:0] node37560;
	wire [4-1:0] node37563;
	wire [4-1:0] node37566;
	wire [4-1:0] node37567;
	wire [4-1:0] node37570;
	wire [4-1:0] node37573;
	wire [4-1:0] node37574;
	wire [4-1:0] node37575;
	wire [4-1:0] node37576;
	wire [4-1:0] node37577;
	wire [4-1:0] node37580;
	wire [4-1:0] node37583;
	wire [4-1:0] node37585;
	wire [4-1:0] node37588;
	wire [4-1:0] node37589;
	wire [4-1:0] node37590;
	wire [4-1:0] node37593;
	wire [4-1:0] node37596;
	wire [4-1:0] node37597;
	wire [4-1:0] node37598;
	wire [4-1:0] node37601;
	wire [4-1:0] node37604;
	wire [4-1:0] node37605;
	wire [4-1:0] node37608;
	wire [4-1:0] node37611;
	wire [4-1:0] node37612;
	wire [4-1:0] node37613;
	wire [4-1:0] node37614;
	wire [4-1:0] node37617;
	wire [4-1:0] node37620;
	wire [4-1:0] node37621;
	wire [4-1:0] node37625;
	wire [4-1:0] node37627;
	wire [4-1:0] node37629;
	wire [4-1:0] node37631;
	wire [4-1:0] node37634;
	wire [4-1:0] node37635;
	wire [4-1:0] node37636;
	wire [4-1:0] node37637;
	wire [4-1:0] node37638;
	wire [4-1:0] node37639;
	wire [4-1:0] node37640;
	wire [4-1:0] node37642;
	wire [4-1:0] node37646;
	wire [4-1:0] node37647;
	wire [4-1:0] node37650;
	wire [4-1:0] node37653;
	wire [4-1:0] node37654;
	wire [4-1:0] node37657;
	wire [4-1:0] node37660;
	wire [4-1:0] node37661;
	wire [4-1:0] node37662;
	wire [4-1:0] node37666;
	wire [4-1:0] node37667;
	wire [4-1:0] node37670;
	wire [4-1:0] node37673;
	wire [4-1:0] node37674;
	wire [4-1:0] node37675;
	wire [4-1:0] node37678;
	wire [4-1:0] node37681;
	wire [4-1:0] node37682;
	wire [4-1:0] node37683;
	wire [4-1:0] node37684;
	wire [4-1:0] node37688;
	wire [4-1:0] node37689;
	wire [4-1:0] node37692;
	wire [4-1:0] node37695;
	wire [4-1:0] node37697;
	wire [4-1:0] node37700;
	wire [4-1:0] node37701;
	wire [4-1:0] node37702;
	wire [4-1:0] node37703;
	wire [4-1:0] node37706;
	wire [4-1:0] node37709;
	wire [4-1:0] node37710;
	wire [4-1:0] node37711;
	wire [4-1:0] node37714;
	wire [4-1:0] node37717;
	wire [4-1:0] node37718;
	wire [4-1:0] node37721;
	wire [4-1:0] node37724;
	wire [4-1:0] node37725;
	wire [4-1:0] node37726;
	wire [4-1:0] node37727;
	wire [4-1:0] node37730;
	wire [4-1:0] node37733;
	wire [4-1:0] node37734;
	wire [4-1:0] node37735;
	wire [4-1:0] node37738;
	wire [4-1:0] node37741;
	wire [4-1:0] node37742;
	wire [4-1:0] node37746;
	wire [4-1:0] node37747;
	wire [4-1:0] node37748;
	wire [4-1:0] node37751;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37756;
	wire [4-1:0] node37758;
	wire [4-1:0] node37762;
	wire [4-1:0] node37763;
	wire [4-1:0] node37767;
	wire [4-1:0] node37768;
	wire [4-1:0] node37769;
	wire [4-1:0] node37773;
	wire [4-1:0] node37774;
	wire [4-1:0] node37778;
	wire [4-1:0] node37779;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37783;
	wire [4-1:0] node37784;
	wire [4-1:0] node37785;
	wire [4-1:0] node37786;
	wire [4-1:0] node37787;
	wire [4-1:0] node37788;
	wire [4-1:0] node37791;
	wire [4-1:0] node37794;
	wire [4-1:0] node37795;
	wire [4-1:0] node37796;
	wire [4-1:0] node37799;
	wire [4-1:0] node37802;
	wire [4-1:0] node37803;
	wire [4-1:0] node37806;
	wire [4-1:0] node37809;
	wire [4-1:0] node37810;
	wire [4-1:0] node37811;
	wire [4-1:0] node37812;
	wire [4-1:0] node37816;
	wire [4-1:0] node37818;
	wire [4-1:0] node37820;
	wire [4-1:0] node37823;
	wire [4-1:0] node37824;
	wire [4-1:0] node37825;
	wire [4-1:0] node37826;
	wire [4-1:0] node37830;
	wire [4-1:0] node37831;
	wire [4-1:0] node37832;
	wire [4-1:0] node37836;
	wire [4-1:0] node37839;
	wire [4-1:0] node37840;
	wire [4-1:0] node37841;
	wire [4-1:0] node37845;
	wire [4-1:0] node37846;
	wire [4-1:0] node37850;
	wire [4-1:0] node37851;
	wire [4-1:0] node37852;
	wire [4-1:0] node37853;
	wire [4-1:0] node37855;
	wire [4-1:0] node37856;
	wire [4-1:0] node37859;
	wire [4-1:0] node37862;
	wire [4-1:0] node37863;
	wire [4-1:0] node37865;
	wire [4-1:0] node37868;
	wire [4-1:0] node37870;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37875;
	wire [4-1:0] node37877;
	wire [4-1:0] node37880;
	wire [4-1:0] node37882;
	wire [4-1:0] node37885;
	wire [4-1:0] node37886;
	wire [4-1:0] node37888;
	wire [4-1:0] node37891;
	wire [4-1:0] node37893;
	wire [4-1:0] node37896;
	wire [4-1:0] node37897;
	wire [4-1:0] node37898;
	wire [4-1:0] node37899;
	wire [4-1:0] node37900;
	wire [4-1:0] node37901;
	wire [4-1:0] node37905;
	wire [4-1:0] node37908;
	wire [4-1:0] node37909;
	wire [4-1:0] node37913;
	wire [4-1:0] node37914;
	wire [4-1:0] node37915;
	wire [4-1:0] node37916;
	wire [4-1:0] node37919;
	wire [4-1:0] node37922;
	wire [4-1:0] node37923;
	wire [4-1:0] node37927;
	wire [4-1:0] node37929;
	wire [4-1:0] node37930;
	wire [4-1:0] node37933;
	wire [4-1:0] node37936;
	wire [4-1:0] node37937;
	wire [4-1:0] node37939;
	wire [4-1:0] node37940;
	wire [4-1:0] node37941;
	wire [4-1:0] node37944;
	wire [4-1:0] node37947;
	wire [4-1:0] node37948;
	wire [4-1:0] node37951;
	wire [4-1:0] node37954;
	wire [4-1:0] node37955;
	wire [4-1:0] node37957;
	wire [4-1:0] node37960;
	wire [4-1:0] node37961;
	wire [4-1:0] node37964;
	wire [4-1:0] node37967;
	wire [4-1:0] node37968;
	wire [4-1:0] node37969;
	wire [4-1:0] node37970;
	wire [4-1:0] node37971;
	wire [4-1:0] node37972;
	wire [4-1:0] node37974;
	wire [4-1:0] node37975;
	wire [4-1:0] node37978;
	wire [4-1:0] node37981;
	wire [4-1:0] node37982;
	wire [4-1:0] node37983;
	wire [4-1:0] node37986;
	wire [4-1:0] node37990;
	wire [4-1:0] node37991;
	wire [4-1:0] node37992;
	wire [4-1:0] node37995;
	wire [4-1:0] node37998;
	wire [4-1:0] node37999;
	wire [4-1:0] node38002;
	wire [4-1:0] node38005;
	wire [4-1:0] node38006;
	wire [4-1:0] node38007;
	wire [4-1:0] node38008;
	wire [4-1:0] node38011;
	wire [4-1:0] node38014;
	wire [4-1:0] node38015;
	wire [4-1:0] node38018;
	wire [4-1:0] node38021;
	wire [4-1:0] node38022;
	wire [4-1:0] node38023;
	wire [4-1:0] node38026;
	wire [4-1:0] node38029;
	wire [4-1:0] node38030;
	wire [4-1:0] node38033;
	wire [4-1:0] node38036;
	wire [4-1:0] node38037;
	wire [4-1:0] node38038;
	wire [4-1:0] node38039;
	wire [4-1:0] node38041;
	wire [4-1:0] node38044;
	wire [4-1:0] node38047;
	wire [4-1:0] node38048;
	wire [4-1:0] node38050;
	wire [4-1:0] node38053;
	wire [4-1:0] node38056;
	wire [4-1:0] node38057;
	wire [4-1:0] node38058;
	wire [4-1:0] node38060;
	wire [4-1:0] node38063;
	wire [4-1:0] node38066;
	wire [4-1:0] node38068;
	wire [4-1:0] node38070;
	wire [4-1:0] node38073;
	wire [4-1:0] node38074;
	wire [4-1:0] node38075;
	wire [4-1:0] node38076;
	wire [4-1:0] node38077;
	wire [4-1:0] node38079;
	wire [4-1:0] node38080;
	wire [4-1:0] node38083;
	wire [4-1:0] node38087;
	wire [4-1:0] node38088;
	wire [4-1:0] node38089;
	wire [4-1:0] node38092;
	wire [4-1:0] node38095;
	wire [4-1:0] node38096;
	wire [4-1:0] node38099;
	wire [4-1:0] node38102;
	wire [4-1:0] node38103;
	wire [4-1:0] node38104;
	wire [4-1:0] node38105;
	wire [4-1:0] node38108;
	wire [4-1:0] node38111;
	wire [4-1:0] node38113;
	wire [4-1:0] node38114;
	wire [4-1:0] node38117;
	wire [4-1:0] node38120;
	wire [4-1:0] node38122;
	wire [4-1:0] node38123;
	wire [4-1:0] node38126;
	wire [4-1:0] node38129;
	wire [4-1:0] node38130;
	wire [4-1:0] node38131;
	wire [4-1:0] node38132;
	wire [4-1:0] node38134;
	wire [4-1:0] node38136;
	wire [4-1:0] node38139;
	wire [4-1:0] node38141;
	wire [4-1:0] node38142;
	wire [4-1:0] node38145;
	wire [4-1:0] node38148;
	wire [4-1:0] node38149;
	wire [4-1:0] node38152;
	wire [4-1:0] node38155;
	wire [4-1:0] node38156;
	wire [4-1:0] node38157;
	wire [4-1:0] node38159;
	wire [4-1:0] node38163;
	wire [4-1:0] node38164;
	wire [4-1:0] node38166;
	wire [4-1:0] node38169;
	wire [4-1:0] node38171;
	wire [4-1:0] node38174;
	wire [4-1:0] node38175;
	wire [4-1:0] node38176;
	wire [4-1:0] node38177;
	wire [4-1:0] node38178;
	wire [4-1:0] node38179;
	wire [4-1:0] node38181;
	wire [4-1:0] node38184;
	wire [4-1:0] node38187;
	wire [4-1:0] node38188;
	wire [4-1:0] node38190;
	wire [4-1:0] node38193;
	wire [4-1:0] node38195;
	wire [4-1:0] node38198;
	wire [4-1:0] node38199;
	wire [4-1:0] node38200;
	wire [4-1:0] node38201;
	wire [4-1:0] node38204;
	wire [4-1:0] node38207;
	wire [4-1:0] node38208;
	wire [4-1:0] node38210;
	wire [4-1:0] node38212;
	wire [4-1:0] node38215;
	wire [4-1:0] node38216;
	wire [4-1:0] node38218;
	wire [4-1:0] node38222;
	wire [4-1:0] node38223;
	wire [4-1:0] node38224;
	wire [4-1:0] node38225;
	wire [4-1:0] node38227;
	wire [4-1:0] node38230;
	wire [4-1:0] node38231;
	wire [4-1:0] node38234;
	wire [4-1:0] node38237;
	wire [4-1:0] node38239;
	wire [4-1:0] node38241;
	wire [4-1:0] node38244;
	wire [4-1:0] node38245;
	wire [4-1:0] node38248;
	wire [4-1:0] node38251;
	wire [4-1:0] node38252;
	wire [4-1:0] node38253;
	wire [4-1:0] node38254;
	wire [4-1:0] node38255;
	wire [4-1:0] node38256;
	wire [4-1:0] node38258;
	wire [4-1:0] node38261;
	wire [4-1:0] node38263;
	wire [4-1:0] node38266;
	wire [4-1:0] node38267;
	wire [4-1:0] node38269;
	wire [4-1:0] node38272;
	wire [4-1:0] node38274;
	wire [4-1:0] node38277;
	wire [4-1:0] node38278;
	wire [4-1:0] node38281;
	wire [4-1:0] node38282;
	wire [4-1:0] node38286;
	wire [4-1:0] node38287;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38291;
	wire [4-1:0] node38294;
	wire [4-1:0] node38295;
	wire [4-1:0] node38298;
	wire [4-1:0] node38301;
	wire [4-1:0] node38302;
	wire [4-1:0] node38306;
	wire [4-1:0] node38307;
	wire [4-1:0] node38308;
	wire [4-1:0] node38310;
	wire [4-1:0] node38314;
	wire [4-1:0] node38315;
	wire [4-1:0] node38318;
	wire [4-1:0] node38321;
	wire [4-1:0] node38322;
	wire [4-1:0] node38323;
	wire [4-1:0] node38325;
	wire [4-1:0] node38326;
	wire [4-1:0] node38328;
	wire [4-1:0] node38331;
	wire [4-1:0] node38333;
	wire [4-1:0] node38336;
	wire [4-1:0] node38337;
	wire [4-1:0] node38338;
	wire [4-1:0] node38341;
	wire [4-1:0] node38344;
	wire [4-1:0] node38346;
	wire [4-1:0] node38348;
	wire [4-1:0] node38351;
	wire [4-1:0] node38352;
	wire [4-1:0] node38353;
	wire [4-1:0] node38356;
	wire [4-1:0] node38359;
	wire [4-1:0] node38360;
	wire [4-1:0] node38361;
	wire [4-1:0] node38365;
	wire [4-1:0] node38366;
	wire [4-1:0] node38369;
	wire [4-1:0] node38372;
	wire [4-1:0] node38373;
	wire [4-1:0] node38374;
	wire [4-1:0] node38375;
	wire [4-1:0] node38376;
	wire [4-1:0] node38378;
	wire [4-1:0] node38381;
	wire [4-1:0] node38383;
	wire [4-1:0] node38386;
	wire [4-1:0] node38387;
	wire [4-1:0] node38389;
	wire [4-1:0] node38392;
	wire [4-1:0] node38394;
	wire [4-1:0] node38397;
	wire [4-1:0] node38398;
	wire [4-1:0] node38399;
	wire [4-1:0] node38400;
	wire [4-1:0] node38401;
	wire [4-1:0] node38402;
	wire [4-1:0] node38407;
	wire [4-1:0] node38408;
	wire [4-1:0] node38410;
	wire [4-1:0] node38413;
	wire [4-1:0] node38415;
	wire [4-1:0] node38418;
	wire [4-1:0] node38419;
	wire [4-1:0] node38421;
	wire [4-1:0] node38423;
	wire [4-1:0] node38426;
	wire [4-1:0] node38428;
	wire [4-1:0] node38429;
	wire [4-1:0] node38433;
	wire [4-1:0] node38434;
	wire [4-1:0] node38435;
	wire [4-1:0] node38437;
	wire [4-1:0] node38440;
	wire [4-1:0] node38442;
	wire [4-1:0] node38445;
	wire [4-1:0] node38446;
	wire [4-1:0] node38448;
	wire [4-1:0] node38451;
	wire [4-1:0] node38454;
	wire [4-1:0] node38455;
	wire [4-1:0] node38456;
	wire [4-1:0] node38457;
	wire [4-1:0] node38458;
	wire [4-1:0] node38459;
	wire [4-1:0] node38463;
	wire [4-1:0] node38464;
	wire [4-1:0] node38465;
	wire [4-1:0] node38469;
	wire [4-1:0] node38472;
	wire [4-1:0] node38473;
	wire [4-1:0] node38474;
	wire [4-1:0] node38475;
	wire [4-1:0] node38479;
	wire [4-1:0] node38482;
	wire [4-1:0] node38484;
	wire [4-1:0] node38485;
	wire [4-1:0] node38489;
	wire [4-1:0] node38490;
	wire [4-1:0] node38491;
	wire [4-1:0] node38492;
	wire [4-1:0] node38495;
	wire [4-1:0] node38498;
	wire [4-1:0] node38499;
	wire [4-1:0] node38502;
	wire [4-1:0] node38505;
	wire [4-1:0] node38506;
	wire [4-1:0] node38509;
	wire [4-1:0] node38510;
	wire [4-1:0] node38513;
	wire [4-1:0] node38516;
	wire [4-1:0] node38517;
	wire [4-1:0] node38518;
	wire [4-1:0] node38520;
	wire [4-1:0] node38521;
	wire [4-1:0] node38525;
	wire [4-1:0] node38527;
	wire [4-1:0] node38528;
	wire [4-1:0] node38532;
	wire [4-1:0] node38533;
	wire [4-1:0] node38534;
	wire [4-1:0] node38537;
	wire [4-1:0] node38538;
	wire [4-1:0] node38539;
	wire [4-1:0] node38543;
	wire [4-1:0] node38544;
	wire [4-1:0] node38548;
	wire [4-1:0] node38549;
	wire [4-1:0] node38550;
	wire [4-1:0] node38553;
	wire [4-1:0] node38556;
	wire [4-1:0] node38558;
	wire [4-1:0] node38561;
	wire [4-1:0] node38562;
	wire [4-1:0] node38563;
	wire [4-1:0] node38564;
	wire [4-1:0] node38565;
	wire [4-1:0] node38566;
	wire [4-1:0] node38567;
	wire [4-1:0] node38570;
	wire [4-1:0] node38572;
	wire [4-1:0] node38573;
	wire [4-1:0] node38577;
	wire [4-1:0] node38578;
	wire [4-1:0] node38579;
	wire [4-1:0] node38580;
	wire [4-1:0] node38584;
	wire [4-1:0] node38586;
	wire [4-1:0] node38589;
	wire [4-1:0] node38590;
	wire [4-1:0] node38592;
	wire [4-1:0] node38595;
	wire [4-1:0] node38596;
	wire [4-1:0] node38599;
	wire [4-1:0] node38600;
	wire [4-1:0] node38604;
	wire [4-1:0] node38605;
	wire [4-1:0] node38606;
	wire [4-1:0] node38609;
	wire [4-1:0] node38611;
	wire [4-1:0] node38612;
	wire [4-1:0] node38615;
	wire [4-1:0] node38618;
	wire [4-1:0] node38619;
	wire [4-1:0] node38620;
	wire [4-1:0] node38622;
	wire [4-1:0] node38624;
	wire [4-1:0] node38629;
	wire [4-1:0] node38630;
	wire [4-1:0] node38631;
	wire [4-1:0] node38632;
	wire [4-1:0] node38635;
	wire [4-1:0] node38636;
	wire [4-1:0] node38638;
	wire [4-1:0] node38641;
	wire [4-1:0] node38642;
	wire [4-1:0] node38646;
	wire [4-1:0] node38647;
	wire [4-1:0] node38648;
	wire [4-1:0] node38650;
	wire [4-1:0] node38651;
	wire [4-1:0] node38655;
	wire [4-1:0] node38656;
	wire [4-1:0] node38657;
	wire [4-1:0] node38660;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38668;
	wire [4-1:0] node38669;
	wire [4-1:0] node38671;
	wire [4-1:0] node38674;
	wire [4-1:0] node38676;
	wire [4-1:0] node38679;
	wire [4-1:0] node38680;
	wire [4-1:0] node38681;
	wire [4-1:0] node38684;
	wire [4-1:0] node38685;
	wire [4-1:0] node38687;
	wire [4-1:0] node38690;
	wire [4-1:0] node38691;
	wire [4-1:0] node38695;
	wire [4-1:0] node38696;
	wire [4-1:0] node38697;
	wire [4-1:0] node38698;
	wire [4-1:0] node38701;
	wire [4-1:0] node38704;
	wire [4-1:0] node38705;
	wire [4-1:0] node38709;
	wire [4-1:0] node38710;
	wire [4-1:0] node38712;
	wire [4-1:0] node38715;
	wire [4-1:0] node38717;
	wire [4-1:0] node38720;
	wire [4-1:0] node38721;
	wire [4-1:0] node38722;
	wire [4-1:0] node38723;
	wire [4-1:0] node38724;
	wire [4-1:0] node38727;
	wire [4-1:0] node38728;
	wire [4-1:0] node38730;
	wire [4-1:0] node38733;
	wire [4-1:0] node38734;
	wire [4-1:0] node38738;
	wire [4-1:0] node38739;
	wire [4-1:0] node38742;
	wire [4-1:0] node38743;
	wire [4-1:0] node38745;
	wire [4-1:0] node38748;
	wire [4-1:0] node38749;
	wire [4-1:0] node38753;
	wire [4-1:0] node38754;
	wire [4-1:0] node38755;
	wire [4-1:0] node38758;
	wire [4-1:0] node38759;
	wire [4-1:0] node38762;
	wire [4-1:0] node38763;
	wire [4-1:0] node38767;
	wire [4-1:0] node38768;
	wire [4-1:0] node38771;
	wire [4-1:0] node38772;
	wire [4-1:0] node38774;
	wire [4-1:0] node38777;
	wire [4-1:0] node38778;
	wire [4-1:0] node38782;
	wire [4-1:0] node38783;
	wire [4-1:0] node38784;
	wire [4-1:0] node38785;
	wire [4-1:0] node38786;
	wire [4-1:0] node38788;
	wire [4-1:0] node38791;
	wire [4-1:0] node38792;
	wire [4-1:0] node38793;
	wire [4-1:0] node38798;
	wire [4-1:0] node38799;
	wire [4-1:0] node38802;
	wire [4-1:0] node38804;
	wire [4-1:0] node38807;
	wire [4-1:0] node38808;
	wire [4-1:0] node38809;
	wire [4-1:0] node38811;
	wire [4-1:0] node38812;
	wire [4-1:0] node38815;
	wire [4-1:0] node38818;
	wire [4-1:0] node38819;
	wire [4-1:0] node38820;
	wire [4-1:0] node38823;
	wire [4-1:0] node38826;
	wire [4-1:0] node38829;
	wire [4-1:0] node38830;
	wire [4-1:0] node38831;
	wire [4-1:0] node38832;
	wire [4-1:0] node38835;
	wire [4-1:0] node38838;
	wire [4-1:0] node38841;
	wire [4-1:0] node38842;
	wire [4-1:0] node38846;
	wire [4-1:0] node38847;
	wire [4-1:0] node38848;
	wire [4-1:0] node38849;
	wire [4-1:0] node38850;
	wire [4-1:0] node38852;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38859;
	wire [4-1:0] node38862;
	wire [4-1:0] node38863;
	wire [4-1:0] node38865;
	wire [4-1:0] node38868;
	wire [4-1:0] node38870;
	wire [4-1:0] node38873;
	wire [4-1:0] node38874;
	wire [4-1:0] node38875;
	wire [4-1:0] node38876;
	wire [4-1:0] node38879;
	wire [4-1:0] node38882;
	wire [4-1:0] node38884;
	wire [4-1:0] node38887;
	wire [4-1:0] node38888;
	wire [4-1:0] node38891;
	wire [4-1:0] node38894;
	wire [4-1:0] node38895;
	wire [4-1:0] node38896;
	wire [4-1:0] node38897;
	wire [4-1:0] node38900;
	wire [4-1:0] node38901;
	wire [4-1:0] node38905;
	wire [4-1:0] node38906;
	wire [4-1:0] node38908;
	wire [4-1:0] node38912;
	wire [4-1:0] node38913;
	wire [4-1:0] node38914;
	wire [4-1:0] node38915;
	wire [4-1:0] node38918;
	wire [4-1:0] node38922;
	wire [4-1:0] node38924;
	wire [4-1:0] node38927;
	wire [4-1:0] node38928;
	wire [4-1:0] node38929;
	wire [4-1:0] node38930;
	wire [4-1:0] node38931;
	wire [4-1:0] node38932;
	wire [4-1:0] node38933;
	wire [4-1:0] node38936;
	wire [4-1:0] node38938;
	wire [4-1:0] node38941;
	wire [4-1:0] node38942;
	wire [4-1:0] node38943;
	wire [4-1:0] node38947;
	wire [4-1:0] node38948;
	wire [4-1:0] node38949;
	wire [4-1:0] node38953;
	wire [4-1:0] node38954;
	wire [4-1:0] node38958;
	wire [4-1:0] node38959;
	wire [4-1:0] node38960;
	wire [4-1:0] node38962;
	wire [4-1:0] node38966;
	wire [4-1:0] node38967;
	wire [4-1:0] node38968;
	wire [4-1:0] node38972;
	wire [4-1:0] node38973;
	wire [4-1:0] node38977;
	wire [4-1:0] node38978;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38981;
	wire [4-1:0] node38983;
	wire [4-1:0] node38986;
	wire [4-1:0] node38987;
	wire [4-1:0] node38990;
	wire [4-1:0] node38993;
	wire [4-1:0] node38994;
	wire [4-1:0] node38998;
	wire [4-1:0] node38999;
	wire [4-1:0] node39001;
	wire [4-1:0] node39002;
	wire [4-1:0] node39005;
	wire [4-1:0] node39008;
	wire [4-1:0] node39009;
	wire [4-1:0] node39011;
	wire [4-1:0] node39014;
	wire [4-1:0] node39015;
	wire [4-1:0] node39019;
	wire [4-1:0] node39020;
	wire [4-1:0] node39021;
	wire [4-1:0] node39025;
	wire [4-1:0] node39027;
	wire [4-1:0] node39030;
	wire [4-1:0] node39031;
	wire [4-1:0] node39032;
	wire [4-1:0] node39035;
	wire [4-1:0] node39036;
	wire [4-1:0] node39038;
	wire [4-1:0] node39040;
	wire [4-1:0] node39043;
	wire [4-1:0] node39044;
	wire [4-1:0] node39048;
	wire [4-1:0] node39049;
	wire [4-1:0] node39050;
	wire [4-1:0] node39051;
	wire [4-1:0] node39052;
	wire [4-1:0] node39053;
	wire [4-1:0] node39057;
	wire [4-1:0] node39059;
	wire [4-1:0] node39062;
	wire [4-1:0] node39063;
	wire [4-1:0] node39067;
	wire [4-1:0] node39068;
	wire [4-1:0] node39069;
	wire [4-1:0] node39073;
	wire [4-1:0] node39074;
	wire [4-1:0] node39077;
	wire [4-1:0] node39078;
	wire [4-1:0] node39082;
	wire [4-1:0] node39083;
	wire [4-1:0] node39085;
	wire [4-1:0] node39088;
	wire [4-1:0] node39089;
	wire [4-1:0] node39093;
	wire [4-1:0] node39094;
	wire [4-1:0] node39095;
	wire [4-1:0] node39096;
	wire [4-1:0] node39099;
	wire [4-1:0] node39100;
	wire [4-1:0] node39102;
	wire [4-1:0] node39105;
	wire [4-1:0] node39106;
	wire [4-1:0] node39110;
	wire [4-1:0] node39111;
	wire [4-1:0] node39112;
	wire [4-1:0] node39113;
	wire [4-1:0] node39116;
	wire [4-1:0] node39119;
	wire [4-1:0] node39120;
	wire [4-1:0] node39121;
	wire [4-1:0] node39124;
	wire [4-1:0] node39127;
	wire [4-1:0] node39129;
	wire [4-1:0] node39132;
	wire [4-1:0] node39133;
	wire [4-1:0] node39134;
	wire [4-1:0] node39138;
	wire [4-1:0] node39139;
	wire [4-1:0] node39143;
	wire [4-1:0] node39144;
	wire [4-1:0] node39145;
	wire [4-1:0] node39148;
	wire [4-1:0] node39149;
	wire [4-1:0] node39151;
	wire [4-1:0] node39154;
	wire [4-1:0] node39155;
	wire [4-1:0] node39159;
	wire [4-1:0] node39160;
	wire [4-1:0] node39161;
	wire [4-1:0] node39162;
	wire [4-1:0] node39164;
	wire [4-1:0] node39165;
	wire [4-1:0] node39168;
	wire [4-1:0] node39171;
	wire [4-1:0] node39172;
	wire [4-1:0] node39175;
	wire [4-1:0] node39178;
	wire [4-1:0] node39179;
	wire [4-1:0] node39181;
	wire [4-1:0] node39184;
	wire [4-1:0] node39185;
	wire [4-1:0] node39188;
	wire [4-1:0] node39191;
	wire [4-1:0] node39192;
	wire [4-1:0] node39194;
	wire [4-1:0] node39197;
	wire [4-1:0] node39198;
	wire [4-1:0] node39202;
	wire [4-1:0] node39203;
	wire [4-1:0] node39204;
	wire [4-1:0] node39205;
	wire [4-1:0] node39206;
	wire [4-1:0] node39207;
	wire [4-1:0] node39208;
	wire [4-1:0] node39209;
	wire [4-1:0] node39210;
	wire [4-1:0] node39213;
	wire [4-1:0] node39216;
	wire [4-1:0] node39217;
	wire [4-1:0] node39219;
	wire [4-1:0] node39222;
	wire [4-1:0] node39224;
	wire [4-1:0] node39227;
	wire [4-1:0] node39228;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39231;
	wire [4-1:0] node39237;
	wire [4-1:0] node39238;
	wire [4-1:0] node39239;
	wire [4-1:0] node39242;
	wire [4-1:0] node39245;
	wire [4-1:0] node39246;
	wire [4-1:0] node39247;
	wire [4-1:0] node39250;
	wire [4-1:0] node39253;
	wire [4-1:0] node39254;
	wire [4-1:0] node39257;
	wire [4-1:0] node39260;
	wire [4-1:0] node39261;
	wire [4-1:0] node39262;
	wire [4-1:0] node39264;
	wire [4-1:0] node39267;
	wire [4-1:0] node39268;
	wire [4-1:0] node39271;
	wire [4-1:0] node39274;
	wire [4-1:0] node39275;
	wire [4-1:0] node39277;
	wire [4-1:0] node39280;
	wire [4-1:0] node39281;
	wire [4-1:0] node39284;
	wire [4-1:0] node39287;
	wire [4-1:0] node39288;
	wire [4-1:0] node39289;
	wire [4-1:0] node39290;
	wire [4-1:0] node39291;
	wire [4-1:0] node39292;
	wire [4-1:0] node39293;
	wire [4-1:0] node39296;
	wire [4-1:0] node39299;
	wire [4-1:0] node39300;
	wire [4-1:0] node39303;
	wire [4-1:0] node39306;
	wire [4-1:0] node39307;
	wire [4-1:0] node39310;
	wire [4-1:0] node39313;
	wire [4-1:0] node39315;
	wire [4-1:0] node39316;
	wire [4-1:0] node39317;
	wire [4-1:0] node39320;
	wire [4-1:0] node39324;
	wire [4-1:0] node39325;
	wire [4-1:0] node39326;
	wire [4-1:0] node39329;
	wire [4-1:0] node39332;
	wire [4-1:0] node39333;
	wire [4-1:0] node39336;
	wire [4-1:0] node39339;
	wire [4-1:0] node39340;
	wire [4-1:0] node39341;
	wire [4-1:0] node39344;
	wire [4-1:0] node39347;
	wire [4-1:0] node39348;
	wire [4-1:0] node39351;
	wire [4-1:0] node39354;
	wire [4-1:0] node39355;
	wire [4-1:0] node39356;
	wire [4-1:0] node39357;
	wire [4-1:0] node39358;
	wire [4-1:0] node39359;
	wire [4-1:0] node39362;
	wire [4-1:0] node39365;
	wire [4-1:0] node39366;
	wire [4-1:0] node39370;
	wire [4-1:0] node39371;
	wire [4-1:0] node39374;
	wire [4-1:0] node39377;
	wire [4-1:0] node39378;
	wire [4-1:0] node39379;
	wire [4-1:0] node39382;
	wire [4-1:0] node39385;
	wire [4-1:0] node39386;
	wire [4-1:0] node39389;
	wire [4-1:0] node39392;
	wire [4-1:0] node39393;
	wire [4-1:0] node39394;
	wire [4-1:0] node39396;
	wire [4-1:0] node39399;
	wire [4-1:0] node39400;
	wire [4-1:0] node39404;
	wire [4-1:0] node39407;
	wire [4-1:0] node39408;
	wire [4-1:0] node39409;
	wire [4-1:0] node39410;
	wire [4-1:0] node39411;
	wire [4-1:0] node39412;
	wire [4-1:0] node39415;
	wire [4-1:0] node39416;
	wire [4-1:0] node39419;
	wire [4-1:0] node39422;
	wire [4-1:0] node39423;
	wire [4-1:0] node39425;
	wire [4-1:0] node39428;
	wire [4-1:0] node39429;
	wire [4-1:0] node39432;
	wire [4-1:0] node39435;
	wire [4-1:0] node39436;
	wire [4-1:0] node39437;
	wire [4-1:0] node39440;
	wire [4-1:0] node39441;
	wire [4-1:0] node39444;
	wire [4-1:0] node39447;
	wire [4-1:0] node39448;
	wire [4-1:0] node39449;
	wire [4-1:0] node39452;
	wire [4-1:0] node39455;
	wire [4-1:0] node39456;
	wire [4-1:0] node39459;
	wire [4-1:0] node39462;
	wire [4-1:0] node39463;
	wire [4-1:0] node39464;
	wire [4-1:0] node39465;
	wire [4-1:0] node39466;
	wire [4-1:0] node39467;
	wire [4-1:0] node39468;
	wire [4-1:0] node39472;
	wire [4-1:0] node39474;
	wire [4-1:0] node39477;
	wire [4-1:0] node39478;
	wire [4-1:0] node39482;
	wire [4-1:0] node39483;
	wire [4-1:0] node39484;
	wire [4-1:0] node39488;
	wire [4-1:0] node39491;
	wire [4-1:0] node39492;
	wire [4-1:0] node39493;
	wire [4-1:0] node39494;
	wire [4-1:0] node39498;
	wire [4-1:0] node39500;
	wire [4-1:0] node39503;
	wire [4-1:0] node39504;
	wire [4-1:0] node39505;
	wire [4-1:0] node39508;
	wire [4-1:0] node39511;
	wire [4-1:0] node39513;
	wire [4-1:0] node39516;
	wire [4-1:0] node39517;
	wire [4-1:0] node39518;
	wire [4-1:0] node39519;
	wire [4-1:0] node39520;
	wire [4-1:0] node39521;
	wire [4-1:0] node39524;
	wire [4-1:0] node39527;
	wire [4-1:0] node39528;
	wire [4-1:0] node39531;
	wire [4-1:0] node39534;
	wire [4-1:0] node39536;
	wire [4-1:0] node39537;
	wire [4-1:0] node39541;
	wire [4-1:0] node39542;
	wire [4-1:0] node39543;
	wire [4-1:0] node39545;
	wire [4-1:0] node39548;
	wire [4-1:0] node39549;
	wire [4-1:0] node39552;
	wire [4-1:0] node39555;
	wire [4-1:0] node39556;
	wire [4-1:0] node39557;
	wire [4-1:0] node39561;
	wire [4-1:0] node39562;
	wire [4-1:0] node39566;
	wire [4-1:0] node39567;
	wire [4-1:0] node39568;
	wire [4-1:0] node39569;
	wire [4-1:0] node39570;
	wire [4-1:0] node39573;
	wire [4-1:0] node39577;
	wire [4-1:0] node39578;
	wire [4-1:0] node39579;
	wire [4-1:0] node39582;
	wire [4-1:0] node39585;
	wire [4-1:0] node39588;
	wire [4-1:0] node39589;
	wire [4-1:0] node39590;
	wire [4-1:0] node39591;
	wire [4-1:0] node39594;
	wire [4-1:0] node39597;
	wire [4-1:0] node39598;
	wire [4-1:0] node39602;
	wire [4-1:0] node39605;
	wire [4-1:0] node39606;
	wire [4-1:0] node39607;
	wire [4-1:0] node39608;
	wire [4-1:0] node39609;
	wire [4-1:0] node39613;
	wire [4-1:0] node39615;
	wire [4-1:0] node39618;
	wire [4-1:0] node39619;
	wire [4-1:0] node39620;
	wire [4-1:0] node39623;
	wire [4-1:0] node39626;
	wire [4-1:0] node39627;
	wire [4-1:0] node39628;
	wire [4-1:0] node39629;
	wire [4-1:0] node39632;
	wire [4-1:0] node39635;
	wire [4-1:0] node39637;
	wire [4-1:0] node39640;
	wire [4-1:0] node39641;
	wire [4-1:0] node39644;
	wire [4-1:0] node39647;
	wire [4-1:0] node39648;
	wire [4-1:0] node39649;
	wire [4-1:0] node39651;
	wire [4-1:0] node39654;
	wire [4-1:0] node39655;
	wire [4-1:0] node39659;
	wire [4-1:0] node39662;
	wire [4-1:0] node39663;
	wire [4-1:0] node39664;
	wire [4-1:0] node39665;
	wire [4-1:0] node39666;
	wire [4-1:0] node39667;
	wire [4-1:0] node39669;
	wire [4-1:0] node39672;
	wire [4-1:0] node39673;
	wire [4-1:0] node39674;
	wire [4-1:0] node39678;
	wire [4-1:0] node39680;
	wire [4-1:0] node39681;
	wire [4-1:0] node39684;
	wire [4-1:0] node39687;
	wire [4-1:0] node39688;
	wire [4-1:0] node39689;
	wire [4-1:0] node39691;
	wire [4-1:0] node39695;
	wire [4-1:0] node39696;
	wire [4-1:0] node39699;
	wire [4-1:0] node39702;
	wire [4-1:0] node39703;
	wire [4-1:0] node39704;
	wire [4-1:0] node39705;
	wire [4-1:0] node39708;
	wire [4-1:0] node39711;
	wire [4-1:0] node39712;
	wire [4-1:0] node39713;
	wire [4-1:0] node39717;
	wire [4-1:0] node39718;
	wire [4-1:0] node39719;
	wire [4-1:0] node39721;
	wire [4-1:0] node39724;
	wire [4-1:0] node39725;
	wire [4-1:0] node39729;
	wire [4-1:0] node39730;
	wire [4-1:0] node39733;
	wire [4-1:0] node39736;
	wire [4-1:0] node39737;
	wire [4-1:0] node39738;
	wire [4-1:0] node39741;
	wire [4-1:0] node39742;
	wire [4-1:0] node39746;
	wire [4-1:0] node39749;
	wire [4-1:0] node39750;
	wire [4-1:0] node39751;
	wire [4-1:0] node39752;
	wire [4-1:0] node39754;
	wire [4-1:0] node39757;
	wire [4-1:0] node39759;
	wire [4-1:0] node39762;
	wire [4-1:0] node39763;
	wire [4-1:0] node39764;
	wire [4-1:0] node39767;
	wire [4-1:0] node39770;
	wire [4-1:0] node39771;
	wire [4-1:0] node39774;
	wire [4-1:0] node39777;
	wire [4-1:0] node39778;
	wire [4-1:0] node39779;
	wire [4-1:0] node39781;
	wire [4-1:0] node39784;
	wire [4-1:0] node39785;
	wire [4-1:0] node39789;
	wire [4-1:0] node39792;
	wire [4-1:0] node39793;
	wire [4-1:0] node39794;
	wire [4-1:0] node39795;
	wire [4-1:0] node39796;
	wire [4-1:0] node39798;
	wire [4-1:0] node39801;
	wire [4-1:0] node39802;
	wire [4-1:0] node39804;
	wire [4-1:0] node39808;
	wire [4-1:0] node39809;
	wire [4-1:0] node39810;
	wire [4-1:0] node39811;
	wire [4-1:0] node39815;
	wire [4-1:0] node39816;
	wire [4-1:0] node39817;
	wire [4-1:0] node39820;
	wire [4-1:0] node39823;
	wire [4-1:0] node39824;
	wire [4-1:0] node39827;
	wire [4-1:0] node39830;
	wire [4-1:0] node39831;
	wire [4-1:0] node39834;
	wire [4-1:0] node39837;
	wire [4-1:0] node39838;
	wire [4-1:0] node39839;
	wire [4-1:0] node39840;
	wire [4-1:0] node39843;
	wire [4-1:0] node39846;
	wire [4-1:0] node39848;
	wire [4-1:0] node39849;
	wire [4-1:0] node39853;
	wire [4-1:0] node39854;
	wire [4-1:0] node39855;
	wire [4-1:0] node39856;
	wire [4-1:0] node39859;
	wire [4-1:0] node39862;
	wire [4-1:0] node39863;
	wire [4-1:0] node39864;
	wire [4-1:0] node39867;
	wire [4-1:0] node39870;
	wire [4-1:0] node39871;
	wire [4-1:0] node39874;
	wire [4-1:0] node39877;
	wire [4-1:0] node39878;
	wire [4-1:0] node39880;
	wire [4-1:0] node39881;
	wire [4-1:0] node39882;
	wire [4-1:0] node39885;
	wire [4-1:0] node39888;
	wire [4-1:0] node39889;
	wire [4-1:0] node39894;
	wire [4-1:0] node39895;
	wire [4-1:0] node39896;
	wire [4-1:0] node39897;
	wire [4-1:0] node39898;
	wire [4-1:0] node39902;
	wire [4-1:0] node39903;
	wire [4-1:0] node39907;
	wire [4-1:0] node39908;
	wire [4-1:0] node39909;
	wire [4-1:0] node39912;
	wire [4-1:0] node39915;
	wire [4-1:0] node39916;
	wire [4-1:0] node39917;
	wire [4-1:0] node39918;
	wire [4-1:0] node39919;
	wire [4-1:0] node39922;
	wire [4-1:0] node39925;
	wire [4-1:0] node39927;
	wire [4-1:0] node39930;
	wire [4-1:0] node39932;
	wire [4-1:0] node39935;
	wire [4-1:0] node39936;
	wire [4-1:0] node39939;
	wire [4-1:0] node39942;
	wire [4-1:0] node39943;
	wire [4-1:0] node39944;
	wire [4-1:0] node39946;
	wire [4-1:0] node39949;
	wire [4-1:0] node39950;
	wire [4-1:0] node39954;
	wire [4-1:0] node39957;
	wire [4-1:0] node39958;
	wire [4-1:0] node39959;
	wire [4-1:0] node39960;
	wire [4-1:0] node39961;
	wire [4-1:0] node39962;
	wire [4-1:0] node39963;
	wire [4-1:0] node39964;
	wire [4-1:0] node39965;
	wire [4-1:0] node39966;
	wire [4-1:0] node39968;
	wire [4-1:0] node39969;
	wire [4-1:0] node39972;
	wire [4-1:0] node39975;
	wire [4-1:0] node39976;
	wire [4-1:0] node39979;
	wire [4-1:0] node39982;
	wire [4-1:0] node39983;
	wire [4-1:0] node39984;
	wire [4-1:0] node39986;
	wire [4-1:0] node39989;
	wire [4-1:0] node39990;
	wire [4-1:0] node39994;
	wire [4-1:0] node39995;
	wire [4-1:0] node39999;
	wire [4-1:0] node40000;
	wire [4-1:0] node40001;
	wire [4-1:0] node40004;
	wire [4-1:0] node40007;
	wire [4-1:0] node40008;
	wire [4-1:0] node40009;
	wire [4-1:0] node40014;
	wire [4-1:0] node40015;
	wire [4-1:0] node40016;
	wire [4-1:0] node40017;
	wire [4-1:0] node40019;
	wire [4-1:0] node40022;
	wire [4-1:0] node40023;
	wire [4-1:0] node40027;
	wire [4-1:0] node40029;
	wire [4-1:0] node40030;
	wire [4-1:0] node40034;
	wire [4-1:0] node40035;
	wire [4-1:0] node40036;
	wire [4-1:0] node40037;
	wire [4-1:0] node40039;
	wire [4-1:0] node40042;
	wire [4-1:0] node40044;
	wire [4-1:0] node40047;
	wire [4-1:0] node40048;
	wire [4-1:0] node40050;
	wire [4-1:0] node40054;
	wire [4-1:0] node40055;
	wire [4-1:0] node40056;
	wire [4-1:0] node40060;
	wire [4-1:0] node40061;
	wire [4-1:0] node40064;
	wire [4-1:0] node40067;
	wire [4-1:0] node40068;
	wire [4-1:0] node40069;
	wire [4-1:0] node40070;
	wire [4-1:0] node40073;
	wire [4-1:0] node40076;
	wire [4-1:0] node40077;
	wire [4-1:0] node40078;
	wire [4-1:0] node40081;
	wire [4-1:0] node40084;
	wire [4-1:0] node40085;
	wire [4-1:0] node40089;
	wire [4-1:0] node40090;
	wire [4-1:0] node40091;
	wire [4-1:0] node40092;
	wire [4-1:0] node40095;
	wire [4-1:0] node40098;
	wire [4-1:0] node40099;
	wire [4-1:0] node40100;
	wire [4-1:0] node40103;
	wire [4-1:0] node40106;
	wire [4-1:0] node40107;
	wire [4-1:0] node40110;
	wire [4-1:0] node40113;
	wire [4-1:0] node40114;
	wire [4-1:0] node40115;
	wire [4-1:0] node40118;
	wire [4-1:0] node40121;
	wire [4-1:0] node40122;
	wire [4-1:0] node40124;
	wire [4-1:0] node40127;
	wire [4-1:0] node40130;
	wire [4-1:0] node40131;
	wire [4-1:0] node40132;
	wire [4-1:0] node40133;
	wire [4-1:0] node40135;
	wire [4-1:0] node40138;
	wire [4-1:0] node40139;
	wire [4-1:0] node40143;
	wire [4-1:0] node40144;
	wire [4-1:0] node40145;
	wire [4-1:0] node40149;
	wire [4-1:0] node40150;
	wire [4-1:0] node40154;
	wire [4-1:0] node40155;
	wire [4-1:0] node40156;
	wire [4-1:0] node40157;
	wire [4-1:0] node40160;
	wire [4-1:0] node40163;
	wire [4-1:0] node40164;
	wire [4-1:0] node40165;
	wire [4-1:0] node40168;
	wire [4-1:0] node40171;
	wire [4-1:0] node40172;
	wire [4-1:0] node40175;
	wire [4-1:0] node40178;
	wire [4-1:0] node40179;
	wire [4-1:0] node40180;
	wire [4-1:0] node40182;
	wire [4-1:0] node40183;
	wire [4-1:0] node40186;
	wire [4-1:0] node40188;
	wire [4-1:0] node40191;
	wire [4-1:0] node40192;
	wire [4-1:0] node40193;
	wire [4-1:0] node40196;
	wire [4-1:0] node40199;
	wire [4-1:0] node40200;
	wire [4-1:0] node40204;
	wire [4-1:0] node40205;
	wire [4-1:0] node40206;
	wire [4-1:0] node40208;
	wire [4-1:0] node40211;
	wire [4-1:0] node40213;
	wire [4-1:0] node40214;
	wire [4-1:0] node40217;
	wire [4-1:0] node40220;
	wire [4-1:0] node40222;
	wire [4-1:0] node40224;
	wire [4-1:0] node40225;
	wire [4-1:0] node40228;
	wire [4-1:0] node40231;
	wire [4-1:0] node40232;
	wire [4-1:0] node40233;
	wire [4-1:0] node40234;
	wire [4-1:0] node40235;
	wire [4-1:0] node40236;
	wire [4-1:0] node40239;
	wire [4-1:0] node40242;
	wire [4-1:0] node40243;
	wire [4-1:0] node40244;
	wire [4-1:0] node40247;
	wire [4-1:0] node40250;
	wire [4-1:0] node40253;
	wire [4-1:0] node40254;
	wire [4-1:0] node40255;
	wire [4-1:0] node40257;
	wire [4-1:0] node40258;
	wire [4-1:0] node40261;
	wire [4-1:0] node40264;
	wire [4-1:0] node40265;
	wire [4-1:0] node40268;
	wire [4-1:0] node40271;
	wire [4-1:0] node40272;
	wire [4-1:0] node40273;
	wire [4-1:0] node40274;
	wire [4-1:0] node40277;
	wire [4-1:0] node40280;
	wire [4-1:0] node40282;
	wire [4-1:0] node40285;
	wire [4-1:0] node40286;
	wire [4-1:0] node40289;
	wire [4-1:0] node40292;
	wire [4-1:0] node40293;
	wire [4-1:0] node40294;
	wire [4-1:0] node40295;
	wire [4-1:0] node40296;
	wire [4-1:0] node40299;
	wire [4-1:0] node40302;
	wire [4-1:0] node40303;
	wire [4-1:0] node40306;
	wire [4-1:0] node40309;
	wire [4-1:0] node40310;
	wire [4-1:0] node40311;
	wire [4-1:0] node40314;
	wire [4-1:0] node40317;
	wire [4-1:0] node40318;
	wire [4-1:0] node40321;
	wire [4-1:0] node40324;
	wire [4-1:0] node40325;
	wire [4-1:0] node40326;
	wire [4-1:0] node40327;
	wire [4-1:0] node40329;
	wire [4-1:0] node40332;
	wire [4-1:0] node40333;
	wire [4-1:0] node40336;
	wire [4-1:0] node40339;
	wire [4-1:0] node40340;
	wire [4-1:0] node40341;
	wire [4-1:0] node40344;
	wire [4-1:0] node40347;
	wire [4-1:0] node40348;
	wire [4-1:0] node40349;
	wire [4-1:0] node40352;
	wire [4-1:0] node40356;
	wire [4-1:0] node40357;
	wire [4-1:0] node40358;
	wire [4-1:0] node40361;
	wire [4-1:0] node40364;
	wire [4-1:0] node40365;
	wire [4-1:0] node40367;
	wire [4-1:0] node40369;
	wire [4-1:0] node40372;
	wire [4-1:0] node40373;
	wire [4-1:0] node40376;
	wire [4-1:0] node40379;
	wire [4-1:0] node40380;
	wire [4-1:0] node40381;
	wire [4-1:0] node40382;
	wire [4-1:0] node40383;
	wire [4-1:0] node40384;
	wire [4-1:0] node40387;
	wire [4-1:0] node40390;
	wire [4-1:0] node40391;
	wire [4-1:0] node40395;
	wire [4-1:0] node40396;
	wire [4-1:0] node40397;
	wire [4-1:0] node40398;
	wire [4-1:0] node40401;
	wire [4-1:0] node40404;
	wire [4-1:0] node40405;
	wire [4-1:0] node40409;
	wire [4-1:0] node40410;
	wire [4-1:0] node40411;
	wire [4-1:0] node40414;
	wire [4-1:0] node40415;
	wire [4-1:0] node40419;
	wire [4-1:0] node40420;
	wire [4-1:0] node40421;
	wire [4-1:0] node40424;
	wire [4-1:0] node40427;
	wire [4-1:0] node40429;
	wire [4-1:0] node40432;
	wire [4-1:0] node40433;
	wire [4-1:0] node40434;
	wire [4-1:0] node40435;
	wire [4-1:0] node40436;
	wire [4-1:0] node40439;
	wire [4-1:0] node40442;
	wire [4-1:0] node40445;
	wire [4-1:0] node40446;
	wire [4-1:0] node40448;
	wire [4-1:0] node40450;
	wire [4-1:0] node40453;
	wire [4-1:0] node40455;
	wire [4-1:0] node40456;
	wire [4-1:0] node40459;
	wire [4-1:0] node40462;
	wire [4-1:0] node40463;
	wire [4-1:0] node40464;
	wire [4-1:0] node40467;
	wire [4-1:0] node40470;
	wire [4-1:0] node40471;
	wire [4-1:0] node40474;
	wire [4-1:0] node40477;
	wire [4-1:0] node40478;
	wire [4-1:0] node40479;
	wire [4-1:0] node40480;
	wire [4-1:0] node40481;
	wire [4-1:0] node40484;
	wire [4-1:0] node40487;
	wire [4-1:0] node40489;
	wire [4-1:0] node40492;
	wire [4-1:0] node40493;
	wire [4-1:0] node40494;
	wire [4-1:0] node40498;
	wire [4-1:0] node40499;
	wire [4-1:0] node40502;
	wire [4-1:0] node40505;
	wire [4-1:0] node40506;
	wire [4-1:0] node40507;
	wire [4-1:0] node40508;
	wire [4-1:0] node40511;
	wire [4-1:0] node40514;
	wire [4-1:0] node40516;
	wire [4-1:0] node40519;
	wire [4-1:0] node40520;
	wire [4-1:0] node40521;
	wire [4-1:0] node40524;
	wire [4-1:0] node40527;
	wire [4-1:0] node40528;
	wire [4-1:0] node40531;
	wire [4-1:0] node40534;
	wire [4-1:0] node40535;
	wire [4-1:0] node40536;
	wire [4-1:0] node40537;
	wire [4-1:0] node40538;
	wire [4-1:0] node40539;
	wire [4-1:0] node40540;
	wire [4-1:0] node40541;
	wire [4-1:0] node40542;
	wire [4-1:0] node40544;
	wire [4-1:0] node40547;
	wire [4-1:0] node40550;
	wire [4-1:0] node40551;
	wire [4-1:0] node40552;
	wire [4-1:0] node40557;
	wire [4-1:0] node40558;
	wire [4-1:0] node40559;
	wire [4-1:0] node40560;
	wire [4-1:0] node40565;
	wire [4-1:0] node40566;
	wire [4-1:0] node40570;
	wire [4-1:0] node40571;
	wire [4-1:0] node40573;
	wire [4-1:0] node40574;
	wire [4-1:0] node40577;
	wire [4-1:0] node40580;
	wire [4-1:0] node40581;
	wire [4-1:0] node40582;
	wire [4-1:0] node40585;
	wire [4-1:0] node40588;
	wire [4-1:0] node40589;
	wire [4-1:0] node40593;
	wire [4-1:0] node40594;
	wire [4-1:0] node40595;
	wire [4-1:0] node40598;
	wire [4-1:0] node40601;
	wire [4-1:0] node40602;
	wire [4-1:0] node40603;
	wire [4-1:0] node40604;
	wire [4-1:0] node40608;
	wire [4-1:0] node40609;
	wire [4-1:0] node40613;
	wire [4-1:0] node40614;
	wire [4-1:0] node40618;
	wire [4-1:0] node40619;
	wire [4-1:0] node40620;
	wire [4-1:0] node40621;
	wire [4-1:0] node40624;
	wire [4-1:0] node40627;
	wire [4-1:0] node40628;
	wire [4-1:0] node40629;
	wire [4-1:0] node40631;
	wire [4-1:0] node40632;
	wire [4-1:0] node40635;
	wire [4-1:0] node40638;
	wire [4-1:0] node40639;
	wire [4-1:0] node40642;
	wire [4-1:0] node40645;
	wire [4-1:0] node40646;
	wire [4-1:0] node40649;
	wire [4-1:0] node40652;
	wire [4-1:0] node40653;
	wire [4-1:0] node40654;
	wire [4-1:0] node40656;
	wire [4-1:0] node40659;
	wire [4-1:0] node40661;
	wire [4-1:0] node40664;
	wire [4-1:0] node40665;
	wire [4-1:0] node40667;
	wire [4-1:0] node40670;
	wire [4-1:0] node40672;
	wire [4-1:0] node40675;
	wire [4-1:0] node40676;
	wire [4-1:0] node40677;
	wire [4-1:0] node40678;
	wire [4-1:0] node40679;
	wire [4-1:0] node40681;
	wire [4-1:0] node40682;
	wire [4-1:0] node40683;
	wire [4-1:0] node40686;
	wire [4-1:0] node40690;
	wire [4-1:0] node40691;
	wire [4-1:0] node40694;
	wire [4-1:0] node40697;
	wire [4-1:0] node40698;
	wire [4-1:0] node40699;
	wire [4-1:0] node40701;
	wire [4-1:0] node40704;
	wire [4-1:0] node40705;
	wire [4-1:0] node40709;
	wire [4-1:0] node40710;
	wire [4-1:0] node40711;
	wire [4-1:0] node40714;
	wire [4-1:0] node40717;
	wire [4-1:0] node40718;
	wire [4-1:0] node40721;
	wire [4-1:0] node40724;
	wire [4-1:0] node40725;
	wire [4-1:0] node40726;
	wire [4-1:0] node40727;
	wire [4-1:0] node40731;
	wire [4-1:0] node40732;
	wire [4-1:0] node40736;
	wire [4-1:0] node40737;
	wire [4-1:0] node40738;
	wire [4-1:0] node40742;
	wire [4-1:0] node40743;
	wire [4-1:0] node40747;
	wire [4-1:0] node40748;
	wire [4-1:0] node40749;
	wire [4-1:0] node40750;
	wire [4-1:0] node40751;
	wire [4-1:0] node40752;
	wire [4-1:0] node40753;
	wire [4-1:0] node40756;
	wire [4-1:0] node40760;
	wire [4-1:0] node40761;
	wire [4-1:0] node40764;
	wire [4-1:0] node40767;
	wire [4-1:0] node40768;
	wire [4-1:0] node40771;
	wire [4-1:0] node40774;
	wire [4-1:0] node40775;
	wire [4-1:0] node40776;
	wire [4-1:0] node40779;
	wire [4-1:0] node40782;
	wire [4-1:0] node40783;
	wire [4-1:0] node40786;
	wire [4-1:0] node40789;
	wire [4-1:0] node40790;
	wire [4-1:0] node40791;
	wire [4-1:0] node40794;
	wire [4-1:0] node40797;
	wire [4-1:0] node40798;
	wire [4-1:0] node40801;
	wire [4-1:0] node40804;
	wire [4-1:0] node40805;
	wire [4-1:0] node40806;
	wire [4-1:0] node40807;
	wire [4-1:0] node40808;
	wire [4-1:0] node40809;
	wire [4-1:0] node40810;
	wire [4-1:0] node40814;
	wire [4-1:0] node40815;
	wire [4-1:0] node40819;
	wire [4-1:0] node40820;
	wire [4-1:0] node40821;
	wire [4-1:0] node40825;
	wire [4-1:0] node40826;
	wire [4-1:0] node40830;
	wire [4-1:0] node40831;
	wire [4-1:0] node40832;
	wire [4-1:0] node40833;
	wire [4-1:0] node40836;
	wire [4-1:0] node40839;
	wire [4-1:0] node40840;
	wire [4-1:0] node40843;
	wire [4-1:0] node40846;
	wire [4-1:0] node40847;
	wire [4-1:0] node40849;
	wire [4-1:0] node40852;
	wire [4-1:0] node40853;
	wire [4-1:0] node40856;
	wire [4-1:0] node40859;
	wire [4-1:0] node40860;
	wire [4-1:0] node40861;
	wire [4-1:0] node40862;
	wire [4-1:0] node40863;
	wire [4-1:0] node40864;
	wire [4-1:0] node40867;
	wire [4-1:0] node40870;
	wire [4-1:0] node40872;
	wire [4-1:0] node40875;
	wire [4-1:0] node40876;
	wire [4-1:0] node40877;
	wire [4-1:0] node40878;
	wire [4-1:0] node40882;
	wire [4-1:0] node40883;
	wire [4-1:0] node40887;
	wire [4-1:0] node40889;
	wire [4-1:0] node40892;
	wire [4-1:0] node40893;
	wire [4-1:0] node40896;
	wire [4-1:0] node40899;
	wire [4-1:0] node40900;
	wire [4-1:0] node40901;
	wire [4-1:0] node40903;
	wire [4-1:0] node40904;
	wire [4-1:0] node40906;
	wire [4-1:0] node40909;
	wire [4-1:0] node40910;
	wire [4-1:0] node40914;
	wire [4-1:0] node40915;
	wire [4-1:0] node40918;
	wire [4-1:0] node40921;
	wire [4-1:0] node40922;
	wire [4-1:0] node40923;
	wire [4-1:0] node40925;
	wire [4-1:0] node40926;
	wire [4-1:0] node40929;
	wire [4-1:0] node40932;
	wire [4-1:0] node40933;
	wire [4-1:0] node40934;
	wire [4-1:0] node40938;
	wire [4-1:0] node40939;
	wire [4-1:0] node40942;
	wire [4-1:0] node40945;
	wire [4-1:0] node40946;
	wire [4-1:0] node40949;
	wire [4-1:0] node40952;
	wire [4-1:0] node40953;
	wire [4-1:0] node40954;
	wire [4-1:0] node40955;
	wire [4-1:0] node40956;
	wire [4-1:0] node40958;
	wire [4-1:0] node40961;
	wire [4-1:0] node40963;
	wire [4-1:0] node40966;
	wire [4-1:0] node40967;
	wire [4-1:0] node40969;
	wire [4-1:0] node40972;
	wire [4-1:0] node40974;
	wire [4-1:0] node40977;
	wire [4-1:0] node40978;
	wire [4-1:0] node40979;
	wire [4-1:0] node40980;
	wire [4-1:0] node40984;
	wire [4-1:0] node40985;
	wire [4-1:0] node40989;
	wire [4-1:0] node40990;
	wire [4-1:0] node40991;
	wire [4-1:0] node40995;
	wire [4-1:0] node40996;
	wire [4-1:0] node41000;
	wire [4-1:0] node41001;
	wire [4-1:0] node41002;
	wire [4-1:0] node41003;
	wire [4-1:0] node41006;
	wire [4-1:0] node41009;
	wire [4-1:0] node41010;
	wire [4-1:0] node41011;
	wire [4-1:0] node41012;
	wire [4-1:0] node41015;
	wire [4-1:0] node41019;
	wire [4-1:0] node41020;
	wire [4-1:0] node41023;
	wire [4-1:0] node41026;
	wire [4-1:0] node41027;
	wire [4-1:0] node41030;
	wire [4-1:0] node41033;
	wire [4-1:0] node41034;
	wire [4-1:0] node41035;
	wire [4-1:0] node41036;
	wire [4-1:0] node41037;
	wire [4-1:0] node41038;
	wire [4-1:0] node41040;
	wire [4-1:0] node41043;
	wire [4-1:0] node41045;
	wire [4-1:0] node41048;
	wire [4-1:0] node41049;
	wire [4-1:0] node41051;
	wire [4-1:0] node41054;
	wire [4-1:0] node41056;
	wire [4-1:0] node41059;
	wire [4-1:0] node41060;
	wire [4-1:0] node41061;
	wire [4-1:0] node41062;
	wire [4-1:0] node41063;
	wire [4-1:0] node41066;
	wire [4-1:0] node41069;
	wire [4-1:0] node41070;
	wire [4-1:0] node41073;
	wire [4-1:0] node41076;
	wire [4-1:0] node41077;
	wire [4-1:0] node41078;
	wire [4-1:0] node41079;
	wire [4-1:0] node41082;
	wire [4-1:0] node41085;
	wire [4-1:0] node41086;
	wire [4-1:0] node41089;
	wire [4-1:0] node41092;
	wire [4-1:0] node41093;
	wire [4-1:0] node41094;
	wire [4-1:0] node41095;
	wire [4-1:0] node41098;
	wire [4-1:0] node41103;
	wire [4-1:0] node41104;
	wire [4-1:0] node41105;
	wire [4-1:0] node41106;
	wire [4-1:0] node41109;
	wire [4-1:0] node41112;
	wire [4-1:0] node41113;
	wire [4-1:0] node41114;
	wire [4-1:0] node41117;
	wire [4-1:0] node41120;
	wire [4-1:0] node41121;
	wire [4-1:0] node41122;
	wire [4-1:0] node41125;
	wire [4-1:0] node41128;
	wire [4-1:0] node41130;
	wire [4-1:0] node41131;
	wire [4-1:0] node41134;
	wire [4-1:0] node41137;
	wire [4-1:0] node41138;
	wire [4-1:0] node41139;
	wire [4-1:0] node41142;
	wire [4-1:0] node41145;
	wire [4-1:0] node41146;
	wire [4-1:0] node41149;
	wire [4-1:0] node41152;
	wire [4-1:0] node41153;
	wire [4-1:0] node41154;
	wire [4-1:0] node41155;
	wire [4-1:0] node41156;
	wire [4-1:0] node41157;
	wire [4-1:0] node41158;
	wire [4-1:0] node41160;
	wire [4-1:0] node41163;
	wire [4-1:0] node41165;
	wire [4-1:0] node41168;
	wire [4-1:0] node41169;
	wire [4-1:0] node41171;
	wire [4-1:0] node41174;
	wire [4-1:0] node41175;
	wire [4-1:0] node41179;
	wire [4-1:0] node41180;
	wire [4-1:0] node41182;
	wire [4-1:0] node41185;
	wire [4-1:0] node41186;
	wire [4-1:0] node41187;
	wire [4-1:0] node41190;
	wire [4-1:0] node41193;
	wire [4-1:0] node41195;
	wire [4-1:0] node41196;
	wire [4-1:0] node41200;
	wire [4-1:0] node41201;
	wire [4-1:0] node41202;
	wire [4-1:0] node41203;
	wire [4-1:0] node41204;
	wire [4-1:0] node41207;
	wire [4-1:0] node41208;
	wire [4-1:0] node41212;
	wire [4-1:0] node41213;
	wire [4-1:0] node41214;
	wire [4-1:0] node41218;
	wire [4-1:0] node41219;
	wire [4-1:0] node41223;
	wire [4-1:0] node41224;
	wire [4-1:0] node41226;
	wire [4-1:0] node41229;
	wire [4-1:0] node41230;
	wire [4-1:0] node41233;
	wire [4-1:0] node41236;
	wire [4-1:0] node41237;
	wire [4-1:0] node41239;
	wire [4-1:0] node41240;
	wire [4-1:0] node41242;
	wire [4-1:0] node41245;
	wire [4-1:0] node41248;
	wire [4-1:0] node41249;
	wire [4-1:0] node41250;
	wire [4-1:0] node41252;
	wire [4-1:0] node41255;
	wire [4-1:0] node41258;
	wire [4-1:0] node41259;
	wire [4-1:0] node41262;
	wire [4-1:0] node41265;
	wire [4-1:0] node41266;
	wire [4-1:0] node41267;
	wire [4-1:0] node41268;
	wire [4-1:0] node41269;
	wire [4-1:0] node41273;
	wire [4-1:0] node41276;
	wire [4-1:0] node41277;
	wire [4-1:0] node41279;
	wire [4-1:0] node41282;
	wire [4-1:0] node41283;
	wire [4-1:0] node41284;
	wire [4-1:0] node41288;
	wire [4-1:0] node41289;
	wire [4-1:0] node41292;
	wire [4-1:0] node41295;
	wire [4-1:0] node41296;
	wire [4-1:0] node41297;
	wire [4-1:0] node41298;
	wire [4-1:0] node41303;
	wire [4-1:0] node41304;
	wire [4-1:0] node41308;
	wire [4-1:0] node41309;
	wire [4-1:0] node41310;
	wire [4-1:0] node41311;
	wire [4-1:0] node41312;
	wire [4-1:0] node41316;
	wire [4-1:0] node41317;
	wire [4-1:0] node41321;
	wire [4-1:0] node41322;
	wire [4-1:0] node41323;
	wire [4-1:0] node41327;
	wire [4-1:0] node41328;
	wire [4-1:0] node41332;
	wire [4-1:0] node41333;
	wire [4-1:0] node41334;
	wire [4-1:0] node41337;
	wire [4-1:0] node41340;
	wire [4-1:0] node41341;
	wire [4-1:0] node41342;
	wire [4-1:0] node41343;
	wire [4-1:0] node41345;
	wire [4-1:0] node41348;
	wire [4-1:0] node41349;
	wire [4-1:0] node41352;
	wire [4-1:0] node41355;
	wire [4-1:0] node41356;
	wire [4-1:0] node41359;
	wire [4-1:0] node41362;
	wire [4-1:0] node41363;
	wire [4-1:0] node41364;
	wire [4-1:0] node41365;
	wire [4-1:0] node41369;
	wire [4-1:0] node41370;
	wire [4-1:0] node41374;
	wire [4-1:0] node41376;
	wire [4-1:0] node41378;
	wire [4-1:0] node41380;
	wire [4-1:0] node41383;
	wire [4-1:0] node41384;
	wire [4-1:0] node41385;
	wire [4-1:0] node41386;
	wire [4-1:0] node41387;
	wire [4-1:0] node41388;
	wire [4-1:0] node41392;
	wire [4-1:0] node41393;
	wire [4-1:0] node41397;
	wire [4-1:0] node41398;
	wire [4-1:0] node41399;
	wire [4-1:0] node41403;
	wire [4-1:0] node41405;
	wire [4-1:0] node41408;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41411;
	wire [4-1:0] node41412;
	wire [4-1:0] node41413;
	wire [4-1:0] node41414;
	wire [4-1:0] node41415;
	wire [4-1:0] node41418;
	wire [4-1:0] node41422;
	wire [4-1:0] node41423;
	wire [4-1:0] node41425;
	wire [4-1:0] node41428;
	wire [4-1:0] node41429;
	wire [4-1:0] node41433;
	wire [4-1:0] node41434;
	wire [4-1:0] node41438;
	wire [4-1:0] node41439;
	wire [4-1:0] node41440;
	wire [4-1:0] node41442;
	wire [4-1:0] node41445;
	wire [4-1:0] node41446;
	wire [4-1:0] node41449;
	wire [4-1:0] node41452;
	wire [4-1:0] node41453;
	wire [4-1:0] node41455;
	wire [4-1:0] node41458;
	wire [4-1:0] node41459;
	wire [4-1:0] node41460;
	wire [4-1:0] node41465;
	wire [4-1:0] node41466;
	wire [4-1:0] node41467;
	wire [4-1:0] node41468;
	wire [4-1:0] node41469;
	wire [4-1:0] node41472;
	wire [4-1:0] node41475;
	wire [4-1:0] node41476;
	wire [4-1:0] node41479;
	wire [4-1:0] node41482;
	wire [4-1:0] node41483;
	wire [4-1:0] node41486;
	wire [4-1:0] node41489;
	wire [4-1:0] node41490;
	wire [4-1:0] node41491;
	wire [4-1:0] node41495;
	wire [4-1:0] node41496;
	wire [4-1:0] node41499;
	wire [4-1:0] node41502;
	wire [4-1:0] node41503;
	wire [4-1:0] node41504;
	wire [4-1:0] node41505;
	wire [4-1:0] node41507;
	wire [4-1:0] node41510;
	wire [4-1:0] node41511;
	wire [4-1:0] node41513;
	wire [4-1:0] node41516;
	wire [4-1:0] node41518;
	wire [4-1:0] node41521;
	wire [4-1:0] node41522;
	wire [4-1:0] node41523;
	wire [4-1:0] node41524;
	wire [4-1:0] node41527;
	wire [4-1:0] node41530;
	wire [4-1:0] node41532;
	wire [4-1:0] node41535;
	wire [4-1:0] node41536;
	wire [4-1:0] node41539;
	wire [4-1:0] node41542;
	wire [4-1:0] node41543;
	wire [4-1:0] node41544;
	wire [4-1:0] node41545;
	wire [4-1:0] node41548;
	wire [4-1:0] node41551;
	wire [4-1:0] node41552;
	wire [4-1:0] node41555;
	wire [4-1:0] node41558;
	wire [4-1:0] node41559;
	wire [4-1:0] node41560;
	wire [4-1:0] node41563;
	wire [4-1:0] node41566;
	wire [4-1:0] node41567;
	wire [4-1:0] node41568;
	wire [4-1:0] node41571;
	wire [4-1:0] node41574;
	wire [4-1:0] node41575;
	wire [4-1:0] node41578;
	wire [4-1:0] node41581;
	wire [4-1:0] node41582;
	wire [4-1:0] node41583;
	wire [4-1:0] node41587;
	wire [4-1:0] node41588;
	wire [4-1:0] node41592;
	wire [4-1:0] node41593;
	wire [4-1:0] node41594;
	wire [4-1:0] node41595;
	wire [4-1:0] node41596;
	wire [4-1:0] node41597;
	wire [4-1:0] node41598;
	wire [4-1:0] node41599;
	wire [4-1:0] node41600;
	wire [4-1:0] node41601;
	wire [4-1:0] node41603;
	wire [4-1:0] node41605;
	wire [4-1:0] node41606;
	wire [4-1:0] node41610;
	wire [4-1:0] node41612;
	wire [4-1:0] node41614;
	wire [4-1:0] node41617;
	wire [4-1:0] node41618;
	wire [4-1:0] node41619;
	wire [4-1:0] node41620;
	wire [4-1:0] node41622;
	wire [4-1:0] node41626;
	wire [4-1:0] node41627;
	wire [4-1:0] node41631;
	wire [4-1:0] node41632;
	wire [4-1:0] node41633;
	wire [4-1:0] node41636;
	wire [4-1:0] node41639;
	wire [4-1:0] node41640;
	wire [4-1:0] node41643;
	wire [4-1:0] node41646;
	wire [4-1:0] node41647;
	wire [4-1:0] node41648;
	wire [4-1:0] node41651;
	wire [4-1:0] node41654;
	wire [4-1:0] node41655;
	wire [4-1:0] node41656;
	wire [4-1:0] node41658;
	wire [4-1:0] node41661;
	wire [4-1:0] node41663;
	wire [4-1:0] node41666;
	wire [4-1:0] node41668;
	wire [4-1:0] node41671;
	wire [4-1:0] node41672;
	wire [4-1:0] node41673;
	wire [4-1:0] node41674;
	wire [4-1:0] node41675;
	wire [4-1:0] node41677;
	wire [4-1:0] node41680;
	wire [4-1:0] node41681;
	wire [4-1:0] node41682;
	wire [4-1:0] node41685;
	wire [4-1:0] node41689;
	wire [4-1:0] node41690;
	wire [4-1:0] node41691;
	wire [4-1:0] node41694;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41701;
	wire [4-1:0] node41704;
	wire [4-1:0] node41705;
	wire [4-1:0] node41706;
	wire [4-1:0] node41707;
	wire [4-1:0] node41710;
	wire [4-1:0] node41713;
	wire [4-1:0] node41714;
	wire [4-1:0] node41717;
	wire [4-1:0] node41720;
	wire [4-1:0] node41721;
	wire [4-1:0] node41722;
	wire [4-1:0] node41724;
	wire [4-1:0] node41727;
	wire [4-1:0] node41728;
	wire [4-1:0] node41731;
	wire [4-1:0] node41734;
	wire [4-1:0] node41735;
	wire [4-1:0] node41736;
	wire [4-1:0] node41739;
	wire [4-1:0] node41743;
	wire [4-1:0] node41744;
	wire [4-1:0] node41745;
	wire [4-1:0] node41747;
	wire [4-1:0] node41749;
	wire [4-1:0] node41752;
	wire [4-1:0] node41753;
	wire [4-1:0] node41755;
	wire [4-1:0] node41758;
	wire [4-1:0] node41761;
	wire [4-1:0] node41762;
	wire [4-1:0] node41763;
	wire [4-1:0] node41766;
	wire [4-1:0] node41768;
	wire [4-1:0] node41771;
	wire [4-1:0] node41772;
	wire [4-1:0] node41775;
	wire [4-1:0] node41777;
	wire [4-1:0] node41780;
	wire [4-1:0] node41781;
	wire [4-1:0] node41782;
	wire [4-1:0] node41783;
	wire [4-1:0] node41784;
	wire [4-1:0] node41785;
	wire [4-1:0] node41786;
	wire [4-1:0] node41787;
	wire [4-1:0] node41790;
	wire [4-1:0] node41793;
	wire [4-1:0] node41794;
	wire [4-1:0] node41797;
	wire [4-1:0] node41800;
	wire [4-1:0] node41802;
	wire [4-1:0] node41803;
	wire [4-1:0] node41806;
	wire [4-1:0] node41809;
	wire [4-1:0] node41810;
	wire [4-1:0] node41811;
	wire [4-1:0] node41812;
	wire [4-1:0] node41815;
	wire [4-1:0] node41819;
	wire [4-1:0] node41820;
	wire [4-1:0] node41821;
	wire [4-1:0] node41824;
	wire [4-1:0] node41828;
	wire [4-1:0] node41829;
	wire [4-1:0] node41831;
	wire [4-1:0] node41832;
	wire [4-1:0] node41833;
	wire [4-1:0] node41836;
	wire [4-1:0] node41840;
	wire [4-1:0] node41842;
	wire [4-1:0] node41843;
	wire [4-1:0] node41845;
	wire [4-1:0] node41848;
	wire [4-1:0] node41850;
	wire [4-1:0] node41853;
	wire [4-1:0] node41854;
	wire [4-1:0] node41855;
	wire [4-1:0] node41856;
	wire [4-1:0] node41857;
	wire [4-1:0] node41859;
	wire [4-1:0] node41863;
	wire [4-1:0] node41865;
	wire [4-1:0] node41866;
	wire [4-1:0] node41869;
	wire [4-1:0] node41872;
	wire [4-1:0] node41874;
	wire [4-1:0] node41876;
	wire [4-1:0] node41877;
	wire [4-1:0] node41881;
	wire [4-1:0] node41882;
	wire [4-1:0] node41884;
	wire [4-1:0] node41885;
	wire [4-1:0] node41886;
	wire [4-1:0] node41890;
	wire [4-1:0] node41891;
	wire [4-1:0] node41895;
	wire [4-1:0] node41896;
	wire [4-1:0] node41898;
	wire [4-1:0] node41901;
	wire [4-1:0] node41902;
	wire [4-1:0] node41904;
	wire [4-1:0] node41907;
	wire [4-1:0] node41909;
	wire [4-1:0] node41912;
	wire [4-1:0] node41913;
	wire [4-1:0] node41914;
	wire [4-1:0] node41915;
	wire [4-1:0] node41917;
	wire [4-1:0] node41918;
	wire [4-1:0] node41922;
	wire [4-1:0] node41924;
	wire [4-1:0] node41925;
	wire [4-1:0] node41929;
	wire [4-1:0] node41930;
	wire [4-1:0] node41932;
	wire [4-1:0] node41933;
	wire [4-1:0] node41937;
	wire [4-1:0] node41938;
	wire [4-1:0] node41940;
	wire [4-1:0] node41944;
	wire [4-1:0] node41945;
	wire [4-1:0] node41946;
	wire [4-1:0] node41947;
	wire [4-1:0] node41948;
	wire [4-1:0] node41949;
	wire [4-1:0] node41953;
	wire [4-1:0] node41954;
	wire [4-1:0] node41958;
	wire [4-1:0] node41960;
	wire [4-1:0] node41961;
	wire [4-1:0] node41965;
	wire [4-1:0] node41966;
	wire [4-1:0] node41967;
	wire [4-1:0] node41972;
	wire [4-1:0] node41973;
	wire [4-1:0] node41974;
	wire [4-1:0] node41976;
	wire [4-1:0] node41979;
	wire [4-1:0] node41981;
	wire [4-1:0] node41984;
	wire [4-1:0] node41986;
	wire [4-1:0] node41988;
	wire [4-1:0] node41991;
	wire [4-1:0] node41992;
	wire [4-1:0] node41993;
	wire [4-1:0] node41994;
	wire [4-1:0] node41995;
	wire [4-1:0] node41996;
	wire [4-1:0] node41997;
	wire [4-1:0] node42000;
	wire [4-1:0] node42003;
	wire [4-1:0] node42004;
	wire [4-1:0] node42007;
	wire [4-1:0] node42008;
	wire [4-1:0] node42009;
	wire [4-1:0] node42013;
	wire [4-1:0] node42015;
	wire [4-1:0] node42018;
	wire [4-1:0] node42019;
	wire [4-1:0] node42020;
	wire [4-1:0] node42021;
	wire [4-1:0] node42024;
	wire [4-1:0] node42027;
	wire [4-1:0] node42028;
	wire [4-1:0] node42029;
	wire [4-1:0] node42033;
	wire [4-1:0] node42035;
	wire [4-1:0] node42038;
	wire [4-1:0] node42039;
	wire [4-1:0] node42040;
	wire [4-1:0] node42041;
	wire [4-1:0] node42045;
	wire [4-1:0] node42047;
	wire [4-1:0] node42050;
	wire [4-1:0] node42051;
	wire [4-1:0] node42055;
	wire [4-1:0] node42056;
	wire [4-1:0] node42057;
	wire [4-1:0] node42058;
	wire [4-1:0] node42059;
	wire [4-1:0] node42061;
	wire [4-1:0] node42064;
	wire [4-1:0] node42066;
	wire [4-1:0] node42069;
	wire [4-1:0] node42070;
	wire [4-1:0] node42074;
	wire [4-1:0] node42075;
	wire [4-1:0] node42076;
	wire [4-1:0] node42078;
	wire [4-1:0] node42083;
	wire [4-1:0] node42084;
	wire [4-1:0] node42086;
	wire [4-1:0] node42089;
	wire [4-1:0] node42090;
	wire [4-1:0] node42093;
	wire [4-1:0] node42094;
	wire [4-1:0] node42098;
	wire [4-1:0] node42099;
	wire [4-1:0] node42100;
	wire [4-1:0] node42101;
	wire [4-1:0] node42102;
	wire [4-1:0] node42103;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42111;
	wire [4-1:0] node42112;
	wire [4-1:0] node42116;
	wire [4-1:0] node42117;
	wire [4-1:0] node42118;
	wire [4-1:0] node42120;
	wire [4-1:0] node42124;
	wire [4-1:0] node42125;
	wire [4-1:0] node42127;
	wire [4-1:0] node42130;
	wire [4-1:0] node42131;
	wire [4-1:0] node42135;
	wire [4-1:0] node42136;
	wire [4-1:0] node42137;
	wire [4-1:0] node42138;
	wire [4-1:0] node42140;
	wire [4-1:0] node42145;
	wire [4-1:0] node42146;
	wire [4-1:0] node42147;
	wire [4-1:0] node42148;
	wire [4-1:0] node42151;
	wire [4-1:0] node42155;
	wire [4-1:0] node42156;
	wire [4-1:0] node42158;
	wire [4-1:0] node42162;
	wire [4-1:0] node42163;
	wire [4-1:0] node42164;
	wire [4-1:0] node42165;
	wire [4-1:0] node42167;
	wire [4-1:0] node42168;
	wire [4-1:0] node42171;
	wire [4-1:0] node42174;
	wire [4-1:0] node42175;
	wire [4-1:0] node42177;
	wire [4-1:0] node42180;
	wire [4-1:0] node42183;
	wire [4-1:0] node42184;
	wire [4-1:0] node42186;
	wire [4-1:0] node42187;
	wire [4-1:0] node42191;
	wire [4-1:0] node42192;
	wire [4-1:0] node42195;
	wire [4-1:0] node42198;
	wire [4-1:0] node42199;
	wire [4-1:0] node42200;
	wire [4-1:0] node42201;
	wire [4-1:0] node42202;
	wire [4-1:0] node42205;
	wire [4-1:0] node42209;
	wire [4-1:0] node42210;
	wire [4-1:0] node42213;
	wire [4-1:0] node42216;
	wire [4-1:0] node42217;
	wire [4-1:0] node42218;
	wire [4-1:0] node42220;
	wire [4-1:0] node42224;
	wire [4-1:0] node42226;
	wire [4-1:0] node42229;
	wire [4-1:0] node42230;
	wire [4-1:0] node42231;
	wire [4-1:0] node42232;
	wire [4-1:0] node42233;
	wire [4-1:0] node42234;
	wire [4-1:0] node42237;
	wire [4-1:0] node42239;
	wire [4-1:0] node42242;
	wire [4-1:0] node42243;
	wire [4-1:0] node42245;
	wire [4-1:0] node42246;
	wire [4-1:0] node42251;
	wire [4-1:0] node42252;
	wire [4-1:0] node42253;
	wire [4-1:0] node42254;
	wire [4-1:0] node42258;
	wire [4-1:0] node42260;
	wire [4-1:0] node42263;
	wire [4-1:0] node42264;
	wire [4-1:0] node42267;
	wire [4-1:0] node42269;
	wire [4-1:0] node42272;
	wire [4-1:0] node42273;
	wire [4-1:0] node42274;
	wire [4-1:0] node42276;
	wire [4-1:0] node42277;
	wire [4-1:0] node42279;
	wire [4-1:0] node42282;
	wire [4-1:0] node42284;
	wire [4-1:0] node42287;
	wire [4-1:0] node42288;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42295;
	wire [4-1:0] node42296;
	wire [4-1:0] node42299;
	wire [4-1:0] node42302;
	wire [4-1:0] node42303;
	wire [4-1:0] node42304;
	wire [4-1:0] node42305;
	wire [4-1:0] node42306;
	wire [4-1:0] node42310;
	wire [4-1:0] node42314;
	wire [4-1:0] node42315;
	wire [4-1:0] node42316;
	wire [4-1:0] node42319;
	wire [4-1:0] node42322;
	wire [4-1:0] node42323;
	wire [4-1:0] node42326;
	wire [4-1:0] node42329;
	wire [4-1:0] node42330;
	wire [4-1:0] node42331;
	wire [4-1:0] node42332;
	wire [4-1:0] node42333;
	wire [4-1:0] node42336;
	wire [4-1:0] node42340;
	wire [4-1:0] node42341;
	wire [4-1:0] node42342;
	wire [4-1:0] node42345;
	wire [4-1:0] node42349;
	wire [4-1:0] node42350;
	wire [4-1:0] node42351;
	wire [4-1:0] node42352;
	wire [4-1:0] node42353;
	wire [4-1:0] node42356;
	wire [4-1:0] node42359;
	wire [4-1:0] node42361;
	wire [4-1:0] node42365;
	wire [4-1:0] node42366;
	wire [4-1:0] node42367;
	wire [4-1:0] node42370;
	wire [4-1:0] node42374;
	wire [4-1:0] node42375;
	wire [4-1:0] node42376;
	wire [4-1:0] node42377;
	wire [4-1:0] node42378;
	wire [4-1:0] node42379;
	wire [4-1:0] node42380;
	wire [4-1:0] node42383;
	wire [4-1:0] node42386;
	wire [4-1:0] node42387;
	wire [4-1:0] node42389;
	wire [4-1:0] node42390;
	wire [4-1:0] node42391;
	wire [4-1:0] node42395;
	wire [4-1:0] node42398;
	wire [4-1:0] node42399;
	wire [4-1:0] node42400;
	wire [4-1:0] node42401;
	wire [4-1:0] node42404;
	wire [4-1:0] node42408;
	wire [4-1:0] node42409;
	wire [4-1:0] node42410;
	wire [4-1:0] node42413;
	wire [4-1:0] node42416;
	wire [4-1:0] node42417;
	wire [4-1:0] node42420;
	wire [4-1:0] node42423;
	wire [4-1:0] node42424;
	wire [4-1:0] node42425;
	wire [4-1:0] node42426;
	wire [4-1:0] node42430;
	wire [4-1:0] node42431;
	wire [4-1:0] node42433;
	wire [4-1:0] node42434;
	wire [4-1:0] node42437;
	wire [4-1:0] node42440;
	wire [4-1:0] node42441;
	wire [4-1:0] node42442;
	wire [4-1:0] node42445;
	wire [4-1:0] node42448;
	wire [4-1:0] node42449;
	wire [4-1:0] node42452;
	wire [4-1:0] node42455;
	wire [4-1:0] node42456;
	wire [4-1:0] node42457;
	wire [4-1:0] node42458;
	wire [4-1:0] node42461;
	wire [4-1:0] node42464;
	wire [4-1:0] node42465;
	wire [4-1:0] node42469;
	wire [4-1:0] node42470;
	wire [4-1:0] node42471;
	wire [4-1:0] node42475;
	wire [4-1:0] node42476;
	wire [4-1:0] node42480;
	wire [4-1:0] node42481;
	wire [4-1:0] node42482;
	wire [4-1:0] node42483;
	wire [4-1:0] node42484;
	wire [4-1:0] node42487;
	wire [4-1:0] node42490;
	wire [4-1:0] node42491;
	wire [4-1:0] node42493;
	wire [4-1:0] node42496;
	wire [4-1:0] node42498;
	wire [4-1:0] node42500;
	wire [4-1:0] node42503;
	wire [4-1:0] node42504;
	wire [4-1:0] node42505;
	wire [4-1:0] node42506;
	wire [4-1:0] node42509;
	wire [4-1:0] node42512;
	wire [4-1:0] node42513;
	wire [4-1:0] node42516;
	wire [4-1:0] node42519;
	wire [4-1:0] node42520;
	wire [4-1:0] node42521;
	wire [4-1:0] node42524;
	wire [4-1:0] node42527;
	wire [4-1:0] node42528;
	wire [4-1:0] node42531;
	wire [4-1:0] node42532;
	wire [4-1:0] node42536;
	wire [4-1:0] node42537;
	wire [4-1:0] node42538;
	wire [4-1:0] node42539;
	wire [4-1:0] node42541;
	wire [4-1:0] node42544;
	wire [4-1:0] node42546;
	wire [4-1:0] node42549;
	wire [4-1:0] node42551;
	wire [4-1:0] node42552;
	wire [4-1:0] node42555;
	wire [4-1:0] node42558;
	wire [4-1:0] node42559;
	wire [4-1:0] node42561;
	wire [4-1:0] node42562;
	wire [4-1:0] node42563;
	wire [4-1:0] node42567;
	wire [4-1:0] node42568;
	wire [4-1:0] node42572;
	wire [4-1:0] node42573;
	wire [4-1:0] node42575;
	wire [4-1:0] node42578;
	wire [4-1:0] node42579;
	wire [4-1:0] node42583;
	wire [4-1:0] node42584;
	wire [4-1:0] node42585;
	wire [4-1:0] node42586;
	wire [4-1:0] node42587;
	wire [4-1:0] node42588;
	wire [4-1:0] node42593;
	wire [4-1:0] node42594;
	wire [4-1:0] node42598;
	wire [4-1:0] node42599;
	wire [4-1:0] node42601;
	wire [4-1:0] node42602;
	wire [4-1:0] node42603;
	wire [4-1:0] node42608;
	wire [4-1:0] node42609;
	wire [4-1:0] node42611;
	wire [4-1:0] node42612;
	wire [4-1:0] node42617;
	wire [4-1:0] node42618;
	wire [4-1:0] node42619;
	wire [4-1:0] node42620;
	wire [4-1:0] node42623;
	wire [4-1:0] node42626;
	wire [4-1:0] node42627;
	wire [4-1:0] node42629;
	wire [4-1:0] node42631;
	wire [4-1:0] node42632;
	wire [4-1:0] node42635;
	wire [4-1:0] node42638;
	wire [4-1:0] node42639;
	wire [4-1:0] node42640;
	wire [4-1:0] node42641;
	wire [4-1:0] node42644;
	wire [4-1:0] node42647;
	wire [4-1:0] node42649;
	wire [4-1:0] node42652;
	wire [4-1:0] node42653;
	wire [4-1:0] node42655;
	wire [4-1:0] node42659;
	wire [4-1:0] node42660;
	wire [4-1:0] node42661;
	wire [4-1:0] node42662;
	wire [4-1:0] node42663;
	wire [4-1:0] node42665;
	wire [4-1:0] node42668;
	wire [4-1:0] node42669;
	wire [4-1:0] node42672;
	wire [4-1:0] node42675;
	wire [4-1:0] node42677;
	wire [4-1:0] node42680;
	wire [4-1:0] node42681;
	wire [4-1:0] node42684;
	wire [4-1:0] node42687;
	wire [4-1:0] node42688;
	wire [4-1:0] node42689;
	wire [4-1:0] node42690;
	wire [4-1:0] node42693;
	wire [4-1:0] node42696;
	wire [4-1:0] node42698;
	wire [4-1:0] node42701;
	wire [4-1:0] node42702;
	wire [4-1:0] node42705;
	wire [4-1:0] node42708;
	wire [4-1:0] node42709;
	wire [4-1:0] node42710;
	wire [4-1:0] node42711;
	wire [4-1:0] node42712;
	wire [4-1:0] node42713;
	wire [4-1:0] node42717;
	wire [4-1:0] node42718;
	wire [4-1:0] node42719;
	wire [4-1:0] node42720;
	wire [4-1:0] node42721;
	wire [4-1:0] node42725;
	wire [4-1:0] node42726;
	wire [4-1:0] node42729;
	wire [4-1:0] node42733;
	wire [4-1:0] node42734;
	wire [4-1:0] node42735;
	wire [4-1:0] node42738;
	wire [4-1:0] node42741;
	wire [4-1:0] node42743;
	wire [4-1:0] node42746;
	wire [4-1:0] node42748;
	wire [4-1:0] node42749;
	wire [4-1:0] node42753;
	wire [4-1:0] node42754;
	wire [4-1:0] node42755;
	wire [4-1:0] node42756;
	wire [4-1:0] node42760;
	wire [4-1:0] node42761;
	wire [4-1:0] node42764;
	wire [4-1:0] node42767;
	wire [4-1:0] node42768;
	wire [4-1:0] node42769;
	wire [4-1:0] node42771;
	wire [4-1:0] node42776;
	wire [4-1:0] node42777;
	wire [4-1:0] node42778;
	wire [4-1:0] node42779;
	wire [4-1:0] node42780;
	wire [4-1:0] node42781;
	wire [4-1:0] node42784;
	wire [4-1:0] node42787;
	wire [4-1:0] node42788;
	wire [4-1:0] node42791;
	wire [4-1:0] node42794;
	wire [4-1:0] node42796;
	wire [4-1:0] node42799;
	wire [4-1:0] node42801;
	wire [4-1:0] node42802;
	wire [4-1:0] node42806;
	wire [4-1:0] node42807;
	wire [4-1:0] node42808;
	wire [4-1:0] node42809;
	wire [4-1:0] node42813;
	wire [4-1:0] node42814;
	wire [4-1:0] node42815;
	wire [4-1:0] node42816;
	wire [4-1:0] node42819;
	wire [4-1:0] node42822;
	wire [4-1:0] node42823;
	wire [4-1:0] node42824;
	wire [4-1:0] node42827;
	wire [4-1:0] node42830;
	wire [4-1:0] node42831;
	wire [4-1:0] node42835;
	wire [4-1:0] node42836;
	wire [4-1:0] node42839;
	wire [4-1:0] node42842;
	wire [4-1:0] node42843;
	wire [4-1:0] node42845;
	wire [4-1:0] node42849;
	wire [4-1:0] node42850;
	wire [4-1:0] node42851;
	wire [4-1:0] node42852;
	wire [4-1:0] node42853;
	wire [4-1:0] node42854;
	wire [4-1:0] node42855;
	wire [4-1:0] node42856;
	wire [4-1:0] node42857;
	wire [4-1:0] node42859;
	wire [4-1:0] node42862;
	wire [4-1:0] node42863;
	wire [4-1:0] node42866;
	wire [4-1:0] node42869;
	wire [4-1:0] node42870;
	wire [4-1:0] node42871;
	wire [4-1:0] node42872;
	wire [4-1:0] node42876;
	wire [4-1:0] node42878;
	wire [4-1:0] node42881;
	wire [4-1:0] node42882;
	wire [4-1:0] node42885;
	wire [4-1:0] node42888;
	wire [4-1:0] node42889;
	wire [4-1:0] node42890;
	wire [4-1:0] node42893;
	wire [4-1:0] node42896;
	wire [4-1:0] node42898;
	wire [4-1:0] node42901;
	wire [4-1:0] node42902;
	wire [4-1:0] node42903;
	wire [4-1:0] node42904;
	wire [4-1:0] node42905;
	wire [4-1:0] node42906;
	wire [4-1:0] node42911;
	wire [4-1:0] node42913;
	wire [4-1:0] node42916;
	wire [4-1:0] node42917;
	wire [4-1:0] node42918;
	wire [4-1:0] node42921;
	wire [4-1:0] node42924;
	wire [4-1:0] node42925;
	wire [4-1:0] node42928;
	wire [4-1:0] node42931;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42938;
	wire [4-1:0] node42939;
	wire [4-1:0] node42940;
	wire [4-1:0] node42941;
	wire [4-1:0] node42942;
	wire [4-1:0] node42943;
	wire [4-1:0] node42947;
	wire [4-1:0] node42948;
	wire [4-1:0] node42952;
	wire [4-1:0] node42953;
	wire [4-1:0] node42956;
	wire [4-1:0] node42959;
	wire [4-1:0] node42960;
	wire [4-1:0] node42963;
	wire [4-1:0] node42966;
	wire [4-1:0] node42967;
	wire [4-1:0] node42968;
	wire [4-1:0] node42971;
	wire [4-1:0] node42974;
	wire [4-1:0] node42975;
	wire [4-1:0] node42976;
	wire [4-1:0] node42977;
	wire [4-1:0] node42978;
	wire [4-1:0] node42981;
	wire [4-1:0] node42984;
	wire [4-1:0] node42985;
	wire [4-1:0] node42989;
	wire [4-1:0] node42990;
	wire [4-1:0] node42991;
	wire [4-1:0] node42994;
	wire [4-1:0] node42997;
	wire [4-1:0] node42999;
	wire [4-1:0] node43002;
	wire [4-1:0] node43003;
	wire [4-1:0] node43004;
	wire [4-1:0] node43005;
	wire [4-1:0] node43010;
	wire [4-1:0] node43011;
	wire [4-1:0] node43014;
	wire [4-1:0] node43017;
	wire [4-1:0] node43018;
	wire [4-1:0] node43019;
	wire [4-1:0] node43020;
	wire [4-1:0] node43024;
	wire [4-1:0] node43025;
	wire [4-1:0] node43029;
	wire [4-1:0] node43030;
	wire [4-1:0] node43032;
	wire [4-1:0] node43035;
	wire [4-1:0] node43036;
	wire [4-1:0] node43040;
	wire [4-1:0] node43041;
	wire [4-1:0] node43042;
	wire [4-1:0] node43043;
	wire [4-1:0] node43046;
	wire [4-1:0] node43049;
	wire [4-1:0] node43050;
	wire [4-1:0] node43051;
	wire [4-1:0] node43052;
	wire [4-1:0] node43053;
	wire [4-1:0] node43056;
	wire [4-1:0] node43059;
	wire [4-1:0] node43060;
	wire [4-1:0] node43063;
	wire [4-1:0] node43066;
	wire [4-1:0] node43067;
	wire [4-1:0] node43068;
	wire [4-1:0] node43071;
	wire [4-1:0] node43074;
	wire [4-1:0] node43075;
	wire [4-1:0] node43078;
	wire [4-1:0] node43081;
	wire [4-1:0] node43082;
	wire [4-1:0] node43083;
	wire [4-1:0] node43086;
	wire [4-1:0] node43089;
	wire [4-1:0] node43090;
	wire [4-1:0] node43091;
	wire [4-1:0] node43094;
	wire [4-1:0] node43097;
	wire [4-1:0] node43099;
	wire [4-1:0] node43100;
	wire [4-1:0] node43103;
	wire [4-1:0] node43106;
	wire [4-1:0] node43107;
	wire [4-1:0] node43108;
	wire [4-1:0] node43111;
	wire [4-1:0] node43114;
	wire [4-1:0] node43115;
	wire [4-1:0] node43116;
	wire [4-1:0] node43117;
	wire [4-1:0] node43118;
	wire [4-1:0] node43122;
	wire [4-1:0] node43123;
	wire [4-1:0] node43124;
	wire [4-1:0] node43126;
	wire [4-1:0] node43129;
	wire [4-1:0] node43130;
	wire [4-1:0] node43134;
	wire [4-1:0] node43135;
	wire [4-1:0] node43136;
	wire [4-1:0] node43139;
	wire [4-1:0] node43143;
	wire [4-1:0] node43144;
	wire [4-1:0] node43145;
	wire [4-1:0] node43146;
	wire [4-1:0] node43149;
	wire [4-1:0] node43152;
	wire [4-1:0] node43153;
	wire [4-1:0] node43156;
	wire [4-1:0] node43159;
	wire [4-1:0] node43160;
	wire [4-1:0] node43161;
	wire [4-1:0] node43165;
	wire [4-1:0] node43167;
	wire [4-1:0] node43170;
	wire [4-1:0] node43171;
	wire [4-1:0] node43172;
	wire [4-1:0] node43173;
	wire [4-1:0] node43176;
	wire [4-1:0] node43179;
	wire [4-1:0] node43180;
	wire [4-1:0] node43181;
	wire [4-1:0] node43184;
	wire [4-1:0] node43187;
	wire [4-1:0] node43188;
	wire [4-1:0] node43191;
	wire [4-1:0] node43194;
	wire [4-1:0] node43195;
	wire [4-1:0] node43196;
	wire [4-1:0] node43199;
	wire [4-1:0] node43202;
	wire [4-1:0] node43203;
	wire [4-1:0] node43206;
	wire [4-1:0] node43209;
	wire [4-1:0] node43210;
	wire [4-1:0] node43211;
	wire [4-1:0] node43212;
	wire [4-1:0] node43213;
	wire [4-1:0] node43214;
	wire [4-1:0] node43215;
	wire [4-1:0] node43216;
	wire [4-1:0] node43217;
	wire [4-1:0] node43220;
	wire [4-1:0] node43223;
	wire [4-1:0] node43224;
	wire [4-1:0] node43227;
	wire [4-1:0] node43230;
	wire [4-1:0] node43231;
	wire [4-1:0] node43232;
	wire [4-1:0] node43236;
	wire [4-1:0] node43237;
	wire [4-1:0] node43240;
	wire [4-1:0] node43243;
	wire [4-1:0] node43244;
	wire [4-1:0] node43245;
	wire [4-1:0] node43247;
	wire [4-1:0] node43248;
	wire [4-1:0] node43251;
	wire [4-1:0] node43254;
	wire [4-1:0] node43257;
	wire [4-1:0] node43258;
	wire [4-1:0] node43259;
	wire [4-1:0] node43262;
	wire [4-1:0] node43266;
	wire [4-1:0] node43267;
	wire [4-1:0] node43268;
	wire [4-1:0] node43269;
	wire [4-1:0] node43270;
	wire [4-1:0] node43273;
	wire [4-1:0] node43276;
	wire [4-1:0] node43277;
	wire [4-1:0] node43281;
	wire [4-1:0] node43282;
	wire [4-1:0] node43283;
	wire [4-1:0] node43286;
	wire [4-1:0] node43289;
	wire [4-1:0] node43290;
	wire [4-1:0] node43293;
	wire [4-1:0] node43296;
	wire [4-1:0] node43297;
	wire [4-1:0] node43298;
	wire [4-1:0] node43300;
	wire [4-1:0] node43303;
	wire [4-1:0] node43304;
	wire [4-1:0] node43305;
	wire [4-1:0] node43308;
	wire [4-1:0] node43311;
	wire [4-1:0] node43312;
	wire [4-1:0] node43316;
	wire [4-1:0] node43317;
	wire [4-1:0] node43319;
	wire [4-1:0] node43321;
	wire [4-1:0] node43324;
	wire [4-1:0] node43325;
	wire [4-1:0] node43326;
	wire [4-1:0] node43331;
	wire [4-1:0] node43332;
	wire [4-1:0] node43333;
	wire [4-1:0] node43334;
	wire [4-1:0] node43335;
	wire [4-1:0] node43336;
	wire [4-1:0] node43340;
	wire [4-1:0] node43341;
	wire [4-1:0] node43344;
	wire [4-1:0] node43347;
	wire [4-1:0] node43348;
	wire [4-1:0] node43349;
	wire [4-1:0] node43350;
	wire [4-1:0] node43354;
	wire [4-1:0] node43358;
	wire [4-1:0] node43359;
	wire [4-1:0] node43360;
	wire [4-1:0] node43363;
	wire [4-1:0] node43366;
	wire [4-1:0] node43367;
	wire [4-1:0] node43369;
	wire [4-1:0] node43372;
	wire [4-1:0] node43373;
	wire [4-1:0] node43374;
	wire [4-1:0] node43377;
	wire [4-1:0] node43380;
	wire [4-1:0] node43381;
	wire [4-1:0] node43385;
	wire [4-1:0] node43386;
	wire [4-1:0] node43389;
	wire [4-1:0] node43392;
	wire [4-1:0] node43393;
	wire [4-1:0] node43394;
	wire [4-1:0] node43395;
	wire [4-1:0] node43398;
	wire [4-1:0] node43401;
	wire [4-1:0] node43402;
	wire [4-1:0] node43405;
	wire [4-1:0] node43408;
	wire [4-1:0] node43409;
	wire [4-1:0] node43410;
	wire [4-1:0] node43411;
	wire [4-1:0] node43412;
	wire [4-1:0] node43413;
	wire [4-1:0] node43414;
	wire [4-1:0] node43417;
	wire [4-1:0] node43420;
	wire [4-1:0] node43421;
	wire [4-1:0] node43425;
	wire [4-1:0] node43426;
	wire [4-1:0] node43429;
	wire [4-1:0] node43432;
	wire [4-1:0] node43433;
	wire [4-1:0] node43436;
	wire [4-1:0] node43439;
	wire [4-1:0] node43440;
	wire [4-1:0] node43441;
	wire [4-1:0] node43444;
	wire [4-1:0] node43447;
	wire [4-1:0] node43448;
	wire [4-1:0] node43451;
	wire [4-1:0] node43454;
	wire [4-1:0] node43455;
	wire [4-1:0] node43456;
	wire [4-1:0] node43459;
	wire [4-1:0] node43462;
	wire [4-1:0] node43463;
	wire [4-1:0] node43466;
	wire [4-1:0] node43469;
	wire [4-1:0] node43470;
	wire [4-1:0] node43471;
	wire [4-1:0] node43472;
	wire [4-1:0] node43473;
	wire [4-1:0] node43477;
	wire [4-1:0] node43478;
	wire [4-1:0] node43483;
	wire [4-1:0] node43484;
	wire [4-1:0] node43485;
	wire [4-1:0] node43486;
	wire [4-1:0] node43490;
	wire [4-1:0] node43491;
	wire [4-1:0] node43496;
	wire [4-1:0] node43497;
	wire [4-1:0] node43498;
	wire [4-1:0] node43499;
	wire [4-1:0] node43500;
	wire [4-1:0] node43501;
	wire [4-1:0] node43502;
	wire [4-1:0] node43503;
	wire [4-1:0] node43504;
	wire [4-1:0] node43507;
	wire [4-1:0] node43510;
	wire [4-1:0] node43511;
	wire [4-1:0] node43512;
	wire [4-1:0] node43515;
	wire [4-1:0] node43518;
	wire [4-1:0] node43519;
	wire [4-1:0] node43520;
	wire [4-1:0] node43524;
	wire [4-1:0] node43526;
	wire [4-1:0] node43529;
	wire [4-1:0] node43530;
	wire [4-1:0] node43531;
	wire [4-1:0] node43534;
	wire [4-1:0] node43537;
	wire [4-1:0] node43538;
	wire [4-1:0] node43539;
	wire [4-1:0] node43541;
	wire [4-1:0] node43542;
	wire [4-1:0] node43545;
	wire [4-1:0] node43548;
	wire [4-1:0] node43549;
	wire [4-1:0] node43552;
	wire [4-1:0] node43555;
	wire [4-1:0] node43556;
	wire [4-1:0] node43557;
	wire [4-1:0] node43558;
	wire [4-1:0] node43562;
	wire [4-1:0] node43563;
	wire [4-1:0] node43568;
	wire [4-1:0] node43569;
	wire [4-1:0] node43570;
	wire [4-1:0] node43572;
	wire [4-1:0] node43575;
	wire [4-1:0] node43577;
	wire [4-1:0] node43580;
	wire [4-1:0] node43581;
	wire [4-1:0] node43583;
	wire [4-1:0] node43586;
	wire [4-1:0] node43588;
	wire [4-1:0] node43591;
	wire [4-1:0] node43592;
	wire [4-1:0] node43593;
	wire [4-1:0] node43594;
	wire [4-1:0] node43595;
	wire [4-1:0] node43596;
	wire [4-1:0] node43597;
	wire [4-1:0] node43598;
	wire [4-1:0] node43601;
	wire [4-1:0] node43604;
	wire [4-1:0] node43605;
	wire [4-1:0] node43609;
	wire [4-1:0] node43611;
	wire [4-1:0] node43613;
	wire [4-1:0] node43616;
	wire [4-1:0] node43617;
	wire [4-1:0] node43620;
	wire [4-1:0] node43623;
	wire [4-1:0] node43624;
	wire [4-1:0] node43625;
	wire [4-1:0] node43626;
	wire [4-1:0] node43629;
	wire [4-1:0] node43632;
	wire [4-1:0] node43633;
	wire [4-1:0] node43634;
	wire [4-1:0] node43638;
	wire [4-1:0] node43639;
	wire [4-1:0] node43643;
	wire [4-1:0] node43644;
	wire [4-1:0] node43647;
	wire [4-1:0] node43650;
	wire [4-1:0] node43651;
	wire [4-1:0] node43654;
	wire [4-1:0] node43657;
	wire [4-1:0] node43658;
	wire [4-1:0] node43661;
	wire [4-1:0] node43664;
	wire [4-1:0] node43665;
	wire [4-1:0] node43666;
	wire [4-1:0] node43667;
	wire [4-1:0] node43668;
	wire [4-1:0] node43671;
	wire [4-1:0] node43675;
	wire [4-1:0] node43676;
	wire [4-1:0] node43677;
	wire [4-1:0] node43678;
	wire [4-1:0] node43679;
	wire [4-1:0] node43680;
	wire [4-1:0] node43683;
	wire [4-1:0] node43686;
	wire [4-1:0] node43687;
	wire [4-1:0] node43690;
	wire [4-1:0] node43693;
	wire [4-1:0] node43694;
	wire [4-1:0] node43697;
	wire [4-1:0] node43700;
	wire [4-1:0] node43701;
	wire [4-1:0] node43702;
	wire [4-1:0] node43703;
	wire [4-1:0] node43705;
	wire [4-1:0] node43708;
	wire [4-1:0] node43710;
	wire [4-1:0] node43713;
	wire [4-1:0] node43714;
	wire [4-1:0] node43716;
	wire [4-1:0] node43720;
	wire [4-1:0] node43721;
	wire [4-1:0] node43722;
	wire [4-1:0] node43725;
	wire [4-1:0] node43728;
	wire [4-1:0] node43729;
	wire [4-1:0] node43732;
	wire [4-1:0] node43733;
	wire [4-1:0] node43738;
	wire [4-1:0] node43739;
	wire [4-1:0] node43740;
	wire [4-1:0] node43744;
	wire [4-1:0] node43745;
	wire [4-1:0] node43749;
	wire [4-1:0] node43750;
	wire [4-1:0] node43751;
	wire [4-1:0] node43752;
	wire [4-1:0] node43755;
	wire [4-1:0] node43758;
	wire [4-1:0] node43759;
	wire [4-1:0] node43760;
	wire [4-1:0] node43763;
	wire [4-1:0] node43766;
	wire [4-1:0] node43767;
	wire [4-1:0] node43768;
	wire [4-1:0] node43771;
	wire [4-1:0] node43774;
	wire [4-1:0] node43775;
	wire [4-1:0] node43776;
	wire [4-1:0] node43777;
	wire [4-1:0] node43780;
	wire [4-1:0] node43783;
	wire [4-1:0] node43784;
	wire [4-1:0] node43786;
	wire [4-1:0] node43789;
	wire [4-1:0] node43791;
	wire [4-1:0] node43793;
	wire [4-1:0] node43796;
	wire [4-1:0] node43797;
	wire [4-1:0] node43798;
	wire [4-1:0] node43800;
	wire [4-1:0] node43803;
	wire [4-1:0] node43804;
	wire [4-1:0] node43808;
	wire [4-1:0] node43809;
	wire [4-1:0] node43810;
	wire [4-1:0] node43814;
	wire [4-1:0] node43815;
	wire [4-1:0] node43816;
	wire [4-1:0] node43820;
	wire [4-1:0] node43822;
	wire [4-1:0] node43825;
	wire [4-1:0] node43826;
	wire [4-1:0] node43827;
	wire [4-1:0] node43831;
	wire [4-1:0] node43832;
	wire [4-1:0] node43836;
	wire [4-1:0] node43837;
	wire [4-1:0] node43838;
	wire [4-1:0] node43839;
	wire [4-1:0] node43840;
	wire [4-1:0] node43841;
	wire [4-1:0] node43842;
	wire [4-1:0] node43843;
	wire [4-1:0] node43844;
	wire [4-1:0] node43847;
	wire [4-1:0] node43851;
	wire [4-1:0] node43852;
	wire [4-1:0] node43853;
	wire [4-1:0] node43855;
	wire [4-1:0] node43856;
	wire [4-1:0] node43859;
	wire [4-1:0] node43862;
	wire [4-1:0] node43864;
	wire [4-1:0] node43865;
	wire [4-1:0] node43868;
	wire [4-1:0] node43872;
	wire [4-1:0] node43873;
	wire [4-1:0] node43874;
	wire [4-1:0] node43878;
	wire [4-1:0] node43879;
	wire [4-1:0] node43883;
	wire [4-1:0] node43884;
	wire [4-1:0] node43885;
	wire [4-1:0] node43886;
	wire [4-1:0] node43887;
	wire [4-1:0] node43889;
	wire [4-1:0] node43890;
	wire [4-1:0] node43893;
	wire [4-1:0] node43896;
	wire [4-1:0] node43898;
	wire [4-1:0] node43899;
	wire [4-1:0] node43902;
	wire [4-1:0] node43905;
	wire [4-1:0] node43906;
	wire [4-1:0] node43908;
	wire [4-1:0] node43911;
	wire [4-1:0] node43913;
	wire [4-1:0] node43914;
	wire [4-1:0] node43917;
	wire [4-1:0] node43920;
	wire [4-1:0] node43921;
	wire [4-1:0] node43922;
	wire [4-1:0] node43925;
	wire [4-1:0] node43928;
	wire [4-1:0] node43929;
	wire [4-1:0] node43932;
	wire [4-1:0] node43935;
	wire [4-1:0] node43936;
	wire [4-1:0] node43937;
	wire [4-1:0] node43938;
	wire [4-1:0] node43939;
	wire [4-1:0] node43943;
	wire [4-1:0] node43944;
	wire [4-1:0] node43945;
	wire [4-1:0] node43949;
	wire [4-1:0] node43952;
	wire [4-1:0] node43953;
	wire [4-1:0] node43955;
	wire [4-1:0] node43956;
	wire [4-1:0] node43959;
	wire [4-1:0] node43962;
	wire [4-1:0] node43963;
	wire [4-1:0] node43965;
	wire [4-1:0] node43969;
	wire [4-1:0] node43970;
	wire [4-1:0] node43971;
	wire [4-1:0] node43973;
	wire [4-1:0] node43974;
	wire [4-1:0] node43978;
	wire [4-1:0] node43979;
	wire [4-1:0] node43981;
	wire [4-1:0] node43984;
	wire [4-1:0] node43987;
	wire [4-1:0] node43988;
	wire [4-1:0] node43989;
	wire [4-1:0] node43993;
	wire [4-1:0] node43994;
	wire [4-1:0] node43998;
	wire [4-1:0] node43999;
	wire [4-1:0] node44000;
	wire [4-1:0] node44001;
	wire [4-1:0] node44003;
	wire [4-1:0] node44006;
	wire [4-1:0] node44008;
	wire [4-1:0] node44011;
	wire [4-1:0] node44012;
	wire [4-1:0] node44014;
	wire [4-1:0] node44017;
	wire [4-1:0] node44018;
	wire [4-1:0] node44022;
	wire [4-1:0] node44023;
	wire [4-1:0] node44024;
	wire [4-1:0] node44026;
	wire [4-1:0] node44029;
	wire [4-1:0] node44030;
	wire [4-1:0] node44033;
	wire [4-1:0] node44036;
	wire [4-1:0] node44037;
	wire [4-1:0] node44038;
	wire [4-1:0] node44041;
	wire [4-1:0] node44044;
	wire [4-1:0] node44045;
	wire [4-1:0] node44048;
	wire [4-1:0] node44051;
	wire [4-1:0] node44052;
	wire [4-1:0] node44053;
	wire [4-1:0] node44057;
	wire [4-1:0] node44058;
	wire [4-1:0] node44062;
	wire [4-1:0] node44063;
	wire [4-1:0] node44064;
	wire [4-1:0] node44065;
	wire [4-1:0] node44066;
	wire [4-1:0] node44067;
	wire [4-1:0] node44071;
	wire [4-1:0] node44072;
	wire [4-1:0] node44077;
	wire [4-1:0] node44078;
	wire [4-1:0] node44082;
	wire [4-1:0] node44083;
	wire [4-1:0] node44084;
	wire [4-1:0] node44085;
	wire [4-1:0] node44086;
	wire [4-1:0] node44091;
	wire [4-1:0] node44092;
	wire [4-1:0] node44093;

	assign outp = (inp[8]) ? node27418 : node1;
		assign node1 = (inp[14]) ? node15391 : node2;
			assign node2 = (inp[6]) ? node8324 : node3;
				assign node3 = (inp[3]) ? node4163 : node4;
					assign node4 = (inp[0]) ? node1906 : node5;
						assign node5 = (inp[9]) ? node957 : node6;
							assign node6 = (inp[10]) ? node466 : node7;
								assign node7 = (inp[4]) ? node219 : node8;
									assign node8 = (inp[13]) ? node114 : node9;
										assign node9 = (inp[1]) ? node49 : node10;
											assign node10 = (inp[2]) ? node28 : node11;
												assign node11 = (inp[7]) ? node15 : node12;
													assign node12 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node15 = (inp[12]) ? node19 : node16;
														assign node16 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node19 = (inp[15]) ? node23 : node20;
															assign node20 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node23 = (inp[5]) ? 4'b0000 : node24;
																assign node24 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node28 = (inp[7]) ? node32 : node29;
													assign node29 = (inp[12]) ? 4'b0110 : 4'b0100;
													assign node32 = (inp[12]) ? node44 : node33;
														assign node33 = (inp[15]) ? node37 : node34;
															assign node34 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node37 = (inp[5]) ? node41 : node38;
																assign node38 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node44 = (inp[11]) ? 4'b0101 : node45;
															assign node45 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node49 = (inp[7]) ? node83 : node50;
												assign node50 = (inp[12]) ? node68 : node51;
													assign node51 = (inp[15]) ? node61 : node52;
														assign node52 = (inp[11]) ? 4'b0100 : node53;
															assign node53 = (inp[5]) ? node57 : node54;
																assign node54 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node57 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node61 = (inp[2]) ? node65 : node62;
															assign node62 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node65 = (inp[5]) ? 4'b0001 : 4'b0100;
													assign node68 = (inp[15]) ? node76 : node69;
														assign node69 = (inp[2]) ? node73 : node70;
															assign node70 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node73 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node76 = (inp[5]) ? node78 : 4'b0010;
															assign node78 = (inp[2]) ? 4'b0010 : node79;
																assign node79 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node83 = (inp[12]) ? node103 : node84;
													assign node84 = (inp[5]) ? node94 : node85;
														assign node85 = (inp[15]) ? node89 : node86;
															assign node86 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node89 = (inp[2]) ? 4'b0011 : node90;
																assign node90 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node94 = (inp[15]) ? node100 : node95;
															assign node95 = (inp[2]) ? node97 : 4'b0111;
																assign node97 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node100 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node103 = (inp[5]) ? 4'b0101 : node104;
														assign node104 = (inp[15]) ? node110 : node105;
															assign node105 = (inp[11]) ? node107 : 4'b0101;
																assign node107 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node110 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node114 = (inp[2]) ? node162 : node115;
											assign node115 = (inp[15]) ? node137 : node116;
												assign node116 = (inp[1]) ? node124 : node117;
													assign node117 = (inp[7]) ? node121 : node118;
														assign node118 = (inp[12]) ? 4'b0110 : 4'b0100;
														assign node121 = (inp[12]) ? 4'b0000 : 4'b0111;
													assign node124 = (inp[5]) ? node132 : node125;
														assign node125 = (inp[11]) ? node127 : 4'b0000;
															assign node127 = (inp[12]) ? 4'b0111 : node128;
																assign node128 = (inp[7]) ? 4'b0110 : 4'b0100;
														assign node132 = (inp[12]) ? node134 : 4'b0001;
															assign node134 = (inp[7]) ? 4'b0001 : 4'b0010;
												assign node137 = (inp[11]) ? node147 : node138;
													assign node138 = (inp[7]) ? node142 : node139;
														assign node139 = (inp[12]) ? 4'b0111 : 4'b0101;
														assign node142 = (inp[5]) ? node144 : 4'b0101;
															assign node144 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node147 = (inp[7]) ? node155 : node148;
														assign node148 = (inp[1]) ? node152 : node149;
															assign node149 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node152 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node155 = (inp[5]) ? node159 : node156;
															assign node156 = (inp[12]) ? 4'b0000 : 4'b0010;
															assign node159 = (inp[12]) ? 4'b0101 : 4'b0111;
											assign node162 = (inp[7]) ? node190 : node163;
												assign node163 = (inp[12]) ? node177 : node164;
													assign node164 = (inp[5]) ? node170 : node165;
														assign node165 = (inp[11]) ? node167 : 4'b0000;
															assign node167 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node170 = (inp[1]) ? 4'b0100 : node171;
															assign node171 = (inp[15]) ? node173 : 4'b0001;
																assign node173 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node177 = (inp[1]) ? node183 : node178;
														assign node178 = (inp[15]) ? node180 : 4'b0011;
															assign node180 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node183 = (inp[5]) ? node185 : 4'b0011;
															assign node185 = (inp[15]) ? 4'b0111 : node186;
																assign node186 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node190 = (inp[12]) ? node208 : node191;
													assign node191 = (inp[15]) ? node199 : node192;
														assign node192 = (inp[5]) ? node196 : node193;
															assign node193 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node196 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node199 = (inp[5]) ? node205 : node200;
															assign node200 = (inp[11]) ? 4'b0110 : node201;
																assign node201 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node205 = (inp[11]) ? 4'b0111 : 4'b0011;
													assign node208 = (inp[15]) ? node214 : node209;
														assign node209 = (inp[1]) ? node211 : 4'b0100;
															assign node211 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node214 = (inp[5]) ? 4'b0001 : node215;
															assign node215 = (inp[1]) ? 4'b0000 : 4'b0100;
									assign node219 = (inp[15]) ? node345 : node220;
										assign node220 = (inp[2]) ? node280 : node221;
											assign node221 = (inp[13]) ? node249 : node222;
												assign node222 = (inp[11]) ? node240 : node223;
													assign node223 = (inp[7]) ? node231 : node224;
														assign node224 = (inp[12]) ? 4'b0010 : node225;
															assign node225 = (inp[1]) ? node227 : 4'b0000;
																assign node227 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node231 = (inp[5]) ? node237 : node232;
															assign node232 = (inp[1]) ? node234 : 4'b0100;
																assign node234 = (inp[12]) ? 4'b0000 : 4'b0010;
															assign node237 = (inp[12]) ? 4'b0001 : 4'b0011;
													assign node240 = (inp[12]) ? node244 : node241;
														assign node241 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node244 = (inp[7]) ? node246 : 4'b0111;
															assign node246 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node249 = (inp[11]) ? node271 : node250;
													assign node250 = (inp[12]) ? node262 : node251;
														assign node251 = (inp[7]) ? node257 : node252;
															assign node252 = (inp[1]) ? node254 : 4'b0100;
																assign node254 = (inp[5]) ? 4'b0001 : 4'b0100;
															assign node257 = (inp[1]) ? node259 : 4'b0111;
																assign node259 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node262 = (inp[7]) ? node266 : node263;
															assign node263 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node266 = (inp[1]) ? node268 : 4'b0001;
																assign node268 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node271 = (inp[7]) ? 4'b0100 : node272;
														assign node272 = (inp[12]) ? 4'b0011 : node273;
															assign node273 = (inp[5]) ? node275 : 4'b0100;
																assign node275 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node280 = (inp[13]) ? node312 : node281;
												assign node281 = (inp[7]) ? node295 : node282;
													assign node282 = (inp[12]) ? node288 : node283;
														assign node283 = (inp[5]) ? node285 : 4'b0101;
															assign node285 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node288 = (inp[11]) ? 4'b0010 : node289;
															assign node289 = (inp[5]) ? 4'b0010 : node290;
																assign node290 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node295 = (inp[12]) ? node303 : node296;
														assign node296 = (inp[1]) ? node300 : node297;
															assign node297 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node300 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node303 = (inp[1]) ? node307 : node304;
															assign node304 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node307 = (inp[5]) ? node309 : 4'b0101;
																assign node309 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node312 = (inp[11]) ? node328 : node313;
													assign node313 = (inp[12]) ? node319 : node314;
														assign node314 = (inp[7]) ? node316 : 4'b0001;
															assign node316 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node319 = (inp[7]) ? node325 : node320;
															assign node320 = (inp[5]) ? 4'b0110 : node321;
																assign node321 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node325 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node328 = (inp[12]) ? node334 : node329;
														assign node329 = (inp[7]) ? node331 : 4'b0000;
															assign node331 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node334 = (inp[7]) ? node338 : node335;
															assign node335 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node338 = (inp[1]) ? node342 : node339;
																assign node339 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node342 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node345 = (inp[12]) ? node399 : node346;
											assign node346 = (inp[7]) ? node366 : node347;
												assign node347 = (inp[2]) ? node357 : node348;
													assign node348 = (inp[11]) ? 4'b0111 : node349;
														assign node349 = (inp[1]) ? node353 : node350;
															assign node350 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node353 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node357 = (inp[13]) ? 4'b0111 : node358;
														assign node358 = (inp[1]) ? node362 : node359;
															assign node359 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node362 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node366 = (inp[1]) ? node382 : node367;
													assign node367 = (inp[11]) ? node373 : node368;
														assign node368 = (inp[5]) ? node370 : 4'b0101;
															assign node370 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node373 = (inp[2]) ? 4'b0001 : node374;
															assign node374 = (inp[13]) ? node378 : node375;
																assign node375 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node378 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node382 = (inp[11]) ? node396 : node383;
														assign node383 = (inp[5]) ? node389 : node384;
															assign node384 = (inp[2]) ? 4'b0100 : node385;
																assign node385 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node389 = (inp[2]) ? node393 : node390;
																assign node390 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node393 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node396 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node399 = (inp[7]) ? node427 : node400;
												assign node400 = (inp[1]) ? node416 : node401;
													assign node401 = (inp[2]) ? node411 : node402;
														assign node402 = (inp[13]) ? node408 : node403;
															assign node403 = (inp[5]) ? 4'b0001 : node404;
																assign node404 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node408 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node411 = (inp[11]) ? 4'b0100 : node412;
															assign node412 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node416 = (inp[5]) ? 4'b0101 : node417;
														assign node417 = (inp[13]) ? node421 : node418;
															assign node418 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node421 = (inp[11]) ? node423 : 4'b0000;
																assign node423 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node427 = (inp[11]) ? node445 : node428;
													assign node428 = (inp[13]) ? node436 : node429;
														assign node429 = (inp[1]) ? node431 : 4'b0010;
															assign node431 = (inp[2]) ? 4'b0111 : node432;
																assign node432 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node436 = (inp[5]) ? node438 : 4'b0111;
															assign node438 = (inp[2]) ? node442 : node439;
																assign node439 = (inp[1]) ? 4'b0111 : 4'b0010;
																assign node442 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node445 = (inp[13]) ? node455 : node446;
														assign node446 = (inp[2]) ? node450 : node447;
															assign node447 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node450 = (inp[1]) ? 4'b0010 : node451;
																assign node451 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node455 = (inp[2]) ? node463 : node456;
															assign node456 = (inp[1]) ? node460 : node457;
																assign node457 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node460 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node463 = (inp[5]) ? 4'b0011 : 4'b0110;
								assign node466 = (inp[2]) ? node704 : node467;
									assign node467 = (inp[13]) ? node587 : node468;
										assign node468 = (inp[4]) ? node502 : node469;
											assign node469 = (inp[7]) ? node479 : node470;
												assign node470 = (inp[12]) ? node472 : 4'b0001;
													assign node472 = (inp[1]) ? node474 : 4'b0011;
														assign node474 = (inp[5]) ? node476 : 4'b0010;
															assign node476 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node479 = (inp[12]) ? node489 : node480;
													assign node480 = (inp[1]) ? node484 : node481;
														assign node481 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node484 = (inp[5]) ? 4'b0011 : node485;
															assign node485 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node489 = (inp[15]) ? node497 : node490;
														assign node490 = (inp[5]) ? node492 : 4'b0101;
															assign node492 = (inp[1]) ? node494 : 4'b0101;
																assign node494 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node497 = (inp[5]) ? 4'b0001 : node498;
															assign node498 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node502 = (inp[11]) ? node554 : node503;
												assign node503 = (inp[1]) ? node529 : node504;
													assign node504 = (inp[12]) ? node518 : node505;
														assign node505 = (inp[5]) ? node513 : node506;
															assign node506 = (inp[7]) ? node510 : node507;
																assign node507 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node510 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node513 = (inp[15]) ? node515 : 4'b0010;
																assign node515 = (inp[7]) ? 4'b0001 : 4'b0111;
														assign node518 = (inp[15]) ? node524 : node519;
															assign node519 = (inp[5]) ? 4'b0001 : node520;
																assign node520 = (inp[7]) ? 4'b0101 : 4'b0111;
															assign node524 = (inp[7]) ? 4'b0111 : node525;
																assign node525 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node529 = (inp[12]) ? node539 : node530;
														assign node530 = (inp[7]) ? node536 : node531;
															assign node531 = (inp[15]) ? node533 : 4'b0101;
																assign node533 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node536 = (inp[5]) ? 4'b0110 : 4'b0000;
														assign node539 = (inp[15]) ? node547 : node540;
															assign node540 = (inp[7]) ? node544 : node541;
																assign node541 = (inp[5]) ? 4'b0011 : 4'b0110;
																assign node544 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node547 = (inp[7]) ? node551 : node548;
																assign node548 = (inp[5]) ? 4'b0101 : 4'b0001;
																assign node551 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node554 = (inp[15]) ? node570 : node555;
													assign node555 = (inp[5]) ? node561 : node556;
														assign node556 = (inp[12]) ? node558 : 4'b0001;
															assign node558 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node561 = (inp[7]) ? node565 : node562;
															assign node562 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node565 = (inp[12]) ? 4'b0001 : node566;
																assign node566 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node570 = (inp[7]) ? node578 : node571;
														assign node571 = (inp[12]) ? node573 : 4'b0110;
															assign node573 = (inp[1]) ? node575 : 4'b0000;
																assign node575 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node578 = (inp[12]) ? node582 : node579;
															assign node579 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node582 = (inp[5]) ? node584 : 4'b0110;
																assign node584 = (inp[1]) ? 4'b0010 : 4'b0110;
										assign node587 = (inp[1]) ? node639 : node588;
											assign node588 = (inp[15]) ? node612 : node589;
												assign node589 = (inp[12]) ? node601 : node590;
													assign node590 = (inp[7]) ? node598 : node591;
														assign node591 = (inp[4]) ? node593 : 4'b0101;
															assign node593 = (inp[11]) ? node595 : 4'b0101;
																assign node595 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node598 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node601 = (inp[7]) ? node605 : node602;
														assign node602 = (inp[4]) ? 4'b0010 : 4'b0111;
														assign node605 = (inp[5]) ? node609 : node606;
															assign node606 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node609 = (inp[11]) ? 4'b0001 : 4'b0101;
												assign node612 = (inp[7]) ? node626 : node613;
													assign node613 = (inp[4]) ? node617 : node614;
														assign node614 = (inp[12]) ? 4'b0110 : 4'b0100;
														assign node617 = (inp[12]) ? node621 : node618;
															assign node618 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node621 = (inp[11]) ? 4'b0101 : node622;
																assign node622 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node626 = (inp[11]) ? node632 : node627;
														assign node627 = (inp[5]) ? 4'b0100 : node628;
															assign node628 = (inp[12]) ? 4'b0011 : 4'b0100;
														assign node632 = (inp[12]) ? node634 : 4'b0010;
															assign node634 = (inp[4]) ? node636 : 4'b0001;
																assign node636 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node639 = (inp[12]) ? node669 : node640;
												assign node640 = (inp[5]) ? node654 : node641;
													assign node641 = (inp[15]) ? node645 : node642;
														assign node642 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node645 = (inp[4]) ? node651 : node646;
															assign node646 = (inp[7]) ? 4'b0011 : node647;
																assign node647 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node651 = (inp[7]) ? 4'b0101 : 4'b0011;
													assign node654 = (inp[7]) ? node662 : node655;
														assign node655 = (inp[4]) ? node657 : 4'b0001;
															assign node657 = (inp[15]) ? node659 : 4'b0000;
																assign node659 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node662 = (inp[15]) ? 4'b0001 : node663;
															assign node663 = (inp[11]) ? 4'b0011 : node664;
																assign node664 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node669 = (inp[7]) ? node687 : node670;
													assign node670 = (inp[4]) ? node678 : node671;
														assign node671 = (inp[5]) ? 4'b0010 : node672;
															assign node672 = (inp[11]) ? 4'b0110 : node673;
																assign node673 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node678 = (inp[15]) ? node684 : node679;
															assign node679 = (inp[5]) ? 4'b0111 : node680;
																assign node680 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node684 = (inp[5]) ? 4'b0001 : 4'b0100;
													assign node687 = (inp[15]) ? node695 : node688;
														assign node688 = (inp[4]) ? node690 : 4'b0001;
															assign node690 = (inp[5]) ? node692 : 4'b0101;
																assign node692 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node695 = (inp[4]) ? node699 : node696;
															assign node696 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node699 = (inp[11]) ? node701 : 4'b0110;
																assign node701 = (inp[5]) ? 4'b0111 : 4'b0011;
									assign node704 = (inp[13]) ? node814 : node705;
										assign node705 = (inp[7]) ? node761 : node706;
											assign node706 = (inp[12]) ? node732 : node707;
												assign node707 = (inp[4]) ? node717 : node708;
													assign node708 = (inp[1]) ? node710 : 4'b0101;
														assign node710 = (inp[5]) ? 4'b0000 : node711;
															assign node711 = (inp[15]) ? node713 : 4'b0101;
																assign node713 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node717 = (inp[15]) ? node723 : node718;
														assign node718 = (inp[11]) ? node720 : 4'b0100;
															assign node720 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node723 = (inp[1]) ? node727 : node724;
															assign node724 = (inp[11]) ? 4'b0011 : 4'b0110;
															assign node727 = (inp[5]) ? node729 : 4'b0011;
																assign node729 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node732 = (inp[15]) ? node752 : node733;
													assign node733 = (inp[1]) ? node741 : node734;
														assign node734 = (inp[4]) ? node736 : 4'b0111;
															assign node736 = (inp[11]) ? 4'b0011 : node737;
																assign node737 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node741 = (inp[4]) ? node747 : node742;
															assign node742 = (inp[5]) ? node744 : 4'b0110;
																assign node744 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node747 = (inp[5]) ? 4'b0110 : node748;
																assign node748 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node752 = (inp[4]) ? node756 : node753;
														assign node753 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node756 = (inp[5]) ? node758 : 4'b0100;
															assign node758 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node761 = (inp[12]) ? node785 : node762;
												assign node762 = (inp[4]) ? node778 : node763;
													assign node763 = (inp[15]) ? node769 : node764;
														assign node764 = (inp[5]) ? node766 : 4'b0111;
															assign node766 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node769 = (inp[5]) ? node775 : node770;
															assign node770 = (inp[11]) ? 4'b0010 : node771;
																assign node771 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node775 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node778 = (inp[15]) ? node782 : node779;
														assign node779 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node782 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node785 = (inp[4]) ? node799 : node786;
													assign node786 = (inp[1]) ? node796 : node787;
														assign node787 = (inp[5]) ? node793 : node788;
															assign node788 = (inp[15]) ? 4'b0000 : node789;
																assign node789 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node793 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node796 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node799 = (inp[15]) ? node809 : node800;
														assign node800 = (inp[5]) ? node804 : node801;
															assign node801 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node804 = (inp[1]) ? node806 : 4'b0100;
																assign node806 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node809 = (inp[5]) ? node811 : 4'b0011;
															assign node811 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node814 = (inp[5]) ? node884 : node815;
											assign node815 = (inp[12]) ? node853 : node816;
												assign node816 = (inp[7]) ? node834 : node817;
													assign node817 = (inp[15]) ? node825 : node818;
														assign node818 = (inp[11]) ? node822 : node819;
															assign node819 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node822 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node825 = (inp[4]) ? node829 : node826;
															assign node826 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node829 = (inp[1]) ? 4'b0110 : node830;
																assign node830 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node834 = (inp[15]) ? node842 : node835;
														assign node835 = (inp[11]) ? node839 : node836;
															assign node836 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node839 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node842 = (inp[4]) ? node848 : node843;
															assign node843 = (inp[11]) ? 4'b0111 : node844;
																assign node844 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node848 = (inp[11]) ? node850 : 4'b0000;
																assign node850 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node853 = (inp[7]) ? node871 : node854;
													assign node854 = (inp[15]) ? node864 : node855;
														assign node855 = (inp[4]) ? node859 : node856;
															assign node856 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node859 = (inp[1]) ? node861 : 4'b0111;
																assign node861 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node864 = (inp[4]) ? node866 : 4'b0010;
															assign node866 = (inp[11]) ? 4'b0000 : node867;
																assign node867 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node871 = (inp[4]) ? node879 : node872;
														assign node872 = (inp[1]) ? node876 : node873;
															assign node873 = (inp[11]) ? 4'b0101 : 4'b0000;
															assign node876 = (inp[11]) ? 4'b0001 : 4'b0101;
														assign node879 = (inp[15]) ? 4'b0110 : node880;
															assign node880 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node884 = (inp[1]) ? node930 : node885;
												assign node885 = (inp[4]) ? node911 : node886;
													assign node886 = (inp[7]) ? node900 : node887;
														assign node887 = (inp[12]) ? node895 : node888;
															assign node888 = (inp[15]) ? node892 : node889;
																assign node889 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node892 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node895 = (inp[11]) ? 4'b0011 : node896;
																assign node896 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node900 = (inp[12]) ? node908 : node901;
															assign node901 = (inp[15]) ? node905 : node902;
																assign node902 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node905 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node908 = (inp[15]) ? 4'b0000 : 4'b0101;
													assign node911 = (inp[11]) ? node923 : node912;
														assign node912 = (inp[7]) ? node916 : node913;
															assign node913 = (inp[12]) ? 4'b0000 : 4'b0110;
															assign node916 = (inp[12]) ? node920 : node917;
																assign node917 = (inp[15]) ? 4'b0001 : 4'b0010;
																assign node920 = (inp[15]) ? 4'b0110 : 4'b0001;
														assign node923 = (inp[12]) ? node927 : node924;
															assign node924 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node927 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node930 = (inp[7]) ? node942 : node931;
													assign node931 = (inp[12]) ? node939 : node932;
														assign node932 = (inp[15]) ? node936 : node933;
															assign node933 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node936 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node939 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node942 = (inp[15]) ? node948 : node943;
														assign node943 = (inp[12]) ? node945 : 4'b0110;
															assign node945 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node948 = (inp[11]) ? node950 : 4'b0010;
															assign node950 = (inp[4]) ? node954 : node951;
																assign node951 = (inp[12]) ? 4'b0000 : 4'b0011;
																assign node954 = (inp[12]) ? 4'b0010 : 4'b0100;
							assign node957 = (inp[10]) ? node1443 : node958;
								assign node958 = (inp[13]) ? node1196 : node959;
									assign node959 = (inp[2]) ? node1081 : node960;
										assign node960 = (inp[5]) ? node1014 : node961;
											assign node961 = (inp[12]) ? node981 : node962;
												assign node962 = (inp[7]) ? node972 : node963;
													assign node963 = (inp[15]) ? node965 : 4'b0001;
														assign node965 = (inp[1]) ? node969 : node966;
															assign node966 = (inp[4]) ? 4'b0011 : 4'b0001;
															assign node969 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node972 = (inp[15]) ? node974 : 4'b0011;
														assign node974 = (inp[4]) ? node978 : node975;
															assign node975 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node978 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node981 = (inp[7]) ? node997 : node982;
													assign node982 = (inp[4]) ? node990 : node983;
														assign node983 = (inp[1]) ? node985 : 4'b0011;
															assign node985 = (inp[11]) ? node987 : 4'b0010;
																assign node987 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node990 = (inp[15]) ? node994 : node991;
															assign node991 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node994 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node997 = (inp[15]) ? node1009 : node998;
														assign node998 = (inp[11]) ? node1004 : node999;
															assign node999 = (inp[4]) ? 4'b0001 : node1000;
																assign node1000 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node1004 = (inp[1]) ? 4'b0001 : node1005;
																assign node1005 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1009 = (inp[4]) ? node1011 : 4'b0001;
															assign node1011 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node1014 = (inp[1]) ? node1048 : node1015;
												assign node1015 = (inp[11]) ? node1031 : node1016;
													assign node1016 = (inp[7]) ? node1020 : node1017;
														assign node1017 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node1020 = (inp[4]) ? node1026 : node1021;
															assign node1021 = (inp[12]) ? node1023 : 4'b0110;
																assign node1023 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node1026 = (inp[15]) ? node1028 : 4'b0001;
																assign node1028 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node1031 = (inp[12]) ? node1045 : node1032;
														assign node1032 = (inp[15]) ? node1038 : node1033;
															assign node1033 = (inp[7]) ? 4'b0010 : node1034;
																assign node1034 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node1038 = (inp[7]) ? node1042 : node1039;
																assign node1039 = (inp[4]) ? 4'b0110 : 4'b0001;
																assign node1042 = (inp[4]) ? 4'b0001 : 4'b0110;
														assign node1045 = (inp[4]) ? 4'b0110 : 4'b0011;
												assign node1048 = (inp[12]) ? node1060 : node1049;
													assign node1049 = (inp[11]) ? node1051 : 4'b0101;
														assign node1051 = (inp[15]) ? node1055 : node1052;
															assign node1052 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node1055 = (inp[4]) ? node1057 : 4'b0100;
																assign node1057 = (inp[7]) ? 4'b0100 : 4'b0110;
													assign node1060 = (inp[4]) ? node1070 : node1061;
														assign node1061 = (inp[7]) ? node1067 : node1062;
															assign node1062 = (inp[11]) ? node1064 : 4'b0110;
																assign node1064 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node1067 = (inp[15]) ? 4'b0000 : 4'b0101;
														assign node1070 = (inp[11]) ? node1076 : node1071;
															assign node1071 = (inp[7]) ? 4'b0011 : node1072;
																assign node1072 = (inp[15]) ? 4'b0101 : 4'b0011;
															assign node1076 = (inp[15]) ? 4'b0010 : node1077;
																assign node1077 = (inp[7]) ? 4'b0001 : 4'b0011;
										assign node1081 = (inp[1]) ? node1131 : node1082;
											assign node1082 = (inp[4]) ? node1100 : node1083;
												assign node1083 = (inp[7]) ? node1087 : node1084;
													assign node1084 = (inp[12]) ? 4'b0111 : 4'b0101;
													assign node1087 = (inp[12]) ? node1093 : node1088;
														assign node1088 = (inp[15]) ? node1090 : 4'b0111;
															assign node1090 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node1093 = (inp[5]) ? node1097 : node1094;
															assign node1094 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node1097 = (inp[15]) ? 4'b0101 : 4'b0001;
												assign node1100 = (inp[12]) ? node1120 : node1101;
													assign node1101 = (inp[11]) ? node1109 : node1102;
														assign node1102 = (inp[7]) ? node1106 : node1103;
															assign node1103 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node1106 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1109 = (inp[15]) ? node1115 : node1110;
															assign node1110 = (inp[7]) ? 4'b0110 : node1111;
																assign node1111 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node1115 = (inp[7]) ? node1117 : 4'b0011;
																assign node1117 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node1120 = (inp[7]) ? node1126 : node1121;
														assign node1121 = (inp[15]) ? node1123 : 4'b0010;
															assign node1123 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node1126 = (inp[15]) ? 4'b0011 : node1127;
															assign node1127 = (inp[5]) ? 4'b0101 : 4'b0001;
											assign node1131 = (inp[5]) ? node1157 : node1132;
												assign node1132 = (inp[4]) ? node1144 : node1133;
													assign node1133 = (inp[12]) ? node1137 : node1134;
														assign node1134 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node1137 = (inp[7]) ? node1139 : 4'b0110;
															assign node1139 = (inp[15]) ? node1141 : 4'b0001;
																assign node1141 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node1144 = (inp[11]) ? 4'b0011 : node1145;
														assign node1145 = (inp[12]) ? node1149 : node1146;
															assign node1146 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node1149 = (inp[15]) ? node1153 : node1150;
																assign node1150 = (inp[7]) ? 4'b0100 : 4'b0011;
																assign node1153 = (inp[7]) ? 4'b0011 : 4'b0100;
												assign node1157 = (inp[12]) ? node1177 : node1158;
													assign node1158 = (inp[7]) ? node1170 : node1159;
														assign node1159 = (inp[15]) ? node1165 : node1160;
															assign node1160 = (inp[11]) ? node1162 : 4'b0001;
																assign node1162 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node1165 = (inp[4]) ? node1167 : 4'b0000;
																assign node1167 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1170 = (inp[15]) ? 4'b0001 : node1171;
															assign node1171 = (inp[11]) ? node1173 : 4'b0010;
																assign node1173 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node1177 = (inp[7]) ? node1185 : node1178;
														assign node1178 = (inp[4]) ? 4'b0110 : node1179;
															assign node1179 = (inp[15]) ? 4'b0011 : node1180;
																assign node1180 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1185 = (inp[4]) ? node1191 : node1186;
															assign node1186 = (inp[15]) ? node1188 : 4'b0000;
																assign node1188 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node1191 = (inp[15]) ? 4'b0110 : node1192;
																assign node1192 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node1196 = (inp[2]) ? node1322 : node1197;
										assign node1197 = (inp[1]) ? node1263 : node1198;
											assign node1198 = (inp[11]) ? node1226 : node1199;
												assign node1199 = (inp[15]) ? node1211 : node1200;
													assign node1200 = (inp[12]) ? node1206 : node1201;
														assign node1201 = (inp[7]) ? node1203 : 4'b0101;
															assign node1203 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node1206 = (inp[7]) ? 4'b0001 : node1207;
															assign node1207 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node1211 = (inp[4]) ? node1219 : node1212;
														assign node1212 = (inp[12]) ? node1216 : node1213;
															assign node1213 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node1216 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node1219 = (inp[12]) ? node1223 : node1220;
															assign node1220 = (inp[5]) ? 4'b0011 : 4'b0100;
															assign node1223 = (inp[7]) ? 4'b0011 : 4'b0101;
												assign node1226 = (inp[12]) ? node1248 : node1227;
													assign node1227 = (inp[15]) ? node1237 : node1228;
														assign node1228 = (inp[7]) ? node1232 : node1229;
															assign node1229 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node1232 = (inp[4]) ? 4'b0111 : node1233;
																assign node1233 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node1237 = (inp[4]) ? node1241 : node1238;
															assign node1238 = (inp[7]) ? 4'b0010 : 4'b0100;
															assign node1241 = (inp[7]) ? node1245 : node1242;
																assign node1242 = (inp[5]) ? 4'b0011 : 4'b0110;
																assign node1245 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node1248 = (inp[7]) ? node1254 : node1249;
														assign node1249 = (inp[4]) ? 4'b0010 : node1250;
															assign node1250 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1254 = (inp[5]) ? 4'b0100 : node1255;
															assign node1255 = (inp[15]) ? node1259 : node1256;
																assign node1256 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node1259 = (inp[4]) ? 4'b0010 : 4'b0001;
											assign node1263 = (inp[5]) ? node1295 : node1264;
												assign node1264 = (inp[7]) ? node1280 : node1265;
													assign node1265 = (inp[12]) ? node1269 : node1266;
														assign node1266 = (inp[4]) ? 4'b0011 : 4'b0101;
														assign node1269 = (inp[15]) ? node1275 : node1270;
															assign node1270 = (inp[4]) ? node1272 : 4'b0110;
																assign node1272 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1275 = (inp[11]) ? node1277 : 4'b0111;
																assign node1277 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node1280 = (inp[4]) ? node1288 : node1281;
														assign node1281 = (inp[12]) ? node1283 : 4'b0011;
															assign node1283 = (inp[15]) ? node1285 : 4'b0001;
																assign node1285 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node1288 = (inp[15]) ? node1292 : node1289;
															assign node1289 = (inp[12]) ? 4'b0101 : 4'b0111;
															assign node1292 = (inp[12]) ? 4'b0011 : 4'b0101;
												assign node1295 = (inp[7]) ? node1307 : node1296;
													assign node1296 = (inp[12]) ? node1302 : node1297;
														assign node1297 = (inp[15]) ? node1299 : 4'b0000;
															assign node1299 = (inp[4]) ? 4'b0010 : 4'b0001;
														assign node1302 = (inp[4]) ? 4'b0001 : node1303;
															assign node1303 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node1307 = (inp[12]) ? node1317 : node1308;
														assign node1308 = (inp[4]) ? node1314 : node1309;
															assign node1309 = (inp[15]) ? 4'b0110 : node1310;
																assign node1310 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1314 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node1317 = (inp[11]) ? 4'b0100 : node1318;
															assign node1318 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node1322 = (inp[5]) ? node1380 : node1323;
											assign node1323 = (inp[7]) ? node1351 : node1324;
												assign node1324 = (inp[12]) ? node1336 : node1325;
													assign node1325 = (inp[15]) ? node1333 : node1326;
														assign node1326 = (inp[11]) ? node1330 : node1327;
															assign node1327 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node1330 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node1333 = (inp[11]) ? 4'b0001 : 4'b0011;
													assign node1336 = (inp[15]) ? node1340 : node1337;
														assign node1337 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node1340 = (inp[4]) ? node1346 : node1341;
															assign node1341 = (inp[1]) ? 4'b0010 : node1342;
																assign node1342 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1346 = (inp[11]) ? 4'b0000 : node1347;
																assign node1347 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node1351 = (inp[12]) ? node1363 : node1352;
													assign node1352 = (inp[4]) ? node1360 : node1353;
														assign node1353 = (inp[15]) ? node1357 : node1354;
															assign node1354 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node1357 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1360 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1363 = (inp[15]) ? node1373 : node1364;
														assign node1364 = (inp[1]) ? node1368 : node1365;
															assign node1365 = (inp[4]) ? 4'b0101 : 4'b0000;
															assign node1368 = (inp[4]) ? node1370 : 4'b0101;
																assign node1370 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node1373 = (inp[4]) ? node1377 : node1374;
															assign node1374 = (inp[11]) ? 4'b0001 : 4'b0101;
															assign node1377 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node1380 = (inp[1]) ? node1410 : node1381;
												assign node1381 = (inp[15]) ? node1397 : node1382;
													assign node1382 = (inp[11]) ? node1390 : node1383;
														assign node1383 = (inp[7]) ? node1387 : node1384;
															assign node1384 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node1387 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1390 = (inp[4]) ? node1394 : node1391;
															assign node1391 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node1394 = (inp[7]) ? 4'b0001 : 4'b0111;
													assign node1397 = (inp[12]) ? node1407 : node1398;
														assign node1398 = (inp[11]) ? 4'b0001 : node1399;
															assign node1399 = (inp[7]) ? node1403 : node1400;
																assign node1400 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node1403 = (inp[4]) ? 4'b0001 : 4'b0111;
														assign node1407 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node1410 = (inp[7]) ? node1422 : node1411;
													assign node1411 = (inp[12]) ? node1417 : node1412;
														assign node1412 = (inp[11]) ? node1414 : 4'b0110;
															assign node1414 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node1417 = (inp[15]) ? 4'b0110 : node1418;
															assign node1418 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node1422 = (inp[12]) ? node1432 : node1423;
														assign node1423 = (inp[4]) ? node1429 : node1424;
															assign node1424 = (inp[11]) ? node1426 : 4'b0010;
																assign node1426 = (inp[15]) ? 4'b0011 : 4'b0111;
															assign node1429 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node1432 = (inp[11]) ? node1438 : node1433;
															assign node1433 = (inp[4]) ? node1435 : 4'b0000;
																assign node1435 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node1438 = (inp[15]) ? 4'b0000 : node1439;
																assign node1439 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node1443 = (inp[2]) ? node1675 : node1444;
									assign node1444 = (inp[13]) ? node1564 : node1445;
										assign node1445 = (inp[5]) ? node1499 : node1446;
											assign node1446 = (inp[12]) ? node1468 : node1447;
												assign node1447 = (inp[7]) ? node1459 : node1448;
													assign node1448 = (inp[4]) ? node1454 : node1449;
														assign node1449 = (inp[11]) ? node1451 : 4'b0000;
															assign node1451 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node1454 = (inp[15]) ? node1456 : 4'b0000;
															assign node1456 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node1459 = (inp[15]) ? node1461 : 4'b0010;
														assign node1461 = (inp[4]) ? node1463 : 4'b0110;
															assign node1463 = (inp[1]) ? 4'b0001 : node1464;
																assign node1464 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node1468 = (inp[7]) ? node1486 : node1469;
													assign node1469 = (inp[15]) ? node1477 : node1470;
														assign node1470 = (inp[4]) ? node1474 : node1471;
															assign node1471 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node1474 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node1477 = (inp[4]) ? node1481 : node1478;
															assign node1478 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node1481 = (inp[11]) ? node1483 : 4'b0000;
																assign node1483 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1486 = (inp[1]) ? node1494 : node1487;
														assign node1487 = (inp[4]) ? node1491 : node1488;
															assign node1488 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node1491 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node1494 = (inp[4]) ? 4'b0000 : node1495;
															assign node1495 = (inp[15]) ? 4'b0000 : 4'b0101;
											assign node1499 = (inp[1]) ? node1535 : node1500;
												assign node1500 = (inp[4]) ? node1512 : node1501;
													assign node1501 = (inp[7]) ? node1505 : node1502;
														assign node1502 = (inp[12]) ? 4'b0010 : 4'b0000;
														assign node1505 = (inp[12]) ? node1507 : 4'b0111;
															assign node1507 = (inp[15]) ? 4'b0000 : node1508;
																assign node1508 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node1512 = (inp[11]) ? node1522 : node1513;
														assign node1513 = (inp[7]) ? node1519 : node1514;
															assign node1514 = (inp[12]) ? node1516 : 4'b0110;
																assign node1516 = (inp[15]) ? 4'b0001 : 4'b0110;
															assign node1519 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node1522 = (inp[7]) ? node1528 : node1523;
															assign node1523 = (inp[12]) ? 4'b0001 : node1524;
																assign node1524 = (inp[15]) ? 4'b0111 : 4'b0001;
															assign node1528 = (inp[12]) ? node1532 : node1529;
																assign node1529 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node1532 = (inp[15]) ? 4'b0111 : 4'b0001;
												assign node1535 = (inp[7]) ? node1551 : node1536;
													assign node1536 = (inp[11]) ? node1546 : node1537;
														assign node1537 = (inp[15]) ? node1541 : node1538;
															assign node1538 = (inp[12]) ? 4'b0010 : 4'b0100;
															assign node1541 = (inp[12]) ? node1543 : 4'b0111;
																assign node1543 = (inp[4]) ? 4'b0100 : 4'b0111;
														assign node1546 = (inp[12]) ? node1548 : 4'b0101;
															assign node1548 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node1551 = (inp[12]) ? node1557 : node1552;
														assign node1552 = (inp[15]) ? node1554 : 4'b0111;
															assign node1554 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node1557 = (inp[4]) ? node1559 : 4'b0100;
															assign node1559 = (inp[15]) ? 4'b0011 : node1560;
																assign node1560 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node1564 = (inp[4]) ? node1624 : node1565;
											assign node1565 = (inp[7]) ? node1593 : node1566;
												assign node1566 = (inp[12]) ? node1578 : node1567;
													assign node1567 = (inp[15]) ? node1573 : node1568;
														assign node1568 = (inp[5]) ? node1570 : 4'b0100;
															assign node1570 = (inp[11]) ? 4'b0001 : 4'b0100;
														assign node1573 = (inp[1]) ? node1575 : 4'b0101;
															assign node1575 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node1578 = (inp[5]) ? node1588 : node1579;
														assign node1579 = (inp[1]) ? node1583 : node1580;
															assign node1580 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node1583 = (inp[11]) ? 4'b0111 : node1584;
																assign node1584 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node1588 = (inp[1]) ? 4'b0011 : node1589;
															assign node1589 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node1593 = (inp[12]) ? node1605 : node1594;
													assign node1594 = (inp[15]) ? node1600 : node1595;
														assign node1595 = (inp[5]) ? node1597 : 4'b0110;
															assign node1597 = (inp[1]) ? 4'b0010 : 4'b0111;
														assign node1600 = (inp[5]) ? node1602 : 4'b0010;
															assign node1602 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node1605 = (inp[15]) ? node1615 : node1606;
														assign node1606 = (inp[1]) ? node1612 : node1607;
															assign node1607 = (inp[5]) ? 4'b0000 : node1608;
																assign node1608 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node1612 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node1615 = (inp[5]) ? node1619 : node1616;
															assign node1616 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node1619 = (inp[1]) ? node1621 : 4'b0101;
																assign node1621 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node1624 = (inp[15]) ? node1646 : node1625;
												assign node1625 = (inp[7]) ? node1637 : node1626;
													assign node1626 = (inp[12]) ? node1630 : node1627;
														assign node1627 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node1630 = (inp[1]) ? node1632 : 4'b0011;
															assign node1632 = (inp[5]) ? 4'b0110 : node1633;
																assign node1633 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1637 = (inp[12]) ? node1641 : node1638;
														assign node1638 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node1641 = (inp[1]) ? 4'b0100 : node1642;
															assign node1642 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1646 = (inp[5]) ? node1662 : node1647;
													assign node1647 = (inp[7]) ? node1655 : node1648;
														assign node1648 = (inp[12]) ? node1652 : node1649;
															assign node1649 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node1652 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node1655 = (inp[12]) ? node1657 : 4'b0100;
															assign node1657 = (inp[1]) ? 4'b0010 : node1658;
																assign node1658 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1662 = (inp[1]) ? node1668 : node1663;
														assign node1663 = (inp[7]) ? 4'b0010 : node1664;
															assign node1664 = (inp[11]) ? 4'b0010 : 4'b0100;
														assign node1668 = (inp[12]) ? node1672 : node1669;
															assign node1669 = (inp[7]) ? 4'b0000 : 4'b0011;
															assign node1672 = (inp[7]) ? 4'b0111 : 4'b0000;
									assign node1675 = (inp[13]) ? node1777 : node1676;
										assign node1676 = (inp[1]) ? node1714 : node1677;
											assign node1677 = (inp[12]) ? node1689 : node1678;
												assign node1678 = (inp[7]) ? node1684 : node1679;
													assign node1679 = (inp[4]) ? node1681 : 4'b0100;
														assign node1681 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node1684 = (inp[15]) ? node1686 : 4'b0111;
														assign node1686 = (inp[4]) ? 4'b0101 : 4'b0011;
												assign node1689 = (inp[7]) ? node1695 : node1690;
													assign node1690 = (inp[4]) ? node1692 : 4'b0110;
														assign node1692 = (inp[15]) ? 4'b0100 : 4'b0010;
													assign node1695 = (inp[5]) ? node1703 : node1696;
														assign node1696 = (inp[4]) ? node1698 : 4'b0001;
															assign node1698 = (inp[15]) ? node1700 : 4'b0000;
																assign node1700 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1703 = (inp[11]) ? node1709 : node1704;
															assign node1704 = (inp[15]) ? node1706 : 4'b0101;
																assign node1706 = (inp[4]) ? 4'b0010 : 4'b0100;
															assign node1709 = (inp[15]) ? 4'b0100 : node1710;
																assign node1710 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node1714 = (inp[5]) ? node1744 : node1715;
												assign node1715 = (inp[11]) ? node1725 : node1716;
													assign node1716 = (inp[4]) ? 4'b0101 : node1717;
														assign node1717 = (inp[7]) ? node1721 : node1718;
															assign node1718 = (inp[12]) ? 4'b0111 : 4'b0100;
															assign node1721 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node1725 = (inp[7]) ? node1737 : node1726;
														assign node1726 = (inp[12]) ? node1734 : node1727;
															assign node1727 = (inp[15]) ? node1731 : node1728;
																assign node1728 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node1731 = (inp[4]) ? 4'b0010 : 4'b0101;
															assign node1734 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node1737 = (inp[4]) ? 4'b0100 : node1738;
															assign node1738 = (inp[12]) ? node1740 : 4'b0011;
																assign node1740 = (inp[15]) ? 4'b0101 : 4'b0000;
												assign node1744 = (inp[7]) ? node1760 : node1745;
													assign node1745 = (inp[12]) ? node1753 : node1746;
														assign node1746 = (inp[4]) ? node1750 : node1747;
															assign node1747 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node1750 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1753 = (inp[15]) ? node1757 : node1754;
															assign node1754 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node1757 = (inp[4]) ? 4'b0000 : 4'b0010;
													assign node1760 = (inp[15]) ? node1768 : node1761;
														assign node1761 = (inp[12]) ? node1765 : node1762;
															assign node1762 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node1765 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node1768 = (inp[12]) ? node1770 : 4'b0110;
															assign node1770 = (inp[11]) ? node1774 : node1771;
																assign node1771 = (inp[4]) ? 4'b0111 : 4'b0101;
																assign node1774 = (inp[4]) ? 4'b0110 : 4'b0100;
										assign node1777 = (inp[15]) ? node1839 : node1778;
											assign node1778 = (inp[12]) ? node1806 : node1779;
												assign node1779 = (inp[7]) ? node1793 : node1780;
													assign node1780 = (inp[11]) ? node1790 : node1781;
														assign node1781 = (inp[4]) ? node1787 : node1782;
															assign node1782 = (inp[5]) ? node1784 : 4'b0000;
																assign node1784 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node1787 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node1790 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node1793 = (inp[4]) ? node1801 : node1794;
														assign node1794 = (inp[11]) ? node1798 : node1795;
															assign node1795 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node1798 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node1801 = (inp[11]) ? node1803 : 4'b0011;
															assign node1803 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node1806 = (inp[7]) ? node1826 : node1807;
													assign node1807 = (inp[4]) ? node1817 : node1808;
														assign node1808 = (inp[1]) ? node1812 : node1809;
															assign node1809 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1812 = (inp[5]) ? node1814 : 4'b0010;
																assign node1814 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node1817 = (inp[5]) ? node1823 : node1818;
															assign node1818 = (inp[11]) ? node1820 : 4'b0110;
																assign node1820 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node1823 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node1826 = (inp[1]) ? node1834 : node1827;
														assign node1827 = (inp[4]) ? node1831 : node1828;
															assign node1828 = (inp[5]) ? 4'b0100 : 4'b0001;
															assign node1831 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node1834 = (inp[4]) ? 4'b0001 : node1835;
															assign node1835 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node1839 = (inp[4]) ? node1873 : node1840;
												assign node1840 = (inp[11]) ? node1858 : node1841;
													assign node1841 = (inp[5]) ? node1851 : node1842;
														assign node1842 = (inp[7]) ? node1848 : node1843;
															assign node1843 = (inp[12]) ? 4'b0011 : node1844;
																assign node1844 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node1848 = (inp[12]) ? 4'b0100 : 4'b0111;
														assign node1851 = (inp[7]) ? node1855 : node1852;
															assign node1852 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node1855 = (inp[12]) ? 4'b0001 : 4'b0011;
													assign node1858 = (inp[12]) ? node1866 : node1859;
														assign node1859 = (inp[7]) ? node1863 : node1860;
															assign node1860 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node1863 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node1866 = (inp[7]) ? 4'b0000 : node1867;
															assign node1867 = (inp[1]) ? node1869 : 4'b0010;
																assign node1869 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node1873 = (inp[5]) ? node1893 : node1874;
													assign node1874 = (inp[11]) ? node1884 : node1875;
														assign node1875 = (inp[7]) ? node1881 : node1876;
															assign node1876 = (inp[12]) ? node1878 : 4'b0111;
																assign node1878 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node1881 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node1884 = (inp[12]) ? node1890 : node1885;
															assign node1885 = (inp[1]) ? 4'b0000 : node1886;
																assign node1886 = (inp[7]) ? 4'b0001 : 4'b0011;
															assign node1890 = (inp[7]) ? 4'b0111 : 4'b0001;
													assign node1893 = (inp[12]) ? node1901 : node1894;
														assign node1894 = (inp[7]) ? 4'b0101 : node1895;
															assign node1895 = (inp[11]) ? node1897 : 4'b0111;
																assign node1897 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node1901 = (inp[7]) ? node1903 : 4'b0000;
															assign node1903 = (inp[1]) ? 4'b0011 : 4'b0111;
						assign node1906 = (inp[9]) ? node2996 : node1907;
							assign node1907 = (inp[13]) ? node2467 : node1908;
								assign node1908 = (inp[2]) ? node2196 : node1909;
									assign node1909 = (inp[1]) ? node2057 : node1910;
										assign node1910 = (inp[7]) ? node1984 : node1911;
											assign node1911 = (inp[12]) ? node1943 : node1912;
												assign node1912 = (inp[15]) ? node1926 : node1913;
													assign node1913 = (inp[11]) ? node1923 : node1914;
														assign node1914 = (inp[10]) ? node1918 : node1915;
															assign node1915 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node1918 = (inp[4]) ? node1920 : 4'b0001;
																assign node1920 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node1923 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1926 = (inp[4]) ? node1932 : node1927;
														assign node1927 = (inp[10]) ? 4'b0000 : node1928;
															assign node1928 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node1932 = (inp[5]) ? node1940 : node1933;
															assign node1933 = (inp[10]) ? node1937 : node1934;
																assign node1934 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node1937 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node1940 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node1943 = (inp[4]) ? node1967 : node1944;
													assign node1944 = (inp[5]) ? node1952 : node1945;
														assign node1945 = (inp[10]) ? node1949 : node1946;
															assign node1946 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1949 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1952 = (inp[15]) ? node1960 : node1953;
															assign node1953 = (inp[11]) ? node1957 : node1954;
																assign node1954 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node1957 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node1960 = (inp[11]) ? node1964 : node1961;
																assign node1961 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node1964 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1967 = (inp[15]) ? node1975 : node1968;
														assign node1968 = (inp[11]) ? 4'b0110 : node1969;
															assign node1969 = (inp[10]) ? 4'b0111 : node1970;
																assign node1970 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1975 = (inp[11]) ? node1979 : node1976;
															assign node1976 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node1979 = (inp[10]) ? 4'b0001 : node1980;
																assign node1980 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node1984 = (inp[12]) ? node2020 : node1985;
												assign node1985 = (inp[15]) ? node2003 : node1986;
													assign node1986 = (inp[11]) ? node1996 : node1987;
														assign node1987 = (inp[4]) ? 4'b0011 : node1988;
															assign node1988 = (inp[10]) ? node1992 : node1989;
																assign node1989 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node1992 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node1996 = (inp[5]) ? node2000 : node1997;
															assign node1997 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node2000 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node2003 = (inp[4]) ? node2011 : node2004;
														assign node2004 = (inp[11]) ? node2006 : 4'b0110;
															assign node2006 = (inp[5]) ? node2008 : 4'b0111;
																assign node2008 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node2011 = (inp[10]) ? node2017 : node2012;
															assign node2012 = (inp[5]) ? node2014 : 4'b0001;
																assign node2014 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node2017 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node2020 = (inp[15]) ? node2038 : node2021;
													assign node2021 = (inp[10]) ? node2031 : node2022;
														assign node2022 = (inp[11]) ? node2024 : 4'b0100;
															assign node2024 = (inp[4]) ? node2028 : node2025;
																assign node2025 = (inp[5]) ? 4'b0100 : 4'b0001;
																assign node2028 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node2031 = (inp[11]) ? 4'b0000 : node2032;
															assign node2032 = (inp[5]) ? 4'b0000 : node2033;
																assign node2033 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2038 = (inp[4]) ? node2048 : node2039;
														assign node2039 = (inp[5]) ? node2043 : node2040;
															assign node2040 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2043 = (inp[10]) ? node2045 : 4'b0001;
																assign node2045 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node2048 = (inp[5]) ? 4'b0110 : node2049;
															assign node2049 = (inp[11]) ? node2053 : node2050;
																assign node2050 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node2053 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node2057 = (inp[5]) ? node2133 : node2058;
											assign node2058 = (inp[15]) ? node2094 : node2059;
												assign node2059 = (inp[12]) ? node2075 : node2060;
													assign node2060 = (inp[7]) ? node2068 : node2061;
														assign node2061 = (inp[10]) ? node2065 : node2062;
															assign node2062 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node2065 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node2068 = (inp[10]) ? node2072 : node2069;
															assign node2069 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node2072 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node2075 = (inp[7]) ? node2087 : node2076;
														assign node2076 = (inp[4]) ? node2082 : node2077;
															assign node2077 = (inp[11]) ? 4'b0011 : node2078;
																assign node2078 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node2082 = (inp[10]) ? 4'b0111 : node2083;
																assign node2083 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node2087 = (inp[4]) ? node2091 : node2088;
															assign node2088 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node2091 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node2094 = (inp[12]) ? node2120 : node2095;
													assign node2095 = (inp[10]) ? node2105 : node2096;
														assign node2096 = (inp[11]) ? node2098 : 4'b0001;
															assign node2098 = (inp[4]) ? node2102 : node2099;
																assign node2099 = (inp[7]) ? 4'b0111 : 4'b0001;
																assign node2102 = (inp[7]) ? 4'b0000 : 4'b0111;
														assign node2105 = (inp[11]) ? node2113 : node2106;
															assign node2106 = (inp[4]) ? node2110 : node2107;
																assign node2107 = (inp[7]) ? 4'b0110 : 4'b0000;
																assign node2110 = (inp[7]) ? 4'b0000 : 4'b0110;
															assign node2113 = (inp[4]) ? node2117 : node2114;
																assign node2114 = (inp[7]) ? 4'b0110 : 4'b0000;
																assign node2117 = (inp[7]) ? 4'b0001 : 4'b0110;
													assign node2120 = (inp[4]) ? node2128 : node2121;
														assign node2121 = (inp[7]) ? node2125 : node2122;
															assign node2122 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2125 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2128 = (inp[11]) ? 4'b0000 : node2129;
															assign node2129 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node2133 = (inp[12]) ? node2165 : node2134;
												assign node2134 = (inp[7]) ? node2148 : node2135;
													assign node2135 = (inp[10]) ? node2141 : node2136;
														assign node2136 = (inp[15]) ? node2138 : 4'b0101;
															assign node2138 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node2141 = (inp[4]) ? node2143 : 4'b0100;
															assign node2143 = (inp[15]) ? node2145 : 4'b0100;
																assign node2145 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node2148 = (inp[15]) ? node2156 : node2149;
														assign node2149 = (inp[10]) ? node2151 : 4'b0110;
															assign node2151 = (inp[4]) ? 4'b0111 : node2152;
																assign node2152 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node2156 = (inp[4]) ? node2162 : node2157;
															assign node2157 = (inp[10]) ? node2159 : 4'b0011;
																assign node2159 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node2162 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node2165 = (inp[7]) ? node2185 : node2166;
													assign node2166 = (inp[4]) ? node2174 : node2167;
														assign node2167 = (inp[15]) ? 4'b0111 : node2168;
															assign node2168 = (inp[10]) ? node2170 : 4'b0111;
																assign node2170 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node2174 = (inp[15]) ? node2182 : node2175;
															assign node2175 = (inp[11]) ? node2179 : node2176;
																assign node2176 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node2179 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node2182 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node2185 = (inp[4]) ? node2189 : node2186;
														assign node2186 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2189 = (inp[15]) ? node2193 : node2190;
															assign node2190 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node2193 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node2196 = (inp[5]) ? node2318 : node2197;
										assign node2197 = (inp[12]) ? node2253 : node2198;
											assign node2198 = (inp[7]) ? node2228 : node2199;
												assign node2199 = (inp[4]) ? node2213 : node2200;
													assign node2200 = (inp[15]) ? node2206 : node2201;
														assign node2201 = (inp[11]) ? node2203 : 4'b0100;
															assign node2203 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node2206 = (inp[11]) ? 4'b0101 : node2207;
															assign node2207 = (inp[10]) ? 4'b0101 : node2208;
																assign node2208 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node2213 = (inp[15]) ? node2221 : node2214;
														assign node2214 = (inp[11]) ? node2218 : node2215;
															assign node2215 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2218 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node2221 = (inp[1]) ? node2223 : 4'b0110;
															assign node2223 = (inp[10]) ? node2225 : 4'b0010;
																assign node2225 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node2228 = (inp[15]) ? node2240 : node2229;
													assign node2229 = (inp[1]) ? node2233 : node2230;
														assign node2230 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node2233 = (inp[11]) ? node2235 : 4'b0110;
															assign node2235 = (inp[4]) ? node2237 : 4'b0111;
																assign node2237 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node2240 = (inp[4]) ? node2246 : node2241;
														assign node2241 = (inp[1]) ? node2243 : 4'b0010;
															assign node2243 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node2246 = (inp[10]) ? node2250 : node2247;
															assign node2247 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2250 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node2253 = (inp[7]) ? node2281 : node2254;
												assign node2254 = (inp[15]) ? node2266 : node2255;
													assign node2255 = (inp[4]) ? node2257 : 4'b0111;
														assign node2257 = (inp[11]) ? node2259 : 4'b0010;
															assign node2259 = (inp[10]) ? node2263 : node2260;
																assign node2260 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node2263 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node2266 = (inp[4]) ? node2272 : node2267;
														assign node2267 = (inp[10]) ? 4'b0111 : node2268;
															assign node2268 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node2272 = (inp[11]) ? node2278 : node2273;
															assign node2273 = (inp[10]) ? 4'b0100 : node2274;
																assign node2274 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2278 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node2281 = (inp[4]) ? node2303 : node2282;
													assign node2282 = (inp[10]) ? node2294 : node2283;
														assign node2283 = (inp[1]) ? node2289 : node2284;
															assign node2284 = (inp[15]) ? node2286 : 4'b0101;
																assign node2286 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node2289 = (inp[15]) ? 4'b0101 : node2290;
																assign node2290 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node2294 = (inp[15]) ? node2298 : node2295;
															assign node2295 = (inp[1]) ? 4'b0001 : 4'b0100;
															assign node2298 = (inp[11]) ? 4'b0001 : node2299;
																assign node2299 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node2303 = (inp[15]) ? node2309 : node2304;
														assign node2304 = (inp[1]) ? 4'b0100 : node2305;
															assign node2305 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2309 = (inp[1]) ? node2311 : 4'b0011;
															assign node2311 = (inp[10]) ? node2315 : node2312;
																assign node2312 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node2315 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node2318 = (inp[1]) ? node2402 : node2319;
											assign node2319 = (inp[4]) ? node2365 : node2320;
												assign node2320 = (inp[7]) ? node2342 : node2321;
													assign node2321 = (inp[12]) ? node2329 : node2322;
														assign node2322 = (inp[15]) ? node2324 : 4'b0100;
															assign node2324 = (inp[10]) ? node2326 : 4'b0101;
																assign node2326 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2329 = (inp[15]) ? node2337 : node2330;
															assign node2330 = (inp[11]) ? node2334 : node2331;
																assign node2331 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node2334 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node2337 = (inp[11]) ? node2339 : 4'b0110;
																assign node2339 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2342 = (inp[12]) ? node2354 : node2343;
														assign node2343 = (inp[15]) ? node2351 : node2344;
															assign node2344 = (inp[11]) ? node2348 : node2345;
																assign node2345 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node2348 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2351 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node2354 = (inp[15]) ? node2360 : node2355;
															assign node2355 = (inp[11]) ? node2357 : 4'b0001;
																assign node2357 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node2360 = (inp[10]) ? 4'b0100 : node2361;
																assign node2361 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node2365 = (inp[7]) ? node2387 : node2366;
													assign node2366 = (inp[15]) ? node2376 : node2367;
														assign node2367 = (inp[12]) ? node2369 : 4'b0101;
															assign node2369 = (inp[11]) ? node2373 : node2370;
																assign node2370 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node2373 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node2376 = (inp[12]) ? node2382 : node2377;
															assign node2377 = (inp[10]) ? node2379 : 4'b0011;
																assign node2379 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node2382 = (inp[11]) ? 4'b0101 : node2383;
																assign node2383 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node2387 = (inp[12]) ? node2395 : node2388;
														assign node2388 = (inp[15]) ? node2390 : 4'b0111;
															assign node2390 = (inp[10]) ? 4'b0100 : node2391;
																assign node2391 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2395 = (inp[15]) ? node2397 : 4'b0101;
															assign node2397 = (inp[11]) ? node2399 : 4'b0011;
																assign node2399 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node2402 = (inp[7]) ? node2440 : node2403;
												assign node2403 = (inp[12]) ? node2423 : node2404;
													assign node2404 = (inp[4]) ? node2414 : node2405;
														assign node2405 = (inp[11]) ? node2407 : 4'b0001;
															assign node2407 = (inp[15]) ? node2411 : node2408;
																assign node2408 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node2411 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2414 = (inp[15]) ? node2420 : node2415;
															assign node2415 = (inp[10]) ? 4'b0000 : node2416;
																assign node2416 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node2420 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node2423 = (inp[15]) ? node2433 : node2424;
														assign node2424 = (inp[4]) ? node2428 : node2425;
															assign node2425 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2428 = (inp[11]) ? node2430 : 4'b0110;
																assign node2430 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node2433 = (inp[4]) ? node2435 : 4'b0011;
															assign node2435 = (inp[10]) ? node2437 : 4'b0001;
																assign node2437 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node2440 = (inp[12]) ? node2454 : node2441;
													assign node2441 = (inp[4]) ? node2445 : node2442;
														assign node2442 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node2445 = (inp[15]) ? node2449 : node2446;
															assign node2446 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2449 = (inp[11]) ? node2451 : 4'b0001;
																assign node2451 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node2454 = (inp[15]) ? node2460 : node2455;
														assign node2455 = (inp[4]) ? node2457 : 4'b0000;
															assign node2457 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node2460 = (inp[10]) ? node2464 : node2461;
															assign node2461 = (inp[4]) ? 4'b0110 : 4'b0100;
															assign node2464 = (inp[4]) ? 4'b0111 : 4'b0101;
								assign node2467 = (inp[2]) ? node2739 : node2468;
									assign node2468 = (inp[11]) ? node2602 : node2469;
										assign node2469 = (inp[10]) ? node2535 : node2470;
											assign node2470 = (inp[5]) ? node2504 : node2471;
												assign node2471 = (inp[12]) ? node2489 : node2472;
													assign node2472 = (inp[7]) ? node2482 : node2473;
														assign node2473 = (inp[4]) ? node2479 : node2474;
															assign node2474 = (inp[1]) ? 4'b0100 : node2475;
																assign node2475 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node2479 = (inp[1]) ? 4'b0010 : 4'b0100;
														assign node2482 = (inp[4]) ? node2486 : node2483;
															assign node2483 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node2486 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node2489 = (inp[15]) ? node2495 : node2490;
														assign node2490 = (inp[4]) ? 4'b0010 : node2491;
															assign node2491 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node2495 = (inp[7]) ? node2501 : node2496;
															assign node2496 = (inp[4]) ? node2498 : 4'b0111;
																assign node2498 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2501 = (inp[1]) ? 4'b0100 : 4'b0011;
												assign node2504 = (inp[1]) ? node2524 : node2505;
													assign node2505 = (inp[15]) ? node2517 : node2506;
														assign node2506 = (inp[12]) ? node2514 : node2507;
															assign node2507 = (inp[7]) ? node2511 : node2508;
																assign node2508 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node2511 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node2514 = (inp[4]) ? 4'b0011 : 4'b0110;
														assign node2517 = (inp[12]) ? node2521 : node2518;
															assign node2518 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node2521 = (inp[7]) ? 4'b0101 : 4'b0111;
													assign node2524 = (inp[15]) ? node2526 : 4'b0001;
														assign node2526 = (inp[7]) ? node2532 : node2527;
															assign node2527 = (inp[4]) ? node2529 : 4'b0000;
																assign node2529 = (inp[12]) ? 4'b0000 : 4'b0011;
															assign node2532 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node2535 = (inp[1]) ? node2567 : node2536;
												assign node2536 = (inp[12]) ? node2548 : node2537;
													assign node2537 = (inp[7]) ? node2541 : node2538;
														assign node2538 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node2541 = (inp[15]) ? node2545 : node2542;
															assign node2542 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node2545 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node2548 = (inp[7]) ? node2556 : node2549;
														assign node2549 = (inp[15]) ? node2553 : node2550;
															assign node2550 = (inp[4]) ? 4'b0010 : 4'b0111;
															assign node2553 = (inp[4]) ? 4'b0101 : 4'b0110;
														assign node2556 = (inp[5]) ? node2562 : node2557;
															assign node2557 = (inp[4]) ? node2559 : 4'b0001;
																assign node2559 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node2562 = (inp[15]) ? 4'b0100 : node2563;
																assign node2563 = (inp[4]) ? 4'b0100 : 4'b0001;
												assign node2567 = (inp[7]) ? node2587 : node2568;
													assign node2568 = (inp[12]) ? node2576 : node2569;
														assign node2569 = (inp[5]) ? node2573 : node2570;
															assign node2570 = (inp[15]) ? 4'b0011 : 4'b0101;
															assign node2573 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node2576 = (inp[4]) ? node2582 : node2577;
															assign node2577 = (inp[15]) ? node2579 : 4'b0011;
																assign node2579 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node2582 = (inp[15]) ? 4'b0001 : node2583;
																assign node2583 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node2587 = (inp[12]) ? node2595 : node2588;
														assign node2588 = (inp[15]) ? node2590 : 4'b0111;
															assign node2590 = (inp[4]) ? node2592 : 4'b0011;
																assign node2592 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node2595 = (inp[5]) ? 4'b0111 : node2596;
															assign node2596 = (inp[15]) ? 4'b0101 : node2597;
																assign node2597 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node2602 = (inp[5]) ? node2672 : node2603;
											assign node2603 = (inp[12]) ? node2633 : node2604;
												assign node2604 = (inp[7]) ? node2620 : node2605;
													assign node2605 = (inp[4]) ? node2613 : node2606;
														assign node2606 = (inp[10]) ? node2610 : node2607;
															assign node2607 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node2610 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node2613 = (inp[15]) ? node2617 : node2614;
															assign node2614 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2617 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node2620 = (inp[15]) ? node2624 : node2621;
														assign node2621 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node2624 = (inp[4]) ? node2630 : node2625;
															assign node2625 = (inp[1]) ? 4'b0011 : node2626;
																assign node2626 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2630 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node2633 = (inp[7]) ? node2653 : node2634;
													assign node2634 = (inp[15]) ? node2644 : node2635;
														assign node2635 = (inp[4]) ? node2639 : node2636;
															assign node2636 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node2639 = (inp[10]) ? 4'b0010 : node2640;
																assign node2640 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node2644 = (inp[4]) ? node2650 : node2645;
															assign node2645 = (inp[1]) ? 4'b0110 : node2646;
																assign node2646 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2650 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node2653 = (inp[1]) ? node2661 : node2654;
														assign node2654 = (inp[15]) ? node2658 : node2655;
															assign node2655 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node2658 = (inp[4]) ? 4'b0010 : 4'b0000;
														assign node2661 = (inp[4]) ? node2667 : node2662;
															assign node2662 = (inp[15]) ? node2664 : 4'b0001;
																assign node2664 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node2667 = (inp[15]) ? 4'b0010 : node2668;
																assign node2668 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node2672 = (inp[1]) ? node2712 : node2673;
												assign node2673 = (inp[4]) ? node2691 : node2674;
													assign node2674 = (inp[10]) ? node2684 : node2675;
														assign node2675 = (inp[15]) ? node2679 : node2676;
															assign node2676 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node2679 = (inp[12]) ? node2681 : 4'b0100;
																assign node2681 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node2684 = (inp[15]) ? node2686 : 4'b0000;
															assign node2686 = (inp[12]) ? node2688 : 4'b0101;
																assign node2688 = (inp[7]) ? 4'b0101 : 4'b0111;
													assign node2691 = (inp[15]) ? node2701 : node2692;
														assign node2692 = (inp[10]) ? node2696 : node2693;
															assign node2693 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node2696 = (inp[12]) ? 4'b0100 : node2697;
																assign node2697 = (inp[7]) ? 4'b0111 : 4'b0100;
														assign node2701 = (inp[10]) ? node2707 : node2702;
															assign node2702 = (inp[12]) ? node2704 : 4'b0100;
																assign node2704 = (inp[7]) ? 4'b0011 : 4'b0101;
															assign node2707 = (inp[12]) ? node2709 : 4'b0010;
																assign node2709 = (inp[7]) ? 4'b0010 : 4'b0100;
												assign node2712 = (inp[7]) ? node2722 : node2713;
													assign node2713 = (inp[15]) ? node2717 : node2714;
														assign node2714 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node2717 = (inp[4]) ? 4'b0010 : node2718;
															assign node2718 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node2722 = (inp[12]) ? node2730 : node2723;
														assign node2723 = (inp[4]) ? node2727 : node2724;
															assign node2724 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2727 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node2730 = (inp[15]) ? node2736 : node2731;
															assign node2731 = (inp[10]) ? 4'b0101 : node2732;
																assign node2732 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node2736 = (inp[4]) ? 4'b0111 : 4'b0101;
									assign node2739 = (inp[5]) ? node2855 : node2740;
										assign node2740 = (inp[12]) ? node2796 : node2741;
											assign node2741 = (inp[7]) ? node2765 : node2742;
												assign node2742 = (inp[15]) ? node2756 : node2743;
													assign node2743 = (inp[11]) ? node2749 : node2744;
														assign node2744 = (inp[4]) ? 4'b0001 : node2745;
															assign node2745 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2749 = (inp[4]) ? node2753 : node2750;
															assign node2750 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node2753 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node2756 = (inp[4]) ? node2760 : node2757;
														assign node2757 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2760 = (inp[1]) ? node2762 : 4'b0010;
															assign node2762 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node2765 = (inp[15]) ? node2781 : node2766;
													assign node2766 = (inp[11]) ? node2772 : node2767;
														assign node2767 = (inp[4]) ? 4'b0010 : node2768;
															assign node2768 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node2772 = (inp[1]) ? node2774 : 4'b0010;
															assign node2774 = (inp[4]) ? node2778 : node2775;
																assign node2775 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node2778 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node2781 = (inp[4]) ? node2785 : node2782;
														assign node2782 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node2785 = (inp[10]) ? node2791 : node2786;
															assign node2786 = (inp[1]) ? 4'b0000 : node2787;
																assign node2787 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node2791 = (inp[1]) ? 4'b0001 : node2792;
																assign node2792 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node2796 = (inp[7]) ? node2828 : node2797;
												assign node2797 = (inp[4]) ? node2815 : node2798;
													assign node2798 = (inp[11]) ? node2806 : node2799;
														assign node2799 = (inp[10]) ? node2801 : 4'b0011;
															assign node2801 = (inp[15]) ? node2803 : 4'b0011;
																assign node2803 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node2806 = (inp[10]) ? node2812 : node2807;
															assign node2807 = (inp[1]) ? 4'b0010 : node2808;
																assign node2808 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node2812 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node2815 = (inp[15]) ? node2821 : node2816;
														assign node2816 = (inp[1]) ? node2818 : 4'b0110;
															assign node2818 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node2821 = (inp[11]) ? node2823 : 4'b0000;
															assign node2823 = (inp[10]) ? node2825 : 4'b0001;
																assign node2825 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node2828 = (inp[15]) ? node2842 : node2829;
													assign node2829 = (inp[1]) ? node2839 : node2830;
														assign node2830 = (inp[4]) ? 4'b0100 : node2831;
															assign node2831 = (inp[11]) ? node2835 : node2832;
																assign node2832 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node2835 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2839 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node2842 = (inp[4]) ? node2852 : node2843;
														assign node2843 = (inp[1]) ? 4'b0000 : node2844;
															assign node2844 = (inp[10]) ? node2848 : node2845;
																assign node2845 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node2848 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2852 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node2855 = (inp[1]) ? node2921 : node2856;
											assign node2856 = (inp[7]) ? node2892 : node2857;
												assign node2857 = (inp[12]) ? node2877 : node2858;
													assign node2858 = (inp[4]) ? node2864 : node2859;
														assign node2859 = (inp[10]) ? 4'b0001 : node2860;
															assign node2860 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node2864 = (inp[15]) ? node2872 : node2865;
															assign node2865 = (inp[11]) ? node2869 : node2866;
																assign node2866 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node2869 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node2872 = (inp[11]) ? 4'b0110 : node2873;
																assign node2873 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2877 = (inp[4]) ? node2885 : node2878;
														assign node2878 = (inp[10]) ? node2882 : node2879;
															assign node2879 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node2882 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node2885 = (inp[15]) ? node2889 : node2886;
															assign node2886 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node2889 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node2892 = (inp[12]) ? node2904 : node2893;
													assign node2893 = (inp[15]) ? node2899 : node2894;
														assign node2894 = (inp[10]) ? 4'b0011 : node2895;
															assign node2895 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node2899 = (inp[4]) ? 4'b0001 : node2900;
															assign node2900 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2904 = (inp[4]) ? node2914 : node2905;
														assign node2905 = (inp[15]) ? node2911 : node2906;
															assign node2906 = (inp[11]) ? node2908 : 4'b0101;
																assign node2908 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2911 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node2914 = (inp[15]) ? 4'b0110 : node2915;
															assign node2915 = (inp[11]) ? node2917 : 4'b0000;
																assign node2917 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node2921 = (inp[12]) ? node2959 : node2922;
												assign node2922 = (inp[7]) ? node2940 : node2923;
													assign node2923 = (inp[4]) ? node2931 : node2924;
														assign node2924 = (inp[10]) ? 4'b0100 : node2925;
															assign node2925 = (inp[11]) ? 4'b0101 : node2926;
																assign node2926 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node2931 = (inp[15]) ? node2937 : node2932;
															assign node2932 = (inp[11]) ? node2934 : 4'b0100;
																assign node2934 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node2937 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node2940 = (inp[15]) ? node2950 : node2941;
														assign node2941 = (inp[10]) ? node2947 : node2942;
															assign node2942 = (inp[11]) ? 4'b0110 : node2943;
																assign node2943 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node2947 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node2950 = (inp[4]) ? node2954 : node2951;
															assign node2951 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2954 = (inp[11]) ? 4'b0101 : node2955;
																assign node2955 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node2959 = (inp[7]) ? node2979 : node2960;
													assign node2960 = (inp[15]) ? node2968 : node2961;
														assign node2961 = (inp[4]) ? node2965 : node2962;
															assign node2962 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2965 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node2968 = (inp[4]) ? node2974 : node2969;
															assign node2969 = (inp[11]) ? 4'b0110 : node2970;
																assign node2970 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node2974 = (inp[10]) ? node2976 : 4'b0100;
																assign node2976 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node2979 = (inp[4]) ? node2989 : node2980;
														assign node2980 = (inp[15]) ? node2986 : node2981;
															assign node2981 = (inp[11]) ? node2983 : 4'b0101;
																assign node2983 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node2986 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node2989 = (inp[15]) ? node2991 : 4'b0000;
															assign node2991 = (inp[10]) ? node2993 : 4'b0011;
																assign node2993 = (inp[11]) ? 4'b0011 : 4'b0010;
							assign node2996 = (inp[10]) ? node3602 : node2997;
								assign node2997 = (inp[11]) ? node3307 : node2998;
									assign node2998 = (inp[15]) ? node3158 : node2999;
										assign node2999 = (inp[5]) ? node3065 : node3000;
											assign node3000 = (inp[2]) ? node3032 : node3001;
												assign node3001 = (inp[13]) ? node3015 : node3002;
													assign node3002 = (inp[12]) ? node3006 : node3003;
														assign node3003 = (inp[7]) ? 4'b0011 : 4'b0001;
														assign node3006 = (inp[7]) ? node3010 : node3007;
															assign node3007 = (inp[4]) ? 4'b0110 : 4'b0011;
															assign node3010 = (inp[1]) ? node3012 : 4'b0000;
																assign node3012 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node3015 = (inp[12]) ? node3019 : node3016;
														assign node3016 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node3019 = (inp[7]) ? node3025 : node3020;
															assign node3020 = (inp[4]) ? 4'b0010 : node3021;
																assign node3021 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node3025 = (inp[1]) ? node3029 : node3026;
																assign node3026 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node3029 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node3032 = (inp[13]) ? node3048 : node3033;
													assign node3033 = (inp[4]) ? node3041 : node3034;
														assign node3034 = (inp[12]) ? node3038 : node3035;
															assign node3035 = (inp[7]) ? 4'b0111 : 4'b0101;
															assign node3038 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node3041 = (inp[12]) ? node3045 : node3042;
															assign node3042 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node3045 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node3048 = (inp[12]) ? node3056 : node3049;
														assign node3049 = (inp[4]) ? node3053 : node3050;
															assign node3050 = (inp[7]) ? 4'b0010 : 4'b0000;
															assign node3053 = (inp[7]) ? 4'b0011 : 4'b0001;
														assign node3056 = (inp[7]) ? node3060 : node3057;
															assign node3057 = (inp[4]) ? 4'b0110 : 4'b0011;
															assign node3060 = (inp[1]) ? 4'b0101 : node3061;
																assign node3061 = (inp[4]) ? 4'b0101 : 4'b0000;
											assign node3065 = (inp[12]) ? node3109 : node3066;
												assign node3066 = (inp[7]) ? node3086 : node3067;
													assign node3067 = (inp[13]) ? node3079 : node3068;
														assign node3068 = (inp[4]) ? node3074 : node3069;
															assign node3069 = (inp[1]) ? node3071 : 4'b0101;
																assign node3071 = (inp[2]) ? 4'b0000 : 4'b0101;
															assign node3074 = (inp[2]) ? node3076 : 4'b0000;
																assign node3076 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node3079 = (inp[4]) ? 4'b0001 : node3080;
															assign node3080 = (inp[2]) ? node3082 : 4'b0000;
																assign node3082 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node3086 = (inp[2]) ? node3096 : node3087;
														assign node3087 = (inp[13]) ? node3091 : node3088;
															assign node3088 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node3091 = (inp[1]) ? 4'b0011 : node3092;
																assign node3092 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node3096 = (inp[4]) ? node3102 : node3097;
															assign node3097 = (inp[1]) ? 4'b0011 : node3098;
																assign node3098 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node3102 = (inp[13]) ? node3106 : node3103;
																assign node3103 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node3106 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node3109 = (inp[7]) ? node3133 : node3110;
													assign node3110 = (inp[2]) ? node3120 : node3111;
														assign node3111 = (inp[1]) ? node3115 : node3112;
															assign node3112 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node3115 = (inp[4]) ? node3117 : 4'b0110;
																assign node3117 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node3120 = (inp[1]) ? node3128 : node3121;
															assign node3121 = (inp[4]) ? node3125 : node3122;
																assign node3122 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node3125 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node3128 = (inp[13]) ? node3130 : 4'b0011;
																assign node3130 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node3133 = (inp[1]) ? node3147 : node3134;
														assign node3134 = (inp[4]) ? node3142 : node3135;
															assign node3135 = (inp[2]) ? node3139 : node3136;
																assign node3136 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node3139 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3142 = (inp[2]) ? 4'b0001 : node3143;
																assign node3143 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node3147 = (inp[2]) ? node3153 : node3148;
															assign node3148 = (inp[4]) ? node3150 : 4'b0100;
																assign node3150 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3153 = (inp[13]) ? 4'b0100 : node3154;
																assign node3154 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node3158 = (inp[2]) ? node3228 : node3159;
											assign node3159 = (inp[13]) ? node3193 : node3160;
												assign node3160 = (inp[4]) ? node3178 : node3161;
													assign node3161 = (inp[12]) ? node3173 : node3162;
														assign node3162 = (inp[7]) ? node3168 : node3163;
															assign node3163 = (inp[1]) ? node3165 : 4'b0001;
																assign node3165 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node3168 = (inp[5]) ? node3170 : 4'b0110;
																assign node3170 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node3173 = (inp[7]) ? node3175 : 4'b0011;
															assign node3175 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node3178 = (inp[5]) ? node3188 : node3179;
														assign node3179 = (inp[7]) ? node3185 : node3180;
															assign node3180 = (inp[12]) ? node3182 : 4'b0110;
																assign node3182 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3185 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node3188 = (inp[12]) ? node3190 : 4'b0110;
															assign node3190 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node3193 = (inp[4]) ? node3215 : node3194;
													assign node3194 = (inp[12]) ? node3204 : node3195;
														assign node3195 = (inp[7]) ? node3199 : node3196;
															assign node3196 = (inp[5]) ? 4'b0001 : 4'b0100;
															assign node3199 = (inp[5]) ? node3201 : 4'b0011;
																assign node3201 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node3204 = (inp[7]) ? node3210 : node3205;
															assign node3205 = (inp[5]) ? node3207 : 4'b0110;
																assign node3207 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node3210 = (inp[5]) ? 4'b0100 : node3211;
																assign node3211 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node3215 = (inp[5]) ? node3219 : node3216;
														assign node3216 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node3219 = (inp[7]) ? node3225 : node3220;
															assign node3220 = (inp[12]) ? node3222 : 4'b0011;
																assign node3222 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node3225 = (inp[12]) ? 4'b0111 : 4'b0100;
											assign node3228 = (inp[1]) ? node3270 : node3229;
												assign node3229 = (inp[13]) ? node3251 : node3230;
													assign node3230 = (inp[7]) ? node3238 : node3231;
														assign node3231 = (inp[12]) ? node3235 : node3232;
															assign node3232 = (inp[4]) ? 4'b0011 : 4'b0101;
															assign node3235 = (inp[4]) ? 4'b0101 : 4'b0111;
														assign node3238 = (inp[4]) ? node3246 : node3239;
															assign node3239 = (inp[5]) ? node3243 : node3240;
																assign node3240 = (inp[12]) ? 4'b0000 : 4'b0010;
																assign node3243 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node3246 = (inp[12]) ? 4'b0011 : node3247;
																assign node3247 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node3251 = (inp[4]) ? node3259 : node3252;
														assign node3252 = (inp[7]) ? node3256 : node3253;
															assign node3253 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node3256 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node3259 = (inp[12]) ? node3263 : node3260;
															assign node3260 = (inp[7]) ? 4'b0000 : 4'b0010;
															assign node3263 = (inp[7]) ? node3267 : node3264;
																assign node3264 = (inp[5]) ? 4'b0001 : 4'b0000;
																assign node3267 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node3270 = (inp[12]) ? node3288 : node3271;
													assign node3271 = (inp[13]) ? node3281 : node3272;
														assign node3272 = (inp[5]) ? node3278 : node3273;
															assign node3273 = (inp[4]) ? 4'b0101 : node3274;
																assign node3274 = (inp[7]) ? 4'b0010 : 4'b0100;
															assign node3278 = (inp[4]) ? 4'b0010 : 4'b0000;
														assign node3281 = (inp[5]) ? node3283 : 4'b0001;
															assign node3283 = (inp[7]) ? 4'b0100 : node3284;
																assign node3284 = (inp[4]) ? 4'b0111 : 4'b0101;
													assign node3288 = (inp[5]) ? node3300 : node3289;
														assign node3289 = (inp[13]) ? node3295 : node3290;
															assign node3290 = (inp[7]) ? node3292 : 4'b0100;
																assign node3292 = (inp[4]) ? 4'b0011 : 4'b0100;
															assign node3295 = (inp[4]) ? 4'b0110 : node3296;
																assign node3296 = (inp[7]) ? 4'b0001 : 4'b0010;
														assign node3300 = (inp[13]) ? node3304 : node3301;
															assign node3301 = (inp[4]) ? 4'b0001 : 4'b0011;
															assign node3304 = (inp[4]) ? 4'b0010 : 4'b0000;
									assign node3307 = (inp[2]) ? node3447 : node3308;
										assign node3308 = (inp[5]) ? node3374 : node3309;
											assign node3309 = (inp[15]) ? node3339 : node3310;
												assign node3310 = (inp[13]) ? node3326 : node3311;
													assign node3311 = (inp[12]) ? node3315 : node3312;
														assign node3312 = (inp[7]) ? 4'b0010 : 4'b0000;
														assign node3315 = (inp[7]) ? node3319 : node3316;
															assign node3316 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node3319 = (inp[1]) ? node3323 : node3320;
																assign node3320 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node3323 = (inp[4]) ? 4'b0000 : 4'b0101;
													assign node3326 = (inp[12]) ? node3330 : node3327;
														assign node3327 = (inp[7]) ? 4'b0110 : 4'b0100;
														assign node3330 = (inp[7]) ? node3334 : node3331;
															assign node3331 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node3334 = (inp[4]) ? 4'b0100 : node3335;
																assign node3335 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node3339 = (inp[1]) ? node3353 : node3340;
													assign node3340 = (inp[7]) ? node3346 : node3341;
														assign node3341 = (inp[4]) ? node3343 : 4'b0111;
															assign node3343 = (inp[12]) ? 4'b0101 : 4'b0111;
														assign node3346 = (inp[4]) ? node3348 : 4'b0100;
															assign node3348 = (inp[12]) ? node3350 : 4'b0101;
																assign node3350 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node3353 = (inp[4]) ? node3367 : node3354;
														assign node3354 = (inp[13]) ? node3360 : node3355;
															assign node3355 = (inp[12]) ? 4'b0000 : node3356;
																assign node3356 = (inp[7]) ? 4'b0110 : 4'b0000;
															assign node3360 = (inp[12]) ? node3364 : node3361;
																assign node3361 = (inp[7]) ? 4'b0010 : 4'b0101;
																assign node3364 = (inp[7]) ? 4'b0101 : 4'b0110;
														assign node3367 = (inp[12]) ? 4'b0010 : node3368;
															assign node3368 = (inp[7]) ? 4'b0100 : node3369;
																assign node3369 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node3374 = (inp[4]) ? node3412 : node3375;
												assign node3375 = (inp[7]) ? node3389 : node3376;
													assign node3376 = (inp[12]) ? node3382 : node3377;
														assign node3377 = (inp[15]) ? node3379 : 4'b0000;
															assign node3379 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node3382 = (inp[1]) ? node3386 : node3383;
															assign node3383 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node3386 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node3389 = (inp[12]) ? node3401 : node3390;
														assign node3390 = (inp[13]) ? node3396 : node3391;
															assign node3391 = (inp[15]) ? 4'b0010 : node3392;
																assign node3392 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node3396 = (inp[1]) ? node3398 : 4'b0111;
																assign node3398 = (inp[15]) ? 4'b0111 : 4'b0011;
														assign node3401 = (inp[15]) ? node3407 : node3402;
															assign node3402 = (inp[13]) ? node3404 : 4'b0101;
																assign node3404 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3407 = (inp[13]) ? node3409 : 4'b0000;
																assign node3409 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node3412 = (inp[12]) ? node3426 : node3413;
													assign node3413 = (inp[13]) ? node3421 : node3414;
														assign node3414 = (inp[1]) ? node3416 : 4'b0000;
															assign node3416 = (inp[7]) ? 4'b0100 : node3417;
																assign node3417 = (inp[15]) ? 4'b0111 : 4'b0100;
														assign node3421 = (inp[15]) ? node3423 : 4'b0001;
															assign node3423 = (inp[7]) ? 4'b0000 : 4'b0010;
													assign node3426 = (inp[7]) ? node3434 : node3427;
														assign node3427 = (inp[15]) ? node3429 : 4'b0110;
															assign node3429 = (inp[13]) ? 4'b0100 : node3430;
																assign node3430 = (inp[1]) ? 4'b0100 : 4'b0001;
														assign node3434 = (inp[15]) ? node3440 : node3435;
															assign node3435 = (inp[13]) ? 4'b0100 : node3436;
																assign node3436 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3440 = (inp[13]) ? node3444 : node3441;
																assign node3441 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node3444 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node3447 = (inp[13]) ? node3531 : node3448;
											assign node3448 = (inp[1]) ? node3486 : node3449;
												assign node3449 = (inp[12]) ? node3469 : node3450;
													assign node3450 = (inp[7]) ? node3458 : node3451;
														assign node3451 = (inp[4]) ? node3453 : 4'b0100;
															assign node3453 = (inp[15]) ? node3455 : 4'b0101;
																assign node3455 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node3458 = (inp[15]) ? node3466 : node3459;
															assign node3459 = (inp[5]) ? node3463 : node3460;
																assign node3460 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node3463 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node3466 = (inp[4]) ? 4'b0101 : 4'b0010;
													assign node3469 = (inp[7]) ? node3475 : node3470;
														assign node3470 = (inp[4]) ? node3472 : 4'b0110;
															assign node3472 = (inp[15]) ? 4'b0100 : 4'b0010;
														assign node3475 = (inp[5]) ? node3481 : node3476;
															assign node3476 = (inp[4]) ? node3478 : 4'b0001;
																assign node3478 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node3481 = (inp[4]) ? 4'b0101 : node3482;
																assign node3482 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node3486 = (inp[5]) ? node3510 : node3487;
													assign node3487 = (inp[12]) ? node3495 : node3488;
														assign node3488 = (inp[7]) ? node3490 : 4'b0100;
															assign node3490 = (inp[4]) ? 4'b0100 : node3491;
																assign node3491 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node3495 = (inp[7]) ? node3503 : node3496;
															assign node3496 = (inp[15]) ? node3500 : node3497;
																assign node3497 = (inp[4]) ? 4'b0010 : 4'b0111;
																assign node3500 = (inp[4]) ? 4'b0101 : 4'b0111;
															assign node3503 = (inp[4]) ? node3507 : node3504;
																assign node3504 = (inp[15]) ? 4'b0100 : 4'b0000;
																assign node3507 = (inp[15]) ? 4'b0010 : 4'b0101;
													assign node3510 = (inp[7]) ? node3520 : node3511;
														assign node3511 = (inp[15]) ? node3515 : node3512;
															assign node3512 = (inp[12]) ? 4'b0011 : 4'b0000;
															assign node3515 = (inp[4]) ? node3517 : 4'b0010;
																assign node3517 = (inp[12]) ? 4'b0000 : 4'b0010;
														assign node3520 = (inp[15]) ? node3524 : node3521;
															assign node3521 = (inp[12]) ? 4'b0001 : 4'b0011;
															assign node3524 = (inp[12]) ? node3528 : node3525;
																assign node3525 = (inp[4]) ? 4'b0000 : 4'b0110;
																assign node3528 = (inp[4]) ? 4'b0111 : 4'b0101;
											assign node3531 = (inp[5]) ? node3565 : node3532;
												assign node3532 = (inp[15]) ? node3550 : node3533;
													assign node3533 = (inp[4]) ? node3543 : node3534;
														assign node3534 = (inp[12]) ? node3538 : node3535;
															assign node3535 = (inp[1]) ? 4'b0000 : 4'b0010;
															assign node3538 = (inp[7]) ? 4'b0001 : node3539;
																assign node3539 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node3543 = (inp[12]) ? node3547 : node3544;
															assign node3544 = (inp[7]) ? 4'b0011 : 4'b0001;
															assign node3547 = (inp[7]) ? 4'b0001 : 4'b0110;
													assign node3550 = (inp[7]) ? node3558 : node3551;
														assign node3551 = (inp[1]) ? node3553 : 4'b0001;
															assign node3553 = (inp[4]) ? node3555 : 4'b0000;
																assign node3555 = (inp[12]) ? 4'b0000 : 4'b0111;
														assign node3558 = (inp[4]) ? 4'b0111 : node3559;
															assign node3559 = (inp[12]) ? 4'b0100 : node3560;
																assign node3560 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node3565 = (inp[1]) ? node3585 : node3566;
													assign node3566 = (inp[15]) ? node3576 : node3567;
														assign node3567 = (inp[12]) ? node3571 : node3568;
															assign node3568 = (inp[7]) ? 4'b0011 : 4'b0000;
															assign node3571 = (inp[7]) ? node3573 : 4'b0110;
																assign node3573 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node3576 = (inp[12]) ? node3582 : node3577;
															assign node3577 = (inp[7]) ? node3579 : 4'b0111;
																assign node3579 = (inp[4]) ? 4'b0000 : 4'b0110;
															assign node3582 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node3585 = (inp[12]) ? node3595 : node3586;
														assign node3586 = (inp[7]) ? node3592 : node3587;
															assign node3587 = (inp[15]) ? node3589 : 4'b0100;
																assign node3589 = (inp[4]) ? 4'b0111 : 4'b0100;
															assign node3592 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node3595 = (inp[7]) ? node3597 : 4'b0111;
															assign node3597 = (inp[4]) ? node3599 : 4'b0001;
																assign node3599 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node3602 = (inp[11]) ? node3888 : node3603;
									assign node3603 = (inp[5]) ? node3737 : node3604;
										assign node3604 = (inp[12]) ? node3658 : node3605;
											assign node3605 = (inp[7]) ? node3627 : node3606;
												assign node3606 = (inp[15]) ? node3618 : node3607;
													assign node3607 = (inp[2]) ? node3611 : node3608;
														assign node3608 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node3611 = (inp[13]) ? node3615 : node3612;
															assign node3612 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node3615 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node3618 = (inp[4]) ? node3622 : node3619;
														assign node3619 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node3622 = (inp[2]) ? node3624 : 4'b0111;
															assign node3624 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node3627 = (inp[13]) ? node3643 : node3628;
													assign node3628 = (inp[1]) ? node3636 : node3629;
														assign node3629 = (inp[15]) ? node3633 : node3630;
															assign node3630 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node3633 = (inp[4]) ? 4'b0100 : 4'b0110;
														assign node3636 = (inp[15]) ? node3640 : node3637;
															assign node3637 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node3640 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node3643 = (inp[2]) ? node3649 : node3644;
														assign node3644 = (inp[15]) ? node3646 : 4'b0110;
															assign node3646 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node3649 = (inp[4]) ? node3653 : node3650;
															assign node3650 = (inp[15]) ? 4'b0110 : 4'b0011;
															assign node3653 = (inp[15]) ? node3655 : 4'b0010;
																assign node3655 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node3658 = (inp[7]) ? node3696 : node3659;
												assign node3659 = (inp[15]) ? node3679 : node3660;
													assign node3660 = (inp[1]) ? node3668 : node3661;
														assign node3661 = (inp[2]) ? 4'b0110 : node3662;
															assign node3662 = (inp[4]) ? node3664 : 4'b0110;
																assign node3664 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node3668 = (inp[13]) ? node3672 : node3669;
															assign node3669 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node3672 = (inp[2]) ? node3676 : node3673;
																assign node3673 = (inp[4]) ? 4'b0010 : 4'b0111;
																assign node3676 = (inp[4]) ? 4'b0111 : 4'b0010;
													assign node3679 = (inp[4]) ? node3689 : node3680;
														assign node3680 = (inp[13]) ? node3684 : node3681;
															assign node3681 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node3684 = (inp[2]) ? node3686 : 4'b0111;
																assign node3686 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node3689 = (inp[1]) ? 4'b0101 : node3690;
															assign node3690 = (inp[2]) ? 4'b0100 : node3691;
																assign node3691 = (inp[13]) ? 4'b0100 : 4'b0001;
												assign node3696 = (inp[4]) ? node3720 : node3697;
													assign node3697 = (inp[13]) ? node3709 : node3698;
														assign node3698 = (inp[15]) ? node3704 : node3699;
															assign node3699 = (inp[1]) ? node3701 : 4'b0001;
																assign node3701 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node3704 = (inp[1]) ? node3706 : 4'b0001;
																assign node3706 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node3709 = (inp[15]) ? node3713 : node3710;
															assign node3710 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node3713 = (inp[1]) ? node3717 : node3714;
																assign node3714 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3717 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node3720 = (inp[15]) ? node3730 : node3721;
														assign node3721 = (inp[1]) ? node3725 : node3722;
															assign node3722 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node3725 = (inp[13]) ? node3727 : 4'b0000;
																assign node3727 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node3730 = (inp[13]) ? node3732 : 4'b0010;
															assign node3732 = (inp[2]) ? 4'b0111 : node3733;
																assign node3733 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node3737 = (inp[7]) ? node3813 : node3738;
											assign node3738 = (inp[12]) ? node3768 : node3739;
												assign node3739 = (inp[15]) ? node3755 : node3740;
													assign node3740 = (inp[1]) ? node3748 : node3741;
														assign node3741 = (inp[13]) ? node3745 : node3742;
															assign node3742 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node3745 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node3748 = (inp[2]) ? node3750 : 4'b0100;
															assign node3750 = (inp[4]) ? 4'b0100 : node3751;
																assign node3751 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node3755 = (inp[4]) ? node3759 : node3756;
														assign node3756 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node3759 = (inp[2]) ? node3763 : node3760;
															assign node3760 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node3763 = (inp[13]) ? node3765 : 4'b0010;
																assign node3765 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node3768 = (inp[4]) ? node3786 : node3769;
													assign node3769 = (inp[13]) ? node3779 : node3770;
														assign node3770 = (inp[2]) ? node3776 : node3771;
															assign node3771 = (inp[1]) ? node3773 : 4'b0010;
																assign node3773 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node3776 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node3779 = (inp[15]) ? node3781 : 4'b0110;
															assign node3781 = (inp[2]) ? 4'b0111 : node3782;
																assign node3782 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node3786 = (inp[15]) ? node3798 : node3787;
														assign node3787 = (inp[2]) ? node3793 : node3788;
															assign node3788 = (inp[1]) ? 4'b0010 : node3789;
																assign node3789 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node3793 = (inp[13]) ? node3795 : 4'b0010;
																assign node3795 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node3798 = (inp[2]) ? node3806 : node3799;
															assign node3799 = (inp[13]) ? node3803 : node3800;
																assign node3800 = (inp[1]) ? 4'b0101 : 4'b0001;
																assign node3803 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node3806 = (inp[13]) ? node3810 : node3807;
																assign node3807 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node3810 = (inp[1]) ? 4'b0101 : 4'b0000;
											assign node3813 = (inp[12]) ? node3855 : node3814;
												assign node3814 = (inp[1]) ? node3830 : node3815;
													assign node3815 = (inp[4]) ? node3823 : node3816;
														assign node3816 = (inp[13]) ? 4'b0111 : node3817;
															assign node3817 = (inp[2]) ? 4'b0111 : node3818;
																assign node3818 = (inp[15]) ? 4'b0111 : 4'b0011;
														assign node3823 = (inp[15]) ? node3827 : node3824;
															assign node3824 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node3827 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3830 = (inp[4]) ? node3844 : node3831;
														assign node3831 = (inp[2]) ? node3839 : node3832;
															assign node3832 = (inp[13]) ? node3836 : node3833;
																assign node3833 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node3836 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node3839 = (inp[15]) ? node3841 : 4'b0010;
																assign node3841 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node3844 = (inp[2]) ? node3850 : node3845;
															assign node3845 = (inp[15]) ? 4'b0000 : node3846;
																assign node3846 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node3850 = (inp[15]) ? 4'b0101 : node3851;
																assign node3851 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node3855 = (inp[15]) ? node3873 : node3856;
													assign node3856 = (inp[1]) ? node3866 : node3857;
														assign node3857 = (inp[2]) ? node3863 : node3858;
															assign node3858 = (inp[4]) ? node3860 : 4'b0000;
																assign node3860 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3863 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node3866 = (inp[13]) ? node3868 : 4'b0101;
															assign node3868 = (inp[2]) ? node3870 : 4'b0001;
																assign node3870 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node3873 = (inp[4]) ? node3881 : node3874;
														assign node3874 = (inp[13]) ? node3876 : 4'b0000;
															assign node3876 = (inp[2]) ? node3878 : 4'b0101;
																assign node3878 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node3881 = (inp[1]) ? node3883 : 4'b0010;
															assign node3883 = (inp[13]) ? node3885 : 4'b0011;
																assign node3885 = (inp[2]) ? 4'b0011 : 4'b0110;
									assign node3888 = (inp[2]) ? node4032 : node3889;
										assign node3889 = (inp[13]) ? node3961 : node3890;
											assign node3890 = (inp[5]) ? node3928 : node3891;
												assign node3891 = (inp[1]) ? node3911 : node3892;
													assign node3892 = (inp[7]) ? node3902 : node3893;
														assign node3893 = (inp[15]) ? node3897 : node3894;
															assign node3894 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node3897 = (inp[12]) ? node3899 : 4'b0011;
																assign node3899 = (inp[4]) ? 4'b0001 : 4'b0011;
														assign node3902 = (inp[12]) ? node3906 : node3903;
															assign node3903 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node3906 = (inp[15]) ? 4'b0101 : node3907;
																assign node3907 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node3911 = (inp[12]) ? node3921 : node3912;
														assign node3912 = (inp[7]) ? node3918 : node3913;
															assign node3913 = (inp[4]) ? node3915 : 4'b0001;
																assign node3915 = (inp[15]) ? 4'b0111 : 4'b0001;
															assign node3918 = (inp[15]) ? 4'b0000 : 4'b0011;
														assign node3921 = (inp[7]) ? node3923 : 4'b0010;
															assign node3923 = (inp[4]) ? 4'b0001 : node3924;
																assign node3924 = (inp[15]) ? 4'b0001 : 4'b0100;
												assign node3928 = (inp[1]) ? node3942 : node3929;
													assign node3929 = (inp[7]) ? node3933 : node3930;
														assign node3930 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node3933 = (inp[4]) ? 4'b0001 : node3934;
															assign node3934 = (inp[12]) ? node3938 : node3935;
																assign node3935 = (inp[15]) ? 4'b0110 : 4'b0010;
																assign node3938 = (inp[15]) ? 4'b0001 : 4'b0100;
													assign node3942 = (inp[12]) ? node3952 : node3943;
														assign node3943 = (inp[7]) ? node3949 : node3944;
															assign node3944 = (inp[4]) ? node3946 : 4'b0101;
																assign node3946 = (inp[15]) ? 4'b0110 : 4'b0101;
															assign node3949 = (inp[15]) ? 4'b0101 : 4'b0110;
														assign node3952 = (inp[7]) ? node3956 : node3953;
															assign node3953 = (inp[4]) ? 4'b0101 : 4'b0110;
															assign node3956 = (inp[15]) ? 4'b0000 : node3957;
																assign node3957 = (inp[4]) ? 4'b0000 : 4'b0101;
											assign node3961 = (inp[15]) ? node3991 : node3962;
												assign node3962 = (inp[5]) ? node3974 : node3963;
													assign node3963 = (inp[12]) ? node3967 : node3964;
														assign node3964 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node3967 = (inp[7]) ? node3969 : 4'b0110;
															assign node3969 = (inp[4]) ? node3971 : 4'b0101;
																assign node3971 = (inp[1]) ? 4'b0101 : 4'b0000;
													assign node3974 = (inp[1]) ? node3982 : node3975;
														assign node3975 = (inp[7]) ? node3979 : node3976;
															assign node3976 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node3979 = (inp[12]) ? 4'b0001 : 4'b0110;
														assign node3982 = (inp[4]) ? node3988 : node3983;
															assign node3983 = (inp[12]) ? 4'b0010 : node3984;
																assign node3984 = (inp[7]) ? 4'b0010 : 4'b0001;
															assign node3988 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node3991 = (inp[1]) ? node4009 : node3992;
													assign node3992 = (inp[4]) ? node4004 : node3993;
														assign node3993 = (inp[7]) ? node3997 : node3994;
															assign node3994 = (inp[12]) ? 4'b0110 : 4'b0100;
															assign node3997 = (inp[12]) ? node4001 : node3998;
																assign node3998 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node4001 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node4004 = (inp[12]) ? 4'b0101 : node4005;
															assign node4005 = (inp[7]) ? 4'b0100 : 4'b0110;
													assign node4009 = (inp[7]) ? node4023 : node4010;
														assign node4010 = (inp[5]) ? node4018 : node4011;
															assign node4011 = (inp[12]) ? node4015 : node4012;
																assign node4012 = (inp[4]) ? 4'b0011 : 4'b0100;
																assign node4015 = (inp[4]) ? 4'b0100 : 4'b0111;
															assign node4018 = (inp[12]) ? node4020 : 4'b0001;
																assign node4020 = (inp[4]) ? 4'b0001 : 4'b0010;
														assign node4023 = (inp[12]) ? node4029 : node4024;
															assign node4024 = (inp[4]) ? 4'b0101 : node4025;
																assign node4025 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node4029 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node4032 = (inp[13]) ? node4100 : node4033;
											assign node4033 = (inp[5]) ? node4063 : node4034;
												assign node4034 = (inp[12]) ? node4050 : node4035;
													assign node4035 = (inp[4]) ? node4039 : node4036;
														assign node4036 = (inp[7]) ? 4'b0111 : 4'b0101;
														assign node4039 = (inp[1]) ? node4045 : node4040;
															assign node4040 = (inp[15]) ? node4042 : 4'b0100;
																assign node4042 = (inp[7]) ? 4'b0100 : 4'b0110;
															assign node4045 = (inp[15]) ? node4047 : 4'b0110;
																assign node4047 = (inp[7]) ? 4'b0101 : 4'b0011;
													assign node4050 = (inp[7]) ? node4058 : node4051;
														assign node4051 = (inp[4]) ? node4055 : node4052;
															assign node4052 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node4055 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node4058 = (inp[15]) ? 4'b0011 : node4059;
															assign node4059 = (inp[4]) ? 4'b0100 : 4'b0001;
												assign node4063 = (inp[12]) ? node4081 : node4064;
													assign node4064 = (inp[7]) ? node4070 : node4065;
														assign node4065 = (inp[4]) ? 4'b0011 : node4066;
															assign node4066 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node4070 = (inp[4]) ? node4076 : node4071;
															assign node4071 = (inp[1]) ? node4073 : 4'b0010;
																assign node4073 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node4076 = (inp[1]) ? node4078 : 4'b0111;
																assign node4078 = (inp[15]) ? 4'b0001 : 4'b0010;
													assign node4081 = (inp[7]) ? node4093 : node4082;
														assign node4082 = (inp[1]) ? node4088 : node4083;
															assign node4083 = (inp[15]) ? 4'b0101 : node4084;
																assign node4084 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node4088 = (inp[4]) ? 4'b0110 : node4089;
																assign node4089 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node4093 = (inp[4]) ? node4095 : 4'b0101;
															assign node4095 = (inp[15]) ? 4'b0110 : node4096;
																assign node4096 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node4100 = (inp[1]) ? node4132 : node4101;
												assign node4101 = (inp[15]) ? node4119 : node4102;
													assign node4102 = (inp[4]) ? node4110 : node4103;
														assign node4103 = (inp[7]) ? node4107 : node4104;
															assign node4104 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node4107 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node4110 = (inp[12]) ? node4112 : 4'b0010;
															assign node4112 = (inp[7]) ? node4116 : node4113;
																assign node4113 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node4116 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node4119 = (inp[12]) ? node4125 : node4120;
														assign node4120 = (inp[5]) ? node4122 : 4'b0011;
															assign node4122 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node4125 = (inp[7]) ? node4129 : node4126;
															assign node4126 = (inp[4]) ? 4'b0000 : 4'b0010;
															assign node4129 = (inp[4]) ? 4'b0110 : 4'b0000;
												assign node4132 = (inp[12]) ? node4148 : node4133;
													assign node4133 = (inp[4]) ? node4137 : node4134;
														assign node4134 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4137 = (inp[5]) ? node4141 : node4138;
															assign node4138 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node4141 = (inp[7]) ? node4145 : node4142;
																assign node4142 = (inp[15]) ? 4'b0110 : 4'b0101;
																assign node4145 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node4148 = (inp[7]) ? node4156 : node4149;
														assign node4149 = (inp[15]) ? 4'b0100 : node4150;
															assign node4150 = (inp[4]) ? 4'b0010 : node4151;
																assign node4151 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node4156 = (inp[15]) ? node4158 : 4'b0000;
															assign node4158 = (inp[4]) ? node4160 : 4'b0000;
																assign node4160 = (inp[5]) ? 4'b0010 : 4'b0110;
					assign node4163 = (inp[11]) ? node6325 : node4164;
						assign node4164 = (inp[12]) ? node5254 : node4165;
							assign node4165 = (inp[7]) ? node4703 : node4166;
								assign node4166 = (inp[15]) ? node4450 : node4167;
									assign node4167 = (inp[4]) ? node4297 : node4168;
										assign node4168 = (inp[0]) ? node4222 : node4169;
											assign node4169 = (inp[5]) ? node4201 : node4170;
												assign node4170 = (inp[1]) ? node4184 : node4171;
													assign node4171 = (inp[9]) ? node4179 : node4172;
														assign node4172 = (inp[10]) ? node4176 : node4173;
															assign node4173 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node4176 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node4179 = (inp[13]) ? 4'b1001 : node4180;
															assign node4180 = (inp[2]) ? 4'b1100 : 4'b1001;
													assign node4184 = (inp[10]) ? node4194 : node4185;
														assign node4185 = (inp[9]) ? node4191 : node4186;
															assign node4186 = (inp[13]) ? node4188 : 4'b1000;
																assign node4188 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node4191 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node4194 = (inp[9]) ? node4196 : 4'b1101;
															assign node4196 = (inp[13]) ? node4198 : 4'b1000;
																assign node4198 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node4201 = (inp[10]) ? node4211 : node4202;
													assign node4202 = (inp[9]) ? node4204 : 4'b1100;
														assign node4204 = (inp[13]) ? node4208 : node4205;
															assign node4205 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node4208 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node4211 = (inp[2]) ? node4217 : node4212;
														assign node4212 = (inp[13]) ? node4214 : 4'b1001;
															assign node4214 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node4217 = (inp[13]) ? node4219 : 4'b1100;
															assign node4219 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node4222 = (inp[13]) ? node4268 : node4223;
												assign node4223 = (inp[2]) ? node4251 : node4224;
													assign node4224 = (inp[1]) ? node4238 : node4225;
														assign node4225 = (inp[5]) ? node4233 : node4226;
															assign node4226 = (inp[10]) ? node4230 : node4227;
																assign node4227 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node4230 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node4233 = (inp[9]) ? 4'b1000 : node4234;
																assign node4234 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node4238 = (inp[5]) ? node4246 : node4239;
															assign node4239 = (inp[9]) ? node4243 : node4240;
																assign node4240 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node4243 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node4246 = (inp[10]) ? node4248 : 4'b1001;
																assign node4248 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node4251 = (inp[1]) ? node4259 : node4252;
														assign node4252 = (inp[10]) ? node4256 : node4253;
															assign node4253 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node4256 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node4259 = (inp[5]) ? node4263 : node4260;
															assign node4260 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node4263 = (inp[9]) ? node4265 : 4'b1101;
																assign node4265 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node4268 = (inp[2]) ? node4288 : node4269;
													assign node4269 = (inp[1]) ? node4279 : node4270;
														assign node4270 = (inp[5]) ? 4'b1101 : node4271;
															assign node4271 = (inp[10]) ? node4275 : node4272;
																assign node4272 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node4275 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node4279 = (inp[5]) ? node4285 : node4280;
															assign node4280 = (inp[9]) ? node4282 : 4'b1001;
																assign node4282 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node4285 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node4288 = (inp[1]) ? node4294 : node4289;
														assign node4289 = (inp[9]) ? 4'b1001 : node4290;
															assign node4290 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node4294 = (inp[5]) ? 4'b1000 : 4'b1101;
										assign node4297 = (inp[1]) ? node4383 : node4298;
											assign node4298 = (inp[5]) ? node4352 : node4299;
												assign node4299 = (inp[0]) ? node4329 : node4300;
													assign node4300 = (inp[2]) ? node4316 : node4301;
														assign node4301 = (inp[13]) ? node4309 : node4302;
															assign node4302 = (inp[10]) ? node4306 : node4303;
																assign node4303 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node4306 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node4309 = (inp[10]) ? node4313 : node4310;
																assign node4310 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node4313 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node4316 = (inp[13]) ? node4324 : node4317;
															assign node4317 = (inp[10]) ? node4321 : node4318;
																assign node4318 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node4321 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node4324 = (inp[10]) ? node4326 : 4'b1010;
																assign node4326 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node4329 = (inp[10]) ? node4345 : node4330;
														assign node4330 = (inp[2]) ? node4338 : node4331;
															assign node4331 = (inp[13]) ? node4335 : node4332;
																assign node4332 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node4335 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node4338 = (inp[13]) ? node4342 : node4339;
																assign node4339 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node4342 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node4345 = (inp[9]) ? 4'b1011 : node4346;
															assign node4346 = (inp[13]) ? 4'b1010 : node4347;
																assign node4347 = (inp[2]) ? 4'b1111 : 4'b1010;
												assign node4352 = (inp[10]) ? node4364 : node4353;
													assign node4353 = (inp[13]) ? node4361 : node4354;
														assign node4354 = (inp[2]) ? node4358 : node4355;
															assign node4355 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node4358 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node4361 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node4364 = (inp[9]) ? node4372 : node4365;
														assign node4365 = (inp[2]) ? node4369 : node4366;
															assign node4366 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node4369 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node4372 = (inp[0]) ? node4380 : node4373;
															assign node4373 = (inp[2]) ? node4377 : node4374;
																assign node4374 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node4377 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node4380 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node4383 = (inp[5]) ? node4417 : node4384;
												assign node4384 = (inp[13]) ? node4398 : node4385;
													assign node4385 = (inp[2]) ? node4391 : node4386;
														assign node4386 = (inp[10]) ? 4'b1111 : node4387;
															assign node4387 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node4391 = (inp[10]) ? node4395 : node4392;
															assign node4392 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node4395 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node4398 = (inp[2]) ? node4406 : node4399;
														assign node4399 = (inp[0]) ? 4'b1010 : node4400;
															assign node4400 = (inp[9]) ? 4'b1010 : node4401;
																assign node4401 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node4406 = (inp[9]) ? node4412 : node4407;
															assign node4407 = (inp[10]) ? node4409 : 4'b1110;
																assign node4409 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node4412 = (inp[10]) ? node4414 : 4'b1111;
																assign node4414 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node4417 = (inp[13]) ? node4429 : node4418;
													assign node4418 = (inp[2]) ? 4'b1110 : node4419;
														assign node4419 = (inp[0]) ? node4421 : 4'b1010;
															assign node4421 = (inp[9]) ? node4425 : node4422;
																assign node4422 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node4425 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node4429 = (inp[2]) ? node4437 : node4430;
														assign node4430 = (inp[10]) ? node4434 : node4431;
															assign node4431 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node4434 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node4437 = (inp[9]) ? node4445 : node4438;
															assign node4438 = (inp[10]) ? node4442 : node4439;
																assign node4439 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node4442 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node4445 = (inp[10]) ? 4'b1010 : node4446;
																assign node4446 = (inp[0]) ? 4'b1011 : 4'b1010;
									assign node4450 = (inp[13]) ? node4574 : node4451;
										assign node4451 = (inp[2]) ? node4509 : node4452;
											assign node4452 = (inp[4]) ? node4480 : node4453;
												assign node4453 = (inp[1]) ? node4475 : node4454;
													assign node4454 = (inp[5]) ? node4468 : node4455;
														assign node4455 = (inp[9]) ? node4463 : node4456;
															assign node4456 = (inp[10]) ? node4460 : node4457;
																assign node4457 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node4460 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node4463 = (inp[0]) ? 4'b1001 : node4464;
																assign node4464 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node4468 = (inp[0]) ? node4470 : 4'b1001;
															assign node4470 = (inp[9]) ? node4472 : 4'b1001;
																assign node4472 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node4475 = (inp[5]) ? node4477 : 4'b1101;
														assign node4477 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node4480 = (inp[1]) ? node4500 : node4481;
													assign node4481 = (inp[9]) ? node4491 : node4482;
														assign node4482 = (inp[5]) ? 4'b1101 : node4483;
															assign node4483 = (inp[0]) ? node4487 : node4484;
																assign node4484 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node4487 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node4491 = (inp[0]) ? node4495 : node4492;
															assign node4492 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node4495 = (inp[10]) ? node4497 : 4'b1100;
																assign node4497 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node4500 = (inp[5]) ? node4504 : node4501;
														assign node4501 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node4504 = (inp[10]) ? 4'b1100 : node4505;
															assign node4505 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node4509 = (inp[4]) ? node4543 : node4510;
												assign node4510 = (inp[1]) ? node4526 : node4511;
													assign node4511 = (inp[9]) ? node4519 : node4512;
														assign node4512 = (inp[10]) ? node4516 : node4513;
															assign node4513 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node4516 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node4519 = (inp[10]) ? node4523 : node4520;
															assign node4520 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node4523 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node4526 = (inp[5]) ? node4536 : node4527;
														assign node4527 = (inp[9]) ? node4529 : 4'b1001;
															assign node4529 = (inp[10]) ? node4533 : node4530;
																assign node4530 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node4533 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node4536 = (inp[10]) ? 4'b1101 : node4537;
															assign node4537 = (inp[0]) ? 4'b1100 : node4538;
																assign node4538 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node4543 = (inp[1]) ? node4559 : node4544;
													assign node4544 = (inp[10]) ? node4550 : node4545;
														assign node4545 = (inp[9]) ? node4547 : 4'b1001;
															assign node4547 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node4550 = (inp[0]) ? 4'b1000 : node4551;
															assign node4551 = (inp[9]) ? node4555 : node4552;
																assign node4552 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node4555 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node4559 = (inp[5]) ? node4569 : node4560;
														assign node4560 = (inp[0]) ? 4'b1101 : node4561;
															assign node4561 = (inp[9]) ? node4565 : node4562;
																assign node4562 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node4565 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node4569 = (inp[9]) ? node4571 : 4'b1000;
															assign node4571 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node4574 = (inp[10]) ? node4622 : node4575;
											assign node4575 = (inp[9]) ? node4595 : node4576;
												assign node4576 = (inp[2]) ? node4588 : node4577;
													assign node4577 = (inp[5]) ? node4583 : node4578;
														assign node4578 = (inp[0]) ? node4580 : 4'b1000;
															assign node4580 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node4583 = (inp[4]) ? node4585 : 4'b1101;
															assign node4585 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node4588 = (inp[5]) ? node4590 : 4'b1001;
														assign node4590 = (inp[4]) ? node4592 : 4'b1000;
															assign node4592 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node4595 = (inp[1]) ? node4609 : node4596;
													assign node4596 = (inp[4]) ? node4602 : node4597;
														assign node4597 = (inp[2]) ? node4599 : 4'b1100;
															assign node4599 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node4602 = (inp[2]) ? node4606 : node4603;
															assign node4603 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node4606 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node4609 = (inp[4]) ? node4617 : node4610;
														assign node4610 = (inp[5]) ? node4614 : node4611;
															assign node4611 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node4614 = (inp[2]) ? 4'b1000 : 4'b1101;
														assign node4617 = (inp[2]) ? node4619 : 4'b1000;
															assign node4619 = (inp[5]) ? 4'b1101 : 4'b1000;
											assign node4622 = (inp[0]) ? node4666 : node4623;
												assign node4623 = (inp[5]) ? node4645 : node4624;
													assign node4624 = (inp[9]) ? node4638 : node4625;
														assign node4625 = (inp[1]) ? node4631 : node4626;
															assign node4626 = (inp[4]) ? node4628 : 4'b1100;
																assign node4628 = (inp[2]) ? 4'b1100 : 4'b1001;
															assign node4631 = (inp[2]) ? node4635 : node4632;
																assign node4632 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node4635 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node4638 = (inp[1]) ? node4640 : 4'b1101;
															assign node4640 = (inp[4]) ? 4'b1100 : node4641;
																assign node4641 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node4645 = (inp[2]) ? node4659 : node4646;
														assign node4646 = (inp[4]) ? node4654 : node4647;
															assign node4647 = (inp[1]) ? node4651 : node4648;
																assign node4648 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node4651 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node4654 = (inp[9]) ? node4656 : 4'b1000;
																assign node4656 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node4659 = (inp[4]) ? node4661 : 4'b1000;
															assign node4661 = (inp[9]) ? 4'b1100 : node4662;
																assign node4662 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node4666 = (inp[1]) ? node4678 : node4667;
													assign node4667 = (inp[9]) ? node4673 : node4668;
														assign node4668 = (inp[4]) ? 4'b1000 : node4669;
															assign node4669 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node4673 = (inp[2]) ? node4675 : 4'b1001;
															assign node4675 = (inp[4]) ? 4'b1100 : 4'b1001;
													assign node4678 = (inp[9]) ? node4690 : node4679;
														assign node4679 = (inp[4]) ? node4683 : node4680;
															assign node4680 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node4683 = (inp[2]) ? node4687 : node4684;
																assign node4684 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node4687 = (inp[5]) ? 4'b1101 : 4'b1000;
														assign node4690 = (inp[4]) ? node4698 : node4691;
															assign node4691 = (inp[2]) ? node4695 : node4692;
																assign node4692 = (inp[5]) ? 4'b1100 : 4'b1000;
																assign node4695 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node4698 = (inp[5]) ? node4700 : 4'b1100;
																assign node4700 = (inp[2]) ? 4'b1100 : 4'b1001;
								assign node4703 = (inp[15]) ? node4967 : node4704;
									assign node4704 = (inp[4]) ? node4842 : node4705;
										assign node4705 = (inp[5]) ? node4785 : node4706;
											assign node4706 = (inp[0]) ? node4750 : node4707;
												assign node4707 = (inp[1]) ? node4727 : node4708;
													assign node4708 = (inp[9]) ? node4716 : node4709;
														assign node4709 = (inp[10]) ? node4713 : node4710;
															assign node4710 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node4713 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node4716 = (inp[10]) ? node4720 : node4717;
															assign node4717 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node4720 = (inp[2]) ? node4724 : node4721;
																assign node4721 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node4724 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node4727 = (inp[9]) ? node4737 : node4728;
														assign node4728 = (inp[2]) ? node4734 : node4729;
															assign node4729 = (inp[13]) ? node4731 : 4'b1011;
																assign node4731 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node4734 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node4737 = (inp[2]) ? node4743 : node4738;
															assign node4738 = (inp[13]) ? node4740 : 4'b1010;
																assign node4740 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node4743 = (inp[13]) ? node4747 : node4744;
																assign node4744 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node4747 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node4750 = (inp[1]) ? node4772 : node4751;
													assign node4751 = (inp[9]) ? node4759 : node4752;
														assign node4752 = (inp[13]) ? 4'b1110 : node4753;
															assign node4753 = (inp[2]) ? node4755 : 4'b1011;
																assign node4755 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node4759 = (inp[2]) ? node4765 : node4760;
															assign node4760 = (inp[13]) ? 4'b1111 : node4761;
																assign node4761 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node4765 = (inp[13]) ? node4769 : node4766;
																assign node4766 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node4769 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node4772 = (inp[2]) ? node4776 : node4773;
														assign node4773 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node4776 = (inp[13]) ? node4780 : node4777;
															assign node4777 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node4780 = (inp[9]) ? node4782 : 4'b1010;
																assign node4782 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node4785 = (inp[10]) ? node4805 : node4786;
												assign node4786 = (inp[9]) ? node4800 : node4787;
													assign node4787 = (inp[13]) ? node4793 : node4788;
														assign node4788 = (inp[1]) ? node4790 : 4'b1011;
															assign node4790 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node4793 = (inp[0]) ? 4'b1011 : node4794;
															assign node4794 = (inp[1]) ? node4796 : 4'b1110;
																assign node4796 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node4800 = (inp[13]) ? node4802 : 4'b1010;
														assign node4802 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node4805 = (inp[1]) ? node4827 : node4806;
													assign node4806 = (inp[9]) ? node4816 : node4807;
														assign node4807 = (inp[2]) ? node4813 : node4808;
															assign node4808 = (inp[13]) ? node4810 : 4'b1110;
																assign node4810 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node4813 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node4816 = (inp[0]) ? node4822 : node4817;
															assign node4817 = (inp[13]) ? node4819 : 4'b1111;
																assign node4819 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node4822 = (inp[2]) ? 4'b1011 : node4823;
																assign node4823 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node4827 = (inp[13]) ? node4833 : node4828;
														assign node4828 = (inp[9]) ? node4830 : 4'b1110;
															assign node4830 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node4833 = (inp[2]) ? node4839 : node4834;
															assign node4834 = (inp[0]) ? 4'b1111 : node4835;
																assign node4835 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node4839 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node4842 = (inp[1]) ? node4890 : node4843;
											assign node4843 = (inp[2]) ? node4867 : node4844;
												assign node4844 = (inp[13]) ? node4858 : node4845;
													assign node4845 = (inp[0]) ? 4'b1101 : node4846;
														assign node4846 = (inp[5]) ? node4852 : node4847;
															assign node4847 = (inp[9]) ? 4'b1101 : node4848;
																assign node4848 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node4852 = (inp[10]) ? 4'b1100 : node4853;
																assign node4853 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node4858 = (inp[5]) ? 4'b1001 : node4859;
														assign node4859 = (inp[9]) ? 4'b1000 : node4860;
															assign node4860 = (inp[0]) ? 4'b1001 : node4861;
																assign node4861 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node4867 = (inp[13]) ? node4879 : node4868;
													assign node4868 = (inp[9]) ? 4'b1000 : node4869;
														assign node4869 = (inp[10]) ? node4873 : node4870;
															assign node4870 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node4873 = (inp[0]) ? node4875 : 4'b1000;
																assign node4875 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node4879 = (inp[0]) ? node4887 : node4880;
														assign node4880 = (inp[9]) ? node4882 : 4'b1100;
															assign node4882 = (inp[10]) ? node4884 : 4'b1100;
																assign node4884 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node4887 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node4890 = (inp[0]) ? node4924 : node4891;
												assign node4891 = (inp[13]) ? node4909 : node4892;
													assign node4892 = (inp[2]) ? node4902 : node4893;
														assign node4893 = (inp[5]) ? node4899 : node4894;
															assign node4894 = (inp[10]) ? node4896 : 4'b1000;
																assign node4896 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node4899 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node4902 = (inp[5]) ? node4904 : 4'b1101;
															assign node4904 = (inp[9]) ? 4'b1001 : node4905;
																assign node4905 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node4909 = (inp[9]) ? node4917 : node4910;
														assign node4910 = (inp[5]) ? node4914 : node4911;
															assign node4911 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node4914 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node4917 = (inp[2]) ? node4921 : node4918;
															assign node4918 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node4921 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node4924 = (inp[9]) ? node4938 : node4925;
													assign node4925 = (inp[10]) ? node4931 : node4926;
														assign node4926 = (inp[5]) ? node4928 : 4'b1000;
															assign node4928 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node4931 = (inp[5]) ? node4935 : node4932;
															assign node4932 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node4935 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node4938 = (inp[13]) ? node4954 : node4939;
														assign node4939 = (inp[10]) ? node4947 : node4940;
															assign node4940 = (inp[2]) ? node4944 : node4941;
																assign node4941 = (inp[5]) ? 4'b1100 : 4'b1001;
																assign node4944 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node4947 = (inp[2]) ? node4951 : node4948;
																assign node4948 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node4951 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node4954 = (inp[10]) ? node4960 : node4955;
															assign node4955 = (inp[5]) ? 4'b1100 : node4956;
																assign node4956 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node4960 = (inp[5]) ? node4964 : node4961;
																assign node4961 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node4964 = (inp[2]) ? 4'b1101 : 4'b1000;
									assign node4967 = (inp[1]) ? node5119 : node4968;
										assign node4968 = (inp[10]) ? node5046 : node4969;
											assign node4969 = (inp[9]) ? node5007 : node4970;
												assign node4970 = (inp[5]) ? node4990 : node4971;
													assign node4971 = (inp[4]) ? node4981 : node4972;
														assign node4972 = (inp[0]) ? node4978 : node4973;
															assign node4973 = (inp[13]) ? node4975 : 4'b1010;
																assign node4975 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node4978 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node4981 = (inp[2]) ? node4987 : node4982;
															assign node4982 = (inp[13]) ? node4984 : 4'b1010;
																assign node4984 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node4987 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node4990 = (inp[4]) ? node5000 : node4991;
														assign node4991 = (inp[2]) ? node4997 : node4992;
															assign node4992 = (inp[0]) ? 4'b1110 : node4993;
																assign node4993 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node4997 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node5000 = (inp[0]) ? node5002 : 4'b1010;
															assign node5002 = (inp[2]) ? node5004 : 4'b1011;
																assign node5004 = (inp[13]) ? 4'b1110 : 4'b1011;
												assign node5007 = (inp[4]) ? node5029 : node5008;
													assign node5008 = (inp[5]) ? node5022 : node5009;
														assign node5009 = (inp[0]) ? node5017 : node5010;
															assign node5010 = (inp[13]) ? node5014 : node5011;
																assign node5011 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node5014 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node5017 = (inp[13]) ? 4'b1110 : node5018;
																assign node5018 = (inp[2]) ? 4'b1011 : 4'b1110;
														assign node5022 = (inp[13]) ? node5026 : node5023;
															assign node5023 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node5026 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5029 = (inp[13]) ? node5033 : node5030;
														assign node5030 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node5033 = (inp[2]) ? node5041 : node5034;
															assign node5034 = (inp[5]) ? node5038 : node5035;
																assign node5035 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node5038 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node5041 = (inp[5]) ? node5043 : 4'b1010;
																assign node5043 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5046 = (inp[9]) ? node5084 : node5047;
												assign node5047 = (inp[5]) ? node5067 : node5048;
													assign node5048 = (inp[13]) ? node5056 : node5049;
														assign node5049 = (inp[2]) ? 4'b1011 : node5050;
															assign node5050 = (inp[4]) ? 4'b1011 : node5051;
																assign node5051 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5056 = (inp[0]) ? node5060 : node5057;
															assign node5057 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node5060 = (inp[4]) ? node5064 : node5061;
																assign node5061 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node5064 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node5067 = (inp[4]) ? node5077 : node5068;
														assign node5068 = (inp[0]) ? 4'b1010 : node5069;
															assign node5069 = (inp[13]) ? node5073 : node5070;
																assign node5070 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node5073 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node5077 = (inp[13]) ? node5079 : 4'b1010;
															assign node5079 = (inp[2]) ? 4'b1111 : node5080;
																assign node5080 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5084 = (inp[5]) ? node5106 : node5085;
													assign node5085 = (inp[0]) ? node5095 : node5086;
														assign node5086 = (inp[13]) ? node5088 : 4'b1010;
															assign node5088 = (inp[2]) ? node5092 : node5089;
																assign node5089 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node5092 = (inp[4]) ? 4'b1011 : 4'b1110;
														assign node5095 = (inp[13]) ? node5103 : node5096;
															assign node5096 = (inp[2]) ? node5100 : node5097;
																assign node5097 = (inp[4]) ? 4'b1010 : 4'b1111;
																assign node5100 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node5103 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node5106 = (inp[2]) ? node5114 : node5107;
														assign node5107 = (inp[4]) ? node5111 : node5108;
															assign node5108 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node5111 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node5114 = (inp[4]) ? 4'b1011 : node5115;
															assign node5115 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node5119 = (inp[13]) ? node5183 : node5120;
											assign node5120 = (inp[9]) ? node5146 : node5121;
												assign node5121 = (inp[4]) ? node5137 : node5122;
													assign node5122 = (inp[2]) ? node5130 : node5123;
														assign node5123 = (inp[5]) ? 4'b1110 : node5124;
															assign node5124 = (inp[0]) ? 4'b1111 : node5125;
																assign node5125 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5130 = (inp[10]) ? node5134 : node5131;
															assign node5131 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node5134 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node5137 = (inp[2]) ? node5141 : node5138;
														assign node5138 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5141 = (inp[10]) ? node5143 : 4'b1110;
															assign node5143 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node5146 = (inp[4]) ? node5166 : node5147;
													assign node5147 = (inp[2]) ? node5161 : node5148;
														assign node5148 = (inp[10]) ? node5154 : node5149;
															assign node5149 = (inp[5]) ? 4'b1110 : node5150;
																assign node5150 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5154 = (inp[5]) ? node5158 : node5155;
																assign node5155 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node5158 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node5161 = (inp[5]) ? node5163 : 4'b1010;
															assign node5163 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node5166 = (inp[2]) ? node5174 : node5167;
														assign node5167 = (inp[10]) ? node5169 : 4'b1010;
															assign node5169 = (inp[5]) ? node5171 : 4'b1011;
																assign node5171 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node5174 = (inp[10]) ? node5180 : node5175;
															assign node5175 = (inp[0]) ? node5177 : 4'b1111;
																assign node5177 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node5180 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5183 = (inp[4]) ? node5221 : node5184;
												assign node5184 = (inp[2]) ? node5198 : node5185;
													assign node5185 = (inp[10]) ? node5191 : node5186;
														assign node5186 = (inp[5]) ? 4'b1010 : node5187;
															assign node5187 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node5191 = (inp[9]) ? 4'b1011 : node5192;
															assign node5192 = (inp[0]) ? 4'b1011 : node5193;
																assign node5193 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node5198 = (inp[10]) ? node5208 : node5199;
														assign node5199 = (inp[9]) ? 4'b1111 : node5200;
															assign node5200 = (inp[0]) ? node5204 : node5201;
																assign node5201 = (inp[5]) ? 4'b1110 : 4'b1111;
																assign node5204 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node5208 = (inp[0]) ? node5216 : node5209;
															assign node5209 = (inp[5]) ? node5213 : node5210;
																assign node5210 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node5213 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node5216 = (inp[5]) ? 4'b1110 : node5217;
																assign node5217 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node5221 = (inp[2]) ? node5235 : node5222;
													assign node5222 = (inp[5]) ? node5228 : node5223;
														assign node5223 = (inp[0]) ? node5225 : 4'b1111;
															assign node5225 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5228 = (inp[10]) ? node5232 : node5229;
															assign node5229 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node5232 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node5235 = (inp[10]) ? node5245 : node5236;
														assign node5236 = (inp[5]) ? node5238 : 4'b1010;
															assign node5238 = (inp[0]) ? node5242 : node5239;
																assign node5239 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node5242 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node5245 = (inp[9]) ? node5251 : node5246;
															assign node5246 = (inp[5]) ? node5248 : 4'b1011;
																assign node5248 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node5251 = (inp[0]) ? 4'b1011 : 4'b1010;
							assign node5254 = (inp[7]) ? node5792 : node5255;
								assign node5255 = (inp[4]) ? node5529 : node5256;
									assign node5256 = (inp[0]) ? node5400 : node5257;
										assign node5257 = (inp[13]) ? node5331 : node5258;
											assign node5258 = (inp[2]) ? node5294 : node5259;
												assign node5259 = (inp[1]) ? node5279 : node5260;
													assign node5260 = (inp[15]) ? node5266 : node5261;
														assign node5261 = (inp[9]) ? node5263 : 4'b1010;
															assign node5263 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node5266 = (inp[5]) ? node5274 : node5267;
															assign node5267 = (inp[9]) ? node5271 : node5268;
																assign node5268 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node5271 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node5274 = (inp[10]) ? 4'b1011 : node5275;
																assign node5275 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node5279 = (inp[5]) ? node5287 : node5280;
														assign node5280 = (inp[15]) ? 4'b1111 : node5281;
															assign node5281 = (inp[10]) ? node5283 : 4'b1110;
																assign node5283 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node5287 = (inp[10]) ? 4'b1011 : node5288;
															assign node5288 = (inp[9]) ? 4'b1010 : node5289;
																assign node5289 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node5294 = (inp[1]) ? node5308 : node5295;
													assign node5295 = (inp[5]) ? node5303 : node5296;
														assign node5296 = (inp[10]) ? node5300 : node5297;
															assign node5297 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node5300 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node5303 = (inp[10]) ? 4'b1111 : node5304;
															assign node5304 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node5308 = (inp[5]) ? node5322 : node5309;
														assign node5309 = (inp[10]) ? node5315 : node5310;
															assign node5310 = (inp[9]) ? node5312 : 4'b1011;
																assign node5312 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node5315 = (inp[15]) ? node5319 : node5316;
																assign node5316 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node5319 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node5322 = (inp[10]) ? node5324 : 4'b1111;
															assign node5324 = (inp[15]) ? node5328 : node5325;
																assign node5325 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node5328 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node5331 = (inp[2]) ? node5371 : node5332;
												assign node5332 = (inp[5]) ? node5350 : node5333;
													assign node5333 = (inp[1]) ? node5341 : node5334;
														assign node5334 = (inp[15]) ? node5336 : 4'b1110;
															assign node5336 = (inp[9]) ? node5338 : 4'b1111;
																assign node5338 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5341 = (inp[9]) ? 4'b1010 : node5342;
															assign node5342 = (inp[15]) ? node5346 : node5343;
																assign node5343 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node5346 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node5350 = (inp[1]) ? node5358 : node5351;
														assign node5351 = (inp[15]) ? node5353 : 4'b1110;
															assign node5353 = (inp[9]) ? node5355 : 4'b1110;
																assign node5355 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5358 = (inp[9]) ? node5366 : node5359;
															assign node5359 = (inp[15]) ? node5363 : node5360;
																assign node5360 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node5363 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node5366 = (inp[15]) ? node5368 : 4'b1111;
																assign node5368 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node5371 = (inp[5]) ? node5385 : node5372;
													assign node5372 = (inp[1]) ? node5378 : node5373;
														assign node5373 = (inp[10]) ? 4'b1010 : node5374;
															assign node5374 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node5378 = (inp[9]) ? node5380 : 4'b1110;
															assign node5380 = (inp[10]) ? node5382 : 4'b1111;
																assign node5382 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node5385 = (inp[1]) ? node5387 : 4'b1011;
														assign node5387 = (inp[15]) ? node5395 : node5388;
															assign node5388 = (inp[10]) ? node5392 : node5389;
																assign node5389 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node5392 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node5395 = (inp[10]) ? node5397 : 4'b1010;
																assign node5397 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node5400 = (inp[9]) ? node5466 : node5401;
											assign node5401 = (inp[10]) ? node5429 : node5402;
												assign node5402 = (inp[15]) ? node5416 : node5403;
													assign node5403 = (inp[1]) ? node5407 : node5404;
														assign node5404 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node5407 = (inp[5]) ? node5413 : node5408;
															assign node5408 = (inp[13]) ? node5410 : 4'b1011;
																assign node5410 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node5413 = (inp[13]) ? 4'b1010 : 4'b1111;
													assign node5416 = (inp[5]) ? 4'b1111 : node5417;
														assign node5417 = (inp[1]) ? node5423 : node5418;
															assign node5418 = (inp[13]) ? node5420 : 4'b1111;
																assign node5420 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node5423 = (inp[13]) ? node5425 : 4'b1011;
																assign node5425 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node5429 = (inp[15]) ? node5449 : node5430;
													assign node5430 = (inp[13]) ? node5442 : node5431;
														assign node5431 = (inp[2]) ? node5437 : node5432;
															assign node5432 = (inp[1]) ? node5434 : 4'b1010;
																assign node5434 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node5437 = (inp[5]) ? 4'b1110 : node5438;
																assign node5438 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node5442 = (inp[2]) ? 4'b1011 : node5443;
															assign node5443 = (inp[1]) ? node5445 : 4'b1111;
																assign node5445 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node5449 = (inp[5]) ? node5459 : node5450;
														assign node5450 = (inp[1]) ? 4'b1110 : node5451;
															assign node5451 = (inp[13]) ? node5455 : node5452;
																assign node5452 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node5455 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node5459 = (inp[2]) ? node5463 : node5460;
															assign node5460 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node5463 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node5466 = (inp[10]) ? node5496 : node5467;
												assign node5467 = (inp[15]) ? node5481 : node5468;
													assign node5468 = (inp[2]) ? node5478 : node5469;
														assign node5469 = (inp[1]) ? node5471 : 4'b1010;
															assign node5471 = (inp[5]) ? node5475 : node5472;
																assign node5472 = (inp[13]) ? 4'b1010 : 4'b1111;
																assign node5475 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node5478 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node5481 = (inp[5]) ? node5489 : node5482;
														assign node5482 = (inp[1]) ? node5484 : 4'b1010;
															assign node5484 = (inp[2]) ? node5486 : 4'b1010;
																assign node5486 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node5489 = (inp[13]) ? node5493 : node5490;
															assign node5490 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node5493 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node5496 = (inp[15]) ? node5512 : node5497;
													assign node5497 = (inp[13]) ? node5505 : node5498;
														assign node5498 = (inp[2]) ? 4'b1111 : node5499;
															assign node5499 = (inp[5]) ? 4'b1011 : node5500;
																assign node5500 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node5505 = (inp[1]) ? node5509 : node5506;
															assign node5506 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node5509 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node5512 = (inp[1]) ? node5520 : node5513;
														assign node5513 = (inp[13]) ? node5517 : node5514;
															assign node5514 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node5517 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node5520 = (inp[13]) ? 4'b1011 : node5521;
															assign node5521 = (inp[2]) ? node5525 : node5522;
																assign node5522 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node5525 = (inp[5]) ? 4'b1111 : 4'b1011;
									assign node5529 = (inp[15]) ? node5669 : node5530;
										assign node5530 = (inp[10]) ? node5604 : node5531;
											assign node5531 = (inp[2]) ? node5561 : node5532;
												assign node5532 = (inp[13]) ? node5546 : node5533;
													assign node5533 = (inp[1]) ? node5541 : node5534;
														assign node5534 = (inp[5]) ? node5536 : 4'b1100;
															assign node5536 = (inp[9]) ? node5538 : 4'b1000;
																assign node5538 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node5541 = (inp[5]) ? 4'b1101 : node5542;
															assign node5542 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node5546 = (inp[5]) ? node5554 : node5547;
														assign node5547 = (inp[9]) ? node5551 : node5548;
															assign node5548 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node5551 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node5554 = (inp[1]) ? node5558 : node5555;
															assign node5555 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node5558 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node5561 = (inp[13]) ? node5585 : node5562;
													assign node5562 = (inp[5]) ? node5574 : node5563;
														assign node5563 = (inp[9]) ? node5569 : node5564;
															assign node5564 = (inp[1]) ? node5566 : 4'b1001;
																assign node5566 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node5569 = (inp[0]) ? node5571 : 4'b1000;
																assign node5571 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node5574 = (inp[1]) ? node5582 : node5575;
															assign node5575 = (inp[0]) ? node5579 : node5576;
																assign node5576 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node5579 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node5582 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node5585 = (inp[1]) ? node5595 : node5586;
														assign node5586 = (inp[5]) ? node5592 : node5587;
															assign node5587 = (inp[9]) ? 4'b1101 : node5588;
																assign node5588 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5592 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node5595 = (inp[9]) ? node5599 : node5596;
															assign node5596 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5599 = (inp[0]) ? 4'b1100 : node5600;
																assign node5600 = (inp[5]) ? 4'b1101 : 4'b1100;
											assign node5604 = (inp[9]) ? node5638 : node5605;
												assign node5605 = (inp[0]) ? node5625 : node5606;
													assign node5606 = (inp[13]) ? node5618 : node5607;
														assign node5607 = (inp[1]) ? node5615 : node5608;
															assign node5608 = (inp[2]) ? node5612 : node5609;
																assign node5609 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node5612 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node5615 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node5618 = (inp[1]) ? node5622 : node5619;
															assign node5619 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node5622 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node5625 = (inp[1]) ? node5633 : node5626;
														assign node5626 = (inp[13]) ? 4'b1100 : node5627;
															assign node5627 = (inp[2]) ? node5629 : 4'b1100;
																assign node5629 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node5633 = (inp[5]) ? node5635 : 4'b1100;
															assign node5635 = (inp[2]) ? 4'b1100 : 4'b1001;
												assign node5638 = (inp[13]) ? node5656 : node5639;
													assign node5639 = (inp[2]) ? node5649 : node5640;
														assign node5640 = (inp[1]) ? 4'b1101 : node5641;
															assign node5641 = (inp[5]) ? node5645 : node5642;
																assign node5642 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node5645 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5649 = (inp[5]) ? 4'b1100 : node5650;
															assign node5650 = (inp[0]) ? node5652 : 4'b1001;
																assign node5652 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node5656 = (inp[2]) ? node5664 : node5657;
														assign node5657 = (inp[1]) ? node5659 : 4'b1101;
															assign node5659 = (inp[5]) ? node5661 : 4'b1000;
																assign node5661 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5664 = (inp[0]) ? node5666 : 4'b1100;
															assign node5666 = (inp[1]) ? 4'b1101 : 4'b1000;
										assign node5669 = (inp[13]) ? node5729 : node5670;
											assign node5670 = (inp[2]) ? node5704 : node5671;
												assign node5671 = (inp[5]) ? node5691 : node5672;
													assign node5672 = (inp[1]) ? node5678 : node5673;
														assign node5673 = (inp[10]) ? node5675 : 4'b1011;
															assign node5675 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node5678 = (inp[9]) ? node5684 : node5679;
															assign node5679 = (inp[0]) ? node5681 : 4'b1110;
																assign node5681 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node5684 = (inp[0]) ? node5688 : node5685;
																assign node5685 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node5688 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5691 = (inp[0]) ? node5697 : node5692;
														assign node5692 = (inp[9]) ? node5694 : 4'b1011;
															assign node5694 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node5697 = (inp[10]) ? node5701 : node5698;
															assign node5698 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node5701 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node5704 = (inp[5]) ? node5714 : node5705;
													assign node5705 = (inp[1]) ? node5709 : node5706;
														assign node5706 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node5709 = (inp[10]) ? 4'b1010 : node5710;
															assign node5710 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node5714 = (inp[10]) ? 4'b1110 : node5715;
														assign node5715 = (inp[1]) ? node5723 : node5716;
															assign node5716 = (inp[0]) ? node5720 : node5717;
																assign node5717 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node5720 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node5723 = (inp[9]) ? 4'b1111 : node5724;
																assign node5724 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5729 = (inp[2]) ? node5763 : node5730;
												assign node5730 = (inp[5]) ? node5748 : node5731;
													assign node5731 = (inp[1]) ? node5741 : node5732;
														assign node5732 = (inp[9]) ? 4'b1110 : node5733;
															assign node5733 = (inp[0]) ? node5737 : node5734;
																assign node5734 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node5737 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5741 = (inp[0]) ? node5745 : node5742;
															assign node5742 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node5745 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node5748 = (inp[0]) ? node5756 : node5749;
														assign node5749 = (inp[9]) ? node5753 : node5750;
															assign node5750 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node5753 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5756 = (inp[9]) ? node5760 : node5757;
															assign node5757 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node5760 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node5763 = (inp[5]) ? node5777 : node5764;
													assign node5764 = (inp[1]) ? node5770 : node5765;
														assign node5765 = (inp[10]) ? node5767 : 4'b1010;
															assign node5767 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node5770 = (inp[10]) ? node5772 : 4'b1110;
															assign node5772 = (inp[0]) ? 4'b1111 : node5773;
																assign node5773 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node5777 = (inp[10]) ? node5785 : node5778;
														assign node5778 = (inp[9]) ? node5782 : node5779;
															assign node5779 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node5782 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node5785 = (inp[9]) ? node5789 : node5786;
															assign node5786 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node5789 = (inp[0]) ? 4'b1011 : 4'b1010;
								assign node5792 = (inp[15]) ? node6050 : node5793;
									assign node5793 = (inp[4]) ? node5901 : node5794;
										assign node5794 = (inp[2]) ? node5850 : node5795;
											assign node5795 = (inp[13]) ? node5823 : node5796;
												assign node5796 = (inp[5]) ? node5810 : node5797;
													assign node5797 = (inp[1]) ? node5803 : node5798;
														assign node5798 = (inp[0]) ? node5800 : 4'b1101;
															assign node5800 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node5803 = (inp[9]) ? node5805 : 4'b1000;
															assign node5805 = (inp[0]) ? 4'b1001 : node5806;
																assign node5806 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node5810 = (inp[9]) ? node5816 : node5811;
														assign node5811 = (inp[10]) ? 4'b1100 : node5812;
															assign node5812 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5816 = (inp[10]) ? 4'b1101 : node5817;
															assign node5817 = (inp[0]) ? node5819 : 4'b1100;
																assign node5819 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node5823 = (inp[5]) ? node5837 : node5824;
													assign node5824 = (inp[1]) ? node5830 : node5825;
														assign node5825 = (inp[10]) ? node5827 : 4'b1001;
															assign node5827 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node5830 = (inp[9]) ? node5834 : node5831;
															assign node5831 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node5834 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node5837 = (inp[1]) ? node5841 : node5838;
														assign node5838 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node5841 = (inp[9]) ? node5843 : 4'b1001;
															assign node5843 = (inp[10]) ? node5847 : node5844;
																assign node5844 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node5847 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node5850 = (inp[13]) ? node5874 : node5851;
												assign node5851 = (inp[1]) ? node5865 : node5852;
													assign node5852 = (inp[9]) ? 4'b1000 : node5853;
														assign node5853 = (inp[10]) ? node5859 : node5854;
															assign node5854 = (inp[5]) ? node5856 : 4'b1000;
																assign node5856 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node5859 = (inp[0]) ? 4'b1001 : node5860;
																assign node5860 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node5865 = (inp[5]) ? node5871 : node5866;
														assign node5866 = (inp[9]) ? 4'b1100 : node5867;
															assign node5867 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node5871 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node5874 = (inp[5]) ? node5884 : node5875;
													assign node5875 = (inp[1]) ? node5881 : node5876;
														assign node5876 = (inp[0]) ? node5878 : 4'b1100;
															assign node5878 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node5881 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node5884 = (inp[9]) ? node5892 : node5885;
														assign node5885 = (inp[10]) ? node5889 : node5886;
															assign node5886 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5889 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node5892 = (inp[10]) ? node5896 : node5893;
															assign node5893 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node5896 = (inp[1]) ? node5898 : 4'b1100;
																assign node5898 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node5901 = (inp[2]) ? node5971 : node5902;
											assign node5902 = (inp[13]) ? node5942 : node5903;
												assign node5903 = (inp[5]) ? node5927 : node5904;
													assign node5904 = (inp[1]) ? node5914 : node5905;
														assign node5905 = (inp[0]) ? 4'b1011 : node5906;
															assign node5906 = (inp[10]) ? node5910 : node5907;
																assign node5907 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node5910 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node5914 = (inp[9]) ? node5920 : node5915;
															assign node5915 = (inp[10]) ? 4'b1111 : node5916;
																assign node5916 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5920 = (inp[0]) ? node5924 : node5921;
																assign node5921 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node5924 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5927 = (inp[1]) ? node5935 : node5928;
														assign node5928 = (inp[0]) ? node5930 : 4'b1010;
															assign node5930 = (inp[9]) ? 4'b1011 : node5931;
																assign node5931 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node5935 = (inp[10]) ? 4'b1010 : node5936;
															assign node5936 = (inp[9]) ? node5938 : 4'b1010;
																assign node5938 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5942 = (inp[5]) ? node5956 : node5943;
													assign node5943 = (inp[1]) ? node5949 : node5944;
														assign node5944 = (inp[9]) ? 4'b1110 : node5945;
															assign node5945 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5949 = (inp[9]) ? 4'b1010 : node5950;
															assign node5950 = (inp[10]) ? node5952 : 4'b1011;
																assign node5952 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node5956 = (inp[10]) ? node5964 : node5957;
														assign node5957 = (inp[9]) ? node5959 : 4'b1110;
															assign node5959 = (inp[1]) ? 4'b1111 : node5960;
																assign node5960 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node5964 = (inp[9]) ? node5966 : 4'b1111;
															assign node5966 = (inp[0]) ? 4'b1110 : node5967;
																assign node5967 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node5971 = (inp[13]) ? node6011 : node5972;
												assign node5972 = (inp[5]) ? node5994 : node5973;
													assign node5973 = (inp[1]) ? node5981 : node5974;
														assign node5974 = (inp[10]) ? node5976 : 4'b1110;
															assign node5976 = (inp[9]) ? 4'b1110 : node5977;
																assign node5977 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5981 = (inp[0]) ? node5989 : node5982;
															assign node5982 = (inp[9]) ? node5986 : node5983;
																assign node5983 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node5986 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node5989 = (inp[10]) ? node5991 : 4'b1011;
																assign node5991 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node5994 = (inp[9]) ? node6000 : node5995;
														assign node5995 = (inp[10]) ? node5997 : 4'b1111;
															assign node5997 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6000 = (inp[10]) ? node6006 : node6001;
															assign node6001 = (inp[1]) ? node6003 : 4'b1110;
																assign node6003 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node6006 = (inp[0]) ? node6008 : 4'b1111;
																assign node6008 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node6011 = (inp[1]) ? node6029 : node6012;
													assign node6012 = (inp[5]) ? node6022 : node6013;
														assign node6013 = (inp[9]) ? 4'b1011 : node6014;
															assign node6014 = (inp[10]) ? node6018 : node6015;
																assign node6015 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node6018 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6022 = (inp[9]) ? node6026 : node6023;
															assign node6023 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node6026 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node6029 = (inp[5]) ? node6041 : node6030;
														assign node6030 = (inp[9]) ? node6036 : node6031;
															assign node6031 = (inp[0]) ? node6033 : 4'b1110;
																assign node6033 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node6036 = (inp[10]) ? 4'b1111 : node6037;
																assign node6037 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node6041 = (inp[0]) ? node6043 : 4'b1011;
															assign node6043 = (inp[9]) ? node6047 : node6044;
																assign node6044 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node6047 = (inp[10]) ? 4'b1011 : 4'b1010;
									assign node6050 = (inp[0]) ? node6196 : node6051;
										assign node6051 = (inp[4]) ? node6119 : node6052;
											assign node6052 = (inp[13]) ? node6088 : node6053;
												assign node6053 = (inp[2]) ? node6069 : node6054;
													assign node6054 = (inp[5]) ? node6064 : node6055;
														assign node6055 = (inp[1]) ? node6057 : 4'b1000;
															assign node6057 = (inp[9]) ? node6061 : node6058;
																assign node6058 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node6061 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6064 = (inp[10]) ? node6066 : 4'b1000;
															assign node6066 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node6069 = (inp[5]) ? node6079 : node6070;
														assign node6070 = (inp[1]) ? node6076 : node6071;
															assign node6071 = (inp[10]) ? 4'b1100 : node6072;
																assign node6072 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node6076 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node6079 = (inp[1]) ? node6081 : 4'b1101;
															assign node6081 = (inp[10]) ? node6085 : node6082;
																assign node6082 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node6085 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node6088 = (inp[2]) ? node6108 : node6089;
													assign node6089 = (inp[10]) ? node6099 : node6090;
														assign node6090 = (inp[5]) ? node6096 : node6091;
															assign node6091 = (inp[1]) ? node6093 : 4'b1100;
																assign node6093 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node6096 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6099 = (inp[1]) ? 4'b1100 : node6100;
															assign node6100 = (inp[9]) ? node6104 : node6101;
																assign node6101 = (inp[5]) ? 4'b1100 : 4'b1101;
																assign node6104 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node6108 = (inp[5]) ? node6114 : node6109;
														assign node6109 = (inp[1]) ? 4'b1100 : node6110;
															assign node6110 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node6114 = (inp[10]) ? 4'b1000 : node6115;
															assign node6115 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node6119 = (inp[2]) ? node6159 : node6120;
												assign node6120 = (inp[13]) ? node6134 : node6121;
													assign node6121 = (inp[5]) ? node6127 : node6122;
														assign node6122 = (inp[10]) ? node6124 : 4'b1001;
															assign node6124 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node6127 = (inp[1]) ? node6129 : 4'b1000;
															assign node6129 = (inp[10]) ? node6131 : 4'b1000;
																assign node6131 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node6134 = (inp[1]) ? node6146 : node6135;
														assign node6135 = (inp[10]) ? node6141 : node6136;
															assign node6136 = (inp[9]) ? node6138 : 4'b1101;
																assign node6138 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node6141 = (inp[5]) ? node6143 : 4'b1100;
																assign node6143 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6146 = (inp[5]) ? node6154 : node6147;
															assign node6147 = (inp[9]) ? node6151 : node6148;
																assign node6148 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node6151 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node6154 = (inp[10]) ? 4'b1100 : node6155;
																assign node6155 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node6159 = (inp[13]) ? node6181 : node6160;
													assign node6160 = (inp[5]) ? node6168 : node6161;
														assign node6161 = (inp[1]) ? node6163 : 4'b1101;
															assign node6163 = (inp[9]) ? 4'b1001 : node6164;
																assign node6164 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node6168 = (inp[1]) ? node6176 : node6169;
															assign node6169 = (inp[10]) ? node6173 : node6170;
																assign node6170 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node6173 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node6176 = (inp[9]) ? 4'b1101 : node6177;
																assign node6177 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6181 = (inp[5]) ? node6189 : node6182;
														assign node6182 = (inp[1]) ? node6184 : 4'b1001;
															assign node6184 = (inp[9]) ? node6186 : 4'b1101;
																assign node6186 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6189 = (inp[1]) ? node6193 : node6190;
															assign node6190 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node6193 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node6196 = (inp[1]) ? node6274 : node6197;
											assign node6197 = (inp[10]) ? node6235 : node6198;
												assign node6198 = (inp[9]) ? node6218 : node6199;
													assign node6199 = (inp[5]) ? node6207 : node6200;
														assign node6200 = (inp[2]) ? node6204 : node6201;
															assign node6201 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node6204 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node6207 = (inp[4]) ? node6213 : node6208;
															assign node6208 = (inp[13]) ? node6210 : 4'b1001;
																assign node6210 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node6213 = (inp[2]) ? 4'b1101 : node6214;
																assign node6214 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node6218 = (inp[5]) ? node6228 : node6219;
														assign node6219 = (inp[4]) ? node6225 : node6220;
															assign node6220 = (inp[13]) ? node6222 : 4'b1001;
																assign node6222 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node6225 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node6228 = (inp[4]) ? 4'b1001 : node6229;
															assign node6229 = (inp[13]) ? node6231 : 4'b1000;
																assign node6231 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node6235 = (inp[13]) ? node6253 : node6236;
													assign node6236 = (inp[2]) ? node6246 : node6237;
														assign node6237 = (inp[4]) ? 4'b1001 : node6238;
															assign node6238 = (inp[9]) ? node6242 : node6239;
																assign node6239 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node6242 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node6246 = (inp[9]) ? node6250 : node6247;
															assign node6247 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node6250 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node6253 = (inp[2]) ? node6265 : node6254;
														assign node6254 = (inp[9]) ? node6260 : node6255;
															assign node6255 = (inp[4]) ? 4'b1101 : node6256;
																assign node6256 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node6260 = (inp[5]) ? node6262 : 4'b1100;
																assign node6262 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node6265 = (inp[4]) ? node6267 : 4'b1000;
															assign node6267 = (inp[9]) ? node6271 : node6268;
																assign node6268 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node6271 = (inp[5]) ? 4'b1001 : 4'b1000;
											assign node6274 = (inp[5]) ? node6302 : node6275;
												assign node6275 = (inp[9]) ? node6289 : node6276;
													assign node6276 = (inp[10]) ? node6282 : node6277;
														assign node6277 = (inp[13]) ? node6279 : 4'b1100;
															assign node6279 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node6282 = (inp[2]) ? node6286 : node6283;
															assign node6283 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node6286 = (inp[13]) ? 4'b1100 : 4'b1001;
													assign node6289 = (inp[10]) ? node6297 : node6290;
														assign node6290 = (inp[4]) ? 4'b1101 : node6291;
															assign node6291 = (inp[2]) ? node6293 : 4'b1001;
																assign node6293 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node6297 = (inp[2]) ? node6299 : 4'b1000;
															assign node6299 = (inp[13]) ? 4'b1101 : 4'b1000;
												assign node6302 = (inp[13]) ? node6314 : node6303;
													assign node6303 = (inp[2]) ? node6307 : node6304;
														assign node6304 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node6307 = (inp[9]) ? node6311 : node6308;
															assign node6308 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node6311 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6314 = (inp[2]) ? node6318 : node6315;
														assign node6315 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node6318 = (inp[10]) ? node6322 : node6319;
															assign node6319 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node6322 = (inp[9]) ? 4'b1001 : 4'b1000;
						assign node6325 = (inp[15]) ? node7329 : node6326;
							assign node6326 = (inp[2]) ? node6836 : node6327;
								assign node6327 = (inp[13]) ? node6575 : node6328;
									assign node6328 = (inp[7]) ? node6446 : node6329;
										assign node6329 = (inp[1]) ? node6381 : node6330;
											assign node6330 = (inp[4]) ? node6352 : node6331;
												assign node6331 = (inp[12]) ? node6339 : node6332;
													assign node6332 = (inp[10]) ? node6336 : node6333;
														assign node6333 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6336 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node6339 = (inp[0]) ? node6345 : node6340;
														assign node6340 = (inp[9]) ? node6342 : 4'b1010;
															assign node6342 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node6345 = (inp[10]) ? node6349 : node6346;
															assign node6346 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node6349 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node6352 = (inp[12]) ? node6366 : node6353;
													assign node6353 = (inp[10]) ? node6361 : node6354;
														assign node6354 = (inp[9]) ? node6356 : 4'b1010;
															assign node6356 = (inp[0]) ? 4'b1011 : node6357;
																assign node6357 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node6361 = (inp[9]) ? node6363 : 4'b1011;
															assign node6363 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node6366 = (inp[5]) ? node6374 : node6367;
														assign node6367 = (inp[0]) ? node6369 : 4'b1100;
															assign node6369 = (inp[9]) ? node6371 : 4'b1101;
																assign node6371 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6374 = (inp[9]) ? node6378 : node6375;
															assign node6375 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node6378 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node6381 = (inp[5]) ? node6405 : node6382;
												assign node6382 = (inp[4]) ? node6392 : node6383;
													assign node6383 = (inp[12]) ? 4'b1111 : node6384;
														assign node6384 = (inp[10]) ? node6388 : node6385;
															assign node6385 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node6388 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node6392 = (inp[12]) ? node6400 : node6393;
														assign node6393 = (inp[10]) ? node6397 : node6394;
															assign node6394 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node6397 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6400 = (inp[0]) ? 4'b1100 : node6401;
															assign node6401 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node6405 = (inp[4]) ? node6433 : node6406;
													assign node6406 = (inp[12]) ? node6420 : node6407;
														assign node6407 = (inp[10]) ? node6415 : node6408;
															assign node6408 = (inp[0]) ? node6412 : node6409;
																assign node6409 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node6412 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node6415 = (inp[0]) ? node6417 : 4'b1000;
																assign node6417 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6420 = (inp[9]) ? node6428 : node6421;
															assign node6421 = (inp[0]) ? node6425 : node6422;
																assign node6422 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node6425 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node6428 = (inp[10]) ? node6430 : 4'b1010;
																assign node6430 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6433 = (inp[12]) ? node6439 : node6434;
														assign node6434 = (inp[10]) ? 4'b1010 : node6435;
															assign node6435 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node6439 = (inp[9]) ? node6443 : node6440;
															assign node6440 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node6443 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node6446 = (inp[1]) ? node6506 : node6447;
											assign node6447 = (inp[12]) ? node6471 : node6448;
												assign node6448 = (inp[4]) ? node6460 : node6449;
													assign node6449 = (inp[5]) ? node6455 : node6450;
														assign node6450 = (inp[10]) ? 4'b1010 : node6451;
															assign node6451 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node6455 = (inp[10]) ? node6457 : 4'b1111;
															assign node6457 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6460 = (inp[9]) ? node6466 : node6461;
														assign node6461 = (inp[10]) ? node6463 : 4'b1100;
															assign node6463 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node6466 = (inp[10]) ? node6468 : 4'b1101;
															assign node6468 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node6471 = (inp[4]) ? node6491 : node6472;
													assign node6472 = (inp[10]) ? node6482 : node6473;
														assign node6473 = (inp[0]) ? node6475 : 4'b1101;
															assign node6475 = (inp[5]) ? node6479 : node6476;
																assign node6476 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node6479 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6482 = (inp[9]) ? node6484 : 4'b1100;
															assign node6484 = (inp[0]) ? node6488 : node6485;
																assign node6485 = (inp[5]) ? 4'b1100 : 4'b1101;
																assign node6488 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node6491 = (inp[9]) ? node6497 : node6492;
														assign node6492 = (inp[5]) ? 4'b1010 : node6493;
															assign node6493 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node6497 = (inp[10]) ? node6501 : node6498;
															assign node6498 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node6501 = (inp[0]) ? node6503 : 4'b1011;
																assign node6503 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node6506 = (inp[5]) ? node6536 : node6507;
												assign node6507 = (inp[4]) ? node6521 : node6508;
													assign node6508 = (inp[12]) ? node6514 : node6509;
														assign node6509 = (inp[0]) ? node6511 : 4'b1010;
															assign node6511 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node6514 = (inp[9]) ? node6518 : node6515;
															assign node6515 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node6518 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node6521 = (inp[12]) ? node6531 : node6522;
														assign node6522 = (inp[9]) ? node6524 : 4'b1000;
															assign node6524 = (inp[0]) ? node6528 : node6525;
																assign node6525 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node6528 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node6531 = (inp[9]) ? node6533 : 4'b1111;
															assign node6533 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node6536 = (inp[4]) ? node6560 : node6537;
													assign node6537 = (inp[12]) ? node6545 : node6538;
														assign node6538 = (inp[9]) ? 4'b1011 : node6539;
															assign node6539 = (inp[10]) ? node6541 : 4'b1010;
																assign node6541 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6545 = (inp[0]) ? node6553 : node6546;
															assign node6546 = (inp[10]) ? node6550 : node6547;
																assign node6547 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node6550 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node6553 = (inp[10]) ? node6557 : node6554;
																assign node6554 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node6557 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node6560 = (inp[12]) ? node6568 : node6561;
														assign node6561 = (inp[0]) ? node6563 : 4'b1100;
															assign node6563 = (inp[9]) ? node6565 : 4'b1100;
																assign node6565 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6568 = (inp[10]) ? node6572 : node6569;
															assign node6569 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node6572 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node6575 = (inp[1]) ? node6703 : node6576;
										assign node6576 = (inp[7]) ? node6650 : node6577;
											assign node6577 = (inp[4]) ? node6607 : node6578;
												assign node6578 = (inp[12]) ? node6596 : node6579;
													assign node6579 = (inp[0]) ? node6589 : node6580;
														assign node6580 = (inp[5]) ? node6582 : 4'b1100;
															assign node6582 = (inp[9]) ? node6586 : node6583;
																assign node6583 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node6586 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6589 = (inp[9]) ? node6593 : node6590;
															assign node6590 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node6593 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node6596 = (inp[5]) ? node6600 : node6597;
														assign node6597 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6600 = (inp[0]) ? node6602 : 4'b1110;
															assign node6602 = (inp[10]) ? 4'b1110 : node6603;
																assign node6603 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node6607 = (inp[12]) ? node6629 : node6608;
													assign node6608 = (inp[0]) ? node6614 : node6609;
														assign node6609 = (inp[10]) ? 4'b1110 : node6610;
															assign node6610 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6614 = (inp[10]) ? node6622 : node6615;
															assign node6615 = (inp[9]) ? node6619 : node6616;
																assign node6616 = (inp[5]) ? 4'b1111 : 4'b1110;
																assign node6619 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node6622 = (inp[9]) ? node6626 : node6623;
																assign node6623 = (inp[5]) ? 4'b1110 : 4'b1111;
																assign node6626 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node6629 = (inp[5]) ? node6639 : node6630;
														assign node6630 = (inp[0]) ? node6634 : node6631;
															assign node6631 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node6634 = (inp[10]) ? node6636 : 4'b1000;
																assign node6636 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6639 = (inp[10]) ? node6645 : node6640;
															assign node6640 = (inp[9]) ? 4'b1100 : node6641;
																assign node6641 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node6645 = (inp[9]) ? 4'b1101 : node6646;
																assign node6646 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node6650 = (inp[10]) ? node6674 : node6651;
												assign node6651 = (inp[5]) ? node6665 : node6652;
													assign node6652 = (inp[4]) ? node6658 : node6653;
														assign node6653 = (inp[12]) ? 4'b1000 : node6654;
															assign node6654 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node6658 = (inp[12]) ? node6660 : 4'b1001;
															assign node6660 = (inp[9]) ? 4'b1111 : node6661;
																assign node6661 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node6665 = (inp[4]) ? node6669 : node6666;
														assign node6666 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node6669 = (inp[12]) ? node6671 : 4'b1000;
															assign node6671 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node6674 = (inp[4]) ? node6692 : node6675;
													assign node6675 = (inp[12]) ? node6683 : node6676;
														assign node6676 = (inp[9]) ? node6680 : node6677;
															assign node6677 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node6680 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node6683 = (inp[9]) ? node6685 : 4'b1001;
															assign node6685 = (inp[0]) ? node6689 : node6686;
																assign node6686 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node6689 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node6692 = (inp[12]) ? node6700 : node6693;
														assign node6693 = (inp[9]) ? 4'b1001 : node6694;
															assign node6694 = (inp[5]) ? node6696 : 4'b1000;
																assign node6696 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6700 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node6703 = (inp[12]) ? node6769 : node6704;
											assign node6704 = (inp[5]) ? node6730 : node6705;
												assign node6705 = (inp[7]) ? node6717 : node6706;
													assign node6706 = (inp[4]) ? node6712 : node6707;
														assign node6707 = (inp[9]) ? 4'b1001 : node6708;
															assign node6708 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6712 = (inp[10]) ? 4'b1011 : node6713;
															assign node6713 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6717 = (inp[4]) ? node6721 : node6718;
														assign node6718 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node6721 = (inp[0]) ? node6723 : 4'b1101;
															assign node6723 = (inp[10]) ? node6727 : node6724;
																assign node6724 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node6727 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node6730 = (inp[7]) ? node6750 : node6731;
													assign node6731 = (inp[4]) ? node6739 : node6732;
														assign node6732 = (inp[9]) ? node6736 : node6733;
															assign node6733 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node6736 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6739 = (inp[0]) ? node6745 : node6740;
															assign node6740 = (inp[10]) ? 4'b1111 : node6741;
																assign node6741 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node6745 = (inp[9]) ? 4'b1110 : node6746;
																assign node6746 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node6750 = (inp[4]) ? node6760 : node6751;
														assign node6751 = (inp[0]) ? node6753 : 4'b1110;
															assign node6753 = (inp[10]) ? node6757 : node6754;
																assign node6754 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node6757 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6760 = (inp[0]) ? 4'b1000 : node6761;
															assign node6761 = (inp[9]) ? node6765 : node6762;
																assign node6762 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node6765 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node6769 = (inp[4]) ? node6805 : node6770;
												assign node6770 = (inp[7]) ? node6788 : node6771;
													assign node6771 = (inp[5]) ? node6779 : node6772;
														assign node6772 = (inp[10]) ? node6776 : node6773;
															assign node6773 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node6776 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node6779 = (inp[0]) ? node6781 : 4'b1111;
															assign node6781 = (inp[10]) ? node6785 : node6782;
																assign node6782 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node6785 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node6788 = (inp[5]) ? node6796 : node6789;
														assign node6789 = (inp[0]) ? 4'b1100 : node6790;
															assign node6790 = (inp[10]) ? node6792 : 4'b1101;
																assign node6792 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node6796 = (inp[0]) ? node6798 : 4'b1001;
															assign node6798 = (inp[10]) ? node6802 : node6799;
																assign node6799 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node6802 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6805 = (inp[7]) ? node6823 : node6806;
													assign node6806 = (inp[10]) ? node6816 : node6807;
														assign node6807 = (inp[9]) ? node6813 : node6808;
															assign node6808 = (inp[5]) ? 4'b1001 : node6809;
																assign node6809 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node6813 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6816 = (inp[9]) ? node6818 : 4'b1000;
															assign node6818 = (inp[0]) ? node6820 : 4'b1001;
																assign node6820 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node6823 = (inp[5]) ? node6831 : node6824;
														assign node6824 = (inp[0]) ? 4'b1010 : node6825;
															assign node6825 = (inp[10]) ? node6827 : 4'b1011;
																assign node6827 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node6831 = (inp[0]) ? 4'b1111 : node6832;
															assign node6832 = (inp[10]) ? 4'b1111 : 4'b1110;
								assign node6836 = (inp[13]) ? node7078 : node6837;
									assign node6837 = (inp[12]) ? node6973 : node6838;
										assign node6838 = (inp[4]) ? node6904 : node6839;
											assign node6839 = (inp[7]) ? node6863 : node6840;
												assign node6840 = (inp[1]) ? node6848 : node6841;
													assign node6841 = (inp[9]) ? node6845 : node6842;
														assign node6842 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6845 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node6848 = (inp[5]) ? node6858 : node6849;
														assign node6849 = (inp[10]) ? 4'b1000 : node6850;
															assign node6850 = (inp[0]) ? node6854 : node6851;
																assign node6851 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node6854 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6858 = (inp[10]) ? 4'b1101 : node6859;
															assign node6859 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6863 = (inp[5]) ? node6885 : node6864;
													assign node6864 = (inp[0]) ? node6878 : node6865;
														assign node6865 = (inp[10]) ? node6871 : node6866;
															assign node6866 = (inp[1]) ? 4'b1111 : node6867;
																assign node6867 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node6871 = (inp[9]) ? node6875 : node6872;
																assign node6872 = (inp[1]) ? 4'b1110 : 4'b1111;
																assign node6875 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node6878 = (inp[9]) ? node6882 : node6879;
															assign node6879 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node6882 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node6885 = (inp[1]) ? node6895 : node6886;
														assign node6886 = (inp[9]) ? node6888 : 4'b1010;
															assign node6888 = (inp[0]) ? node6892 : node6889;
																assign node6889 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node6892 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node6895 = (inp[10]) ? node6897 : 4'b1110;
															assign node6897 = (inp[9]) ? node6901 : node6898;
																assign node6898 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node6901 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node6904 = (inp[7]) ? node6940 : node6905;
												assign node6905 = (inp[5]) ? node6925 : node6906;
													assign node6906 = (inp[1]) ? node6918 : node6907;
														assign node6907 = (inp[0]) ? node6913 : node6908;
															assign node6908 = (inp[9]) ? 4'b1110 : node6909;
																assign node6909 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node6913 = (inp[10]) ? 4'b1111 : node6914;
																assign node6914 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node6918 = (inp[9]) ? 4'b1010 : node6919;
															assign node6919 = (inp[10]) ? node6921 : 4'b1011;
																assign node6921 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6925 = (inp[9]) ? node6931 : node6926;
														assign node6926 = (inp[10]) ? node6928 : 4'b1110;
															assign node6928 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node6931 = (inp[10]) ? node6935 : node6932;
															assign node6932 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node6935 = (inp[0]) ? node6937 : 4'b1110;
																assign node6937 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node6940 = (inp[5]) ? node6954 : node6941;
													assign node6941 = (inp[1]) ? node6945 : node6942;
														assign node6942 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node6945 = (inp[9]) ? 4'b1100 : node6946;
															assign node6946 = (inp[0]) ? node6950 : node6947;
																assign node6947 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node6950 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node6954 = (inp[0]) ? node6966 : node6955;
														assign node6955 = (inp[1]) ? node6961 : node6956;
															assign node6956 = (inp[10]) ? 4'b1000 : node6957;
																assign node6957 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node6961 = (inp[9]) ? 4'b1001 : node6962;
																assign node6962 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node6966 = (inp[1]) ? node6968 : 4'b1001;
															assign node6968 = (inp[10]) ? 4'b1001 : node6969;
																assign node6969 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node6973 = (inp[5]) ? node7023 : node6974;
											assign node6974 = (inp[4]) ? node6998 : node6975;
												assign node6975 = (inp[7]) ? node6989 : node6976;
													assign node6976 = (inp[1]) ? node6982 : node6977;
														assign node6977 = (inp[10]) ? 4'b1111 : node6978;
															assign node6978 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node6982 = (inp[10]) ? 4'b1010 : node6983;
															assign node6983 = (inp[9]) ? 4'b1011 : node6984;
																assign node6984 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6989 = (inp[1]) ? node6995 : node6990;
														assign node6990 = (inp[10]) ? 4'b1001 : node6991;
															assign node6991 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6995 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node6998 = (inp[7]) ? node7016 : node6999;
													assign node6999 = (inp[0]) ? node7007 : node7000;
														assign node7000 = (inp[10]) ? 4'b1000 : node7001;
															assign node7001 = (inp[1]) ? node7003 : 4'b1000;
																assign node7003 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node7007 = (inp[1]) ? 4'b1001 : node7008;
															assign node7008 = (inp[9]) ? node7012 : node7009;
																assign node7009 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node7012 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node7016 = (inp[1]) ? node7018 : 4'b1110;
														assign node7018 = (inp[10]) ? 4'b1010 : node7019;
															assign node7019 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node7023 = (inp[4]) ? node7043 : node7024;
												assign node7024 = (inp[7]) ? node7038 : node7025;
													assign node7025 = (inp[1]) ? node7027 : 4'b1110;
														assign node7027 = (inp[9]) ? node7033 : node7028;
															assign node7028 = (inp[0]) ? 4'b1111 : node7029;
																assign node7029 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node7033 = (inp[10]) ? node7035 : 4'b1110;
																assign node7035 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node7038 = (inp[1]) ? 4'b1000 : node7039;
														assign node7039 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node7043 = (inp[7]) ? node7063 : node7044;
													assign node7044 = (inp[1]) ? node7052 : node7045;
														assign node7045 = (inp[0]) ? node7049 : node7046;
															assign node7046 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node7049 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node7052 = (inp[0]) ? node7058 : node7053;
															assign node7053 = (inp[10]) ? 4'b1000 : node7054;
																assign node7054 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node7058 = (inp[10]) ? 4'b1001 : node7059;
																assign node7059 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7063 = (inp[0]) ? node7071 : node7064;
														assign node7064 = (inp[1]) ? node7066 : 4'b1111;
															assign node7066 = (inp[10]) ? 4'b1111 : node7067;
																assign node7067 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node7071 = (inp[10]) ? node7075 : node7072;
															assign node7072 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node7075 = (inp[9]) ? 4'b1111 : 4'b1110;
									assign node7078 = (inp[12]) ? node7196 : node7079;
										assign node7079 = (inp[4]) ? node7141 : node7080;
											assign node7080 = (inp[7]) ? node7110 : node7081;
												assign node7081 = (inp[5]) ? node7093 : node7082;
													assign node7082 = (inp[1]) ? node7088 : node7083;
														assign node7083 = (inp[9]) ? node7085 : 4'b1000;
															assign node7085 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node7088 = (inp[9]) ? 4'b1100 : node7089;
															assign node7089 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node7093 = (inp[1]) ? node7101 : node7094;
														assign node7094 = (inp[10]) ? node7098 : node7095;
															assign node7095 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node7098 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node7101 = (inp[10]) ? node7103 : 4'b1000;
															assign node7103 = (inp[0]) ? node7107 : node7104;
																assign node7104 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node7107 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node7110 = (inp[5]) ? node7132 : node7111;
													assign node7111 = (inp[1]) ? node7119 : node7112;
														assign node7112 = (inp[0]) ? node7114 : 4'b1011;
															assign node7114 = (inp[9]) ? node7116 : 4'b1010;
																assign node7116 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node7119 = (inp[10]) ? node7125 : node7120;
															assign node7120 = (inp[0]) ? node7122 : 4'b1010;
																assign node7122 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node7125 = (inp[0]) ? node7129 : node7126;
																assign node7126 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node7129 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node7132 = (inp[1]) ? node7134 : 4'b1110;
														assign node7134 = (inp[9]) ? node7136 : 4'b1010;
															assign node7136 = (inp[0]) ? 4'b1010 : node7137;
																assign node7137 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node7141 = (inp[7]) ? node7167 : node7142;
												assign node7142 = (inp[1]) ? node7156 : node7143;
													assign node7143 = (inp[9]) ? node7147 : node7144;
														assign node7144 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node7147 = (inp[5]) ? node7149 : 4'b1011;
															assign node7149 = (inp[0]) ? node7153 : node7150;
																assign node7150 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node7153 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node7156 = (inp[5]) ? node7162 : node7157;
														assign node7157 = (inp[9]) ? 4'b1110 : node7158;
															assign node7158 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node7162 = (inp[9]) ? 4'b1010 : node7163;
															assign node7163 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node7167 = (inp[1]) ? node7179 : node7168;
													assign node7168 = (inp[5]) ? node7170 : 4'b1100;
														assign node7170 = (inp[9]) ? 4'b1100 : node7171;
															assign node7171 = (inp[0]) ? node7175 : node7172;
																assign node7172 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node7175 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node7179 = (inp[5]) ? node7189 : node7180;
														assign node7180 = (inp[10]) ? 4'b1001 : node7181;
															assign node7181 = (inp[0]) ? node7185 : node7182;
																assign node7182 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node7185 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node7189 = (inp[9]) ? node7193 : node7190;
															assign node7190 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node7193 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node7196 = (inp[1]) ? node7264 : node7197;
											assign node7197 = (inp[4]) ? node7229 : node7198;
												assign node7198 = (inp[7]) ? node7206 : node7199;
													assign node7199 = (inp[9]) ? node7203 : node7200;
														assign node7200 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node7203 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node7206 = (inp[5]) ? node7220 : node7207;
														assign node7207 = (inp[0]) ? node7213 : node7208;
															assign node7208 = (inp[10]) ? 4'b1101 : node7209;
																assign node7209 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node7213 = (inp[9]) ? node7217 : node7214;
																assign node7214 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node7217 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node7220 = (inp[9]) ? 4'b1100 : node7221;
															assign node7221 = (inp[10]) ? node7225 : node7222;
																assign node7222 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node7225 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node7229 = (inp[7]) ? node7239 : node7230;
													assign node7230 = (inp[5]) ? 4'b1001 : node7231;
														assign node7231 = (inp[9]) ? node7235 : node7232;
															assign node7232 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node7235 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node7239 = (inp[0]) ? node7255 : node7240;
														assign node7240 = (inp[5]) ? node7248 : node7241;
															assign node7241 = (inp[9]) ? node7245 : node7242;
																assign node7242 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node7245 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node7248 = (inp[10]) ? node7252 : node7249;
																assign node7249 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node7252 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node7255 = (inp[10]) ? 4'b1010 : node7256;
															assign node7256 = (inp[9]) ? node7260 : node7257;
																assign node7257 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node7260 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node7264 = (inp[7]) ? node7296 : node7265;
												assign node7265 = (inp[4]) ? node7277 : node7266;
													assign node7266 = (inp[5]) ? node7272 : node7267;
														assign node7267 = (inp[10]) ? 4'b1110 : node7268;
															assign node7268 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node7272 = (inp[0]) ? 4'b1010 : node7273;
															assign node7273 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node7277 = (inp[9]) ? node7287 : node7278;
														assign node7278 = (inp[10]) ? node7284 : node7279;
															assign node7279 = (inp[5]) ? 4'b1100 : node7280;
																assign node7280 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7284 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node7287 = (inp[10]) ? node7293 : node7288;
															assign node7288 = (inp[5]) ? 4'b1101 : node7289;
																assign node7289 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7293 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node7296 = (inp[4]) ? node7318 : node7297;
													assign node7297 = (inp[5]) ? node7311 : node7298;
														assign node7298 = (inp[0]) ? node7304 : node7299;
															assign node7299 = (inp[10]) ? 4'b1000 : node7300;
																assign node7300 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node7304 = (inp[9]) ? node7308 : node7305;
																assign node7305 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node7308 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node7311 = (inp[9]) ? node7315 : node7312;
															assign node7312 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node7315 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node7318 = (inp[5]) ? node7324 : node7319;
														assign node7319 = (inp[9]) ? 4'b1110 : node7320;
															assign node7320 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node7324 = (inp[9]) ? 4'b1011 : node7325;
															assign node7325 = (inp[10]) ? 4'b1011 : 4'b1010;
							assign node7329 = (inp[9]) ? node7815 : node7330;
								assign node7330 = (inp[10]) ? node7596 : node7331;
									assign node7331 = (inp[2]) ? node7487 : node7332;
										assign node7332 = (inp[13]) ? node7410 : node7333;
											assign node7333 = (inp[1]) ? node7377 : node7334;
												assign node7334 = (inp[12]) ? node7356 : node7335;
													assign node7335 = (inp[7]) ? node7343 : node7336;
														assign node7336 = (inp[4]) ? node7338 : 4'b1000;
															assign node7338 = (inp[0]) ? 4'b1100 : node7339;
																assign node7339 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node7343 = (inp[0]) ? node7351 : node7344;
															assign node7344 = (inp[5]) ? node7348 : node7345;
																assign node7345 = (inp[4]) ? 4'b1011 : 4'b1110;
																assign node7348 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node7351 = (inp[4]) ? node7353 : 4'b1011;
																assign node7353 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node7356 = (inp[7]) ? node7364 : node7357;
														assign node7357 = (inp[4]) ? node7359 : 4'b1010;
															assign node7359 = (inp[0]) ? node7361 : 4'b1011;
																assign node7361 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node7364 = (inp[0]) ? node7372 : node7365;
															assign node7365 = (inp[5]) ? node7369 : node7366;
																assign node7366 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node7369 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node7372 = (inp[4]) ? 4'b1001 : node7373;
																assign node7373 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node7377 = (inp[5]) ? node7395 : node7378;
													assign node7378 = (inp[12]) ? node7388 : node7379;
														assign node7379 = (inp[4]) ? node7383 : node7380;
															assign node7380 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7383 = (inp[7]) ? node7385 : 4'b1001;
																assign node7385 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7388 = (inp[7]) ? node7390 : 4'b1110;
															assign node7390 = (inp[0]) ? node7392 : 4'b1101;
																assign node7392 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node7395 = (inp[4]) ? node7401 : node7396;
														assign node7396 = (inp[7]) ? 4'b1110 : node7397;
															assign node7397 = (inp[12]) ? 4'b1010 : 4'b1001;
														assign node7401 = (inp[7]) ? node7407 : node7402;
															assign node7402 = (inp[12]) ? 4'b1011 : node7403;
																assign node7403 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7407 = (inp[12]) ? 4'b1001 : 4'b1011;
											assign node7410 = (inp[1]) ? node7446 : node7411;
												assign node7411 = (inp[12]) ? node7427 : node7412;
													assign node7412 = (inp[7]) ? node7420 : node7413;
														assign node7413 = (inp[4]) ? node7417 : node7414;
															assign node7414 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7417 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node7420 = (inp[5]) ? node7424 : node7421;
															assign node7421 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node7424 = (inp[4]) ? 4'b1010 : 4'b1111;
													assign node7427 = (inp[7]) ? node7435 : node7428;
														assign node7428 = (inp[0]) ? node7432 : node7429;
															assign node7429 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node7432 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node7435 = (inp[5]) ? node7441 : node7436;
															assign node7436 = (inp[0]) ? node7438 : 4'b1101;
																assign node7438 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node7441 = (inp[4]) ? 4'b1100 : node7442;
																assign node7442 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node7446 = (inp[5]) ? node7466 : node7447;
													assign node7447 = (inp[12]) ? node7455 : node7448;
														assign node7448 = (inp[7]) ? node7452 : node7449;
															assign node7449 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node7452 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node7455 = (inp[7]) ? node7461 : node7456;
															assign node7456 = (inp[4]) ? 4'b1010 : node7457;
																assign node7457 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node7461 = (inp[0]) ? node7463 : 4'b1001;
																assign node7463 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node7466 = (inp[12]) ? node7476 : node7467;
														assign node7467 = (inp[7]) ? node7473 : node7468;
															assign node7468 = (inp[4]) ? 4'b1001 : node7469;
																assign node7469 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7473 = (inp[4]) ? 4'b1111 : 4'b1010;
														assign node7476 = (inp[7]) ? node7480 : node7477;
															assign node7477 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node7480 = (inp[0]) ? node7484 : node7481;
																assign node7481 = (inp[4]) ? 4'b1101 : 4'b1100;
																assign node7484 = (inp[4]) ? 4'b1100 : 4'b1101;
										assign node7487 = (inp[13]) ? node7539 : node7488;
											assign node7488 = (inp[5]) ? node7522 : node7489;
												assign node7489 = (inp[1]) ? node7505 : node7490;
													assign node7490 = (inp[12]) ? node7496 : node7491;
														assign node7491 = (inp[7]) ? 4'b1010 : node7492;
															assign node7492 = (inp[0]) ? 4'b1001 : 4'b1100;
														assign node7496 = (inp[7]) ? node7502 : node7497;
															assign node7497 = (inp[4]) ? node7499 : 4'b1110;
																assign node7499 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node7502 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node7505 = (inp[4]) ? node7511 : node7506;
														assign node7506 = (inp[12]) ? node7508 : 4'b1001;
															assign node7508 = (inp[7]) ? 4'b1001 : 4'b1010;
														assign node7511 = (inp[12]) ? node7517 : node7512;
															assign node7512 = (inp[7]) ? node7514 : 4'b1100;
																assign node7514 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node7517 = (inp[7]) ? node7519 : 4'b1010;
																assign node7519 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7522 = (inp[12]) ? node7536 : node7523;
													assign node7523 = (inp[7]) ? node7531 : node7524;
														assign node7524 = (inp[1]) ? node7528 : node7525;
															assign node7525 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node7528 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node7531 = (inp[1]) ? 4'b1110 : node7532;
															assign node7532 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node7536 = (inp[7]) ? 4'b1100 : 4'b1110;
											assign node7539 = (inp[5]) ? node7577 : node7540;
												assign node7540 = (inp[4]) ? node7556 : node7541;
													assign node7541 = (inp[1]) ? node7549 : node7542;
														assign node7542 = (inp[7]) ? node7546 : node7543;
															assign node7543 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node7546 = (inp[12]) ? 4'b1001 : 4'b1110;
														assign node7549 = (inp[7]) ? node7553 : node7550;
															assign node7550 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node7553 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node7556 = (inp[7]) ? node7564 : node7557;
														assign node7557 = (inp[12]) ? node7561 : node7558;
															assign node7558 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node7561 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node7564 = (inp[12]) ? node7572 : node7565;
															assign node7565 = (inp[1]) ? node7569 : node7566;
																assign node7566 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node7569 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node7572 = (inp[1]) ? 4'b1100 : node7573;
																assign node7573 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7577 = (inp[12]) ? node7593 : node7578;
													assign node7578 = (inp[7]) ? node7584 : node7579;
														assign node7579 = (inp[4]) ? 4'b1100 : node7580;
															assign node7580 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node7584 = (inp[0]) ? node7590 : node7585;
															assign node7585 = (inp[4]) ? 4'b1111 : node7586;
																assign node7586 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node7590 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node7593 = (inp[7]) ? 4'b1000 : 4'b1010;
									assign node7596 = (inp[5]) ? node7726 : node7597;
										assign node7597 = (inp[7]) ? node7669 : node7598;
											assign node7598 = (inp[12]) ? node7634 : node7599;
												assign node7599 = (inp[2]) ? node7615 : node7600;
													assign node7600 = (inp[1]) ? node7608 : node7601;
														assign node7601 = (inp[0]) ? node7603 : 4'b1101;
															assign node7603 = (inp[4]) ? 4'b1001 : node7604;
																assign node7604 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node7608 = (inp[4]) ? node7612 : node7609;
															assign node7609 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7612 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node7615 = (inp[0]) ? node7625 : node7616;
														assign node7616 = (inp[13]) ? 4'b1001 : node7617;
															assign node7617 = (inp[1]) ? node7621 : node7618;
																assign node7618 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node7621 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node7625 = (inp[13]) ? node7627 : 4'b1000;
															assign node7627 = (inp[1]) ? node7631 : node7628;
																assign node7628 = (inp[4]) ? 4'b1100 : 4'b1001;
																assign node7631 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node7634 = (inp[0]) ? node7648 : node7635;
													assign node7635 = (inp[2]) ? node7643 : node7636;
														assign node7636 = (inp[1]) ? node7640 : node7637;
															assign node7637 = (inp[13]) ? 4'b1111 : 4'b1010;
															assign node7640 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node7643 = (inp[13]) ? 4'b1011 : node7644;
															assign node7644 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node7648 = (inp[13]) ? node7658 : node7649;
														assign node7649 = (inp[2]) ? node7653 : node7650;
															assign node7650 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node7653 = (inp[1]) ? 4'b1011 : node7654;
																assign node7654 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node7658 = (inp[2]) ? node7666 : node7659;
															assign node7659 = (inp[1]) ? node7663 : node7660;
																assign node7660 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node7663 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node7666 = (inp[1]) ? 4'b1110 : 4'b1010;
											assign node7669 = (inp[12]) ? node7699 : node7670;
												assign node7670 = (inp[1]) ? node7684 : node7671;
													assign node7671 = (inp[13]) ? node7677 : node7672;
														assign node7672 = (inp[2]) ? node7674 : 4'b1111;
															assign node7674 = (inp[0]) ? 4'b1110 : 4'b1010;
														assign node7677 = (inp[4]) ? node7681 : node7678;
															assign node7678 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node7681 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7684 = (inp[13]) ? node7692 : node7685;
														assign node7685 = (inp[2]) ? node7689 : node7686;
															assign node7686 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node7689 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7692 = (inp[4]) ? node7696 : node7693;
															assign node7693 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node7696 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node7699 = (inp[0]) ? node7717 : node7700;
													assign node7700 = (inp[4]) ? node7706 : node7701;
														assign node7701 = (inp[2]) ? node7703 : 4'b1000;
															assign node7703 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node7706 = (inp[2]) ? node7714 : node7707;
															assign node7707 = (inp[13]) ? node7711 : node7708;
																assign node7708 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node7711 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node7714 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node7717 = (inp[4]) ? node7723 : node7718;
														assign node7718 = (inp[13]) ? 4'b1101 : node7719;
															assign node7719 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node7723 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node7726 = (inp[2]) ? node7778 : node7727;
											assign node7727 = (inp[13]) ? node7753 : node7728;
												assign node7728 = (inp[12]) ? node7746 : node7729;
													assign node7729 = (inp[7]) ? node7739 : node7730;
														assign node7730 = (inp[4]) ? node7734 : node7731;
															assign node7731 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node7734 = (inp[1]) ? 4'b1101 : node7735;
																assign node7735 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7739 = (inp[1]) ? 4'b1111 : node7740;
															assign node7740 = (inp[4]) ? 4'b1111 : node7741;
																assign node7741 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7746 = (inp[4]) ? node7750 : node7747;
														assign node7747 = (inp[7]) ? 4'b1001 : 4'b1011;
														assign node7750 = (inp[7]) ? 4'b1000 : 4'b1010;
												assign node7753 = (inp[12]) ? node7767 : node7754;
													assign node7754 = (inp[7]) ? node7762 : node7755;
														assign node7755 = (inp[4]) ? 4'b1000 : node7756;
															assign node7756 = (inp[1]) ? node7758 : 4'b1101;
																assign node7758 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7762 = (inp[1]) ? 4'b1011 : node7763;
															assign node7763 = (inp[4]) ? 4'b1011 : 4'b1110;
													assign node7767 = (inp[7]) ? node7771 : node7768;
														assign node7768 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node7771 = (inp[4]) ? node7775 : node7772;
															assign node7772 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7775 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node7778 = (inp[13]) ? node7796 : node7779;
												assign node7779 = (inp[12]) ? node7793 : node7780;
													assign node7780 = (inp[7]) ? node7786 : node7781;
														assign node7781 = (inp[4]) ? node7783 : 4'b1101;
															assign node7783 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7786 = (inp[0]) ? node7790 : node7787;
															assign node7787 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node7790 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node7793 = (inp[7]) ? 4'b1101 : 4'b1111;
												assign node7796 = (inp[12]) ? node7812 : node7797;
													assign node7797 = (inp[7]) ? node7803 : node7798;
														assign node7798 = (inp[4]) ? 4'b1101 : node7799;
															assign node7799 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7803 = (inp[1]) ? node7809 : node7804;
															assign node7804 = (inp[4]) ? 4'b1110 : node7805;
																assign node7805 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node7809 = (inp[0]) ? 4'b1111 : 4'b1011;
													assign node7812 = (inp[7]) ? 4'b1001 : 4'b1011;
								assign node7815 = (inp[10]) ? node8075 : node7816;
									assign node7816 = (inp[7]) ? node7932 : node7817;
										assign node7817 = (inp[12]) ? node7883 : node7818;
											assign node7818 = (inp[1]) ? node7846 : node7819;
												assign node7819 = (inp[4]) ? node7831 : node7820;
													assign node7820 = (inp[5]) ? node7826 : node7821;
														assign node7821 = (inp[13]) ? node7823 : 4'b1001;
															assign node7823 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node7826 = (inp[13]) ? 4'b1100 : node7827;
															assign node7827 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node7831 = (inp[13]) ? node7839 : node7832;
														assign node7832 = (inp[2]) ? node7836 : node7833;
															assign node7833 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7836 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node7839 = (inp[2]) ? node7843 : node7840;
															assign node7840 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node7843 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node7846 = (inp[5]) ? node7862 : node7847;
													assign node7847 = (inp[4]) ? node7855 : node7848;
														assign node7848 = (inp[2]) ? node7852 : node7849;
															assign node7849 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node7852 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node7855 = (inp[2]) ? node7859 : node7856;
															assign node7856 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node7859 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node7862 = (inp[2]) ? node7874 : node7863;
														assign node7863 = (inp[13]) ? node7867 : node7864;
															assign node7864 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7867 = (inp[4]) ? node7871 : node7868;
																assign node7868 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node7871 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node7874 = (inp[0]) ? node7880 : node7875;
															assign node7875 = (inp[4]) ? 4'b1100 : node7876;
																assign node7876 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node7880 = (inp[13]) ? 4'b1101 : 4'b1000;
											assign node7883 = (inp[4]) ? node7907 : node7884;
												assign node7884 = (inp[13]) ? node7896 : node7885;
													assign node7885 = (inp[2]) ? node7891 : node7886;
														assign node7886 = (inp[5]) ? 4'b1011 : node7887;
															assign node7887 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node7891 = (inp[1]) ? node7893 : 4'b1111;
															assign node7893 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node7896 = (inp[2]) ? node7902 : node7897;
														assign node7897 = (inp[0]) ? node7899 : 4'b1011;
															assign node7899 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node7902 = (inp[1]) ? node7904 : 4'b1011;
															assign node7904 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node7907 = (inp[13]) ? node7921 : node7908;
													assign node7908 = (inp[2]) ? node7914 : node7909;
														assign node7909 = (inp[5]) ? 4'b1010 : node7910;
															assign node7910 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node7914 = (inp[5]) ? 4'b1111 : node7915;
															assign node7915 = (inp[1]) ? 4'b1011 : node7916;
																assign node7916 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7921 = (inp[2]) ? node7927 : node7922;
														assign node7922 = (inp[1]) ? node7924 : 4'b1111;
															assign node7924 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node7927 = (inp[5]) ? 4'b1011 : node7928;
															assign node7928 = (inp[1]) ? 4'b1110 : 4'b1010;
										assign node7932 = (inp[12]) ? node8012 : node7933;
											assign node7933 = (inp[1]) ? node7965 : node7934;
												assign node7934 = (inp[5]) ? node7946 : node7935;
													assign node7935 = (inp[13]) ? node7937 : 4'b1111;
														assign node7937 = (inp[4]) ? node7941 : node7938;
															assign node7938 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node7941 = (inp[2]) ? node7943 : 4'b1111;
																assign node7943 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7946 = (inp[4]) ? node7960 : node7947;
														assign node7947 = (inp[0]) ? node7953 : node7948;
															assign node7948 = (inp[2]) ? node7950 : 4'b1110;
																assign node7950 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node7953 = (inp[13]) ? node7957 : node7954;
																assign node7954 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node7957 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node7960 = (inp[2]) ? 4'b1110 : node7961;
															assign node7961 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node7965 = (inp[5]) ? node7989 : node7966;
													assign node7966 = (inp[2]) ? node7974 : node7967;
														assign node7967 = (inp[13]) ? 4'b1110 : node7968;
															assign node7968 = (inp[4]) ? node7970 : 4'b1110;
																assign node7970 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node7974 = (inp[0]) ? node7982 : node7975;
															assign node7975 = (inp[4]) ? node7979 : node7976;
																assign node7976 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node7979 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node7982 = (inp[4]) ? node7986 : node7983;
																assign node7983 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node7986 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node7989 = (inp[0]) ? node8003 : node7990;
														assign node7990 = (inp[2]) ? node7996 : node7991;
															assign node7991 = (inp[4]) ? node7993 : 4'b1111;
																assign node7993 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node7996 = (inp[4]) ? node8000 : node7997;
																assign node7997 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node8000 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node8003 = (inp[4]) ? 4'b1111 : node8004;
															assign node8004 = (inp[2]) ? node8008 : node8005;
																assign node8005 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node8008 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node8012 = (inp[2]) ? node8042 : node8013;
												assign node8013 = (inp[13]) ? node8023 : node8014;
													assign node8014 = (inp[5]) ? 4'b1000 : node8015;
														assign node8015 = (inp[1]) ? node8019 : node8016;
															assign node8016 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8019 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node8023 = (inp[1]) ? node8033 : node8024;
														assign node8024 = (inp[0]) ? node8026 : 4'b1100;
															assign node8026 = (inp[5]) ? node8030 : node8027;
																assign node8027 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node8030 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node8033 = (inp[5]) ? node8039 : node8034;
															assign node8034 = (inp[0]) ? node8036 : 4'b1000;
																assign node8036 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node8039 = (inp[4]) ? 4'b1100 : 4'b1101;
												assign node8042 = (inp[5]) ? node8072 : node8043;
													assign node8043 = (inp[4]) ? node8059 : node8044;
														assign node8044 = (inp[0]) ? node8052 : node8045;
															assign node8045 = (inp[13]) ? node8049 : node8046;
																assign node8046 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node8049 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node8052 = (inp[1]) ? node8056 : node8053;
																assign node8053 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node8056 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node8059 = (inp[0]) ? node8067 : node8060;
															assign node8060 = (inp[1]) ? node8064 : node8061;
																assign node8061 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node8064 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node8067 = (inp[13]) ? 4'b1101 : node8068;
																assign node8068 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node8072 = (inp[13]) ? 4'b1001 : 4'b1101;
									assign node8075 = (inp[5]) ? node8235 : node8076;
										assign node8076 = (inp[1]) ? node8154 : node8077;
											assign node8077 = (inp[12]) ? node8113 : node8078;
												assign node8078 = (inp[7]) ? node8094 : node8079;
													assign node8079 = (inp[13]) ? node8089 : node8080;
														assign node8080 = (inp[0]) ? node8082 : 4'b1000;
															assign node8082 = (inp[2]) ? node8086 : node8083;
																assign node8083 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node8086 = (inp[4]) ? 4'b1001 : 4'b1100;
														assign node8089 = (inp[4]) ? 4'b1101 : node8090;
															assign node8090 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node8094 = (inp[0]) ? node8104 : node8095;
														assign node8095 = (inp[13]) ? node8097 : 4'b1110;
															assign node8097 = (inp[4]) ? node8101 : node8098;
																assign node8098 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node8101 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node8104 = (inp[2]) ? node8106 : 4'b1010;
															assign node8106 = (inp[4]) ? node8110 : node8107;
																assign node8107 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node8110 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node8113 = (inp[7]) ? node8129 : node8114;
													assign node8114 = (inp[2]) ? node8122 : node8115;
														assign node8115 = (inp[13]) ? 4'b1110 : node8116;
															assign node8116 = (inp[0]) ? 4'b1010 : node8117;
																assign node8117 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node8122 = (inp[13]) ? 4'b1010 : node8123;
															assign node8123 = (inp[0]) ? node8125 : 4'b1110;
																assign node8125 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node8129 = (inp[4]) ? node8143 : node8130;
														assign node8130 = (inp[0]) ? node8138 : node8131;
															assign node8131 = (inp[2]) ? node8135 : node8132;
																assign node8132 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node8135 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node8138 = (inp[2]) ? node8140 : 4'b1100;
																assign node8140 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node8143 = (inp[2]) ? node8149 : node8144;
															assign node8144 = (inp[0]) ? node8146 : 4'b1000;
																assign node8146 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node8149 = (inp[13]) ? node8151 : 4'b1101;
																assign node8151 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node8154 = (inp[7]) ? node8196 : node8155;
												assign node8155 = (inp[12]) ? node8183 : node8156;
													assign node8156 = (inp[13]) ? node8170 : node8157;
														assign node8157 = (inp[0]) ? node8165 : node8158;
															assign node8158 = (inp[2]) ? node8162 : node8159;
																assign node8159 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node8162 = (inp[4]) ? 4'b1100 : 4'b1001;
															assign node8165 = (inp[4]) ? 4'b1001 : node8166;
																assign node8166 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node8170 = (inp[0]) ? node8176 : node8171;
															assign node8171 = (inp[2]) ? 4'b1000 : node8172;
																assign node8172 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node8176 = (inp[4]) ? node8180 : node8177;
																assign node8177 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node8180 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node8183 = (inp[2]) ? node8191 : node8184;
														assign node8184 = (inp[13]) ? node8188 : node8185;
															assign node8185 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node8188 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8191 = (inp[13]) ? 4'b1111 : node8192;
															assign node8192 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node8196 = (inp[12]) ? node8218 : node8197;
													assign node8197 = (inp[13]) ? node8209 : node8198;
														assign node8198 = (inp[0]) ? node8204 : node8199;
															assign node8199 = (inp[2]) ? 4'b1010 : node8200;
																assign node8200 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node8204 = (inp[2]) ? 4'b1011 : node8205;
																assign node8205 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node8209 = (inp[0]) ? 4'b1111 : node8210;
															assign node8210 = (inp[2]) ? node8214 : node8211;
																assign node8211 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node8214 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node8218 = (inp[0]) ? node8228 : node8219;
														assign node8219 = (inp[4]) ? 4'b1001 : node8220;
															assign node8220 = (inp[13]) ? node8224 : node8221;
																assign node8221 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node8224 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node8228 = (inp[4]) ? node8230 : 4'b1100;
															assign node8230 = (inp[2]) ? 4'b1000 : node8231;
																assign node8231 = (inp[13]) ? 4'b1001 : 4'b1101;
										assign node8235 = (inp[12]) ? node8293 : node8236;
											assign node8236 = (inp[7]) ? node8264 : node8237;
												assign node8237 = (inp[1]) ? node8249 : node8238;
													assign node8238 = (inp[4]) ? node8242 : node8239;
														assign node8239 = (inp[0]) ? 4'b1101 : 4'b1000;
														assign node8242 = (inp[0]) ? node8246 : node8243;
															assign node8243 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node8246 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node8249 = (inp[2]) ? node8259 : node8250;
														assign node8250 = (inp[4]) ? node8254 : node8251;
															assign node8251 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node8254 = (inp[13]) ? 4'b1001 : node8255;
																assign node8255 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8259 = (inp[0]) ? 4'b1001 : node8260;
															assign node8260 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node8264 = (inp[13]) ? node8276 : node8265;
													assign node8265 = (inp[1]) ? node8271 : node8266;
														assign node8266 = (inp[4]) ? node8268 : 4'b1011;
															assign node8268 = (inp[2]) ? 4'b1011 : 4'b1110;
														assign node8271 = (inp[4]) ? 4'b1011 : node8272;
															assign node8272 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node8276 = (inp[0]) ? node8278 : 4'b1010;
														assign node8278 = (inp[1]) ? node8286 : node8279;
															assign node8279 = (inp[2]) ? node8283 : node8280;
																assign node8280 = (inp[4]) ? 4'b1010 : 4'b1111;
																assign node8283 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node8286 = (inp[2]) ? node8290 : node8287;
																assign node8287 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node8290 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node8293 = (inp[7]) ? node8307 : node8294;
												assign node8294 = (inp[2]) ? node8304 : node8295;
													assign node8295 = (inp[13]) ? node8299 : node8296;
														assign node8296 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node8299 = (inp[0]) ? 4'b1110 : node8300;
															assign node8300 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node8304 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node8307 = (inp[2]) ? node8321 : node8308;
													assign node8308 = (inp[13]) ? node8312 : node8309;
														assign node8309 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node8312 = (inp[1]) ? node8316 : node8313;
															assign node8313 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8316 = (inp[0]) ? node8318 : 4'b1100;
																assign node8318 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node8321 = (inp[13]) ? 4'b1000 : 4'b1100;
				assign node8324 = (inp[7]) ? node12186 : node8325;
					assign node8325 = (inp[15]) ? node10247 : node8326;
						assign node8326 = (inp[10]) ? node9300 : node8327;
							assign node8327 = (inp[5]) ? node8789 : node8328;
								assign node8328 = (inp[13]) ? node8564 : node8329;
									assign node8329 = (inp[1]) ? node8451 : node8330;
										assign node8330 = (inp[12]) ? node8404 : node8331;
											assign node8331 = (inp[2]) ? node8365 : node8332;
												assign node8332 = (inp[0]) ? node8348 : node8333;
													assign node8333 = (inp[4]) ? node8341 : node8334;
														assign node8334 = (inp[3]) ? 4'b1001 : node8335;
															assign node8335 = (inp[9]) ? 4'b1001 : node8336;
																assign node8336 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node8341 = (inp[11]) ? node8345 : node8342;
															assign node8342 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node8345 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8348 = (inp[9]) ? node8354 : node8349;
														assign node8349 = (inp[3]) ? node8351 : 4'b1000;
															assign node8351 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8354 = (inp[4]) ? node8360 : node8355;
															assign node8355 = (inp[11]) ? 4'b1000 : node8356;
																assign node8356 = (inp[3]) ? 4'b1000 : 4'b1001;
															assign node8360 = (inp[3]) ? node8362 : 4'b1001;
																assign node8362 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node8365 = (inp[3]) ? node8389 : node8366;
													assign node8366 = (inp[11]) ? node8376 : node8367;
														assign node8367 = (inp[4]) ? node8369 : 4'b1001;
															assign node8369 = (inp[9]) ? node8373 : node8370;
																assign node8370 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node8373 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node8376 = (inp[4]) ? node8382 : node8377;
															assign node8377 = (inp[0]) ? node8379 : 4'b1000;
																assign node8379 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node8382 = (inp[0]) ? node8386 : node8383;
																assign node8383 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node8386 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8389 = (inp[9]) ? node8397 : node8390;
														assign node8390 = (inp[0]) ? node8392 : 4'b1001;
															assign node8392 = (inp[11]) ? 4'b1000 : node8393;
																assign node8393 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node8397 = (inp[0]) ? node8399 : 4'b1000;
															assign node8399 = (inp[4]) ? node8401 : 4'b1000;
																assign node8401 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node8404 = (inp[3]) ? node8434 : node8405;
												assign node8405 = (inp[4]) ? node8419 : node8406;
													assign node8406 = (inp[11]) ? 4'b1001 : node8407;
														assign node8407 = (inp[9]) ? node8413 : node8408;
															assign node8408 = (inp[2]) ? node8410 : 4'b1000;
																assign node8410 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node8413 = (inp[2]) ? node8415 : 4'b1001;
																assign node8415 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node8419 = (inp[11]) ? node8429 : node8420;
														assign node8420 = (inp[9]) ? node8424 : node8421;
															assign node8421 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8424 = (inp[0]) ? 4'b1101 : node8425;
																assign node8425 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node8429 = (inp[9]) ? 4'b1100 : node8430;
															assign node8430 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8434 = (inp[11]) ? node8444 : node8435;
													assign node8435 = (inp[9]) ? node8439 : node8436;
														assign node8436 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node8439 = (inp[0]) ? node8441 : 4'b1001;
															assign node8441 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node8444 = (inp[9]) ? 4'b1000 : node8445;
														assign node8445 = (inp[2]) ? node8447 : 4'b1001;
															assign node8447 = (inp[4]) ? 4'b1000 : 4'b1001;
										assign node8451 = (inp[3]) ? node8501 : node8452;
											assign node8452 = (inp[4]) ? node8476 : node8453;
												assign node8453 = (inp[12]) ? node8467 : node8454;
													assign node8454 = (inp[2]) ? node8460 : node8455;
														assign node8455 = (inp[11]) ? 4'b1000 : node8456;
															assign node8456 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8460 = (inp[11]) ? 4'b1001 : node8461;
															assign node8461 = (inp[0]) ? 4'b1000 : node8462;
																assign node8462 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node8467 = (inp[9]) ? node8473 : node8468;
														assign node8468 = (inp[2]) ? node8470 : 4'b1101;
															assign node8470 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8473 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node8476 = (inp[9]) ? node8486 : node8477;
													assign node8477 = (inp[11]) ? node8479 : 4'b1001;
														assign node8479 = (inp[2]) ? 4'b1000 : node8480;
															assign node8480 = (inp[12]) ? node8482 : 4'b1001;
																assign node8482 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node8486 = (inp[11]) ? node8494 : node8487;
														assign node8487 = (inp[2]) ? 4'b1000 : node8488;
															assign node8488 = (inp[12]) ? node8490 : 4'b1001;
																assign node8490 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node8494 = (inp[12]) ? 4'b1001 : node8495;
															assign node8495 = (inp[0]) ? 4'b1000 : node8496;
																assign node8496 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node8501 = (inp[11]) ? node8539 : node8502;
												assign node8502 = (inp[4]) ? node8526 : node8503;
													assign node8503 = (inp[12]) ? node8515 : node8504;
														assign node8504 = (inp[9]) ? node8510 : node8505;
															assign node8505 = (inp[0]) ? node8507 : 4'b1100;
																assign node8507 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node8510 = (inp[2]) ? 4'b1101 : node8511;
																assign node8511 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8515 = (inp[9]) ? node8521 : node8516;
															assign node8516 = (inp[0]) ? 4'b1001 : node8517;
																assign node8517 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node8521 = (inp[2]) ? node8523 : 4'b1000;
																assign node8523 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node8526 = (inp[12]) ? node8532 : node8527;
														assign node8527 = (inp[9]) ? node8529 : 4'b1000;
															assign node8529 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8532 = (inp[2]) ? node8534 : 4'b1100;
															assign node8534 = (inp[9]) ? node8536 : 4'b1100;
																assign node8536 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8539 = (inp[2]) ? node8553 : node8540;
													assign node8540 = (inp[12]) ? node8550 : node8541;
														assign node8541 = (inp[4]) ? 4'b1001 : node8542;
															assign node8542 = (inp[9]) ? node8546 : node8543;
																assign node8543 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node8546 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8550 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node8553 = (inp[4]) ? node8559 : node8554;
														assign node8554 = (inp[12]) ? node8556 : 4'b1100;
															assign node8556 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8559 = (inp[0]) ? 4'b1001 : node8560;
															assign node8560 = (inp[9]) ? 4'b1101 : 4'b1100;
									assign node8564 = (inp[1]) ? node8670 : node8565;
										assign node8565 = (inp[3]) ? node8617 : node8566;
											assign node8566 = (inp[12]) ? node8594 : node8567;
												assign node8567 = (inp[9]) ? node8581 : node8568;
													assign node8568 = (inp[11]) ? node8574 : node8569;
														assign node8569 = (inp[2]) ? node8571 : 4'b1100;
															assign node8571 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8574 = (inp[2]) ? node8576 : 4'b1101;
															assign node8576 = (inp[4]) ? 4'b1100 : node8577;
																assign node8577 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node8581 = (inp[0]) ? node8587 : node8582;
														assign node8582 = (inp[11]) ? node8584 : 4'b1101;
															assign node8584 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node8587 = (inp[4]) ? node8591 : node8588;
															assign node8588 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node8591 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node8594 = (inp[4]) ? node8606 : node8595;
													assign node8595 = (inp[2]) ? node8597 : 4'b1101;
														assign node8597 = (inp[0]) ? 4'b1101 : node8598;
															assign node8598 = (inp[9]) ? node8602 : node8599;
																assign node8599 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node8602 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node8606 = (inp[11]) ? node8614 : node8607;
														assign node8607 = (inp[2]) ? 4'b1001 : node8608;
															assign node8608 = (inp[0]) ? 4'b1000 : node8609;
																assign node8609 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8614 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node8617 = (inp[11]) ? node8645 : node8618;
												assign node8618 = (inp[9]) ? node8634 : node8619;
													assign node8619 = (inp[0]) ? node8629 : node8620;
														assign node8620 = (inp[12]) ? node8624 : node8621;
															assign node8621 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node8624 = (inp[2]) ? 4'b1101 : node8625;
																assign node8625 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node8629 = (inp[2]) ? node8631 : 4'b1100;
															assign node8631 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node8634 = (inp[0]) ? 4'b1101 : node8635;
														assign node8635 = (inp[4]) ? node8639 : node8636;
															assign node8636 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node8639 = (inp[2]) ? 4'b1101 : node8640;
																assign node8640 = (inp[12]) ? 4'b1100 : 4'b1101;
												assign node8645 = (inp[9]) ? node8657 : node8646;
													assign node8646 = (inp[2]) ? node8648 : 4'b1101;
														assign node8648 = (inp[4]) ? node8652 : node8649;
															assign node8649 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node8652 = (inp[0]) ? node8654 : 4'b1101;
																assign node8654 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node8657 = (inp[2]) ? node8659 : 4'b1100;
														assign node8659 = (inp[12]) ? node8665 : node8660;
															assign node8660 = (inp[4]) ? 4'b1101 : node8661;
																assign node8661 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8665 = (inp[4]) ? 4'b1100 : node8666;
																assign node8666 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node8670 = (inp[3]) ? node8724 : node8671;
											assign node8671 = (inp[4]) ? node8695 : node8672;
												assign node8672 = (inp[12]) ? node8686 : node8673;
													assign node8673 = (inp[9]) ? node8679 : node8674;
														assign node8674 = (inp[11]) ? node8676 : 4'b1100;
															assign node8676 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node8679 = (inp[11]) ? node8681 : 4'b1101;
															assign node8681 = (inp[0]) ? node8683 : 4'b1100;
																assign node8683 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node8686 = (inp[11]) ? node8690 : node8687;
														assign node8687 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8690 = (inp[9]) ? 4'b1000 : node8691;
															assign node8691 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node8695 = (inp[9]) ? node8709 : node8696;
													assign node8696 = (inp[11]) ? node8704 : node8697;
														assign node8697 = (inp[2]) ? 4'b1101 : node8698;
															assign node8698 = (inp[12]) ? node8700 : 4'b1100;
																assign node8700 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8704 = (inp[0]) ? 4'b1101 : node8705;
															assign node8705 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node8709 = (inp[11]) ? node8717 : node8710;
														assign node8710 = (inp[12]) ? 4'b1100 : node8711;
															assign node8711 = (inp[2]) ? node8713 : 4'b1101;
																assign node8713 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8717 = (inp[2]) ? 4'b1101 : node8718;
															assign node8718 = (inp[0]) ? 4'b1100 : node8719;
																assign node8719 = (inp[12]) ? 4'b1101 : 4'b1100;
											assign node8724 = (inp[4]) ? node8760 : node8725;
												assign node8725 = (inp[12]) ? node8745 : node8726;
													assign node8726 = (inp[9]) ? node8734 : node8727;
														assign node8727 = (inp[11]) ? node8729 : 4'b1001;
															assign node8729 = (inp[0]) ? node8731 : 4'b1000;
																assign node8731 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node8734 = (inp[11]) ? node8740 : node8735;
															assign node8735 = (inp[2]) ? 4'b1000 : node8736;
																assign node8736 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node8740 = (inp[2]) ? 4'b1001 : node8741;
																assign node8741 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node8745 = (inp[9]) ? node8753 : node8746;
														assign node8746 = (inp[11]) ? node8748 : 4'b1100;
															assign node8748 = (inp[2]) ? 4'b1101 : node8749;
																assign node8749 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8753 = (inp[0]) ? node8755 : 4'b1101;
															assign node8755 = (inp[11]) ? 4'b1101 : node8756;
																assign node8756 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node8760 = (inp[12]) ? node8774 : node8761;
													assign node8761 = (inp[0]) ? node8769 : node8762;
														assign node8762 = (inp[11]) ? node8764 : 4'b1100;
															assign node8764 = (inp[2]) ? 4'b1100 : node8765;
																assign node8765 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node8769 = (inp[11]) ? 4'b1101 : node8770;
															assign node8770 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node8774 = (inp[11]) ? node8784 : node8775;
														assign node8775 = (inp[9]) ? node8781 : node8776;
															assign node8776 = (inp[2]) ? node8778 : 4'b1000;
																assign node8778 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node8781 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node8784 = (inp[9]) ? 4'b1000 : node8785;
															assign node8785 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node8789 = (inp[13]) ? node9037 : node8790;
									assign node8790 = (inp[1]) ? node8888 : node8791;
										assign node8791 = (inp[3]) ? node8845 : node8792;
											assign node8792 = (inp[4]) ? node8812 : node8793;
												assign node8793 = (inp[11]) ? node8803 : node8794;
													assign node8794 = (inp[9]) ? node8798 : node8795;
														assign node8795 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8798 = (inp[2]) ? node8800 : 4'b1101;
															assign node8800 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node8803 = (inp[9]) ? node8807 : node8804;
														assign node8804 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node8807 = (inp[2]) ? node8809 : 4'b1100;
															assign node8809 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8812 = (inp[12]) ? node8824 : node8813;
													assign node8813 = (inp[2]) ? node8821 : node8814;
														assign node8814 = (inp[11]) ? 4'b1100 : node8815;
															assign node8815 = (inp[9]) ? 4'b1101 : node8816;
																assign node8816 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node8821 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node8824 = (inp[2]) ? node8830 : node8825;
														assign node8825 = (inp[11]) ? node8827 : 4'b1000;
															assign node8827 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8830 = (inp[9]) ? node8838 : node8831;
															assign node8831 = (inp[0]) ? node8835 : node8832;
																assign node8832 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node8835 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node8838 = (inp[0]) ? node8842 : node8839;
																assign node8839 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node8842 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node8845 = (inp[2]) ? node8869 : node8846;
												assign node8846 = (inp[4]) ? node8860 : node8847;
													assign node8847 = (inp[0]) ? node8855 : node8848;
														assign node8848 = (inp[11]) ? node8852 : node8849;
															assign node8849 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node8852 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node8855 = (inp[11]) ? node8857 : 4'b1101;
															assign node8857 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node8860 = (inp[0]) ? node8862 : 4'b1101;
														assign node8862 = (inp[9]) ? node8866 : node8863;
															assign node8863 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node8866 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node8869 = (inp[11]) ? node8879 : node8870;
													assign node8870 = (inp[9]) ? 4'b1101 : node8871;
														assign node8871 = (inp[4]) ? node8873 : 4'b1100;
															assign node8873 = (inp[0]) ? node8875 : 4'b1100;
																assign node8875 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node8879 = (inp[9]) ? 4'b1100 : node8880;
														assign node8880 = (inp[12]) ? 4'b1101 : node8881;
															assign node8881 = (inp[0]) ? node8883 : 4'b1101;
																assign node8883 = (inp[4]) ? 4'b1100 : 4'b1101;
										assign node8888 = (inp[4]) ? node8964 : node8889;
											assign node8889 = (inp[3]) ? node8921 : node8890;
												assign node8890 = (inp[12]) ? node8900 : node8891;
													assign node8891 = (inp[9]) ? 4'b1100 : node8892;
														assign node8892 = (inp[2]) ? node8894 : 4'b1101;
															assign node8894 = (inp[0]) ? node8896 : 4'b1100;
																assign node8896 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node8900 = (inp[2]) ? node8914 : node8901;
														assign node8901 = (inp[9]) ? node8907 : node8902;
															assign node8902 = (inp[0]) ? 4'b1001 : node8903;
																assign node8903 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node8907 = (inp[0]) ? node8911 : node8908;
																assign node8908 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node8911 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8914 = (inp[11]) ? node8918 : node8915;
															assign node8915 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node8918 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node8921 = (inp[12]) ? node8943 : node8922;
													assign node8922 = (inp[0]) ? node8932 : node8923;
														assign node8923 = (inp[2]) ? 4'b1000 : node8924;
															assign node8924 = (inp[9]) ? node8928 : node8925;
																assign node8925 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node8928 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8932 = (inp[2]) ? node8938 : node8933;
															assign node8933 = (inp[11]) ? 4'b1000 : node8934;
																assign node8934 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node8938 = (inp[11]) ? node8940 : 4'b1001;
																assign node8940 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8943 = (inp[2]) ? node8949 : node8944;
														assign node8944 = (inp[11]) ? node8946 : 4'b1100;
															assign node8946 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node8949 = (inp[9]) ? node8957 : node8950;
															assign node8950 = (inp[11]) ? node8954 : node8951;
																assign node8951 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node8954 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8957 = (inp[11]) ? node8961 : node8958;
																assign node8958 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node8961 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node8964 = (inp[3]) ? node9002 : node8965;
												assign node8965 = (inp[2]) ? node8983 : node8966;
													assign node8966 = (inp[0]) ? node8974 : node8967;
														assign node8967 = (inp[9]) ? node8971 : node8968;
															assign node8968 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node8971 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node8974 = (inp[11]) ? node8976 : 4'b1101;
															assign node8976 = (inp[9]) ? node8980 : node8977;
																assign node8977 = (inp[12]) ? 4'b1101 : 4'b1100;
																assign node8980 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node8983 = (inp[12]) ? node8997 : node8984;
														assign node8984 = (inp[0]) ? node8990 : node8985;
															assign node8985 = (inp[9]) ? node8987 : 4'b1101;
																assign node8987 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node8990 = (inp[11]) ? node8994 : node8991;
																assign node8991 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node8994 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node8997 = (inp[11]) ? 4'b1101 : node8998;
															assign node8998 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node9002 = (inp[12]) ? node9016 : node9003;
													assign node9003 = (inp[11]) ? node9005 : 4'b1101;
														assign node9005 = (inp[9]) ? node9011 : node9006;
															assign node9006 = (inp[0]) ? 4'b1101 : node9007;
																assign node9007 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9011 = (inp[2]) ? 4'b1100 : node9012;
																assign node9012 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node9016 = (inp[0]) ? node9024 : node9017;
														assign node9017 = (inp[11]) ? node9021 : node9018;
															assign node9018 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9021 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node9024 = (inp[11]) ? node9030 : node9025;
															assign node9025 = (inp[2]) ? node9027 : 4'b1001;
																assign node9027 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9030 = (inp[2]) ? node9034 : node9031;
																assign node9031 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node9034 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node9037 = (inp[1]) ? node9161 : node9038;
										assign node9038 = (inp[3]) ? node9094 : node9039;
											assign node9039 = (inp[4]) ? node9069 : node9040;
												assign node9040 = (inp[2]) ? node9062 : node9041;
													assign node9041 = (inp[12]) ? node9055 : node9042;
														assign node9042 = (inp[0]) ? node9048 : node9043;
															assign node9043 = (inp[11]) ? 4'b1001 : node9044;
																assign node9044 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9048 = (inp[9]) ? node9052 : node9049;
																assign node9049 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node9052 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9055 = (inp[11]) ? node9057 : 4'b1001;
															assign node9057 = (inp[9]) ? node9059 : 4'b1001;
																assign node9059 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node9062 = (inp[9]) ? node9066 : node9063;
														assign node9063 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9066 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node9069 = (inp[12]) ? node9083 : node9070;
													assign node9070 = (inp[2]) ? node9078 : node9071;
														assign node9071 = (inp[9]) ? node9075 : node9072;
															assign node9072 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9075 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9078 = (inp[9]) ? 4'b1000 : node9079;
															assign node9079 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9083 = (inp[11]) ? node9089 : node9084;
														assign node9084 = (inp[9]) ? 4'b1100 : node9085;
															assign node9085 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node9089 = (inp[9]) ? 4'b1101 : node9090;
															assign node9090 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node9094 = (inp[12]) ? node9124 : node9095;
												assign node9095 = (inp[11]) ? node9107 : node9096;
													assign node9096 = (inp[9]) ? node9102 : node9097;
														assign node9097 = (inp[4]) ? node9099 : 4'b1001;
															assign node9099 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node9102 = (inp[2]) ? node9104 : 4'b1000;
															assign node9104 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node9107 = (inp[9]) ? node9115 : node9108;
														assign node9108 = (inp[0]) ? node9110 : 4'b1000;
															assign node9110 = (inp[2]) ? node9112 : 4'b1001;
																assign node9112 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node9115 = (inp[0]) ? node9117 : 4'b1001;
															assign node9117 = (inp[2]) ? node9121 : node9118;
																assign node9118 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node9121 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node9124 = (inp[11]) ? node9142 : node9125;
													assign node9125 = (inp[9]) ? node9135 : node9126;
														assign node9126 = (inp[2]) ? 4'b1001 : node9127;
															assign node9127 = (inp[4]) ? node9131 : node9128;
																assign node9128 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node9131 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node9135 = (inp[2]) ? 4'b1000 : node9136;
															assign node9136 = (inp[4]) ? 4'b1001 : node9137;
																assign node9137 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node9142 = (inp[9]) ? node9152 : node9143;
														assign node9143 = (inp[2]) ? 4'b1000 : node9144;
															assign node9144 = (inp[0]) ? node9148 : node9145;
																assign node9145 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node9148 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node9152 = (inp[2]) ? 4'b1001 : node9153;
															assign node9153 = (inp[0]) ? node9157 : node9154;
																assign node9154 = (inp[4]) ? 4'b1000 : 4'b1001;
																assign node9157 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node9161 = (inp[3]) ? node9215 : node9162;
											assign node9162 = (inp[4]) ? node9192 : node9163;
												assign node9163 = (inp[12]) ? node9179 : node9164;
													assign node9164 = (inp[0]) ? node9172 : node9165;
														assign node9165 = (inp[11]) ? 4'b1000 : node9166;
															assign node9166 = (inp[2]) ? 4'b1001 : node9167;
																assign node9167 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node9172 = (inp[11]) ? node9176 : node9173;
															assign node9173 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9176 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node9179 = (inp[9]) ? node9185 : node9180;
														assign node9180 = (inp[11]) ? 4'b1101 : node9181;
															assign node9181 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node9185 = (inp[11]) ? node9189 : node9186;
															assign node9186 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9189 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node9192 = (inp[12]) ? node9200 : node9193;
													assign node9193 = (inp[11]) ? node9195 : 4'b1001;
														assign node9195 = (inp[9]) ? node9197 : 4'b1000;
															assign node9197 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node9200 = (inp[9]) ? node9206 : node9201;
														assign node9201 = (inp[11]) ? node9203 : 4'b1000;
															assign node9203 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node9206 = (inp[11]) ? node9212 : node9207;
															assign node9207 = (inp[0]) ? node9209 : 4'b1001;
																assign node9209 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node9212 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node9215 = (inp[0]) ? node9265 : node9216;
												assign node9216 = (inp[12]) ? node9238 : node9217;
													assign node9217 = (inp[4]) ? node9231 : node9218;
														assign node9218 = (inp[2]) ? node9224 : node9219;
															assign node9219 = (inp[9]) ? node9221 : 4'b1100;
																assign node9221 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node9224 = (inp[11]) ? node9228 : node9225;
																assign node9225 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node9228 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node9231 = (inp[9]) ? node9233 : 4'b1000;
															assign node9233 = (inp[2]) ? node9235 : 4'b1001;
																assign node9235 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9238 = (inp[4]) ? node9252 : node9239;
														assign node9239 = (inp[11]) ? node9245 : node9240;
															assign node9240 = (inp[2]) ? node9242 : 4'b1001;
																assign node9242 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9245 = (inp[9]) ? node9249 : node9246;
																assign node9246 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node9249 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9252 = (inp[9]) ? node9258 : node9253;
															assign node9253 = (inp[11]) ? node9255 : 4'b1101;
																assign node9255 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9258 = (inp[11]) ? node9262 : node9259;
																assign node9259 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node9262 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node9265 = (inp[2]) ? node9289 : node9266;
													assign node9266 = (inp[11]) ? node9280 : node9267;
														assign node9267 = (inp[9]) ? node9273 : node9268;
															assign node9268 = (inp[4]) ? 4'b1001 : node9269;
																assign node9269 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node9273 = (inp[12]) ? node9277 : node9274;
																assign node9274 = (inp[4]) ? 4'b1000 : 4'b1101;
																assign node9277 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9280 = (inp[9]) ? node9284 : node9281;
															assign node9281 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node9284 = (inp[12]) ? node9286 : 4'b1100;
																assign node9286 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9289 = (inp[9]) ? 4'b1001 : node9290;
														assign node9290 = (inp[12]) ? node9294 : node9291;
															assign node9291 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9294 = (inp[4]) ? 4'b1101 : node9295;
																assign node9295 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node9300 = (inp[3]) ? node9798 : node9301;
								assign node9301 = (inp[0]) ? node9547 : node9302;
									assign node9302 = (inp[9]) ? node9414 : node9303;
										assign node9303 = (inp[11]) ? node9361 : node9304;
											assign node9304 = (inp[4]) ? node9326 : node9305;
												assign node9305 = (inp[1]) ? node9315 : node9306;
													assign node9306 = (inp[5]) ? node9310 : node9307;
														assign node9307 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node9310 = (inp[13]) ? node9312 : 4'b1100;
															assign node9312 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node9315 = (inp[12]) ? node9323 : node9316;
														assign node9316 = (inp[2]) ? node9318 : 4'b1000;
															assign node9318 = (inp[5]) ? 4'b1100 : node9319;
																assign node9319 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node9323 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node9326 = (inp[1]) ? node9348 : node9327;
													assign node9327 = (inp[13]) ? node9339 : node9328;
														assign node9328 = (inp[12]) ? node9334 : node9329;
															assign node9329 = (inp[5]) ? 4'b1100 : node9330;
																assign node9330 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node9334 = (inp[5]) ? node9336 : 4'b1100;
																assign node9336 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node9339 = (inp[5]) ? node9343 : node9340;
															assign node9340 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node9343 = (inp[2]) ? node9345 : 4'b1101;
																assign node9345 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node9348 = (inp[5]) ? node9356 : node9349;
														assign node9349 = (inp[13]) ? node9351 : 4'b1001;
															assign node9351 = (inp[12]) ? 4'b1101 : node9352;
																assign node9352 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node9356 = (inp[13]) ? 4'b1000 : node9357;
															assign node9357 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node9361 = (inp[4]) ? node9383 : node9362;
												assign node9362 = (inp[1]) ? node9372 : node9363;
													assign node9363 = (inp[5]) ? node9367 : node9364;
														assign node9364 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node9367 = (inp[13]) ? node9369 : 4'b1101;
															assign node9369 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node9372 = (inp[12]) ? node9380 : node9373;
														assign node9373 = (inp[5]) ? node9377 : node9374;
															assign node9374 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node9377 = (inp[2]) ? 4'b1000 : 4'b1101;
														assign node9380 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node9383 = (inp[2]) ? node9403 : node9384;
													assign node9384 = (inp[12]) ? node9392 : node9385;
														assign node9385 = (inp[13]) ? node9389 : node9386;
															assign node9386 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node9389 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node9392 = (inp[1]) ? node9400 : node9393;
															assign node9393 = (inp[5]) ? node9397 : node9394;
																assign node9394 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node9397 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node9400 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node9403 = (inp[5]) ? node9409 : node9404;
														assign node9404 = (inp[13]) ? node9406 : 4'b1000;
															assign node9406 = (inp[12]) ? 4'b1001 : 4'b1100;
														assign node9409 = (inp[13]) ? 4'b1001 : node9410;
															assign node9410 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node9414 = (inp[11]) ? node9478 : node9415;
											assign node9415 = (inp[1]) ? node9439 : node9416;
												assign node9416 = (inp[4]) ? node9426 : node9417;
													assign node9417 = (inp[13]) ? node9421 : node9418;
														assign node9418 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node9421 = (inp[5]) ? node9423 : 4'b1101;
															assign node9423 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node9426 = (inp[13]) ? node9432 : node9427;
														assign node9427 = (inp[2]) ? node9429 : 4'b1101;
															assign node9429 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node9432 = (inp[12]) ? node9436 : node9433;
															assign node9433 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node9436 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node9439 = (inp[12]) ? node9461 : node9440;
													assign node9440 = (inp[2]) ? node9452 : node9441;
														assign node9441 = (inp[4]) ? node9447 : node9442;
															assign node9442 = (inp[5]) ? 4'b1101 : node9443;
																assign node9443 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node9447 = (inp[13]) ? node9449 : 4'b1101;
																assign node9449 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node9452 = (inp[5]) ? node9458 : node9453;
															assign node9453 = (inp[13]) ? node9455 : 4'b1000;
																assign node9455 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node9458 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node9461 = (inp[5]) ? node9467 : node9462;
														assign node9462 = (inp[13]) ? node9464 : 4'b1100;
															assign node9464 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9467 = (inp[13]) ? node9473 : node9468;
															assign node9468 = (inp[4]) ? 4'b1100 : node9469;
																assign node9469 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node9473 = (inp[4]) ? 4'b1001 : node9474;
																assign node9474 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node9478 = (inp[4]) ? node9518 : node9479;
												assign node9479 = (inp[12]) ? node9499 : node9480;
													assign node9480 = (inp[1]) ? node9492 : node9481;
														assign node9481 = (inp[2]) ? node9489 : node9482;
															assign node9482 = (inp[5]) ? node9486 : node9483;
																assign node9483 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node9486 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node9489 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node9492 = (inp[5]) ? node9496 : node9493;
															assign node9493 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node9496 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node9499 = (inp[1]) ? node9511 : node9500;
														assign node9500 = (inp[2]) ? node9506 : node9501;
															assign node9501 = (inp[5]) ? node9503 : 4'b1100;
																assign node9503 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node9506 = (inp[5]) ? 4'b1100 : node9507;
																assign node9507 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node9511 = (inp[13]) ? 4'b1100 : node9512;
															assign node9512 = (inp[5]) ? node9514 : 4'b1101;
																assign node9514 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node9518 = (inp[1]) ? node9538 : node9519;
													assign node9519 = (inp[5]) ? node9529 : node9520;
														assign node9520 = (inp[2]) ? 4'b1001 : node9521;
															assign node9521 = (inp[13]) ? node9525 : node9522;
																assign node9522 = (inp[12]) ? 4'b1100 : 4'b1000;
																assign node9525 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node9529 = (inp[2]) ? node9535 : node9530;
															assign node9530 = (inp[12]) ? node9532 : 4'b1001;
																assign node9532 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node9535 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node9538 = (inp[5]) ? node9544 : node9539;
														assign node9539 = (inp[13]) ? 4'b1101 : node9540;
															assign node9540 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9544 = (inp[13]) ? 4'b1000 : 4'b1100;
									assign node9547 = (inp[13]) ? node9685 : node9548;
										assign node9548 = (inp[5]) ? node9610 : node9549;
											assign node9549 = (inp[12]) ? node9567 : node9550;
												assign node9550 = (inp[11]) ? node9562 : node9551;
													assign node9551 = (inp[9]) ? node9557 : node9552;
														assign node9552 = (inp[4]) ? 4'b1000 : node9553;
															assign node9553 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9557 = (inp[4]) ? 4'b1001 : node9558;
															assign node9558 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node9562 = (inp[9]) ? 4'b1000 : node9563;
														assign node9563 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node9567 = (inp[11]) ? node9589 : node9568;
													assign node9568 = (inp[9]) ? node9576 : node9569;
														assign node9569 = (inp[4]) ? 4'b1100 : node9570;
															assign node9570 = (inp[1]) ? 4'b1100 : node9571;
																assign node9571 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9576 = (inp[1]) ? node9582 : node9577;
															assign node9577 = (inp[4]) ? 4'b1101 : node9578;
																assign node9578 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node9582 = (inp[4]) ? node9586 : node9583;
																assign node9583 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node9586 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node9589 = (inp[9]) ? node9601 : node9590;
														assign node9590 = (inp[2]) ? node9596 : node9591;
															assign node9591 = (inp[4]) ? node9593 : 4'b1001;
																assign node9593 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node9596 = (inp[4]) ? 4'b1101 : node9597;
																assign node9597 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node9601 = (inp[2]) ? 4'b1001 : node9602;
															assign node9602 = (inp[1]) ? node9606 : node9603;
																assign node9603 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node9606 = (inp[4]) ? 4'b1000 : 4'b1101;
											assign node9610 = (inp[12]) ? node9646 : node9611;
												assign node9611 = (inp[11]) ? node9627 : node9612;
													assign node9612 = (inp[2]) ? node9618 : node9613;
														assign node9613 = (inp[9]) ? node9615 : 4'b1100;
															assign node9615 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node9618 = (inp[1]) ? node9624 : node9619;
															assign node9619 = (inp[4]) ? 4'b1100 : node9620;
																assign node9620 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node9624 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node9627 = (inp[2]) ? node9633 : node9628;
														assign node9628 = (inp[9]) ? node9630 : 4'b1101;
															assign node9630 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node9633 = (inp[1]) ? node9639 : node9634;
															assign node9634 = (inp[4]) ? 4'b1100 : node9635;
																assign node9635 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node9639 = (inp[4]) ? node9643 : node9640;
																assign node9640 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node9643 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node9646 = (inp[1]) ? node9668 : node9647;
													assign node9647 = (inp[4]) ? node9655 : node9648;
														assign node9648 = (inp[9]) ? 4'b1100 : node9649;
															assign node9649 = (inp[11]) ? 4'b1100 : node9650;
																assign node9650 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node9655 = (inp[2]) ? node9663 : node9656;
															assign node9656 = (inp[11]) ? node9660 : node9657;
																assign node9657 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node9660 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node9663 = (inp[11]) ? 4'b1000 : node9664;
																assign node9664 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node9668 = (inp[4]) ? node9676 : node9669;
														assign node9669 = (inp[2]) ? node9671 : 4'b1001;
															assign node9671 = (inp[9]) ? node9673 : 4'b1000;
																assign node9673 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9676 = (inp[2]) ? node9678 : 4'b1101;
															assign node9678 = (inp[11]) ? node9682 : node9679;
																assign node9679 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node9682 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node9685 = (inp[5]) ? node9745 : node9686;
											assign node9686 = (inp[12]) ? node9704 : node9687;
												assign node9687 = (inp[9]) ? node9697 : node9688;
													assign node9688 = (inp[11]) ? node9694 : node9689;
														assign node9689 = (inp[4]) ? 4'b1100 : node9690;
															assign node9690 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node9694 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node9697 = (inp[11]) ? node9699 : 4'b1101;
														assign node9699 = (inp[4]) ? 4'b1100 : node9700;
															assign node9700 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node9704 = (inp[9]) ? node9720 : node9705;
													assign node9705 = (inp[4]) ? node9717 : node9706;
														assign node9706 = (inp[1]) ? node9714 : node9707;
															assign node9707 = (inp[11]) ? node9711 : node9708;
																assign node9708 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node9711 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node9714 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node9717 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node9720 = (inp[11]) ? node9734 : node9721;
														assign node9721 = (inp[4]) ? node9727 : node9722;
															assign node9722 = (inp[1]) ? 4'b1001 : node9723;
																assign node9723 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node9727 = (inp[1]) ? node9731 : node9728;
																assign node9728 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node9731 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node9734 = (inp[2]) ? node9738 : node9735;
															assign node9735 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node9738 = (inp[4]) ? node9742 : node9739;
																assign node9739 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node9742 = (inp[1]) ? 4'b1101 : 4'b1000;
											assign node9745 = (inp[12]) ? node9765 : node9746;
												assign node9746 = (inp[4]) ? node9760 : node9747;
													assign node9747 = (inp[2]) ? node9753 : node9748;
														assign node9748 = (inp[11]) ? node9750 : 4'b1001;
															assign node9750 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node9753 = (inp[11]) ? node9757 : node9754;
															assign node9754 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9757 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node9760 = (inp[9]) ? node9762 : 4'b1001;
														assign node9762 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node9765 = (inp[1]) ? node9781 : node9766;
													assign node9766 = (inp[4]) ? node9774 : node9767;
														assign node9767 = (inp[11]) ? node9771 : node9768;
															assign node9768 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node9771 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node9774 = (inp[11]) ? node9778 : node9775;
															assign node9775 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node9778 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node9781 = (inp[4]) ? node9789 : node9782;
														assign node9782 = (inp[9]) ? node9786 : node9783;
															assign node9783 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node9786 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node9789 = (inp[9]) ? 4'b1000 : node9790;
															assign node9790 = (inp[11]) ? node9794 : node9791;
																assign node9791 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node9794 = (inp[2]) ? 4'b1001 : 4'b1000;
								assign node9798 = (inp[9]) ? node10024 : node9799;
									assign node9799 = (inp[11]) ? node9909 : node9800;
										assign node9800 = (inp[5]) ? node9848 : node9801;
											assign node9801 = (inp[13]) ? node9825 : node9802;
												assign node9802 = (inp[1]) ? node9812 : node9803;
													assign node9803 = (inp[12]) ? 4'b1000 : node9804;
														assign node9804 = (inp[0]) ? 4'b1001 : node9805;
															assign node9805 = (inp[2]) ? node9807 : 4'b1000;
																assign node9807 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node9812 = (inp[0]) ? node9818 : node9813;
														assign node9813 = (inp[4]) ? 4'b1000 : node9814;
															assign node9814 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node9818 = (inp[4]) ? 4'b1100 : node9819;
															assign node9819 = (inp[12]) ? 4'b1001 : node9820;
																assign node9820 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node9825 = (inp[1]) ? node9835 : node9826;
													assign node9826 = (inp[2]) ? node9828 : 4'b1100;
														assign node9828 = (inp[0]) ? node9832 : node9829;
															assign node9829 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node9832 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node9835 = (inp[4]) ? node9845 : node9836;
														assign node9836 = (inp[12]) ? node9840 : node9837;
															assign node9837 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node9840 = (inp[0]) ? node9842 : 4'b1100;
																assign node9842 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node9845 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node9848 = (inp[13]) ? node9888 : node9849;
												assign node9849 = (inp[1]) ? node9867 : node9850;
													assign node9850 = (inp[0]) ? node9856 : node9851;
														assign node9851 = (inp[12]) ? node9853 : 4'b1100;
															assign node9853 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node9856 = (inp[12]) ? node9862 : node9857;
															assign node9857 = (inp[2]) ? 4'b1101 : node9858;
																assign node9858 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node9862 = (inp[4]) ? 4'b1100 : node9863;
																assign node9863 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node9867 = (inp[12]) ? node9879 : node9868;
														assign node9868 = (inp[4]) ? node9874 : node9869;
															assign node9869 = (inp[2]) ? node9871 : 4'b1000;
																assign node9871 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node9874 = (inp[0]) ? 4'b1100 : node9875;
																assign node9875 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node9879 = (inp[4]) ? node9885 : node9880;
															assign node9880 = (inp[2]) ? node9882 : 4'b1101;
																assign node9882 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node9885 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node9888 = (inp[1]) ? node9894 : node9889;
													assign node9889 = (inp[0]) ? node9891 : 4'b1001;
														assign node9891 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node9894 = (inp[12]) ? node9902 : node9895;
														assign node9895 = (inp[4]) ? node9897 : 4'b1101;
															assign node9897 = (inp[0]) ? 4'b1001 : node9898;
																assign node9898 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9902 = (inp[4]) ? 4'b1101 : node9903;
															assign node9903 = (inp[0]) ? 4'b1000 : node9904;
																assign node9904 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node9909 = (inp[5]) ? node9971 : node9910;
											assign node9910 = (inp[13]) ? node9938 : node9911;
												assign node9911 = (inp[0]) ? node9921 : node9912;
													assign node9912 = (inp[1]) ? node9918 : node9913;
														assign node9913 = (inp[2]) ? node9915 : 4'b1001;
															assign node9915 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node9918 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node9921 = (inp[1]) ? node9927 : node9922;
														assign node9922 = (inp[12]) ? node9924 : 4'b1000;
															assign node9924 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node9927 = (inp[12]) ? node9933 : node9928;
															assign node9928 = (inp[4]) ? 4'b1001 : node9929;
																assign node9929 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9933 = (inp[4]) ? node9935 : 4'b1000;
																assign node9935 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node9938 = (inp[1]) ? node9956 : node9939;
													assign node9939 = (inp[2]) ? node9945 : node9940;
														assign node9940 = (inp[4]) ? node9942 : 4'b1101;
															assign node9942 = (inp[12]) ? 4'b1100 : 4'b1101;
														assign node9945 = (inp[12]) ? node9951 : node9946;
															assign node9946 = (inp[4]) ? node9948 : 4'b1100;
																assign node9948 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node9951 = (inp[0]) ? 4'b1101 : node9952;
																assign node9952 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node9956 = (inp[4]) ? node9964 : node9957;
														assign node9957 = (inp[12]) ? node9959 : 4'b1000;
															assign node9959 = (inp[2]) ? 4'b1101 : node9960;
																assign node9960 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node9964 = (inp[12]) ? node9968 : node9965;
															assign node9965 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9968 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node9971 = (inp[13]) ? node9995 : node9972;
												assign node9972 = (inp[1]) ? node9984 : node9973;
													assign node9973 = (inp[0]) ? node9975 : 4'b1101;
														assign node9975 = (inp[4]) ? node9979 : node9976;
															assign node9976 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node9979 = (inp[2]) ? node9981 : 4'b1101;
																assign node9981 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node9984 = (inp[12]) ? node9990 : node9985;
														assign node9985 = (inp[4]) ? 4'b1100 : node9986;
															assign node9986 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node9990 = (inp[4]) ? 4'b1000 : node9991;
															assign node9991 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node9995 = (inp[1]) ? node10003 : node9996;
													assign node9996 = (inp[0]) ? node9998 : 4'b1000;
														assign node9998 = (inp[2]) ? 4'b1000 : node9999;
															assign node9999 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node10003 = (inp[0]) ? node10017 : node10004;
														assign node10004 = (inp[2]) ? node10010 : node10005;
															assign node10005 = (inp[4]) ? node10007 : 4'b1001;
																assign node10007 = (inp[12]) ? 4'b1100 : 4'b1001;
															assign node10010 = (inp[12]) ? node10014 : node10011;
																assign node10011 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node10014 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node10017 = (inp[12]) ? node10021 : node10018;
															assign node10018 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node10021 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node10024 = (inp[11]) ? node10142 : node10025;
										assign node10025 = (inp[5]) ? node10077 : node10026;
											assign node10026 = (inp[13]) ? node10050 : node10027;
												assign node10027 = (inp[1]) ? node10037 : node10028;
													assign node10028 = (inp[4]) ? node10030 : 4'b1001;
														assign node10030 = (inp[12]) ? node10032 : 4'b1000;
															assign node10032 = (inp[0]) ? node10034 : 4'b1001;
																assign node10034 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10037 = (inp[12]) ? node10041 : node10038;
														assign node10038 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node10041 = (inp[4]) ? node10045 : node10042;
															assign node10042 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node10045 = (inp[0]) ? node10047 : 4'b1100;
																assign node10047 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node10050 = (inp[1]) ? node10056 : node10051;
													assign node10051 = (inp[2]) ? node10053 : 4'b1101;
														assign node10053 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node10056 = (inp[0]) ? node10064 : node10057;
														assign node10057 = (inp[12]) ? 4'b1101 : node10058;
															assign node10058 = (inp[4]) ? node10060 : 4'b1000;
																assign node10060 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node10064 = (inp[2]) ? node10072 : node10065;
															assign node10065 = (inp[4]) ? node10069 : node10066;
																assign node10066 = (inp[12]) ? 4'b1100 : 4'b1001;
																assign node10069 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node10072 = (inp[12]) ? node10074 : 4'b1000;
																assign node10074 = (inp[4]) ? 4'b1000 : 4'b1101;
											assign node10077 = (inp[13]) ? node10109 : node10078;
												assign node10078 = (inp[1]) ? node10094 : node10079;
													assign node10079 = (inp[2]) ? node10089 : node10080;
														assign node10080 = (inp[4]) ? node10084 : node10081;
															assign node10081 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node10084 = (inp[12]) ? node10086 : 4'b1101;
																assign node10086 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node10089 = (inp[12]) ? 4'b1101 : node10090;
															assign node10090 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node10094 = (inp[2]) ? node10100 : node10095;
														assign node10095 = (inp[4]) ? node10097 : 4'b1100;
															assign node10097 = (inp[12]) ? 4'b1001 : 4'b1100;
														assign node10100 = (inp[12]) ? node10104 : node10101;
															assign node10101 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node10104 = (inp[4]) ? 4'b1000 : node10105;
																assign node10105 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node10109 = (inp[1]) ? node10125 : node10110;
													assign node10110 = (inp[2]) ? node10120 : node10111;
														assign node10111 = (inp[0]) ? node10117 : node10112;
															assign node10112 = (inp[4]) ? node10114 : 4'b1000;
																assign node10114 = (inp[12]) ? 4'b1001 : 4'b1000;
															assign node10117 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node10120 = (inp[12]) ? 4'b1000 : node10121;
															assign node10121 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node10125 = (inp[2]) ? node10137 : node10126;
														assign node10126 = (inp[12]) ? node10132 : node10127;
															assign node10127 = (inp[4]) ? node10129 : 4'b1100;
																assign node10129 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node10132 = (inp[4]) ? node10134 : 4'b1001;
																assign node10134 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node10137 = (inp[4]) ? 4'b1000 : node10138;
															assign node10138 = (inp[12]) ? 4'b1000 : 4'b1100;
										assign node10142 = (inp[13]) ? node10196 : node10143;
											assign node10143 = (inp[5]) ? node10175 : node10144;
												assign node10144 = (inp[1]) ? node10158 : node10145;
													assign node10145 = (inp[0]) ? node10151 : node10146;
														assign node10146 = (inp[2]) ? node10148 : 4'b1000;
															assign node10148 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node10151 = (inp[2]) ? node10155 : node10152;
															assign node10152 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node10155 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node10158 = (inp[0]) ? node10168 : node10159;
														assign node10159 = (inp[12]) ? node10163 : node10160;
															assign node10160 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node10163 = (inp[4]) ? 4'b1101 : node10164;
																assign node10164 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node10168 = (inp[4]) ? node10172 : node10169;
															assign node10169 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node10172 = (inp[12]) ? 4'b1100 : 4'b1001;
												assign node10175 = (inp[1]) ? node10183 : node10176;
													assign node10176 = (inp[12]) ? 4'b1100 : node10177;
														assign node10177 = (inp[4]) ? node10179 : 4'b1100;
															assign node10179 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node10183 = (inp[4]) ? node10191 : node10184;
														assign node10184 = (inp[12]) ? node10188 : node10185;
															assign node10185 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node10188 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node10191 = (inp[12]) ? 4'b1000 : node10192;
															assign node10192 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node10196 = (inp[5]) ? node10228 : node10197;
												assign node10197 = (inp[1]) ? node10209 : node10198;
													assign node10198 = (inp[0]) ? 4'b1100 : node10199;
														assign node10199 = (inp[2]) ? node10205 : node10200;
															assign node10200 = (inp[4]) ? node10202 : 4'b1100;
																assign node10202 = (inp[12]) ? 4'b1101 : 4'b1100;
															assign node10205 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node10209 = (inp[0]) ? node10217 : node10210;
														assign node10210 = (inp[12]) ? node10214 : node10211;
															assign node10211 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node10214 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node10217 = (inp[4]) ? node10223 : node10218;
															assign node10218 = (inp[12]) ? node10220 : 4'b1001;
																assign node10220 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node10223 = (inp[12]) ? node10225 : 4'b1100;
																assign node10225 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node10228 = (inp[0]) ? node10232 : node10229;
													assign node10229 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node10232 = (inp[1]) ? node10238 : node10233;
														assign node10233 = (inp[2]) ? node10235 : 4'b1000;
															assign node10235 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node10238 = (inp[12]) ? node10244 : node10239;
															assign node10239 = (inp[4]) ? 4'b1001 : node10240;
																assign node10240 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node10244 = (inp[4]) ? 4'b1100 : 4'b1000;
						assign node10247 = (inp[10]) ? node11183 : node10248;
							assign node10248 = (inp[9]) ? node10760 : node10249;
								assign node10249 = (inp[11]) ? node10491 : node10250;
									assign node10250 = (inp[5]) ? node10366 : node10251;
										assign node10251 = (inp[13]) ? node10315 : node10252;
											assign node10252 = (inp[1]) ? node10284 : node10253;
												assign node10253 = (inp[3]) ? node10271 : node10254;
													assign node10254 = (inp[2]) ? node10262 : node10255;
														assign node10255 = (inp[12]) ? node10257 : 4'b1010;
															assign node10257 = (inp[4]) ? node10259 : 4'b1010;
																assign node10259 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node10262 = (inp[0]) ? node10268 : node10263;
															assign node10263 = (inp[12]) ? 4'b1010 : node10264;
																assign node10264 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node10268 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node10271 = (inp[12]) ? node10279 : node10272;
														assign node10272 = (inp[4]) ? node10274 : 4'b1010;
															assign node10274 = (inp[0]) ? 4'b1111 : node10275;
																assign node10275 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node10279 = (inp[4]) ? 4'b1010 : node10280;
															assign node10280 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node10284 = (inp[12]) ? node10302 : node10285;
													assign node10285 = (inp[3]) ? node10295 : node10286;
														assign node10286 = (inp[4]) ? node10292 : node10287;
															assign node10287 = (inp[0]) ? 4'b1011 : node10288;
																assign node10288 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node10292 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10295 = (inp[4]) ? 4'b1010 : node10296;
															assign node10296 = (inp[2]) ? node10298 : 4'b1110;
																assign node10298 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node10302 = (inp[4]) ? node10312 : node10303;
														assign node10303 = (inp[3]) ? node10309 : node10304;
															assign node10304 = (inp[0]) ? 4'b1110 : node10305;
																assign node10305 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node10309 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node10312 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node10315 = (inp[12]) ? node10341 : node10316;
												assign node10316 = (inp[1]) ? node10324 : node10317;
													assign node10317 = (inp[3]) ? node10319 : 4'b1111;
														assign node10319 = (inp[4]) ? 4'b1010 : node10320;
															assign node10320 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node10324 = (inp[2]) ? node10334 : node10325;
														assign node10325 = (inp[3]) ? node10331 : node10326;
															assign node10326 = (inp[4]) ? 4'b1010 : node10327;
																assign node10327 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node10331 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node10334 = (inp[3]) ? node10338 : node10335;
															assign node10335 = (inp[4]) ? 4'b1011 : 4'b1110;
															assign node10338 = (inp[0]) ? 4'b1111 : 4'b1011;
												assign node10341 = (inp[3]) ? node10357 : node10342;
													assign node10342 = (inp[2]) ? node10352 : node10343;
														assign node10343 = (inp[4]) ? node10347 : node10344;
															assign node10344 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node10347 = (inp[1]) ? 4'b1111 : node10348;
																assign node10348 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node10352 = (inp[4]) ? 4'b1111 : node10353;
															assign node10353 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node10357 = (inp[0]) ? 4'b1111 : node10358;
														assign node10358 = (inp[2]) ? node10362 : node10359;
															assign node10359 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node10362 = (inp[4]) ? 4'b1111 : 4'b1110;
										assign node10366 = (inp[13]) ? node10426 : node10367;
											assign node10367 = (inp[1]) ? node10389 : node10368;
												assign node10368 = (inp[2]) ? node10378 : node10369;
													assign node10369 = (inp[0]) ? 4'b1111 : node10370;
														assign node10370 = (inp[4]) ? node10372 : 4'b1110;
															assign node10372 = (inp[3]) ? node10374 : 4'b1110;
																assign node10374 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node10378 = (inp[12]) ? node10384 : node10379;
														assign node10379 = (inp[3]) ? node10381 : 4'b1110;
															assign node10381 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node10384 = (inp[0]) ? node10386 : 4'b1110;
															assign node10386 = (inp[3]) ? 4'b1110 : 4'b1111;
												assign node10389 = (inp[12]) ? node10411 : node10390;
													assign node10390 = (inp[0]) ? node10404 : node10391;
														assign node10391 = (inp[2]) ? node10397 : node10392;
															assign node10392 = (inp[3]) ? node10394 : 4'b1011;
																assign node10394 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node10397 = (inp[4]) ? node10401 : node10398;
																assign node10398 = (inp[3]) ? 4'b1011 : 4'b1111;
																assign node10401 = (inp[3]) ? 4'b1111 : 4'b1011;
														assign node10404 = (inp[2]) ? 4'b1011 : node10405;
															assign node10405 = (inp[4]) ? 4'b1111 : node10406;
																assign node10406 = (inp[3]) ? 4'b1010 : 4'b1111;
													assign node10411 = (inp[4]) ? node10419 : node10412;
														assign node10412 = (inp[3]) ? node10416 : node10413;
															assign node10413 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node10416 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10419 = (inp[2]) ? 4'b1110 : node10420;
															assign node10420 = (inp[0]) ? node10422 : 4'b1111;
																assign node10422 = (inp[3]) ? 4'b1110 : 4'b1111;
											assign node10426 = (inp[12]) ? node10464 : node10427;
												assign node10427 = (inp[1]) ? node10445 : node10428;
													assign node10428 = (inp[4]) ? node10438 : node10429;
														assign node10429 = (inp[2]) ? 4'b1010 : node10430;
															assign node10430 = (inp[0]) ? node10434 : node10431;
																assign node10431 = (inp[3]) ? 4'b1010 : 4'b1011;
																assign node10434 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node10438 = (inp[3]) ? node10440 : 4'b1010;
															assign node10440 = (inp[0]) ? node10442 : 4'b1110;
																assign node10442 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node10445 = (inp[2]) ? node10455 : node10446;
														assign node10446 = (inp[4]) ? node10450 : node10447;
															assign node10447 = (inp[3]) ? 4'b1110 : 4'b1010;
															assign node10450 = (inp[3]) ? 4'b1011 : node10451;
																assign node10451 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node10455 = (inp[0]) ? node10459 : node10456;
															assign node10456 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node10459 = (inp[3]) ? node10461 : 4'b1110;
																assign node10461 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node10464 = (inp[3]) ? node10482 : node10465;
													assign node10465 = (inp[4]) ? node10473 : node10466;
														assign node10466 = (inp[1]) ? node10468 : 4'b1011;
															assign node10468 = (inp[2]) ? node10470 : 4'b1111;
																assign node10470 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node10473 = (inp[2]) ? node10477 : node10474;
															assign node10474 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node10477 = (inp[0]) ? 4'b1010 : node10478;
																assign node10478 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node10482 = (inp[2]) ? 4'b1010 : node10483;
														assign node10483 = (inp[4]) ? node10487 : node10484;
															assign node10484 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10487 = (inp[0]) ? 4'b1010 : 4'b1011;
									assign node10491 = (inp[5]) ? node10623 : node10492;
										assign node10492 = (inp[13]) ? node10554 : node10493;
											assign node10493 = (inp[1]) ? node10519 : node10494;
												assign node10494 = (inp[0]) ? node10504 : node10495;
													assign node10495 = (inp[4]) ? node10497 : 4'b1011;
														assign node10497 = (inp[3]) ? node10501 : node10498;
															assign node10498 = (inp[12]) ? 4'b1011 : 4'b1010;
															assign node10501 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node10504 = (inp[2]) ? node10514 : node10505;
														assign node10505 = (inp[12]) ? node10509 : node10506;
															assign node10506 = (inp[3]) ? 4'b1110 : 4'b1011;
															assign node10509 = (inp[4]) ? node10511 : 4'b1010;
																assign node10511 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node10514 = (inp[3]) ? 4'b1011 : node10515;
															assign node10515 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node10519 = (inp[12]) ? node10537 : node10520;
													assign node10520 = (inp[4]) ? node10530 : node10521;
														assign node10521 = (inp[3]) ? node10527 : node10522;
															assign node10522 = (inp[0]) ? 4'b1010 : node10523;
																assign node10523 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node10527 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10530 = (inp[3]) ? 4'b1011 : node10531;
															assign node10531 = (inp[2]) ? 4'b1111 : node10532;
																assign node10532 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node10537 = (inp[4]) ? node10547 : node10538;
														assign node10538 = (inp[3]) ? node10544 : node10539;
															assign node10539 = (inp[0]) ? 4'b1111 : node10540;
																assign node10540 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node10544 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10547 = (inp[0]) ? 4'b1011 : node10548;
															assign node10548 = (inp[3]) ? 4'b1011 : node10549;
																assign node10549 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node10554 = (inp[1]) ? node10588 : node10555;
												assign node10555 = (inp[4]) ? node10573 : node10556;
													assign node10556 = (inp[2]) ? node10558 : 4'b1110;
														assign node10558 = (inp[12]) ? node10566 : node10559;
															assign node10559 = (inp[0]) ? node10563 : node10560;
																assign node10560 = (inp[3]) ? 4'b1111 : 4'b1110;
																assign node10563 = (inp[3]) ? 4'b1110 : 4'b1111;
															assign node10566 = (inp[0]) ? node10570 : node10567;
																assign node10567 = (inp[3]) ? 4'b1111 : 4'b1110;
																assign node10570 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node10573 = (inp[12]) ? node10579 : node10574;
														assign node10574 = (inp[3]) ? node10576 : 4'b1110;
															assign node10576 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node10579 = (inp[2]) ? 4'b1110 : node10580;
															assign node10580 = (inp[3]) ? node10584 : node10581;
																assign node10581 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node10584 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node10588 = (inp[12]) ? node10608 : node10589;
													assign node10589 = (inp[2]) ? node10597 : node10590;
														assign node10590 = (inp[4]) ? node10594 : node10591;
															assign node10591 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node10594 = (inp[3]) ? 4'b1111 : 4'b1011;
														assign node10597 = (inp[4]) ? node10601 : node10598;
															assign node10598 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10601 = (inp[3]) ? node10605 : node10602;
																assign node10602 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node10605 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node10608 = (inp[3]) ? node10616 : node10609;
														assign node10609 = (inp[4]) ? 4'b1110 : node10610;
															assign node10610 = (inp[0]) ? node10612 : 4'b1010;
																assign node10612 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node10616 = (inp[0]) ? 4'b1110 : node10617;
															assign node10617 = (inp[4]) ? 4'b1110 : node10618;
																assign node10618 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node10623 = (inp[13]) ? node10695 : node10624;
											assign node10624 = (inp[12]) ? node10662 : node10625;
												assign node10625 = (inp[1]) ? node10639 : node10626;
													assign node10626 = (inp[0]) ? node10632 : node10627;
														assign node10627 = (inp[3]) ? node10629 : 4'b1111;
															assign node10629 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node10632 = (inp[3]) ? node10634 : 4'b1110;
															assign node10634 = (inp[4]) ? 4'b1011 : node10635;
																assign node10635 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node10639 = (inp[2]) ? node10653 : node10640;
														assign node10640 = (inp[0]) ? node10646 : node10641;
															assign node10641 = (inp[3]) ? 4'b1010 : node10642;
																assign node10642 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node10646 = (inp[4]) ? node10650 : node10647;
																assign node10647 = (inp[3]) ? 4'b1011 : 4'b1110;
																assign node10650 = (inp[3]) ? 4'b1110 : 4'b1011;
														assign node10653 = (inp[0]) ? node10659 : node10654;
															assign node10654 = (inp[3]) ? 4'b1110 : node10655;
																assign node10655 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node10659 = (inp[3]) ? 4'b1010 : 4'b1110;
												assign node10662 = (inp[2]) ? node10684 : node10663;
													assign node10663 = (inp[1]) ? node10673 : node10664;
														assign node10664 = (inp[0]) ? node10666 : 4'b1110;
															assign node10666 = (inp[3]) ? node10670 : node10667;
																assign node10667 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node10670 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node10673 = (inp[0]) ? node10679 : node10674;
															assign node10674 = (inp[4]) ? 4'b1111 : node10675;
																assign node10675 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node10679 = (inp[3]) ? 4'b1110 : node10680;
																assign node10680 = (inp[4]) ? 4'b1110 : 4'b1011;
													assign node10684 = (inp[3]) ? 4'b1111 : node10685;
														assign node10685 = (inp[0]) ? node10691 : node10686;
															assign node10686 = (inp[1]) ? node10688 : 4'b1111;
																assign node10688 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node10691 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node10695 = (inp[12]) ? node10729 : node10696;
												assign node10696 = (inp[3]) ? node10712 : node10697;
													assign node10697 = (inp[4]) ? node10707 : node10698;
														assign node10698 = (inp[1]) ? node10702 : node10699;
															assign node10699 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10702 = (inp[0]) ? node10704 : 4'b1011;
																assign node10704 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node10707 = (inp[1]) ? 4'b1111 : node10708;
															assign node10708 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node10712 = (inp[1]) ? node10718 : node10713;
														assign node10713 = (inp[4]) ? 4'b1111 : node10714;
															assign node10714 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10718 = (inp[4]) ? node10724 : node10719;
															assign node10719 = (inp[0]) ? 4'b1111 : node10720;
																assign node10720 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node10724 = (inp[2]) ? node10726 : 4'b1010;
																assign node10726 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node10729 = (inp[2]) ? node10749 : node10730;
													assign node10730 = (inp[4]) ? node10744 : node10731;
														assign node10731 = (inp[1]) ? node10739 : node10732;
															assign node10732 = (inp[3]) ? node10736 : node10733;
																assign node10733 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node10736 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node10739 = (inp[3]) ? node10741 : 4'b1110;
																assign node10741 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10744 = (inp[1]) ? 4'b1011 : node10745;
															assign node10745 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node10749 = (inp[4]) ? node10753 : node10750;
														assign node10750 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node10753 = (inp[0]) ? 4'b1011 : node10754;
															assign node10754 = (inp[1]) ? node10756 : 4'b1011;
																assign node10756 = (inp[3]) ? 4'b1011 : 4'b1010;
								assign node10760 = (inp[11]) ? node10944 : node10761;
									assign node10761 = (inp[13]) ? node10855 : node10762;
										assign node10762 = (inp[5]) ? node10804 : node10763;
											assign node10763 = (inp[12]) ? node10787 : node10764;
												assign node10764 = (inp[3]) ? node10772 : node10765;
													assign node10765 = (inp[4]) ? node10769 : node10766;
														assign node10766 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10769 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node10772 = (inp[1]) ? node10780 : node10773;
														assign node10773 = (inp[0]) ? node10777 : node10774;
															assign node10774 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node10777 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node10780 = (inp[4]) ? 4'b1011 : node10781;
															assign node10781 = (inp[2]) ? node10783 : 4'b1111;
																assign node10783 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node10787 = (inp[3]) ? node10797 : node10788;
													assign node10788 = (inp[1]) ? node10794 : node10789;
														assign node10789 = (inp[2]) ? node10791 : 4'b1011;
															assign node10791 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node10794 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node10797 = (inp[2]) ? 4'b1011 : node10798;
														assign node10798 = (inp[4]) ? 4'b1011 : node10799;
															assign node10799 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node10804 = (inp[1]) ? node10826 : node10805;
												assign node10805 = (inp[0]) ? node10813 : node10806;
													assign node10806 = (inp[3]) ? node10808 : 4'b1111;
														assign node10808 = (inp[4]) ? node10810 : 4'b1111;
															assign node10810 = (inp[12]) ? 4'b1110 : 4'b1011;
													assign node10813 = (inp[4]) ? node10821 : node10814;
														assign node10814 = (inp[3]) ? node10818 : node10815;
															assign node10815 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node10818 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node10821 = (inp[2]) ? node10823 : 4'b1110;
															assign node10823 = (inp[3]) ? 4'b1011 : 4'b1111;
												assign node10826 = (inp[12]) ? node10844 : node10827;
													assign node10827 = (inp[0]) ? node10835 : node10828;
														assign node10828 = (inp[4]) ? node10832 : node10829;
															assign node10829 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node10832 = (inp[3]) ? 4'b1110 : 4'b1010;
														assign node10835 = (inp[4]) ? node10839 : node10836;
															assign node10836 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node10839 = (inp[3]) ? 4'b1111 : node10840;
																assign node10840 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node10844 = (inp[2]) ? 4'b1111 : node10845;
														assign node10845 = (inp[3]) ? node10849 : node10846;
															assign node10846 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node10849 = (inp[4]) ? node10851 : 4'b1110;
																assign node10851 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node10855 = (inp[5]) ? node10905 : node10856;
											assign node10856 = (inp[12]) ? node10886 : node10857;
												assign node10857 = (inp[1]) ? node10875 : node10858;
													assign node10858 = (inp[3]) ? node10868 : node10859;
														assign node10859 = (inp[2]) ? node10861 : 4'b1110;
															assign node10861 = (inp[0]) ? node10865 : node10862;
																assign node10862 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node10865 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node10868 = (inp[4]) ? node10872 : node10869;
															assign node10869 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node10872 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node10875 = (inp[0]) ? node10881 : node10876;
														assign node10876 = (inp[3]) ? 4'b1111 : node10877;
															assign node10877 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node10881 = (inp[4]) ? 4'b1011 : node10882;
															assign node10882 = (inp[3]) ? 4'b1011 : 4'b1111;
												assign node10886 = (inp[4]) ? node10898 : node10887;
													assign node10887 = (inp[2]) ? node10893 : node10888;
														assign node10888 = (inp[1]) ? node10890 : 4'b1110;
															assign node10890 = (inp[0]) ? 4'b1110 : 4'b1010;
														assign node10893 = (inp[0]) ? node10895 : 4'b1111;
															assign node10895 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node10898 = (inp[2]) ? 4'b1110 : node10899;
														assign node10899 = (inp[3]) ? node10901 : 4'b1110;
															assign node10901 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node10905 = (inp[12]) ? node10927 : node10906;
												assign node10906 = (inp[4]) ? node10912 : node10907;
													assign node10907 = (inp[1]) ? node10909 : 4'b1011;
														assign node10909 = (inp[3]) ? 4'b1111 : 4'b1011;
													assign node10912 = (inp[0]) ? node10920 : node10913;
														assign node10913 = (inp[1]) ? node10917 : node10914;
															assign node10914 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node10917 = (inp[3]) ? 4'b1010 : 4'b1111;
														assign node10920 = (inp[1]) ? node10924 : node10921;
															assign node10921 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node10924 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node10927 = (inp[1]) ? node10935 : node10928;
													assign node10928 = (inp[2]) ? 4'b1011 : node10929;
														assign node10929 = (inp[4]) ? node10931 : 4'b1011;
															assign node10931 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node10935 = (inp[4]) ? node10939 : node10936;
														assign node10936 = (inp[3]) ? 4'b1011 : 4'b1110;
														assign node10939 = (inp[0]) ? 4'b1011 : node10940;
															assign node10940 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node10944 = (inp[5]) ? node11060 : node10945;
										assign node10945 = (inp[13]) ? node11007 : node10946;
											assign node10946 = (inp[1]) ? node10972 : node10947;
												assign node10947 = (inp[12]) ? node10961 : node10948;
													assign node10948 = (inp[4]) ? node10952 : node10949;
														assign node10949 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node10952 = (inp[3]) ? node10956 : node10953;
															assign node10953 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node10956 = (inp[2]) ? 4'b1111 : node10957;
																assign node10957 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node10961 = (inp[0]) ? node10963 : 4'b1010;
														assign node10963 = (inp[4]) ? 4'b1010 : node10964;
															assign node10964 = (inp[2]) ? node10968 : node10965;
																assign node10965 = (inp[3]) ? 4'b1011 : 4'b1010;
																assign node10968 = (inp[3]) ? 4'b1010 : 4'b1011;
												assign node10972 = (inp[3]) ? node10992 : node10973;
													assign node10973 = (inp[12]) ? node10985 : node10974;
														assign node10974 = (inp[4]) ? node10980 : node10975;
															assign node10975 = (inp[2]) ? 4'b1011 : node10976;
																assign node10976 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10980 = (inp[0]) ? node10982 : 4'b1110;
																assign node10982 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node10985 = (inp[4]) ? 4'b1010 : node10986;
															assign node10986 = (inp[2]) ? 4'b1110 : node10987;
																assign node10987 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node10992 = (inp[2]) ? node11000 : node10993;
														assign node10993 = (inp[4]) ? node10997 : node10994;
															assign node10994 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node10997 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node11000 = (inp[12]) ? node11004 : node11001;
															assign node11001 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node11004 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node11007 = (inp[12]) ? node11039 : node11008;
												assign node11008 = (inp[1]) ? node11026 : node11009;
													assign node11009 = (inp[4]) ? node11019 : node11010;
														assign node11010 = (inp[2]) ? node11012 : 4'b1111;
															assign node11012 = (inp[3]) ? node11016 : node11013;
																assign node11013 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node11016 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11019 = (inp[3]) ? node11021 : 4'b1111;
															assign node11021 = (inp[2]) ? 4'b1011 : node11022;
																assign node11022 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node11026 = (inp[0]) ? node11030 : node11027;
														assign node11027 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11030 = (inp[3]) ? node11034 : node11031;
															assign node11031 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node11034 = (inp[2]) ? 4'b1111 : node11035;
																assign node11035 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node11039 = (inp[3]) ? node11051 : node11040;
													assign node11040 = (inp[0]) ? node11042 : 4'b1111;
														assign node11042 = (inp[1]) ? 4'b1111 : node11043;
															assign node11043 = (inp[2]) ? node11047 : node11044;
																assign node11044 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node11047 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node11051 = (inp[0]) ? 4'b1111 : node11052;
														assign node11052 = (inp[4]) ? node11056 : node11053;
															assign node11053 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node11056 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node11060 = (inp[13]) ? node11126 : node11061;
											assign node11061 = (inp[12]) ? node11097 : node11062;
												assign node11062 = (inp[4]) ? node11082 : node11063;
													assign node11063 = (inp[3]) ? node11075 : node11064;
														assign node11064 = (inp[2]) ? node11070 : node11065;
															assign node11065 = (inp[1]) ? node11067 : 4'b1110;
																assign node11067 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11070 = (inp[1]) ? 4'b1111 : node11071;
																assign node11071 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11075 = (inp[1]) ? node11079 : node11076;
															assign node11076 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node11079 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node11082 = (inp[2]) ? node11090 : node11083;
														assign node11083 = (inp[0]) ? node11085 : 4'b1011;
															assign node11085 = (inp[1]) ? node11087 : 4'b1111;
																assign node11087 = (inp[3]) ? 4'b1111 : 4'b1010;
														assign node11090 = (inp[1]) ? node11094 : node11091;
															assign node11091 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node11094 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node11097 = (inp[0]) ? node11109 : node11098;
													assign node11098 = (inp[4]) ? node11104 : node11099;
														assign node11099 = (inp[3]) ? 4'b1110 : node11100;
															assign node11100 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node11104 = (inp[2]) ? 4'b1110 : node11105;
															assign node11105 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node11109 = (inp[3]) ? node11121 : node11110;
														assign node11110 = (inp[1]) ? node11116 : node11111;
															assign node11111 = (inp[2]) ? 4'b1111 : node11112;
																assign node11112 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node11116 = (inp[4]) ? node11118 : 4'b1011;
																assign node11118 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11121 = (inp[4]) ? 4'b1110 : node11122;
															assign node11122 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node11126 = (inp[1]) ? node11154 : node11127;
												assign node11127 = (inp[12]) ? node11145 : node11128;
													assign node11128 = (inp[4]) ? node11136 : node11129;
														assign node11129 = (inp[2]) ? 4'b1010 : node11130;
															assign node11130 = (inp[3]) ? node11132 : 4'b1010;
																assign node11132 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11136 = (inp[3]) ? node11142 : node11137;
															assign node11137 = (inp[2]) ? node11139 : 4'b1010;
																assign node11139 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node11142 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node11145 = (inp[2]) ? 4'b1010 : node11146;
														assign node11146 = (inp[3]) ? node11148 : 4'b1010;
															assign node11148 = (inp[4]) ? 4'b1010 : node11149;
																assign node11149 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node11154 = (inp[12]) ? node11168 : node11155;
													assign node11155 = (inp[3]) ? node11163 : node11156;
														assign node11156 = (inp[4]) ? node11158 : 4'b1010;
															assign node11158 = (inp[0]) ? node11160 : 4'b1110;
																assign node11160 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11163 = (inp[2]) ? node11165 : 4'b1110;
															assign node11165 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node11168 = (inp[3]) ? node11176 : node11169;
														assign node11169 = (inp[4]) ? node11171 : 4'b1111;
															assign node11171 = (inp[2]) ? node11173 : 4'b1010;
																assign node11173 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node11176 = (inp[2]) ? 4'b1010 : node11177;
															assign node11177 = (inp[0]) ? 4'b1010 : node11178;
																assign node11178 = (inp[4]) ? 4'b1011 : 4'b1010;
							assign node11183 = (inp[4]) ? node11647 : node11184;
								assign node11184 = (inp[13]) ? node11392 : node11185;
									assign node11185 = (inp[5]) ? node11295 : node11186;
										assign node11186 = (inp[1]) ? node11242 : node11187;
											assign node11187 = (inp[0]) ? node11203 : node11188;
												assign node11188 = (inp[2]) ? node11196 : node11189;
													assign node11189 = (inp[9]) ? node11193 : node11190;
														assign node11190 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11193 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11196 = (inp[11]) ? node11200 : node11197;
														assign node11197 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node11200 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node11203 = (inp[12]) ? node11231 : node11204;
													assign node11204 = (inp[11]) ? node11218 : node11205;
														assign node11205 = (inp[9]) ? node11213 : node11206;
															assign node11206 = (inp[2]) ? node11210 : node11207;
																assign node11207 = (inp[3]) ? 4'b1011 : 4'b1010;
																assign node11210 = (inp[3]) ? 4'b1010 : 4'b1011;
															assign node11213 = (inp[3]) ? node11215 : 4'b1010;
																assign node11215 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node11218 = (inp[2]) ? node11226 : node11219;
															assign node11219 = (inp[3]) ? node11223 : node11220;
																assign node11220 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node11223 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11226 = (inp[9]) ? node11228 : 4'b1010;
																assign node11228 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node11231 = (inp[2]) ? 4'b1010 : node11232;
														assign node11232 = (inp[11]) ? 4'b1010 : node11233;
															assign node11233 = (inp[3]) ? node11237 : node11234;
																assign node11234 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node11237 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node11242 = (inp[11]) ? node11268 : node11243;
												assign node11243 = (inp[9]) ? node11259 : node11244;
													assign node11244 = (inp[3]) ? node11256 : node11245;
														assign node11245 = (inp[12]) ? node11251 : node11246;
															assign node11246 = (inp[2]) ? 4'b1011 : node11247;
																assign node11247 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11251 = (inp[2]) ? 4'b1110 : node11252;
																assign node11252 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node11256 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node11259 = (inp[0]) ? node11261 : 4'b1011;
														assign node11261 = (inp[12]) ? node11263 : 4'b1010;
															assign node11263 = (inp[3]) ? node11265 : 4'b1111;
																assign node11265 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node11268 = (inp[9]) ? node11284 : node11269;
													assign node11269 = (inp[12]) ? node11275 : node11270;
														assign node11270 = (inp[3]) ? node11272 : 4'b1010;
															assign node11272 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11275 = (inp[3]) ? node11279 : node11276;
															assign node11276 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node11279 = (inp[0]) ? node11281 : 4'b1011;
																assign node11281 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node11284 = (inp[12]) ? node11290 : node11285;
														assign node11285 = (inp[3]) ? node11287 : 4'b1011;
															assign node11287 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node11290 = (inp[3]) ? node11292 : 4'b1110;
															assign node11292 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node11295 = (inp[1]) ? node11335 : node11296;
											assign node11296 = (inp[3]) ? node11318 : node11297;
												assign node11297 = (inp[9]) ? node11307 : node11298;
													assign node11298 = (inp[11]) ? node11304 : node11299;
														assign node11299 = (inp[2]) ? node11301 : 4'b1110;
															assign node11301 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11304 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node11307 = (inp[11]) ? node11313 : node11308;
														assign node11308 = (inp[2]) ? node11310 : 4'b1111;
															assign node11310 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node11313 = (inp[0]) ? node11315 : 4'b1110;
															assign node11315 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node11318 = (inp[0]) ? node11326 : node11319;
													assign node11319 = (inp[9]) ? node11323 : node11320;
														assign node11320 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11323 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node11326 = (inp[9]) ? 4'b1111 : node11327;
														assign node11327 = (inp[11]) ? node11331 : node11328;
															assign node11328 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node11331 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node11335 = (inp[11]) ? node11363 : node11336;
												assign node11336 = (inp[9]) ? node11352 : node11337;
													assign node11337 = (inp[2]) ? node11347 : node11338;
														assign node11338 = (inp[3]) ? node11342 : node11339;
															assign node11339 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node11342 = (inp[12]) ? 4'b1111 : node11343;
																assign node11343 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node11347 = (inp[12]) ? 4'b1110 : node11348;
															assign node11348 = (inp[3]) ? 4'b1011 : 4'b1111;
													assign node11352 = (inp[12]) ? node11356 : node11353;
														assign node11353 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11356 = (inp[3]) ? 4'b1111 : node11357;
															assign node11357 = (inp[2]) ? node11359 : 4'b1011;
																assign node11359 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node11363 = (inp[0]) ? node11377 : node11364;
													assign node11364 = (inp[9]) ? node11370 : node11365;
														assign node11365 = (inp[12]) ? 4'b1011 : node11366;
															assign node11366 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node11370 = (inp[12]) ? node11374 : node11371;
															assign node11371 = (inp[3]) ? 4'b1011 : 4'b1110;
															assign node11374 = (inp[3]) ? 4'b1110 : 4'b1010;
													assign node11377 = (inp[9]) ? node11385 : node11378;
														assign node11378 = (inp[12]) ? node11382 : node11379;
															assign node11379 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node11382 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node11385 = (inp[12]) ? node11389 : node11386;
															assign node11386 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node11389 = (inp[2]) ? 4'b1110 : 4'b1111;
									assign node11392 = (inp[5]) ? node11500 : node11393;
										assign node11393 = (inp[1]) ? node11435 : node11394;
											assign node11394 = (inp[9]) ? node11416 : node11395;
												assign node11395 = (inp[11]) ? node11409 : node11396;
													assign node11396 = (inp[2]) ? node11398 : 4'b1111;
														assign node11398 = (inp[12]) ? node11404 : node11399;
															assign node11399 = (inp[0]) ? node11401 : 4'b1111;
																assign node11401 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node11404 = (inp[3]) ? node11406 : 4'b1111;
																assign node11406 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node11409 = (inp[2]) ? node11411 : 4'b1110;
														assign node11411 = (inp[0]) ? node11413 : 4'b1111;
															assign node11413 = (inp[3]) ? 4'b1110 : 4'b1111;
												assign node11416 = (inp[11]) ? node11428 : node11417;
													assign node11417 = (inp[2]) ? node11419 : 4'b1110;
														assign node11419 = (inp[12]) ? node11423 : node11420;
															assign node11420 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node11423 = (inp[0]) ? node11425 : 4'b1110;
																assign node11425 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node11428 = (inp[2]) ? node11430 : 4'b1111;
														assign node11430 = (inp[0]) ? 4'b1111 : node11431;
															assign node11431 = (inp[3]) ? 4'b1110 : 4'b1111;
											assign node11435 = (inp[3]) ? node11465 : node11436;
												assign node11436 = (inp[12]) ? node11452 : node11437;
													assign node11437 = (inp[11]) ? node11445 : node11438;
														assign node11438 = (inp[9]) ? node11440 : 4'b1110;
															assign node11440 = (inp[2]) ? 4'b1111 : node11441;
																assign node11441 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11445 = (inp[9]) ? 4'b1110 : node11446;
															assign node11446 = (inp[0]) ? 4'b1111 : node11447;
																assign node11447 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node11452 = (inp[2]) ? node11460 : node11453;
														assign node11453 = (inp[9]) ? node11457 : node11454;
															assign node11454 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11457 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11460 = (inp[9]) ? node11462 : 4'b1010;
															assign node11462 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node11465 = (inp[12]) ? node11485 : node11466;
													assign node11466 = (inp[2]) ? node11474 : node11467;
														assign node11467 = (inp[9]) ? node11471 : node11468;
															assign node11468 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11471 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11474 = (inp[9]) ? node11480 : node11475;
															assign node11475 = (inp[0]) ? 4'b1010 : node11476;
																assign node11476 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11480 = (inp[11]) ? 4'b1011 : node11481;
																assign node11481 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node11485 = (inp[9]) ? node11491 : node11486;
														assign node11486 = (inp[11]) ? node11488 : 4'b1111;
															assign node11488 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node11491 = (inp[11]) ? node11497 : node11492;
															assign node11492 = (inp[0]) ? 4'b1110 : node11493;
																assign node11493 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node11497 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node11500 = (inp[1]) ? node11584 : node11501;
											assign node11501 = (inp[0]) ? node11543 : node11502;
												assign node11502 = (inp[2]) ? node11530 : node11503;
													assign node11503 = (inp[11]) ? node11517 : node11504;
														assign node11504 = (inp[12]) ? node11512 : node11505;
															assign node11505 = (inp[3]) ? node11509 : node11506;
																assign node11506 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node11509 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11512 = (inp[9]) ? node11514 : 4'b1010;
																assign node11514 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node11517 = (inp[12]) ? node11523 : node11518;
															assign node11518 = (inp[9]) ? node11520 : 4'b1011;
																assign node11520 = (inp[3]) ? 4'b1010 : 4'b1011;
															assign node11523 = (inp[9]) ? node11527 : node11524;
																assign node11524 = (inp[3]) ? 4'b1011 : 4'b1010;
																assign node11527 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node11530 = (inp[3]) ? node11538 : node11531;
														assign node11531 = (inp[12]) ? 4'b1011 : node11532;
															assign node11532 = (inp[9]) ? node11534 : 4'b1010;
																assign node11534 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11538 = (inp[9]) ? node11540 : 4'b1011;
															assign node11540 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11543 = (inp[2]) ? node11565 : node11544;
													assign node11544 = (inp[9]) ? node11550 : node11545;
														assign node11545 = (inp[11]) ? node11547 : 4'b1011;
															assign node11547 = (inp[3]) ? 4'b1010 : 4'b1011;
														assign node11550 = (inp[12]) ? node11558 : node11551;
															assign node11551 = (inp[3]) ? node11555 : node11552;
																assign node11552 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node11555 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11558 = (inp[3]) ? node11562 : node11559;
																assign node11559 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node11562 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11565 = (inp[3]) ? node11577 : node11566;
														assign node11566 = (inp[12]) ? node11572 : node11567;
															assign node11567 = (inp[9]) ? 4'b1010 : node11568;
																assign node11568 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11572 = (inp[9]) ? node11574 : 4'b1010;
																assign node11574 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11577 = (inp[11]) ? node11581 : node11578;
															assign node11578 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node11581 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node11584 = (inp[11]) ? node11616 : node11585;
												assign node11585 = (inp[9]) ? node11599 : node11586;
													assign node11586 = (inp[0]) ? node11588 : 4'b1010;
														assign node11588 = (inp[12]) ? node11594 : node11589;
															assign node11589 = (inp[3]) ? 4'b1110 : node11590;
																assign node11590 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node11594 = (inp[3]) ? 4'b1011 : node11595;
																assign node11595 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node11599 = (inp[12]) ? node11611 : node11600;
														assign node11600 = (inp[3]) ? node11606 : node11601;
															assign node11601 = (inp[0]) ? node11603 : 4'b1011;
																assign node11603 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node11606 = (inp[0]) ? 4'b1111 : node11607;
																assign node11607 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11611 = (inp[3]) ? node11613 : 4'b1110;
															assign node11613 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node11616 = (inp[9]) ? node11634 : node11617;
													assign node11617 = (inp[12]) ? node11625 : node11618;
														assign node11618 = (inp[3]) ? 4'b1111 : node11619;
															assign node11619 = (inp[0]) ? node11621 : 4'b1011;
																assign node11621 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node11625 = (inp[3]) ? node11631 : node11626;
															assign node11626 = (inp[2]) ? node11628 : 4'b1110;
																assign node11628 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node11631 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node11634 = (inp[12]) ? node11640 : node11635;
														assign node11635 = (inp[3]) ? node11637 : 4'b1010;
															assign node11637 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node11640 = (inp[3]) ? node11642 : 4'b1111;
															assign node11642 = (inp[0]) ? node11644 : 4'b1010;
																assign node11644 = (inp[2]) ? 4'b1010 : 4'b1011;
								assign node11647 = (inp[12]) ? node11915 : node11648;
									assign node11648 = (inp[11]) ? node11786 : node11649;
										assign node11649 = (inp[1]) ? node11713 : node11650;
											assign node11650 = (inp[5]) ? node11684 : node11651;
												assign node11651 = (inp[9]) ? node11661 : node11652;
													assign node11652 = (inp[3]) ? node11658 : node11653;
														assign node11653 = (inp[13]) ? node11655 : 4'b1010;
															assign node11655 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node11658 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node11661 = (inp[13]) ? node11673 : node11662;
														assign node11662 = (inp[3]) ? node11668 : node11663;
															assign node11663 = (inp[0]) ? 4'b1011 : node11664;
																assign node11664 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node11668 = (inp[0]) ? 4'b1110 : node11669;
																assign node11669 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11673 = (inp[3]) ? node11679 : node11674;
															assign node11674 = (inp[2]) ? node11676 : 4'b1110;
																assign node11676 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node11679 = (inp[0]) ? 4'b1010 : node11680;
																assign node11680 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node11684 = (inp[9]) ? node11694 : node11685;
													assign node11685 = (inp[3]) ? node11691 : node11686;
														assign node11686 = (inp[13]) ? node11688 : 4'b1110;
															assign node11688 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node11691 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node11694 = (inp[2]) ? node11704 : node11695;
														assign node11695 = (inp[13]) ? node11701 : node11696;
															assign node11696 = (inp[3]) ? node11698 : 4'b1110;
																assign node11698 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11701 = (inp[3]) ? 4'b1111 : 4'b1011;
														assign node11704 = (inp[3]) ? node11710 : node11705;
															assign node11705 = (inp[13]) ? node11707 : 4'b1111;
																assign node11707 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11710 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node11713 = (inp[2]) ? node11755 : node11714;
												assign node11714 = (inp[13]) ? node11734 : node11715;
													assign node11715 = (inp[9]) ? node11723 : node11716;
														assign node11716 = (inp[0]) ? 4'b1010 : node11717;
															assign node11717 = (inp[5]) ? node11719 : 4'b1011;
																assign node11719 = (inp[3]) ? 4'b1111 : 4'b1011;
														assign node11723 = (inp[5]) ? node11731 : node11724;
															assign node11724 = (inp[3]) ? node11728 : node11725;
																assign node11725 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node11728 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11731 = (inp[0]) ? 4'b1110 : 4'b1010;
													assign node11734 = (inp[0]) ? node11744 : node11735;
														assign node11735 = (inp[9]) ? node11741 : node11736;
															assign node11736 = (inp[3]) ? 4'b1110 : node11737;
																assign node11737 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node11741 = (inp[5]) ? 4'b1010 : 4'b1111;
														assign node11744 = (inp[9]) ? node11752 : node11745;
															assign node11745 = (inp[5]) ? node11749 : node11746;
																assign node11746 = (inp[3]) ? 4'b1110 : 4'b1010;
																assign node11749 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node11752 = (inp[3]) ? 4'b1010 : 4'b1011;
												assign node11755 = (inp[5]) ? node11771 : node11756;
													assign node11756 = (inp[9]) ? node11762 : node11757;
														assign node11757 = (inp[3]) ? 4'b1010 : node11758;
															assign node11758 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node11762 = (inp[13]) ? node11766 : node11763;
															assign node11763 = (inp[0]) ? 4'b1111 : 4'b1011;
															assign node11766 = (inp[3]) ? 4'b1111 : node11767;
																assign node11767 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node11771 = (inp[9]) ? node11779 : node11772;
														assign node11772 = (inp[13]) ? node11776 : node11773;
															assign node11773 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node11776 = (inp[3]) ? 4'b1011 : 4'b1110;
														assign node11779 = (inp[13]) ? node11781 : 4'b1010;
															assign node11781 = (inp[3]) ? node11783 : 4'b1111;
																assign node11783 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node11786 = (inp[13]) ? node11854 : node11787;
											assign node11787 = (inp[2]) ? node11825 : node11788;
												assign node11788 = (inp[0]) ? node11806 : node11789;
													assign node11789 = (inp[9]) ? node11799 : node11790;
														assign node11790 = (inp[1]) ? node11794 : node11791;
															assign node11791 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node11794 = (inp[5]) ? node11796 : 4'b1010;
																assign node11796 = (inp[3]) ? 4'b1110 : 4'b1010;
														assign node11799 = (inp[1]) ? 4'b1011 : node11800;
															assign node11800 = (inp[3]) ? 4'b1011 : node11801;
																assign node11801 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node11806 = (inp[1]) ? node11818 : node11807;
														assign node11807 = (inp[5]) ? node11811 : node11808;
															assign node11808 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node11811 = (inp[3]) ? node11815 : node11812;
																assign node11812 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node11815 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11818 = (inp[9]) ? 4'b1111 : node11819;
															assign node11819 = (inp[3]) ? 4'b1110 : node11820;
																assign node11820 = (inp[5]) ? 4'b1011 : 4'b1110;
												assign node11825 = (inp[9]) ? node11841 : node11826;
													assign node11826 = (inp[3]) ? node11834 : node11827;
														assign node11827 = (inp[5]) ? 4'b1010 : node11828;
															assign node11828 = (inp[1]) ? 4'b1111 : node11829;
																assign node11829 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node11834 = (inp[5]) ? node11836 : 4'b1110;
															assign node11836 = (inp[1]) ? node11838 : 4'b1011;
																assign node11838 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node11841 = (inp[3]) ? node11847 : node11842;
														assign node11842 = (inp[1]) ? 4'b1110 : node11843;
															assign node11843 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node11847 = (inp[1]) ? node11851 : node11848;
															assign node11848 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node11851 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node11854 = (inp[9]) ? node11892 : node11855;
												assign node11855 = (inp[1]) ? node11875 : node11856;
													assign node11856 = (inp[5]) ? node11866 : node11857;
														assign node11857 = (inp[3]) ? node11863 : node11858;
															assign node11858 = (inp[0]) ? 4'b1110 : node11859;
																assign node11859 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node11863 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node11866 = (inp[3]) ? node11870 : node11867;
															assign node11867 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node11870 = (inp[2]) ? node11872 : 4'b1111;
																assign node11872 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node11875 = (inp[0]) ? node11883 : node11876;
														assign node11876 = (inp[5]) ? 4'b1111 : node11877;
															assign node11877 = (inp[3]) ? 4'b1111 : node11878;
																assign node11878 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node11883 = (inp[5]) ? node11887 : node11884;
															assign node11884 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node11887 = (inp[3]) ? node11889 : 4'b1110;
																assign node11889 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node11892 = (inp[1]) ? node11908 : node11893;
													assign node11893 = (inp[0]) ? node11903 : node11894;
														assign node11894 = (inp[3]) ? node11900 : node11895;
															assign node11895 = (inp[5]) ? 4'b1011 : node11896;
																assign node11896 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node11900 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node11903 = (inp[5]) ? 4'b1010 : node11904;
															assign node11904 = (inp[3]) ? 4'b1011 : 4'b1111;
													assign node11908 = (inp[5]) ? 4'b1110 : node11909;
														assign node11909 = (inp[3]) ? 4'b1110 : node11910;
															assign node11910 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node11915 = (inp[0]) ? node12049 : node11916;
										assign node11916 = (inp[2]) ? node11990 : node11917;
											assign node11917 = (inp[3]) ? node11955 : node11918;
												assign node11918 = (inp[1]) ? node11926 : node11919;
													assign node11919 = (inp[13]) ? node11923 : node11920;
														assign node11920 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node11923 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11926 = (inp[9]) ? node11942 : node11927;
														assign node11927 = (inp[11]) ? node11935 : node11928;
															assign node11928 = (inp[13]) ? node11932 : node11929;
																assign node11929 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node11932 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node11935 = (inp[13]) ? node11939 : node11936;
																assign node11936 = (inp[5]) ? 4'b1111 : 4'b1011;
																assign node11939 = (inp[5]) ? 4'b1011 : 4'b1110;
														assign node11942 = (inp[11]) ? node11948 : node11943;
															assign node11943 = (inp[5]) ? node11945 : 4'b1011;
																assign node11945 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node11948 = (inp[13]) ? node11952 : node11949;
																assign node11949 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node11952 = (inp[5]) ? 4'b1010 : 4'b1111;
												assign node11955 = (inp[9]) ? node11971 : node11956;
													assign node11956 = (inp[13]) ? node11964 : node11957;
														assign node11957 = (inp[5]) ? node11961 : node11958;
															assign node11958 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11961 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node11964 = (inp[5]) ? node11968 : node11965;
															assign node11965 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11968 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11971 = (inp[1]) ? node11981 : node11972;
														assign node11972 = (inp[5]) ? node11976 : node11973;
															assign node11973 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node11976 = (inp[11]) ? node11978 : 4'b1110;
																assign node11978 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node11981 = (inp[5]) ? node11987 : node11982;
															assign node11982 = (inp[13]) ? 4'b1110 : node11983;
																assign node11983 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11987 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node11990 = (inp[11]) ? node12022 : node11991;
												assign node11991 = (inp[9]) ? node12009 : node11992;
													assign node11992 = (inp[13]) ? node12000 : node11993;
														assign node11993 = (inp[5]) ? 4'b1110 : node11994;
															assign node11994 = (inp[1]) ? node11996 : 4'b1010;
																assign node11996 = (inp[3]) ? 4'b1010 : 4'b1011;
														assign node12000 = (inp[5]) ? node12006 : node12001;
															assign node12001 = (inp[3]) ? 4'b1111 : node12002;
																assign node12002 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node12006 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node12009 = (inp[13]) ? node12017 : node12010;
														assign node12010 = (inp[5]) ? 4'b1111 : node12011;
															assign node12011 = (inp[1]) ? node12013 : 4'b1011;
																assign node12013 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node12017 = (inp[5]) ? 4'b1010 : node12018;
															assign node12018 = (inp[3]) ? 4'b1110 : 4'b1111;
												assign node12022 = (inp[9]) ? node12034 : node12023;
													assign node12023 = (inp[13]) ? node12029 : node12024;
														assign node12024 = (inp[5]) ? 4'b1111 : node12025;
															assign node12025 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node12029 = (inp[5]) ? node12031 : 4'b1110;
															assign node12031 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node12034 = (inp[13]) ? node12038 : node12035;
														assign node12035 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node12038 = (inp[5]) ? node12044 : node12039;
															assign node12039 = (inp[1]) ? node12041 : 4'b1111;
																assign node12041 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node12044 = (inp[3]) ? 4'b1010 : node12045;
																assign node12045 = (inp[1]) ? 4'b1011 : 4'b1010;
										assign node12049 = (inp[1]) ? node12135 : node12050;
											assign node12050 = (inp[5]) ? node12100 : node12051;
												assign node12051 = (inp[13]) ? node12079 : node12052;
													assign node12052 = (inp[2]) ? node12066 : node12053;
														assign node12053 = (inp[3]) ? node12061 : node12054;
															assign node12054 = (inp[11]) ? node12058 : node12055;
																assign node12055 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node12058 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node12061 = (inp[9]) ? node12063 : 4'b1011;
																assign node12063 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12066 = (inp[9]) ? node12072 : node12067;
															assign node12067 = (inp[3]) ? 4'b1010 : node12068;
																assign node12068 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node12072 = (inp[11]) ? node12076 : node12073;
																assign node12073 = (inp[3]) ? 4'b1010 : 4'b1011;
																assign node12076 = (inp[3]) ? 4'b1011 : 4'b1010;
													assign node12079 = (inp[11]) ? node12091 : node12080;
														assign node12080 = (inp[9]) ? node12086 : node12081;
															assign node12081 = (inp[2]) ? 4'b1111 : node12082;
																assign node12082 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node12086 = (inp[2]) ? 4'b1110 : node12087;
																assign node12087 = (inp[3]) ? 4'b1110 : 4'b1111;
														assign node12091 = (inp[9]) ? node12095 : node12092;
															assign node12092 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node12095 = (inp[3]) ? 4'b1111 : node12096;
																assign node12096 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node12100 = (inp[13]) ? node12122 : node12101;
													assign node12101 = (inp[9]) ? node12115 : node12102;
														assign node12102 = (inp[2]) ? node12108 : node12103;
															assign node12103 = (inp[11]) ? node12105 : 4'b1111;
																assign node12105 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node12108 = (inp[11]) ? node12112 : node12109;
																assign node12109 = (inp[3]) ? 4'b1110 : 4'b1111;
																assign node12112 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node12115 = (inp[11]) ? node12119 : node12116;
															assign node12116 = (inp[3]) ? 4'b1111 : 4'b1110;
															assign node12119 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node12122 = (inp[11]) ? node12132 : node12123;
														assign node12123 = (inp[2]) ? node12129 : node12124;
															assign node12124 = (inp[9]) ? node12126 : 4'b1011;
																assign node12126 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node12129 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node12132 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node12135 = (inp[2]) ? node12155 : node12136;
												assign node12136 = (inp[13]) ? node12150 : node12137;
													assign node12137 = (inp[5]) ? node12139 : 4'b1011;
														assign node12139 = (inp[11]) ? node12145 : node12140;
															assign node12140 = (inp[3]) ? 4'b1110 : node12141;
																assign node12141 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12145 = (inp[9]) ? node12147 : 4'b1111;
																assign node12147 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node12150 = (inp[5]) ? node12152 : 4'b1110;
														assign node12152 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node12155 = (inp[9]) ? node12171 : node12156;
													assign node12156 = (inp[11]) ? node12164 : node12157;
														assign node12157 = (inp[5]) ? node12161 : node12158;
															assign node12158 = (inp[13]) ? 4'b1111 : 4'b1010;
															assign node12161 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node12164 = (inp[5]) ? 4'b1011 : node12165;
															assign node12165 = (inp[3]) ? node12167 : 4'b1011;
																assign node12167 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node12171 = (inp[11]) ? node12177 : node12172;
														assign node12172 = (inp[13]) ? 4'b1110 : node12173;
															assign node12173 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node12177 = (inp[5]) ? node12183 : node12178;
															assign node12178 = (inp[13]) ? 4'b1111 : node12179;
																assign node12179 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node12183 = (inp[13]) ? 4'b1010 : 4'b1110;
					assign node12186 = (inp[15]) ? node13804 : node12187;
						assign node12187 = (inp[2]) ? node13011 : node12188;
							assign node12188 = (inp[1]) ? node12604 : node12189;
								assign node12189 = (inp[9]) ? node12389 : node12190;
									assign node12190 = (inp[11]) ? node12274 : node12191;
										assign node12191 = (inp[12]) ? node12229 : node12192;
											assign node12192 = (inp[5]) ? node12208 : node12193;
												assign node12193 = (inp[13]) ? node12203 : node12194;
													assign node12194 = (inp[3]) ? node12196 : 4'b1010;
														assign node12196 = (inp[4]) ? node12200 : node12197;
															assign node12197 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12200 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node12203 = (inp[3]) ? node12205 : 4'b1110;
														assign node12205 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node12208 = (inp[13]) ? node12222 : node12209;
													assign node12209 = (inp[3]) ? node12215 : node12210;
														assign node12210 = (inp[0]) ? node12212 : 4'b1111;
															assign node12212 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node12215 = (inp[4]) ? node12219 : node12216;
															assign node12216 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12219 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12222 = (inp[4]) ? node12226 : node12223;
														assign node12223 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node12226 = (inp[3]) ? 4'b1110 : 4'b1010;
											assign node12229 = (inp[4]) ? node12257 : node12230;
												assign node12230 = (inp[0]) ? node12244 : node12231;
													assign node12231 = (inp[13]) ? node12237 : node12232;
														assign node12232 = (inp[3]) ? 4'b1010 : node12233;
															assign node12233 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node12237 = (inp[5]) ? node12241 : node12238;
															assign node12238 = (inp[3]) ? 4'b1011 : 4'b1110;
															assign node12241 = (inp[3]) ? 4'b1110 : 4'b1010;
													assign node12244 = (inp[5]) ? node12252 : node12245;
														assign node12245 = (inp[13]) ? node12249 : node12246;
															assign node12246 = (inp[3]) ? 4'b1110 : 4'b1011;
															assign node12249 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node12252 = (inp[13]) ? node12254 : 4'b1011;
															assign node12254 = (inp[3]) ? 4'b1110 : 4'b1010;
												assign node12257 = (inp[13]) ? node12267 : node12258;
													assign node12258 = (inp[5]) ? node12264 : node12259;
														assign node12259 = (inp[3]) ? node12261 : 4'b1110;
															assign node12261 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12264 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12267 = (inp[5]) ? node12271 : node12268;
														assign node12268 = (inp[3]) ? 4'b1111 : 4'b1011;
														assign node12271 = (inp[3]) ? 4'b1011 : 4'b1111;
										assign node12274 = (inp[12]) ? node12332 : node12275;
											assign node12275 = (inp[3]) ? node12293 : node12276;
												assign node12276 = (inp[0]) ? node12284 : node12277;
													assign node12277 = (inp[5]) ? node12281 : node12278;
														assign node12278 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node12281 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node12284 = (inp[5]) ? node12288 : node12285;
														assign node12285 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node12288 = (inp[13]) ? 4'b1011 : node12289;
															assign node12289 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node12293 = (inp[4]) ? node12319 : node12294;
													assign node12294 = (inp[10]) ? node12306 : node12295;
														assign node12295 = (inp[0]) ? node12299 : node12296;
															assign node12296 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node12299 = (inp[5]) ? node12303 : node12300;
																assign node12300 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node12303 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node12306 = (inp[13]) ? node12314 : node12307;
															assign node12307 = (inp[5]) ? node12311 : node12308;
																assign node12308 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node12311 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12314 = (inp[5]) ? node12316 : 4'b1111;
																assign node12316 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12319 = (inp[0]) ? node12327 : node12320;
														assign node12320 = (inp[5]) ? node12324 : node12321;
															assign node12321 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node12324 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node12327 = (inp[13]) ? node12329 : 4'b1010;
															assign node12329 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node12332 = (inp[4]) ? node12360 : node12333;
												assign node12333 = (inp[0]) ? node12347 : node12334;
													assign node12334 = (inp[3]) ? node12340 : node12335;
														assign node12335 = (inp[13]) ? node12337 : 4'b1011;
															assign node12337 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node12340 = (inp[5]) ? node12344 : node12341;
															assign node12341 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node12344 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node12347 = (inp[5]) ? node12353 : node12348;
														assign node12348 = (inp[13]) ? node12350 : 4'b1111;
															assign node12350 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node12353 = (inp[10]) ? node12355 : 4'b1111;
															assign node12355 = (inp[3]) ? 4'b1010 : node12356;
																assign node12356 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node12360 = (inp[13]) ? node12374 : node12361;
													assign node12361 = (inp[5]) ? node12369 : node12362;
														assign node12362 = (inp[3]) ? node12366 : node12363;
															assign node12363 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12366 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12369 = (inp[3]) ? 4'b1111 : node12370;
															assign node12370 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node12374 = (inp[10]) ? node12382 : node12375;
														assign node12375 = (inp[5]) ? node12379 : node12376;
															assign node12376 = (inp[3]) ? 4'b1110 : 4'b1010;
															assign node12379 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node12382 = (inp[5]) ? node12386 : node12383;
															assign node12383 = (inp[3]) ? 4'b1110 : 4'b1010;
															assign node12386 = (inp[3]) ? 4'b1010 : 4'b1111;
									assign node12389 = (inp[11]) ? node12501 : node12390;
										assign node12390 = (inp[12]) ? node12438 : node12391;
											assign node12391 = (inp[3]) ? node12407 : node12392;
												assign node12392 = (inp[5]) ? node12396 : node12393;
													assign node12393 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node12396 = (inp[13]) ? node12402 : node12397;
														assign node12397 = (inp[0]) ? node12399 : 4'b1110;
															assign node12399 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node12402 = (inp[4]) ? 4'b1011 : node12403;
															assign node12403 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node12407 = (inp[13]) ? node12423 : node12408;
													assign node12408 = (inp[0]) ? node12416 : node12409;
														assign node12409 = (inp[5]) ? node12413 : node12410;
															assign node12410 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node12413 = (inp[4]) ? 4'b1011 : 4'b1110;
														assign node12416 = (inp[4]) ? node12420 : node12417;
															assign node12417 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node12420 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node12423 = (inp[10]) ? node12429 : node12424;
														assign node12424 = (inp[5]) ? 4'b1111 : node12425;
															assign node12425 = (inp[0]) ? 4'b1011 : 4'b1111;
														assign node12429 = (inp[4]) ? node12433 : node12430;
															assign node12430 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node12433 = (inp[5]) ? 4'b1111 : node12434;
																assign node12434 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node12438 = (inp[0]) ? node12470 : node12439;
												assign node12439 = (inp[5]) ? node12457 : node12440;
													assign node12440 = (inp[13]) ? node12448 : node12441;
														assign node12441 = (inp[3]) ? node12445 : node12442;
															assign node12442 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node12445 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node12448 = (inp[10]) ? node12450 : 4'b1010;
															assign node12450 = (inp[3]) ? node12454 : node12451;
																assign node12451 = (inp[4]) ? 4'b1010 : 4'b1111;
																assign node12454 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node12457 = (inp[13]) ? node12463 : node12458;
														assign node12458 = (inp[3]) ? 4'b1011 : node12459;
															assign node12459 = (inp[4]) ? 4'b1011 : 4'b1110;
														assign node12463 = (inp[4]) ? node12467 : node12464;
															assign node12464 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node12467 = (inp[3]) ? 4'b1010 : 4'b1111;
												assign node12470 = (inp[13]) ? node12484 : node12471;
													assign node12471 = (inp[3]) ? node12479 : node12472;
														assign node12472 = (inp[5]) ? node12476 : node12473;
															assign node12473 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node12476 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node12479 = (inp[10]) ? node12481 : 4'b1111;
															assign node12481 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node12484 = (inp[4]) ? node12490 : node12485;
														assign node12485 = (inp[5]) ? 4'b1011 : node12486;
															assign node12486 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node12490 = (inp[10]) ? node12496 : node12491;
															assign node12491 = (inp[3]) ? 4'b1110 : node12492;
																assign node12492 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node12496 = (inp[3]) ? 4'b1010 : node12497;
																assign node12497 = (inp[5]) ? 4'b1110 : 4'b1010;
										assign node12501 = (inp[12]) ? node12547 : node12502;
											assign node12502 = (inp[5]) ? node12520 : node12503;
												assign node12503 = (inp[13]) ? node12513 : node12504;
													assign node12504 = (inp[4]) ? node12510 : node12505;
														assign node12505 = (inp[0]) ? node12507 : 4'b1010;
															assign node12507 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node12510 = (inp[0]) ? 4'b1010 : 4'b1110;
													assign node12513 = (inp[3]) ? node12515 : 4'b1110;
														assign node12515 = (inp[4]) ? node12517 : 4'b1110;
															assign node12517 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node12520 = (inp[13]) ? node12530 : node12521;
													assign node12521 = (inp[4]) ? node12523 : 4'b1111;
														assign node12523 = (inp[3]) ? node12527 : node12524;
															assign node12524 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12527 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12530 = (inp[4]) ? node12544 : node12531;
														assign node12531 = (inp[10]) ? node12539 : node12532;
															assign node12532 = (inp[0]) ? node12536 : node12533;
																assign node12533 = (inp[3]) ? 4'b1010 : 4'b1011;
																assign node12536 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node12539 = (inp[3]) ? node12541 : 4'b1010;
																assign node12541 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12544 = (inp[3]) ? 4'b1110 : 4'b1010;
											assign node12547 = (inp[5]) ? node12573 : node12548;
												assign node12548 = (inp[13]) ? node12562 : node12549;
													assign node12549 = (inp[4]) ? node12555 : node12550;
														assign node12550 = (inp[3]) ? 4'b1110 : node12551;
															assign node12551 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12555 = (inp[3]) ? node12559 : node12556;
															assign node12556 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12559 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12562 = (inp[10]) ? 4'b1011 : node12563;
														assign node12563 = (inp[0]) ? 4'b1111 : node12564;
															assign node12564 = (inp[3]) ? node12568 : node12565;
																assign node12565 = (inp[4]) ? 4'b1011 : 4'b1110;
																assign node12568 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node12573 = (inp[0]) ? node12589 : node12574;
													assign node12574 = (inp[4]) ? node12582 : node12575;
														assign node12575 = (inp[3]) ? node12579 : node12576;
															assign node12576 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node12579 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node12582 = (inp[13]) ? node12586 : node12583;
															assign node12583 = (inp[3]) ? 4'b1110 : 4'b1010;
															assign node12586 = (inp[3]) ? 4'b1011 : 4'b1110;
													assign node12589 = (inp[4]) ? node12597 : node12590;
														assign node12590 = (inp[3]) ? node12594 : node12591;
															assign node12591 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node12594 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node12597 = (inp[3]) ? node12601 : node12598;
															assign node12598 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node12601 = (inp[13]) ? 4'b1011 : 4'b1110;
								assign node12604 = (inp[5]) ? node12804 : node12605;
									assign node12605 = (inp[13]) ? node12687 : node12606;
										assign node12606 = (inp[12]) ? node12642 : node12607;
											assign node12607 = (inp[10]) ? node12615 : node12608;
												assign node12608 = (inp[11]) ? node12612 : node12609;
													assign node12609 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12612 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node12615 = (inp[4]) ? node12631 : node12616;
													assign node12616 = (inp[0]) ? node12624 : node12617;
														assign node12617 = (inp[3]) ? 4'b1011 : node12618;
															assign node12618 = (inp[9]) ? 4'b1010 : node12619;
																assign node12619 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12624 = (inp[9]) ? node12628 : node12625;
															assign node12625 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node12628 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12631 = (inp[3]) ? 4'b1011 : node12632;
														assign node12632 = (inp[0]) ? 4'b1011 : node12633;
															assign node12633 = (inp[11]) ? node12637 : node12634;
																assign node12634 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node12637 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node12642 = (inp[3]) ? node12664 : node12643;
												assign node12643 = (inp[4]) ? node12657 : node12644;
													assign node12644 = (inp[9]) ? node12650 : node12645;
														assign node12645 = (inp[11]) ? node12647 : 4'b1111;
															assign node12647 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node12650 = (inp[11]) ? node12654 : node12651;
															assign node12651 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12654 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node12657 = (inp[9]) ? node12661 : node12658;
														assign node12658 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12661 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node12664 = (inp[9]) ? node12676 : node12665;
													assign node12665 = (inp[11]) ? node12671 : node12666;
														assign node12666 = (inp[4]) ? 4'b1010 : node12667;
															assign node12667 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12671 = (inp[4]) ? 4'b1011 : node12672;
															assign node12672 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12676 = (inp[11]) ? node12682 : node12677;
														assign node12677 = (inp[4]) ? 4'b1011 : node12678;
															assign node12678 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12682 = (inp[4]) ? 4'b1010 : node12683;
															assign node12683 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node12687 = (inp[3]) ? node12727 : node12688;
											assign node12688 = (inp[4]) ? node12704 : node12689;
												assign node12689 = (inp[12]) ? node12697 : node12690;
													assign node12690 = (inp[11]) ? node12694 : node12691;
														assign node12691 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12694 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12697 = (inp[11]) ? node12701 : node12698;
														assign node12698 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node12701 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node12704 = (inp[12]) ? node12720 : node12705;
													assign node12705 = (inp[10]) ? node12711 : node12706;
														assign node12706 = (inp[9]) ? 4'b1110 : node12707;
															assign node12707 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12711 = (inp[0]) ? node12717 : node12712;
															assign node12712 = (inp[11]) ? 4'b1111 : node12713;
																assign node12713 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node12717 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12720 = (inp[9]) ? node12724 : node12721;
														assign node12721 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12724 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node12727 = (inp[10]) ? node12765 : node12728;
												assign node12728 = (inp[4]) ? node12744 : node12729;
													assign node12729 = (inp[12]) ? node12739 : node12730;
														assign node12730 = (inp[11]) ? node12732 : 4'b1111;
															assign node12732 = (inp[0]) ? node12736 : node12733;
																assign node12733 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node12736 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node12739 = (inp[9]) ? 4'b1111 : node12740;
															assign node12740 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12744 = (inp[12]) ? node12754 : node12745;
														assign node12745 = (inp[9]) ? 4'b1111 : node12746;
															assign node12746 = (inp[0]) ? node12750 : node12747;
																assign node12747 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12750 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12754 = (inp[9]) ? node12760 : node12755;
															assign node12755 = (inp[0]) ? node12757 : 4'b1111;
																assign node12757 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12760 = (inp[0]) ? node12762 : 4'b1110;
																assign node12762 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12765 = (inp[12]) ? node12789 : node12766;
													assign node12766 = (inp[11]) ? node12782 : node12767;
														assign node12767 = (inp[4]) ? node12775 : node12768;
															assign node12768 = (inp[9]) ? node12772 : node12769;
																assign node12769 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node12772 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12775 = (inp[0]) ? node12779 : node12776;
																assign node12776 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12779 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12782 = (inp[0]) ? node12786 : node12783;
															assign node12783 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node12786 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12789 = (inp[11]) ? node12797 : node12790;
														assign node12790 = (inp[9]) ? node12794 : node12791;
															assign node12791 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node12794 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node12797 = (inp[9]) ? 4'b1110 : node12798;
															assign node12798 = (inp[0]) ? 4'b1111 : node12799;
																assign node12799 = (inp[4]) ? 4'b1110 : 4'b1111;
									assign node12804 = (inp[13]) ? node12914 : node12805;
										assign node12805 = (inp[4]) ? node12851 : node12806;
											assign node12806 = (inp[12]) ? node12830 : node12807;
												assign node12807 = (inp[0]) ? node12823 : node12808;
													assign node12808 = (inp[3]) ? node12814 : node12809;
														assign node12809 = (inp[11]) ? node12811 : 4'b1111;
															assign node12811 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12814 = (inp[10]) ? node12816 : 4'b1110;
															assign node12816 = (inp[11]) ? node12820 : node12817;
																assign node12817 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node12820 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12823 = (inp[9]) ? node12827 : node12824;
														assign node12824 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12827 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12830 = (inp[3]) ? node12838 : node12831;
													assign node12831 = (inp[9]) ? node12835 : node12832;
														assign node12832 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12835 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node12838 = (inp[11]) ? node12846 : node12839;
														assign node12839 = (inp[0]) ? node12843 : node12840;
															assign node12840 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12843 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12846 = (inp[0]) ? node12848 : 4'b1111;
															assign node12848 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node12851 = (inp[10]) ? node12883 : node12852;
												assign node12852 = (inp[12]) ? node12866 : node12853;
													assign node12853 = (inp[0]) ? node12861 : node12854;
														assign node12854 = (inp[9]) ? node12856 : 4'b1111;
															assign node12856 = (inp[11]) ? node12858 : 4'b1110;
																assign node12858 = (inp[3]) ? 4'b1110 : 4'b1111;
														assign node12861 = (inp[9]) ? node12863 : 4'b1110;
															assign node12863 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12866 = (inp[0]) ? node12876 : node12867;
														assign node12867 = (inp[3]) ? node12869 : 4'b1110;
															assign node12869 = (inp[9]) ? node12873 : node12870;
																assign node12870 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node12873 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12876 = (inp[3]) ? 4'b1111 : node12877;
															assign node12877 = (inp[11]) ? node12879 : 4'b1111;
																assign node12879 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node12883 = (inp[3]) ? node12897 : node12884;
													assign node12884 = (inp[0]) ? node12886 : 4'b1111;
														assign node12886 = (inp[12]) ? node12892 : node12887;
															assign node12887 = (inp[11]) ? node12889 : 4'b1111;
																assign node12889 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12892 = (inp[9]) ? 4'b1111 : node12893;
																assign node12893 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12897 = (inp[0]) ? node12905 : node12898;
														assign node12898 = (inp[12]) ? 4'b1110 : node12899;
															assign node12899 = (inp[11]) ? node12901 : 4'b1111;
																assign node12901 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node12905 = (inp[12]) ? 4'b1111 : node12906;
															assign node12906 = (inp[9]) ? node12910 : node12907;
																assign node12907 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12910 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node12914 = (inp[12]) ? node12952 : node12915;
											assign node12915 = (inp[4]) ? node12933 : node12916;
												assign node12916 = (inp[11]) ? node12928 : node12917;
													assign node12917 = (inp[9]) ? node12923 : node12918;
														assign node12918 = (inp[0]) ? 4'b1010 : node12919;
															assign node12919 = (inp[3]) ? 4'b1010 : 4'b1011;
														assign node12923 = (inp[3]) ? 4'b1011 : node12924;
															assign node12924 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12928 = (inp[9]) ? 4'b1010 : node12929;
														assign node12929 = (inp[3]) ? 4'b1011 : 4'b1010;
												assign node12933 = (inp[9]) ? node12945 : node12934;
													assign node12934 = (inp[11]) ? node12940 : node12935;
														assign node12935 = (inp[0]) ? 4'b1010 : node12936;
															assign node12936 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node12940 = (inp[0]) ? 4'b1011 : node12941;
															assign node12941 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node12945 = (inp[11]) ? 4'b1010 : node12946;
														assign node12946 = (inp[3]) ? node12948 : 4'b1011;
															assign node12948 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node12952 = (inp[4]) ? node12984 : node12953;
												assign node12953 = (inp[3]) ? node12967 : node12954;
													assign node12954 = (inp[10]) ? node12960 : node12955;
														assign node12955 = (inp[9]) ? node12957 : 4'b1110;
															assign node12957 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12960 = (inp[0]) ? node12962 : 4'b1110;
															assign node12962 = (inp[11]) ? 4'b1110 : node12963;
																assign node12963 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12967 = (inp[9]) ? node12975 : node12968;
														assign node12968 = (inp[11]) ? node12972 : node12969;
															assign node12969 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12972 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12975 = (inp[10]) ? node12981 : node12976;
															assign node12976 = (inp[11]) ? node12978 : 4'b1011;
																assign node12978 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12981 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node12984 = (inp[10]) ? node12996 : node12985;
													assign node12985 = (inp[9]) ? node12993 : node12986;
														assign node12986 = (inp[11]) ? node12988 : 4'b1010;
															assign node12988 = (inp[3]) ? node12990 : 4'b1011;
																assign node12990 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node12993 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12996 = (inp[9]) ? node13006 : node12997;
														assign node12997 = (inp[11]) ? node13003 : node12998;
															assign node12998 = (inp[0]) ? 4'b1010 : node12999;
																assign node12999 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node13003 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node13006 = (inp[11]) ? 4'b1010 : node13007;
															assign node13007 = (inp[3]) ? 4'b1010 : 4'b1011;
							assign node13011 = (inp[4]) ? node13355 : node13012;
								assign node13012 = (inp[11]) ? node13178 : node13013;
									assign node13013 = (inp[9]) ? node13091 : node13014;
										assign node13014 = (inp[13]) ? node13050 : node13015;
											assign node13015 = (inp[5]) ? node13033 : node13016;
												assign node13016 = (inp[12]) ? node13024 : node13017;
													assign node13017 = (inp[0]) ? node13021 : node13018;
														assign node13018 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node13021 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node13024 = (inp[1]) ? node13030 : node13025;
														assign node13025 = (inp[3]) ? node13027 : 4'b1011;
															assign node13027 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13030 = (inp[3]) ? 4'b1010 : 4'b1110;
												assign node13033 = (inp[12]) ? node13041 : node13034;
													assign node13034 = (inp[3]) ? node13038 : node13035;
														assign node13035 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13038 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node13041 = (inp[1]) ? node13045 : node13042;
														assign node13042 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node13045 = (inp[3]) ? 4'b1111 : node13046;
															assign node13046 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node13050 = (inp[5]) ? node13072 : node13051;
												assign node13051 = (inp[12]) ? node13059 : node13052;
													assign node13052 = (inp[0]) ? node13056 : node13053;
														assign node13053 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node13056 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node13059 = (inp[0]) ? node13069 : node13060;
														assign node13060 = (inp[10]) ? node13062 : 4'b1111;
															assign node13062 = (inp[3]) ? node13066 : node13063;
																assign node13063 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node13066 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node13069 = (inp[3]) ? 4'b1110 : 4'b1111;
												assign node13072 = (inp[12]) ? node13078 : node13073;
													assign node13073 = (inp[3]) ? node13075 : 4'b1010;
														assign node13075 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node13078 = (inp[1]) ? node13086 : node13079;
														assign node13079 = (inp[3]) ? node13083 : node13080;
															assign node13080 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node13083 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13086 = (inp[0]) ? node13088 : 4'b1111;
															assign node13088 = (inp[3]) ? 4'b1010 : 4'b1110;
										assign node13091 = (inp[5]) ? node13135 : node13092;
											assign node13092 = (inp[13]) ? node13112 : node13093;
												assign node13093 = (inp[3]) ? node13101 : node13094;
													assign node13094 = (inp[1]) ? node13096 : 4'b1010;
														assign node13096 = (inp[12]) ? 4'b1111 : node13097;
															assign node13097 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node13101 = (inp[12]) ? node13107 : node13102;
														assign node13102 = (inp[1]) ? node13104 : 4'b1011;
															assign node13104 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node13107 = (inp[1]) ? 4'b1011 : node13108;
															assign node13108 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node13112 = (inp[12]) ? node13122 : node13113;
													assign node13113 = (inp[0]) ? node13117 : node13114;
														assign node13114 = (inp[3]) ? 4'b1110 : 4'b1111;
														assign node13117 = (inp[3]) ? node13119 : 4'b1110;
															assign node13119 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node13122 = (inp[0]) ? node13130 : node13123;
														assign node13123 = (inp[3]) ? node13127 : node13124;
															assign node13124 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node13127 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node13130 = (inp[3]) ? node13132 : 4'b1010;
															assign node13132 = (inp[1]) ? 4'b1111 : 4'b1010;
											assign node13135 = (inp[13]) ? node13155 : node13136;
												assign node13136 = (inp[12]) ? node13146 : node13137;
													assign node13137 = (inp[1]) ? node13141 : node13138;
														assign node13138 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node13141 = (inp[0]) ? node13143 : 4'b1111;
															assign node13143 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node13146 = (inp[1]) ? node13150 : node13147;
														assign node13147 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node13150 = (inp[3]) ? 4'b1110 : node13151;
															assign node13151 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node13155 = (inp[12]) ? node13157 : 4'b1011;
													assign node13157 = (inp[0]) ? node13171 : node13158;
														assign node13158 = (inp[10]) ? node13164 : node13159;
															assign node13159 = (inp[1]) ? node13161 : 4'b1110;
																assign node13161 = (inp[3]) ? 4'b1011 : 4'b1110;
															assign node13164 = (inp[3]) ? node13168 : node13165;
																assign node13165 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node13168 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node13171 = (inp[1]) ? node13175 : node13172;
															assign node13172 = (inp[3]) ? 4'b1111 : 4'b1010;
															assign node13175 = (inp[3]) ? 4'b1011 : 4'b1111;
									assign node13178 = (inp[9]) ? node13274 : node13179;
										assign node13179 = (inp[1]) ? node13227 : node13180;
											assign node13180 = (inp[5]) ? node13210 : node13181;
												assign node13181 = (inp[12]) ? node13199 : node13182;
													assign node13182 = (inp[13]) ? node13190 : node13183;
														assign node13183 = (inp[10]) ? 4'b1011 : node13184;
															assign node13184 = (inp[3]) ? 4'b1011 : node13185;
																assign node13185 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node13190 = (inp[10]) ? node13192 : 4'b1111;
															assign node13192 = (inp[0]) ? node13196 : node13193;
																assign node13193 = (inp[3]) ? 4'b1110 : 4'b1111;
																assign node13196 = (inp[3]) ? 4'b1111 : 4'b1110;
													assign node13199 = (inp[3]) ? node13203 : node13200;
														assign node13200 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node13203 = (inp[13]) ? node13207 : node13204;
															assign node13204 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node13207 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node13210 = (inp[13]) ? node13220 : node13211;
													assign node13211 = (inp[12]) ? node13217 : node13212;
														assign node13212 = (inp[0]) ? node13214 : 4'b1110;
															assign node13214 = (inp[3]) ? 4'b1110 : 4'b1111;
														assign node13217 = (inp[3]) ? 4'b1011 : 4'b1111;
													assign node13220 = (inp[12]) ? node13222 : 4'b1011;
														assign node13222 = (inp[3]) ? 4'b1110 : node13223;
															assign node13223 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node13227 = (inp[3]) ? node13255 : node13228;
												assign node13228 = (inp[12]) ? node13244 : node13229;
													assign node13229 = (inp[0]) ? node13237 : node13230;
														assign node13230 = (inp[10]) ? node13232 : 4'b1011;
															assign node13232 = (inp[5]) ? 4'b1011 : node13233;
																assign node13233 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node13237 = (inp[5]) ? node13241 : node13238;
															assign node13238 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node13241 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node13244 = (inp[5]) ? node13248 : node13245;
														assign node13245 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node13248 = (inp[13]) ? node13252 : node13249;
															assign node13249 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node13252 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node13255 = (inp[12]) ? node13269 : node13256;
													assign node13256 = (inp[0]) ? node13260 : node13257;
														assign node13257 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node13260 = (inp[10]) ? node13266 : node13261;
															assign node13261 = (inp[5]) ? 4'b1110 : node13262;
																assign node13262 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node13266 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node13269 = (inp[13]) ? 4'b1011 : node13270;
														assign node13270 = (inp[5]) ? 4'b1110 : 4'b1011;
										assign node13274 = (inp[5]) ? node13318 : node13275;
											assign node13275 = (inp[13]) ? node13295 : node13276;
												assign node13276 = (inp[12]) ? node13288 : node13277;
													assign node13277 = (inp[1]) ? node13283 : node13278;
														assign node13278 = (inp[3]) ? 4'b1010 : node13279;
															assign node13279 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node13283 = (inp[3]) ? 4'b1011 : node13284;
															assign node13284 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node13288 = (inp[1]) ? node13292 : node13289;
														assign node13289 = (inp[3]) ? 4'b1110 : 4'b1011;
														assign node13292 = (inp[3]) ? 4'b1010 : 4'b1110;
												assign node13295 = (inp[12]) ? node13307 : node13296;
													assign node13296 = (inp[1]) ? node13302 : node13297;
														assign node13297 = (inp[0]) ? 4'b1110 : node13298;
															assign node13298 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node13302 = (inp[0]) ? 4'b1111 : node13303;
															assign node13303 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node13307 = (inp[1]) ? node13311 : node13308;
														assign node13308 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node13311 = (inp[3]) ? node13315 : node13312;
															assign node13312 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node13315 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node13318 = (inp[13]) ? node13338 : node13319;
												assign node13319 = (inp[12]) ? node13333 : node13320;
													assign node13320 = (inp[1]) ? node13326 : node13321;
														assign node13321 = (inp[0]) ? node13323 : 4'b1111;
															assign node13323 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node13326 = (inp[10]) ? 4'b1110 : node13327;
															assign node13327 = (inp[0]) ? 4'b1111 : node13328;
																assign node13328 = (inp[3]) ? 4'b1110 : 4'b1111;
													assign node13333 = (inp[3]) ? 4'b1010 : node13334;
														assign node13334 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node13338 = (inp[12]) ? node13346 : node13339;
													assign node13339 = (inp[1]) ? node13341 : 4'b1010;
														assign node13341 = (inp[0]) ? 4'b1010 : node13342;
															assign node13342 = (inp[3]) ? 4'b1011 : 4'b1010;
													assign node13346 = (inp[0]) ? node13352 : node13347;
														assign node13347 = (inp[3]) ? 4'b1111 : node13348;
															assign node13348 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node13352 = (inp[1]) ? 4'b1010 : 4'b1110;
								assign node13355 = (inp[0]) ? node13629 : node13356;
									assign node13356 = (inp[1]) ? node13474 : node13357;
										assign node13357 = (inp[5]) ? node13419 : node13358;
											assign node13358 = (inp[12]) ? node13390 : node13359;
												assign node13359 = (inp[3]) ? node13381 : node13360;
													assign node13360 = (inp[13]) ? node13368 : node13361;
														assign node13361 = (inp[9]) ? node13365 : node13362;
															assign node13362 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node13365 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node13368 = (inp[10]) ? node13376 : node13369;
															assign node13369 = (inp[11]) ? node13373 : node13370;
																assign node13370 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node13373 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node13376 = (inp[9]) ? node13378 : 4'b1110;
																assign node13378 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node13381 = (inp[13]) ? 4'b1011 : node13382;
														assign node13382 = (inp[11]) ? node13386 : node13383;
															assign node13383 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node13386 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node13390 = (inp[11]) ? node13404 : node13391;
													assign node13391 = (inp[9]) ? node13397 : node13392;
														assign node13392 = (inp[13]) ? 4'b1010 : node13393;
															assign node13393 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node13397 = (inp[13]) ? node13401 : node13398;
															assign node13398 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node13401 = (inp[3]) ? 4'b1110 : 4'b1011;
													assign node13404 = (inp[9]) ? node13412 : node13405;
														assign node13405 = (inp[3]) ? node13409 : node13406;
															assign node13406 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node13409 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node13412 = (inp[13]) ? node13416 : node13413;
															assign node13413 = (inp[3]) ? 4'b1010 : 4'b1110;
															assign node13416 = (inp[3]) ? 4'b1111 : 4'b1010;
											assign node13419 = (inp[12]) ? node13449 : node13420;
												assign node13420 = (inp[11]) ? node13436 : node13421;
													assign node13421 = (inp[9]) ? node13431 : node13422;
														assign node13422 = (inp[10]) ? 4'b1011 : node13423;
															assign node13423 = (inp[3]) ? node13427 : node13424;
																assign node13424 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node13427 = (inp[13]) ? 4'b1110 : 4'b1011;
														assign node13431 = (inp[13]) ? node13433 : 4'b1010;
															assign node13433 = (inp[3]) ? 4'b1111 : 4'b1010;
													assign node13436 = (inp[9]) ? node13444 : node13437;
														assign node13437 = (inp[3]) ? node13441 : node13438;
															assign node13438 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node13441 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node13444 = (inp[3]) ? node13446 : 4'b1011;
															assign node13446 = (inp[13]) ? 4'b1110 : 4'b1011;
												assign node13449 = (inp[11]) ? node13463 : node13450;
													assign node13450 = (inp[9]) ? node13456 : node13451;
														assign node13451 = (inp[3]) ? node13453 : 4'b1110;
															assign node13453 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node13456 = (inp[13]) ? node13460 : node13457;
															assign node13457 = (inp[3]) ? 4'b1111 : 4'b1011;
															assign node13460 = (inp[3]) ? 4'b1010 : 4'b1111;
													assign node13463 = (inp[9]) ? node13467 : node13464;
														assign node13464 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node13467 = (inp[3]) ? node13471 : node13468;
															assign node13468 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node13471 = (inp[13]) ? 4'b1011 : 4'b1110;
										assign node13474 = (inp[10]) ? node13536 : node13475;
											assign node13475 = (inp[12]) ? node13507 : node13476;
												assign node13476 = (inp[9]) ? node13494 : node13477;
													assign node13477 = (inp[11]) ? node13485 : node13478;
														assign node13478 = (inp[13]) ? node13480 : 4'b1111;
															assign node13480 = (inp[5]) ? node13482 : 4'b1110;
																assign node13482 = (inp[3]) ? 4'b1010 : 4'b1011;
														assign node13485 = (inp[5]) ? node13491 : node13486;
															assign node13486 = (inp[13]) ? 4'b1110 : node13487;
																assign node13487 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node13491 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node13494 = (inp[5]) ? node13502 : node13495;
														assign node13495 = (inp[13]) ? node13497 : 4'b1010;
															assign node13497 = (inp[3]) ? node13499 : 4'b1110;
																assign node13499 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node13502 = (inp[13]) ? 4'b1010 : node13503;
															assign node13503 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node13507 = (inp[11]) ? node13527 : node13508;
													assign node13508 = (inp[5]) ? node13520 : node13509;
														assign node13509 = (inp[13]) ? node13517 : node13510;
															assign node13510 = (inp[3]) ? node13514 : node13511;
																assign node13511 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node13514 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node13517 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node13520 = (inp[13]) ? node13524 : node13521;
															assign node13521 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node13524 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node13527 = (inp[9]) ? node13531 : node13528;
														assign node13528 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node13531 = (inp[3]) ? node13533 : 4'b1111;
															assign node13533 = (inp[5]) ? 4'b1111 : 4'b1010;
											assign node13536 = (inp[12]) ? node13584 : node13537;
												assign node13537 = (inp[9]) ? node13565 : node13538;
													assign node13538 = (inp[11]) ? node13552 : node13539;
														assign node13539 = (inp[3]) ? node13547 : node13540;
															assign node13540 = (inp[13]) ? node13544 : node13541;
																assign node13541 = (inp[5]) ? 4'b1111 : 4'b1011;
																assign node13544 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node13547 = (inp[13]) ? 4'b1010 : node13548;
																assign node13548 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node13552 = (inp[3]) ? node13558 : node13553;
															assign node13553 = (inp[5]) ? node13555 : 4'b1110;
																assign node13555 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node13558 = (inp[5]) ? node13562 : node13559;
																assign node13559 = (inp[13]) ? 4'b1111 : 4'b1011;
																assign node13562 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node13565 = (inp[11]) ? node13573 : node13566;
														assign node13566 = (inp[13]) ? node13570 : node13567;
															assign node13567 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node13570 = (inp[3]) ? 4'b1111 : 4'b1110;
														assign node13573 = (inp[3]) ? node13581 : node13574;
															assign node13574 = (inp[13]) ? node13578 : node13575;
																assign node13575 = (inp[5]) ? 4'b1111 : 4'b1011;
																assign node13578 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node13581 = (inp[13]) ? 4'b1010 : 4'b1111;
												assign node13584 = (inp[3]) ? node13608 : node13585;
													assign node13585 = (inp[5]) ? node13595 : node13586;
														assign node13586 = (inp[13]) ? node13588 : 4'b1010;
															assign node13588 = (inp[9]) ? node13592 : node13589;
																assign node13589 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node13592 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node13595 = (inp[13]) ? node13601 : node13596;
															assign node13596 = (inp[11]) ? node13598 : 4'b1110;
																assign node13598 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node13601 = (inp[9]) ? node13605 : node13602;
																assign node13602 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node13605 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node13608 = (inp[11]) ? node13614 : node13609;
														assign node13609 = (inp[9]) ? node13611 : 4'b1010;
															assign node13611 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node13614 = (inp[9]) ? node13622 : node13615;
															assign node13615 = (inp[13]) ? node13619 : node13616;
																assign node13616 = (inp[5]) ? 4'b1110 : 4'b1011;
																assign node13619 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node13622 = (inp[5]) ? node13626 : node13623;
																assign node13623 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node13626 = (inp[13]) ? 4'b1010 : 4'b1111;
									assign node13629 = (inp[13]) ? node13723 : node13630;
										assign node13630 = (inp[5]) ? node13676 : node13631;
											assign node13631 = (inp[1]) ? node13657 : node13632;
												assign node13632 = (inp[9]) ? node13644 : node13633;
													assign node13633 = (inp[11]) ? node13639 : node13634;
														assign node13634 = (inp[12]) ? node13636 : 4'b1010;
															assign node13636 = (inp[3]) ? 4'b1010 : 4'b1110;
														assign node13639 = (inp[12]) ? node13641 : 4'b1110;
															assign node13641 = (inp[3]) ? 4'b1011 : 4'b1111;
													assign node13644 = (inp[11]) ? node13650 : node13645;
														assign node13645 = (inp[3]) ? 4'b1110 : node13646;
															assign node13646 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node13650 = (inp[12]) ? node13654 : node13651;
															assign node13651 = (inp[3]) ? 4'b1111 : 4'b1010;
															assign node13654 = (inp[3]) ? 4'b1010 : 4'b1110;
												assign node13657 = (inp[9]) ? node13671 : node13658;
													assign node13658 = (inp[12]) ? node13666 : node13659;
														assign node13659 = (inp[11]) ? node13663 : node13660;
															assign node13660 = (inp[3]) ? 4'b1011 : 4'b1010;
															assign node13663 = (inp[3]) ? 4'b1010 : 4'b1011;
														assign node13666 = (inp[11]) ? 4'b1011 : node13667;
															assign node13667 = (inp[3]) ? 4'b1011 : 4'b1010;
													assign node13671 = (inp[3]) ? 4'b1010 : node13672;
														assign node13672 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node13676 = (inp[1]) ? node13716 : node13677;
												assign node13677 = (inp[10]) ? node13701 : node13678;
													assign node13678 = (inp[11]) ? node13692 : node13679;
														assign node13679 = (inp[9]) ? node13687 : node13680;
															assign node13680 = (inp[12]) ? node13684 : node13681;
																assign node13681 = (inp[3]) ? 4'b1011 : 4'b1111;
																assign node13684 = (inp[3]) ? 4'b1111 : 4'b1010;
															assign node13687 = (inp[3]) ? node13689 : 4'b1110;
																assign node13689 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node13692 = (inp[9]) ? node13698 : node13693;
															assign node13693 = (inp[3]) ? node13695 : 4'b1110;
																assign node13695 = (inp[12]) ? 4'b1110 : 4'b1010;
															assign node13698 = (inp[3]) ? 4'b1011 : 4'b1010;
													assign node13701 = (inp[11]) ? node13713 : node13702;
														assign node13702 = (inp[9]) ? node13708 : node13703;
															assign node13703 = (inp[3]) ? 4'b1111 : node13704;
																assign node13704 = (inp[12]) ? 4'b1010 : 4'b1111;
															assign node13708 = (inp[3]) ? node13710 : 4'b1110;
																assign node13710 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node13713 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node13716 = (inp[9]) ? node13720 : node13717;
													assign node13717 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node13720 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node13723 = (inp[5]) ? node13755 : node13724;
											assign node13724 = (inp[1]) ? node13748 : node13725;
												assign node13725 = (inp[9]) ? node13735 : node13726;
													assign node13726 = (inp[12]) ? node13730 : node13727;
														assign node13727 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node13730 = (inp[3]) ? 4'b1111 : node13731;
															assign node13731 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13735 = (inp[3]) ? node13743 : node13736;
														assign node13736 = (inp[12]) ? node13740 : node13737;
															assign node13737 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13740 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node13743 = (inp[11]) ? 4'b1110 : node13744;
															assign node13744 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node13748 = (inp[11]) ? node13752 : node13749;
													assign node13749 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node13752 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node13755 = (inp[1]) ? node13783 : node13756;
												assign node13756 = (inp[9]) ? node13770 : node13757;
													assign node13757 = (inp[11]) ? node13763 : node13758;
														assign node13758 = (inp[3]) ? 4'b1010 : node13759;
															assign node13759 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node13763 = (inp[10]) ? node13767 : node13764;
															assign node13764 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node13767 = (inp[3]) ? 4'b1110 : 4'b1011;
													assign node13770 = (inp[3]) ? node13778 : node13771;
														assign node13771 = (inp[12]) ? node13775 : node13772;
															assign node13772 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node13775 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node13778 = (inp[12]) ? 4'b1011 : node13779;
															assign node13779 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node13783 = (inp[12]) ? node13791 : node13784;
													assign node13784 = (inp[11]) ? node13788 : node13785;
														assign node13785 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node13788 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node13791 = (inp[10]) ? node13799 : node13792;
														assign node13792 = (inp[9]) ? node13796 : node13793;
															assign node13793 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node13796 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node13799 = (inp[3]) ? node13801 : 4'b1011;
															assign node13801 = (inp[9]) ? 4'b1011 : 4'b1010;
						assign node13804 = (inp[5]) ? node14606 : node13805;
							assign node13805 = (inp[13]) ? node14253 : node13806;
								assign node13806 = (inp[12]) ? node14082 : node13807;
									assign node13807 = (inp[4]) ? node13953 : node13808;
										assign node13808 = (inp[10]) ? node13874 : node13809;
											assign node13809 = (inp[0]) ? node13843 : node13810;
												assign node13810 = (inp[3]) ? node13826 : node13811;
													assign node13811 = (inp[1]) ? 4'b1001 : node13812;
														assign node13812 = (inp[2]) ? node13818 : node13813;
															assign node13813 = (inp[11]) ? 4'b1100 : node13814;
																assign node13814 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node13818 = (inp[9]) ? node13822 : node13819;
																assign node13819 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node13822 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13826 = (inp[1]) ? node13834 : node13827;
														assign node13827 = (inp[9]) ? 4'b1000 : node13828;
															assign node13828 = (inp[2]) ? 4'b1001 : node13829;
																assign node13829 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13834 = (inp[2]) ? node13836 : 4'b1100;
															assign node13836 = (inp[11]) ? node13840 : node13837;
																assign node13837 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node13840 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node13843 = (inp[9]) ? node13867 : node13844;
													assign node13844 = (inp[11]) ? node13856 : node13845;
														assign node13845 = (inp[3]) ? node13851 : node13846;
															assign node13846 = (inp[1]) ? node13848 : 4'b1101;
																assign node13848 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node13851 = (inp[1]) ? node13853 : 4'b1000;
																assign node13853 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node13856 = (inp[3]) ? node13862 : node13857;
															assign node13857 = (inp[1]) ? 4'b1000 : node13858;
																assign node13858 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node13862 = (inp[1]) ? node13864 : 4'b1001;
																assign node13864 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node13867 = (inp[2]) ? 4'b1000 : node13868;
														assign node13868 = (inp[3]) ? 4'b1101 : node13869;
															assign node13869 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node13874 = (inp[9]) ? node13918 : node13875;
												assign node13875 = (inp[2]) ? node13891 : node13876;
													assign node13876 = (inp[11]) ? node13882 : node13877;
														assign node13877 = (inp[1]) ? node13879 : 4'b1000;
															assign node13879 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node13882 = (inp[1]) ? node13886 : node13883;
															assign node13883 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node13886 = (inp[3]) ? node13888 : 4'b1000;
																assign node13888 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13891 = (inp[0]) ? node13903 : node13892;
														assign node13892 = (inp[11]) ? node13898 : node13893;
															assign node13893 = (inp[1]) ? node13895 : 4'b1100;
																assign node13895 = (inp[3]) ? 4'b1101 : 4'b1001;
															assign node13898 = (inp[3]) ? node13900 : 4'b1101;
																assign node13900 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node13903 = (inp[11]) ? node13911 : node13904;
															assign node13904 = (inp[3]) ? node13908 : node13905;
																assign node13905 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node13908 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node13911 = (inp[3]) ? node13915 : node13912;
																assign node13912 = (inp[1]) ? 4'b1001 : 4'b1100;
																assign node13915 = (inp[1]) ? 4'b1100 : 4'b1001;
												assign node13918 = (inp[0]) ? node13928 : node13919;
													assign node13919 = (inp[1]) ? 4'b1101 : node13920;
														assign node13920 = (inp[3]) ? node13922 : 4'b1101;
															assign node13922 = (inp[2]) ? node13924 : 4'b1001;
																assign node13924 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node13928 = (inp[1]) ? node13938 : node13929;
														assign node13929 = (inp[3]) ? 4'b1001 : node13930;
															assign node13930 = (inp[2]) ? node13934 : node13931;
																assign node13931 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13934 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13938 = (inp[3]) ? node13946 : node13939;
															assign node13939 = (inp[11]) ? node13943 : node13940;
																assign node13940 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node13943 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node13946 = (inp[2]) ? node13950 : node13947;
																assign node13947 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node13950 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node13953 = (inp[3]) ? node14025 : node13954;
											assign node13954 = (inp[0]) ? node13982 : node13955;
												assign node13955 = (inp[1]) ? node13969 : node13956;
													assign node13956 = (inp[10]) ? node13962 : node13957;
														assign node13957 = (inp[11]) ? node13959 : 4'b1001;
															assign node13959 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node13962 = (inp[2]) ? 4'b1001 : node13963;
															assign node13963 = (inp[9]) ? 4'b1000 : node13964;
																assign node13964 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node13969 = (inp[2]) ? node13975 : node13970;
														assign node13970 = (inp[11]) ? node13972 : 4'b1000;
															assign node13972 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node13975 = (inp[11]) ? node13979 : node13976;
															assign node13976 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node13979 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node13982 = (inp[2]) ? node13998 : node13983;
													assign node13983 = (inp[1]) ? node13989 : node13984;
														assign node13984 = (inp[9]) ? node13986 : 4'b1000;
															assign node13986 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13989 = (inp[10]) ? node13991 : 4'b1001;
															assign node13991 = (inp[9]) ? node13995 : node13992;
																assign node13992 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node13995 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node13998 = (inp[1]) ? node14012 : node13999;
														assign node13999 = (inp[10]) ? node14005 : node14000;
															assign node14000 = (inp[11]) ? 4'b1001 : node14001;
																assign node14001 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node14005 = (inp[11]) ? node14009 : node14006;
																assign node14006 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node14009 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node14012 = (inp[10]) ? node14018 : node14013;
															assign node14013 = (inp[9]) ? node14015 : 4'b1000;
																assign node14015 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node14018 = (inp[9]) ? node14022 : node14019;
																assign node14019 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node14022 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node14025 = (inp[1]) ? node14057 : node14026;
												assign node14026 = (inp[9]) ? node14038 : node14027;
													assign node14027 = (inp[2]) ? node14029 : 4'b1101;
														assign node14029 = (inp[10]) ? node14035 : node14030;
															assign node14030 = (inp[0]) ? 4'b1101 : node14031;
																assign node14031 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14035 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node14038 = (inp[10]) ? node14048 : node14039;
														assign node14039 = (inp[2]) ? node14043 : node14040;
															assign node14040 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node14043 = (inp[11]) ? node14045 : 4'b1100;
																assign node14045 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14048 = (inp[11]) ? node14054 : node14049;
															assign node14049 = (inp[0]) ? node14051 : 4'b1101;
																assign node14051 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node14054 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node14057 = (inp[9]) ? node14073 : node14058;
													assign node14058 = (inp[10]) ? node14068 : node14059;
														assign node14059 = (inp[11]) ? node14065 : node14060;
															assign node14060 = (inp[0]) ? node14062 : 4'b1001;
																assign node14062 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node14065 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node14068 = (inp[0]) ? 4'b1000 : node14069;
															assign node14069 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node14073 = (inp[11]) ? node14077 : node14074;
														assign node14074 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node14077 = (inp[2]) ? node14079 : 4'b1001;
															assign node14079 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node14082 = (inp[4]) ? node14184 : node14083;
										assign node14083 = (inp[0]) ? node14141 : node14084;
											assign node14084 = (inp[1]) ? node14102 : node14085;
												assign node14085 = (inp[10]) ? node14095 : node14086;
													assign node14086 = (inp[3]) ? node14088 : 4'b1000;
														assign node14088 = (inp[9]) ? node14092 : node14089;
															assign node14089 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node14092 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14095 = (inp[9]) ? node14099 : node14096;
														assign node14096 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node14099 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node14102 = (inp[3]) ? node14126 : node14103;
													assign node14103 = (inp[10]) ? node14117 : node14104;
														assign node14104 = (inp[11]) ? node14110 : node14105;
															assign node14105 = (inp[2]) ? node14107 : 4'b1000;
																assign node14107 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node14110 = (inp[2]) ? node14114 : node14111;
																assign node14111 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node14114 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14117 = (inp[11]) ? 4'b1000 : node14118;
															assign node14118 = (inp[9]) ? node14122 : node14119;
																assign node14119 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node14122 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node14126 = (inp[10]) ? node14134 : node14127;
														assign node14127 = (inp[11]) ? node14131 : node14128;
															assign node14128 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node14131 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14134 = (inp[11]) ? node14138 : node14135;
															assign node14135 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node14138 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node14141 = (inp[3]) ? node14159 : node14142;
												assign node14142 = (inp[9]) ? node14152 : node14143;
													assign node14143 = (inp[11]) ? node14147 : node14144;
														assign node14144 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node14147 = (inp[2]) ? node14149 : 4'b1000;
															assign node14149 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node14152 = (inp[11]) ? 4'b1001 : node14153;
														assign node14153 = (inp[2]) ? node14155 : 4'b1000;
															assign node14155 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node14159 = (inp[11]) ? node14173 : node14160;
													assign node14160 = (inp[10]) ? node14168 : node14161;
														assign node14161 = (inp[9]) ? node14165 : node14162;
															assign node14162 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node14165 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14168 = (inp[2]) ? 4'b1001 : node14169;
															assign node14169 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node14173 = (inp[1]) ? node14179 : node14174;
														assign node14174 = (inp[9]) ? 4'b1001 : node14175;
															assign node14175 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14179 = (inp[9]) ? node14181 : 4'b1001;
															assign node14181 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node14184 = (inp[3]) ? node14232 : node14185;
											assign node14185 = (inp[1]) ? node14209 : node14186;
												assign node14186 = (inp[10]) ? node14198 : node14187;
													assign node14187 = (inp[2]) ? 4'b1100 : node14188;
														assign node14188 = (inp[0]) ? node14190 : 4'b1100;
															assign node14190 = (inp[9]) ? node14194 : node14191;
																assign node14191 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node14194 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node14198 = (inp[0]) ? 4'b1101 : node14199;
														assign node14199 = (inp[9]) ? node14201 : 4'b1101;
															assign node14201 = (inp[11]) ? node14205 : node14202;
																assign node14202 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node14205 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node14209 = (inp[0]) ? node14227 : node14210;
													assign node14210 = (inp[11]) ? node14220 : node14211;
														assign node14211 = (inp[10]) ? node14213 : 4'b1000;
															assign node14213 = (inp[2]) ? node14217 : node14214;
																assign node14214 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node14217 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14220 = (inp[2]) ? node14224 : node14221;
															assign node14221 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node14224 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node14227 = (inp[9]) ? node14229 : 4'b1001;
														assign node14229 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node14232 = (inp[11]) ? node14242 : node14233;
												assign node14233 = (inp[9]) ? node14237 : node14234;
													assign node14234 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node14237 = (inp[2]) ? node14239 : 4'b1000;
														assign node14239 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node14242 = (inp[9]) ? node14248 : node14243;
													assign node14243 = (inp[0]) ? node14245 : 4'b1000;
														assign node14245 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node14248 = (inp[2]) ? node14250 : 4'b1001;
														assign node14250 = (inp[0]) ? 4'b1000 : 4'b1001;
								assign node14253 = (inp[12]) ? node14445 : node14254;
									assign node14254 = (inp[4]) ? node14350 : node14255;
										assign node14255 = (inp[11]) ? node14313 : node14256;
											assign node14256 = (inp[0]) ? node14282 : node14257;
												assign node14257 = (inp[2]) ? node14269 : node14258;
													assign node14258 = (inp[3]) ? node14266 : node14259;
														assign node14259 = (inp[1]) ? node14263 : node14260;
															assign node14260 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node14263 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node14266 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node14269 = (inp[9]) ? node14277 : node14270;
														assign node14270 = (inp[1]) ? node14274 : node14271;
															assign node14271 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node14274 = (inp[3]) ? 4'b1001 : 4'b1100;
														assign node14277 = (inp[3]) ? 4'b1000 : node14278;
															assign node14278 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node14282 = (inp[10]) ? node14302 : node14283;
													assign node14283 = (inp[1]) ? node14295 : node14284;
														assign node14284 = (inp[3]) ? node14288 : node14285;
															assign node14285 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node14288 = (inp[9]) ? node14292 : node14289;
																assign node14289 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node14292 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14295 = (inp[3]) ? 4'b1000 : node14296;
															assign node14296 = (inp[9]) ? 4'b1100 : node14297;
																assign node14297 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node14302 = (inp[3]) ? node14306 : node14303;
														assign node14303 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node14306 = (inp[1]) ? node14308 : 4'b1100;
															assign node14308 = (inp[2]) ? node14310 : 4'b1000;
																assign node14310 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node14313 = (inp[9]) ? node14327 : node14314;
												assign node14314 = (inp[3]) ? node14318 : node14315;
													assign node14315 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node14318 = (inp[1]) ? node14324 : node14319;
														assign node14319 = (inp[0]) ? node14321 : 4'b1101;
															assign node14321 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14324 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node14327 = (inp[1]) ? node14339 : node14328;
													assign node14328 = (inp[3]) ? node14334 : node14329;
														assign node14329 = (inp[0]) ? 4'b1000 : node14330;
															assign node14330 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14334 = (inp[0]) ? node14336 : 4'b1100;
															assign node14336 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node14339 = (inp[3]) ? node14345 : node14340;
														assign node14340 = (inp[0]) ? node14342 : 4'b1100;
															assign node14342 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14345 = (inp[0]) ? node14347 : 4'b1001;
															assign node14347 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node14350 = (inp[3]) ? node14400 : node14351;
											assign node14351 = (inp[11]) ? node14379 : node14352;
												assign node14352 = (inp[10]) ? node14364 : node14353;
													assign node14353 = (inp[9]) ? node14359 : node14354;
														assign node14354 = (inp[0]) ? 4'b1100 : node14355;
															assign node14355 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14359 = (inp[0]) ? 4'b1101 : node14360;
															assign node14360 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node14364 = (inp[2]) ? node14372 : node14365;
														assign node14365 = (inp[1]) ? 4'b1100 : node14366;
															assign node14366 = (inp[9]) ? 4'b1100 : node14367;
																assign node14367 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node14372 = (inp[1]) ? node14374 : 4'b1100;
															assign node14374 = (inp[0]) ? 4'b1101 : node14375;
																assign node14375 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node14379 = (inp[1]) ? node14391 : node14380;
													assign node14380 = (inp[9]) ? node14386 : node14381;
														assign node14381 = (inp[0]) ? node14383 : 4'b1100;
															assign node14383 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node14386 = (inp[0]) ? node14388 : 4'b1101;
															assign node14388 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node14391 = (inp[2]) ? node14393 : 4'b1101;
														assign node14393 = (inp[0]) ? node14397 : node14394;
															assign node14394 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14397 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node14400 = (inp[1]) ? node14424 : node14401;
												assign node14401 = (inp[11]) ? node14413 : node14402;
													assign node14402 = (inp[9]) ? node14408 : node14403;
														assign node14403 = (inp[10]) ? node14405 : 4'b1000;
															assign node14405 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node14408 = (inp[2]) ? node14410 : 4'b1001;
															assign node14410 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node14413 = (inp[9]) ? node14419 : node14414;
														assign node14414 = (inp[2]) ? node14416 : 4'b1001;
															assign node14416 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14419 = (inp[0]) ? node14421 : 4'b1000;
															assign node14421 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node14424 = (inp[2]) ? node14438 : node14425;
													assign node14425 = (inp[9]) ? node14433 : node14426;
														assign node14426 = (inp[10]) ? node14430 : node14427;
															assign node14427 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14430 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14433 = (inp[11]) ? 4'b1101 : node14434;
															assign node14434 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node14438 = (inp[11]) ? node14442 : node14439;
														assign node14439 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node14442 = (inp[9]) ? 4'b1100 : 4'b1101;
									assign node14445 = (inp[4]) ? node14507 : node14446;
										assign node14446 = (inp[11]) ? node14478 : node14447;
											assign node14447 = (inp[9]) ? node14461 : node14448;
												assign node14448 = (inp[2]) ? node14454 : node14449;
													assign node14449 = (inp[1]) ? node14451 : 4'b1100;
														assign node14451 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node14454 = (inp[1]) ? 4'b1100 : node14455;
														assign node14455 = (inp[0]) ? 4'b1101 : node14456;
															assign node14456 = (inp[3]) ? 4'b1101 : 4'b1100;
												assign node14461 = (inp[2]) ? node14469 : node14462;
													assign node14462 = (inp[3]) ? 4'b1101 : node14463;
														assign node14463 = (inp[0]) ? 4'b1101 : node14464;
															assign node14464 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node14469 = (inp[3]) ? node14475 : node14470;
														assign node14470 = (inp[0]) ? node14472 : 4'b1101;
															assign node14472 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node14475 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node14478 = (inp[9]) ? node14494 : node14479;
												assign node14479 = (inp[0]) ? node14489 : node14480;
													assign node14480 = (inp[3]) ? node14486 : node14481;
														assign node14481 = (inp[2]) ? 4'b1101 : node14482;
															assign node14482 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node14486 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node14489 = (inp[1]) ? 4'b1101 : node14490;
														assign node14490 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node14494 = (inp[0]) ? node14502 : node14495;
													assign node14495 = (inp[2]) ? node14499 : node14496;
														assign node14496 = (inp[3]) ? 4'b1100 : 4'b1101;
														assign node14499 = (inp[3]) ? 4'b1101 : 4'b1100;
													assign node14502 = (inp[3]) ? 4'b1100 : node14503;
														assign node14503 = (inp[1]) ? 4'b1100 : 4'b1101;
										assign node14507 = (inp[3]) ? node14555 : node14508;
											assign node14508 = (inp[1]) ? node14526 : node14509;
												assign node14509 = (inp[11]) ? node14515 : node14510;
													assign node14510 = (inp[9]) ? 4'b1001 : node14511;
														assign node14511 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node14515 = (inp[9]) ? node14521 : node14516;
														assign node14516 = (inp[2]) ? 4'b1001 : node14517;
															assign node14517 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node14521 = (inp[0]) ? node14523 : 4'b1000;
															assign node14523 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node14526 = (inp[2]) ? node14542 : node14527;
													assign node14527 = (inp[0]) ? node14535 : node14528;
														assign node14528 = (inp[10]) ? 4'b1100 : node14529;
															assign node14529 = (inp[9]) ? node14531 : 4'b1100;
																assign node14531 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14535 = (inp[11]) ? node14539 : node14536;
															assign node14536 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14539 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node14542 = (inp[0]) ? node14548 : node14543;
														assign node14543 = (inp[11]) ? 4'b1100 : node14544;
															assign node14544 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14548 = (inp[10]) ? node14550 : 4'b1101;
															assign node14550 = (inp[11]) ? 4'b1101 : node14551;
																assign node14551 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node14555 = (inp[2]) ? node14577 : node14556;
												assign node14556 = (inp[0]) ? node14564 : node14557;
													assign node14557 = (inp[9]) ? node14561 : node14558;
														assign node14558 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14561 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node14564 = (inp[1]) ? node14570 : node14565;
														assign node14565 = (inp[11]) ? node14567 : 4'b1101;
															assign node14567 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14570 = (inp[9]) ? node14574 : node14571;
															assign node14571 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14574 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node14577 = (inp[1]) ? node14593 : node14578;
													assign node14578 = (inp[0]) ? node14586 : node14579;
														assign node14579 = (inp[11]) ? node14583 : node14580;
															assign node14580 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14583 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node14586 = (inp[11]) ? node14590 : node14587;
															assign node14587 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14590 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node14593 = (inp[10]) ? node14601 : node14594;
														assign node14594 = (inp[9]) ? node14598 : node14595;
															assign node14595 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14598 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14601 = (inp[11]) ? node14603 : 4'b1100;
															assign node14603 = (inp[0]) ? 4'b1101 : 4'b1100;
							assign node14606 = (inp[13]) ? node14958 : node14607;
								assign node14607 = (inp[1]) ? node14785 : node14608;
									assign node14608 = (inp[12]) ? node14696 : node14609;
										assign node14609 = (inp[9]) ? node14651 : node14610;
											assign node14610 = (inp[11]) ? node14630 : node14611;
												assign node14611 = (inp[4]) ? node14623 : node14612;
													assign node14612 = (inp[3]) ? node14618 : node14613;
														assign node14613 = (inp[0]) ? 4'b1000 : node14614;
															assign node14614 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14618 = (inp[10]) ? 4'b1101 : node14619;
															assign node14619 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node14623 = (inp[3]) ? 4'b1000 : node14624;
														assign node14624 = (inp[0]) ? 4'b1100 : node14625;
															assign node14625 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node14630 = (inp[2]) ? node14640 : node14631;
													assign node14631 = (inp[0]) ? 4'b1001 : node14632;
														assign node14632 = (inp[4]) ? node14636 : node14633;
															assign node14633 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node14636 = (inp[3]) ? 4'b1001 : 4'b1101;
													assign node14640 = (inp[3]) ? node14646 : node14641;
														assign node14641 = (inp[4]) ? node14643 : 4'b1001;
															assign node14643 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14646 = (inp[4]) ? node14648 : 4'b1100;
															assign node14648 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node14651 = (inp[4]) ? node14673 : node14652;
												assign node14652 = (inp[3]) ? node14662 : node14653;
													assign node14653 = (inp[11]) ? node14659 : node14654;
														assign node14654 = (inp[2]) ? 4'b1001 : node14655;
															assign node14655 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node14659 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node14662 = (inp[11]) ? node14668 : node14663;
														assign node14663 = (inp[2]) ? node14665 : 4'b1100;
															assign node14665 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node14668 = (inp[2]) ? node14670 : 4'b1101;
															assign node14670 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node14673 = (inp[3]) ? node14685 : node14674;
													assign node14674 = (inp[11]) ? node14680 : node14675;
														assign node14675 = (inp[10]) ? 4'b1101 : node14676;
															assign node14676 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14680 = (inp[2]) ? node14682 : 4'b1100;
															assign node14682 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node14685 = (inp[11]) ? node14691 : node14686;
														assign node14686 = (inp[0]) ? node14688 : 4'b1001;
															assign node14688 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14691 = (inp[0]) ? node14693 : 4'b1000;
															assign node14693 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node14696 = (inp[3]) ? node14734 : node14697;
											assign node14697 = (inp[4]) ? node14717 : node14698;
												assign node14698 = (inp[9]) ? node14710 : node14699;
													assign node14699 = (inp[11]) ? node14705 : node14700;
														assign node14700 = (inp[2]) ? node14702 : 4'b1100;
															assign node14702 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14705 = (inp[0]) ? node14707 : 4'b1101;
															assign node14707 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node14710 = (inp[11]) ? 4'b1100 : node14711;
														assign node14711 = (inp[0]) ? node14713 : 4'b1101;
															assign node14713 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node14717 = (inp[2]) ? node14725 : node14718;
													assign node14718 = (inp[9]) ? node14722 : node14719;
														assign node14719 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node14722 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14725 = (inp[9]) ? 4'b1001 : node14726;
														assign node14726 = (inp[11]) ? node14730 : node14727;
															assign node14727 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node14730 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node14734 = (inp[9]) ? node14756 : node14735;
												assign node14735 = (inp[11]) ? node14745 : node14736;
													assign node14736 = (inp[2]) ? 4'b1100 : node14737;
														assign node14737 = (inp[0]) ? node14741 : node14738;
															assign node14738 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node14741 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node14745 = (inp[2]) ? 4'b1101 : node14746;
														assign node14746 = (inp[10]) ? 4'b1100 : node14747;
															assign node14747 = (inp[0]) ? node14751 : node14748;
																assign node14748 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node14751 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node14756 = (inp[11]) ? node14774 : node14757;
													assign node14757 = (inp[2]) ? 4'b1101 : node14758;
														assign node14758 = (inp[10]) ? node14766 : node14759;
															assign node14759 = (inp[4]) ? node14763 : node14760;
																assign node14760 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node14763 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node14766 = (inp[0]) ? node14770 : node14767;
																assign node14767 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node14770 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node14774 = (inp[2]) ? 4'b1100 : node14775;
														assign node14775 = (inp[10]) ? 4'b1101 : node14776;
															assign node14776 = (inp[0]) ? node14780 : node14777;
																assign node14777 = (inp[4]) ? 4'b1101 : 4'b1100;
																assign node14780 = (inp[4]) ? 4'b1100 : 4'b1101;
									assign node14785 = (inp[12]) ? node14877 : node14786;
										assign node14786 = (inp[4]) ? node14830 : node14787;
											assign node14787 = (inp[3]) ? node14811 : node14788;
												assign node14788 = (inp[10]) ? node14798 : node14789;
													assign node14789 = (inp[0]) ? 4'b1101 : node14790;
														assign node14790 = (inp[11]) ? node14794 : node14791;
															assign node14791 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14794 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node14798 = (inp[2]) ? node14804 : node14799;
														assign node14799 = (inp[11]) ? node14801 : 4'b1100;
															assign node14801 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14804 = (inp[9]) ? node14806 : 4'b1100;
															assign node14806 = (inp[11]) ? 4'b1100 : node14807;
																assign node14807 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node14811 = (inp[9]) ? node14825 : node14812;
													assign node14812 = (inp[10]) ? 4'b1000 : node14813;
														assign node14813 = (inp[11]) ? node14819 : node14814;
															assign node14814 = (inp[2]) ? node14816 : 4'b1000;
																assign node14816 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node14819 = (inp[2]) ? node14821 : 4'b1001;
																assign node14821 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14825 = (inp[11]) ? node14827 : 4'b1001;
														assign node14827 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node14830 = (inp[2]) ? node14858 : node14831;
												assign node14831 = (inp[3]) ? node14849 : node14832;
													assign node14832 = (inp[0]) ? node14840 : node14833;
														assign node14833 = (inp[11]) ? node14837 : node14834;
															assign node14834 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node14837 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node14840 = (inp[10]) ? 4'b1101 : node14841;
															assign node14841 = (inp[9]) ? node14845 : node14842;
																assign node14842 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node14845 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node14849 = (inp[11]) ? 4'b1100 : node14850;
														assign node14850 = (inp[0]) ? node14854 : node14851;
															assign node14851 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node14854 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node14858 = (inp[10]) ? node14866 : node14859;
													assign node14859 = (inp[9]) ? node14863 : node14860;
														assign node14860 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14863 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node14866 = (inp[0]) ? node14872 : node14867;
														assign node14867 = (inp[9]) ? 4'b1100 : node14868;
															assign node14868 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14872 = (inp[9]) ? 4'b1101 : node14873;
															assign node14873 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node14877 = (inp[11]) ? node14915 : node14878;
											assign node14878 = (inp[9]) ? node14898 : node14879;
												assign node14879 = (inp[2]) ? 4'b1100 : node14880;
													assign node14880 = (inp[0]) ? node14890 : node14881;
														assign node14881 = (inp[10]) ? 4'b1100 : node14882;
															assign node14882 = (inp[3]) ? node14886 : node14883;
																assign node14883 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node14886 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node14890 = (inp[4]) ? node14894 : node14891;
															assign node14891 = (inp[3]) ? 4'b1101 : 4'b1100;
															assign node14894 = (inp[3]) ? 4'b1100 : 4'b1101;
												assign node14898 = (inp[2]) ? 4'b1101 : node14899;
													assign node14899 = (inp[0]) ? 4'b1101 : node14900;
														assign node14900 = (inp[10]) ? node14908 : node14901;
															assign node14901 = (inp[3]) ? node14905 : node14902;
																assign node14902 = (inp[4]) ? 4'b1101 : 4'b1100;
																assign node14905 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node14908 = (inp[3]) ? 4'b1101 : node14909;
																assign node14909 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node14915 = (inp[9]) ? node14935 : node14916;
												assign node14916 = (inp[2]) ? 4'b1101 : node14917;
													assign node14917 = (inp[0]) ? node14927 : node14918;
														assign node14918 = (inp[10]) ? node14920 : 4'b1100;
															assign node14920 = (inp[4]) ? node14924 : node14921;
																assign node14921 = (inp[3]) ? 4'b1101 : 4'b1100;
																assign node14924 = (inp[3]) ? 4'b1100 : 4'b1101;
														assign node14927 = (inp[3]) ? node14931 : node14928;
															assign node14928 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node14931 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node14935 = (inp[2]) ? 4'b1100 : node14936;
													assign node14936 = (inp[3]) ? node14944 : node14937;
														assign node14937 = (inp[4]) ? node14941 : node14938;
															assign node14938 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node14941 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node14944 = (inp[10]) ? node14950 : node14945;
															assign node14945 = (inp[4]) ? 4'b1100 : node14946;
																assign node14946 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node14950 = (inp[4]) ? node14954 : node14951;
																assign node14951 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node14954 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node14958 = (inp[12]) ? node15176 : node14959;
									assign node14959 = (inp[1]) ? node15065 : node14960;
										assign node14960 = (inp[9]) ? node15010 : node14961;
											assign node14961 = (inp[11]) ? node14983 : node14962;
												assign node14962 = (inp[0]) ? node14976 : node14963;
													assign node14963 = (inp[3]) ? node14969 : node14964;
														assign node14964 = (inp[4]) ? 4'b1001 : node14965;
															assign node14965 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node14969 = (inp[4]) ? node14973 : node14970;
															assign node14970 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node14973 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node14976 = (inp[3]) ? node14980 : node14977;
														assign node14977 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node14980 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node14983 = (inp[0]) ? node14997 : node14984;
													assign node14984 = (inp[2]) ? node14990 : node14985;
														assign node14985 = (inp[3]) ? node14987 : 4'b1101;
															assign node14987 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node14990 = (inp[3]) ? node14994 : node14991;
															assign node14991 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node14994 = (inp[4]) ? 4'b1100 : 4'b1001;
													assign node14997 = (inp[10]) ? node15005 : node14998;
														assign node14998 = (inp[2]) ? 4'b1100 : node14999;
															assign node14999 = (inp[4]) ? 4'b1100 : node15000;
																assign node15000 = (inp[3]) ? 4'b1000 : 4'b1100;
														assign node15005 = (inp[3]) ? 4'b1000 : node15006;
															assign node15006 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node15010 = (inp[11]) ? node15042 : node15011;
												assign node15011 = (inp[0]) ? node15027 : node15012;
													assign node15012 = (inp[10]) ? node15016 : node15013;
														assign node15013 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node15016 = (inp[3]) ? node15020 : node15017;
															assign node15017 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node15020 = (inp[4]) ? node15024 : node15021;
																assign node15021 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node15024 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node15027 = (inp[2]) ? node15035 : node15028;
														assign node15028 = (inp[4]) ? node15032 : node15029;
															assign node15029 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node15032 = (inp[3]) ? 4'b1100 : 4'b1001;
														assign node15035 = (inp[10]) ? node15037 : 4'b1000;
															assign node15037 = (inp[4]) ? 4'b1000 : node15038;
																assign node15038 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node15042 = (inp[0]) ? node15056 : node15043;
													assign node15043 = (inp[3]) ? node15049 : node15044;
														assign node15044 = (inp[4]) ? 4'b1001 : node15045;
															assign node15045 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15049 = (inp[4]) ? node15053 : node15050;
															assign node15050 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node15053 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node15056 = (inp[4]) ? node15060 : node15057;
														assign node15057 = (inp[3]) ? 4'b1001 : 4'b1101;
														assign node15060 = (inp[3]) ? 4'b1101 : node15061;
															assign node15061 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node15065 = (inp[3]) ? node15121 : node15066;
											assign node15066 = (inp[4]) ? node15092 : node15067;
												assign node15067 = (inp[2]) ? node15085 : node15068;
													assign node15068 = (inp[10]) ? node15076 : node15069;
														assign node15069 = (inp[11]) ? node15071 : 4'b1001;
															assign node15071 = (inp[9]) ? 4'b1000 : node15072;
																assign node15072 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15076 = (inp[11]) ? 4'b1001 : node15077;
															assign node15077 = (inp[9]) ? node15081 : node15078;
																assign node15078 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node15081 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15085 = (inp[11]) ? node15089 : node15086;
														assign node15086 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15089 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node15092 = (inp[2]) ? node15106 : node15093;
													assign node15093 = (inp[10]) ? node15099 : node15094;
														assign node15094 = (inp[11]) ? node15096 : 4'b1000;
															assign node15096 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node15099 = (inp[11]) ? node15103 : node15100;
															assign node15100 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15103 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15106 = (inp[10]) ? node15116 : node15107;
														assign node15107 = (inp[9]) ? 4'b1001 : node15108;
															assign node15108 = (inp[11]) ? node15112 : node15109;
																assign node15109 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node15112 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15116 = (inp[11]) ? node15118 : 4'b1000;
															assign node15118 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node15121 = (inp[4]) ? node15149 : node15122;
												assign node15122 = (inp[10]) ? node15132 : node15123;
													assign node15123 = (inp[2]) ? node15125 : 4'b1100;
														assign node15125 = (inp[11]) ? node15129 : node15126;
															assign node15126 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node15129 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node15132 = (inp[0]) ? node15140 : node15133;
														assign node15133 = (inp[2]) ? node15135 : 4'b1101;
															assign node15135 = (inp[9]) ? node15137 : 4'b1100;
																assign node15137 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node15140 = (inp[2]) ? node15142 : 4'b1100;
															assign node15142 = (inp[9]) ? node15146 : node15143;
																assign node15143 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node15146 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node15149 = (inp[2]) ? node15169 : node15150;
													assign node15150 = (inp[10]) ? node15164 : node15151;
														assign node15151 = (inp[9]) ? node15157 : node15152;
															assign node15152 = (inp[0]) ? node15154 : 4'b1000;
																assign node15154 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node15157 = (inp[0]) ? node15161 : node15158;
																assign node15158 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node15161 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node15164 = (inp[11]) ? 4'b1001 : node15165;
															assign node15165 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node15169 = (inp[9]) ? node15173 : node15170;
														assign node15170 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15173 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node15176 = (inp[4]) ? node15292 : node15177;
										assign node15177 = (inp[10]) ? node15235 : node15178;
											assign node15178 = (inp[3]) ? node15208 : node15179;
												assign node15179 = (inp[1]) ? node15195 : node15180;
													assign node15180 = (inp[11]) ? node15190 : node15181;
														assign node15181 = (inp[2]) ? node15187 : node15182;
															assign node15182 = (inp[9]) ? 4'b1000 : node15183;
																assign node15183 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15187 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15190 = (inp[9]) ? 4'b1000 : node15191;
															assign node15191 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15195 = (inp[9]) ? node15203 : node15196;
														assign node15196 = (inp[0]) ? node15198 : 4'b1001;
															assign node15198 = (inp[11]) ? node15200 : 4'b1000;
																assign node15200 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node15203 = (inp[11]) ? 4'b1001 : node15204;
															assign node15204 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node15208 = (inp[1]) ? node15224 : node15209;
													assign node15209 = (inp[0]) ? node15217 : node15210;
														assign node15210 = (inp[11]) ? node15214 : node15211;
															assign node15211 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15214 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node15217 = (inp[11]) ? node15219 : 4'b1000;
															assign node15219 = (inp[9]) ? 4'b1000 : node15220;
																assign node15220 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node15224 = (inp[0]) ? node15226 : 4'b1000;
														assign node15226 = (inp[11]) ? 4'b1000 : node15227;
															assign node15227 = (inp[9]) ? node15231 : node15228;
																assign node15228 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node15231 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node15235 = (inp[0]) ? node15259 : node15236;
												assign node15236 = (inp[11]) ? node15246 : node15237;
													assign node15237 = (inp[9]) ? node15241 : node15238;
														assign node15238 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node15241 = (inp[3]) ? 4'b1001 : node15242;
															assign node15242 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node15246 = (inp[9]) ? node15252 : node15247;
														assign node15247 = (inp[3]) ? 4'b1001 : node15248;
															assign node15248 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node15252 = (inp[3]) ? 4'b1000 : node15253;
															assign node15253 = (inp[2]) ? node15255 : 4'b1001;
																assign node15255 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node15259 = (inp[9]) ? node15275 : node15260;
													assign node15260 = (inp[1]) ? node15270 : node15261;
														assign node15261 = (inp[2]) ? node15267 : node15262;
															assign node15262 = (inp[3]) ? node15264 : 4'b1001;
																assign node15264 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node15267 = (inp[3]) ? 4'b1001 : 4'b1000;
														assign node15270 = (inp[11]) ? node15272 : 4'b1000;
															assign node15272 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node15275 = (inp[3]) ? node15287 : node15276;
														assign node15276 = (inp[11]) ? node15282 : node15277;
															assign node15277 = (inp[1]) ? node15279 : 4'b1001;
																assign node15279 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node15282 = (inp[2]) ? 4'b1000 : node15283;
																assign node15283 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node15287 = (inp[11]) ? 4'b1001 : node15288;
															assign node15288 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node15292 = (inp[3]) ? node15334 : node15293;
											assign node15293 = (inp[1]) ? node15313 : node15294;
												assign node15294 = (inp[0]) ? node15306 : node15295;
													assign node15295 = (inp[11]) ? node15301 : node15296;
														assign node15296 = (inp[9]) ? 4'b1101 : node15297;
															assign node15297 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node15301 = (inp[2]) ? 4'b1100 : node15302;
															assign node15302 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node15306 = (inp[9]) ? node15310 : node15307;
														assign node15307 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node15310 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node15313 = (inp[2]) ? node15321 : node15314;
													assign node15314 = (inp[11]) ? node15318 : node15315;
														assign node15315 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15318 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15321 = (inp[9]) ? node15323 : 4'b1000;
														assign node15323 = (inp[10]) ? node15329 : node15324;
															assign node15324 = (inp[11]) ? 4'b1000 : node15325;
																assign node15325 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node15329 = (inp[11]) ? node15331 : 4'b1000;
																assign node15331 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node15334 = (inp[2]) ? node15364 : node15335;
												assign node15335 = (inp[1]) ? node15357 : node15336;
													assign node15336 = (inp[11]) ? node15344 : node15337;
														assign node15337 = (inp[0]) ? node15341 : node15338;
															assign node15338 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node15341 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15344 = (inp[10]) ? node15350 : node15345;
															assign node15345 = (inp[0]) ? node15347 : 4'b1000;
																assign node15347 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node15350 = (inp[9]) ? node15354 : node15351;
																assign node15351 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node15354 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node15357 = (inp[11]) ? node15359 : 4'b1001;
														assign node15359 = (inp[9]) ? 4'b1001 : node15360;
															assign node15360 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node15364 = (inp[0]) ? node15372 : node15365;
													assign node15365 = (inp[11]) ? node15369 : node15366;
														assign node15366 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15369 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15372 = (inp[1]) ? node15384 : node15373;
														assign node15373 = (inp[10]) ? node15379 : node15374;
															assign node15374 = (inp[11]) ? node15376 : 4'b1001;
																assign node15376 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node15379 = (inp[9]) ? 4'b1001 : node15380;
																assign node15380 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15384 = (inp[11]) ? node15388 : node15385;
															assign node15385 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15388 = (inp[9]) ? 4'b1000 : 4'b1001;
			assign node15391 = (inp[6]) ? node23763 : node15392;
				assign node15392 = (inp[3]) ? node19608 : node15393;
					assign node15393 = (inp[12]) ? node17447 : node15394;
						assign node15394 = (inp[7]) ? node16390 : node15395;
							assign node15395 = (inp[4]) ? node15893 : node15396;
								assign node15396 = (inp[15]) ? node15658 : node15397;
									assign node15397 = (inp[5]) ? node15517 : node15398;
										assign node15398 = (inp[1]) ? node15456 : node15399;
											assign node15399 = (inp[9]) ? node15427 : node15400;
												assign node15400 = (inp[10]) ? node15412 : node15401;
													assign node15401 = (inp[11]) ? node15403 : 4'b1100;
														assign node15403 = (inp[13]) ? node15407 : node15404;
															assign node15404 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node15407 = (inp[2]) ? node15409 : 4'b1100;
																assign node15409 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15412 = (inp[11]) ? node15420 : node15413;
														assign node15413 = (inp[2]) ? node15415 : 4'b1101;
															assign node15415 = (inp[13]) ? 4'b1000 : node15416;
																assign node15416 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15420 = (inp[0]) ? 4'b1101 : node15421;
															assign node15421 = (inp[2]) ? 4'b1101 : node15422;
																assign node15422 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node15427 = (inp[13]) ? node15443 : node15428;
													assign node15428 = (inp[2]) ? node15434 : node15429;
														assign node15429 = (inp[10]) ? 4'b1000 : node15430;
															assign node15430 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node15434 = (inp[11]) ? 4'b1100 : node15435;
															assign node15435 = (inp[0]) ? node15439 : node15436;
																assign node15436 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node15439 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node15443 = (inp[2]) ? node15449 : node15444;
														assign node15444 = (inp[10]) ? node15446 : 4'b1101;
															assign node15446 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node15449 = (inp[10]) ? node15451 : 4'b1000;
															assign node15451 = (inp[11]) ? node15453 : 4'b1001;
																assign node15453 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node15456 = (inp[10]) ? node15482 : node15457;
												assign node15457 = (inp[9]) ? node15467 : node15458;
													assign node15458 = (inp[13]) ? node15464 : node15459;
														assign node15459 = (inp[2]) ? 4'b1100 : node15460;
															assign node15460 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15464 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node15467 = (inp[13]) ? node15475 : node15468;
														assign node15468 = (inp[2]) ? node15472 : node15469;
															assign node15469 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node15472 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15475 = (inp[2]) ? 4'b1001 : node15476;
															assign node15476 = (inp[0]) ? 4'b1101 : node15477;
																assign node15477 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node15482 = (inp[9]) ? node15500 : node15483;
													assign node15483 = (inp[13]) ? node15491 : node15484;
														assign node15484 = (inp[2]) ? node15486 : 4'b1001;
															assign node15486 = (inp[0]) ? node15488 : 4'b1101;
																assign node15488 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node15491 = (inp[2]) ? node15497 : node15492;
															assign node15492 = (inp[0]) ? 4'b1101 : node15493;
																assign node15493 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node15497 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node15500 = (inp[2]) ? node15510 : node15501;
														assign node15501 = (inp[13]) ? node15507 : node15502;
															assign node15502 = (inp[0]) ? 4'b1000 : node15503;
																assign node15503 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node15507 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15510 = (inp[13]) ? node15514 : node15511;
															assign node15511 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node15514 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node15517 = (inp[13]) ? node15587 : node15518;
											assign node15518 = (inp[1]) ? node15558 : node15519;
												assign node15519 = (inp[2]) ? node15537 : node15520;
													assign node15520 = (inp[10]) ? node15530 : node15521;
														assign node15521 = (inp[9]) ? node15525 : node15522;
															assign node15522 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node15525 = (inp[11]) ? node15527 : 4'b1101;
																assign node15527 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node15530 = (inp[9]) ? 4'b1100 : node15531;
															assign node15531 = (inp[11]) ? node15533 : 4'b1101;
																assign node15533 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node15537 = (inp[0]) ? node15547 : node15538;
														assign node15538 = (inp[10]) ? 4'b1000 : node15539;
															assign node15539 = (inp[11]) ? node15543 : node15540;
																assign node15540 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node15543 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node15547 = (inp[11]) ? node15553 : node15548;
															assign node15548 = (inp[10]) ? node15550 : 4'b1001;
																assign node15550 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node15553 = (inp[10]) ? 4'b1001 : node15554;
																assign node15554 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node15558 = (inp[2]) ? node15576 : node15559;
													assign node15559 = (inp[9]) ? node15567 : node15560;
														assign node15560 = (inp[10]) ? node15562 : 4'b1000;
															assign node15562 = (inp[0]) ? node15564 : 4'b1001;
																assign node15564 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15567 = (inp[10]) ? node15573 : node15568;
															assign node15568 = (inp[0]) ? node15570 : 4'b1001;
																assign node15570 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node15573 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15576 = (inp[9]) ? node15582 : node15577;
														assign node15577 = (inp[11]) ? 4'b1101 : node15578;
															assign node15578 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node15582 = (inp[0]) ? 4'b1100 : node15583;
															assign node15583 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node15587 = (inp[9]) ? node15619 : node15588;
												assign node15588 = (inp[2]) ? node15600 : node15589;
													assign node15589 = (inp[1]) ? node15595 : node15590;
														assign node15590 = (inp[10]) ? 4'b1001 : node15591;
															assign node15591 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15595 = (inp[10]) ? 4'b1101 : node15596;
															assign node15596 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node15600 = (inp[1]) ? node15612 : node15601;
														assign node15601 = (inp[10]) ? node15607 : node15602;
															assign node15602 = (inp[11]) ? node15604 : 4'b1101;
																assign node15604 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node15607 = (inp[0]) ? 4'b1100 : node15608;
																assign node15608 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node15612 = (inp[10]) ? node15616 : node15613;
															assign node15613 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15616 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node15619 = (inp[0]) ? node15637 : node15620;
													assign node15620 = (inp[11]) ? node15628 : node15621;
														assign node15621 = (inp[1]) ? node15625 : node15622;
															assign node15622 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node15625 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node15628 = (inp[10]) ? node15630 : 4'b1001;
															assign node15630 = (inp[2]) ? node15634 : node15631;
																assign node15631 = (inp[1]) ? 4'b1100 : 4'b1000;
																assign node15634 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node15637 = (inp[10]) ? node15649 : node15638;
														assign node15638 = (inp[11]) ? node15644 : node15639;
															assign node15639 = (inp[1]) ? 4'b1100 : node15640;
																assign node15640 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node15644 = (inp[2]) ? node15646 : 4'b1001;
																assign node15646 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node15649 = (inp[1]) ? node15653 : node15650;
															assign node15650 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node15653 = (inp[2]) ? node15655 : 4'b1101;
																assign node15655 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node15658 = (inp[9]) ? node15762 : node15659;
										assign node15659 = (inp[13]) ? node15709 : node15660;
											assign node15660 = (inp[2]) ? node15682 : node15661;
												assign node15661 = (inp[5]) ? node15675 : node15662;
													assign node15662 = (inp[10]) ? node15668 : node15663;
														assign node15663 = (inp[0]) ? 4'b1010 : node15664;
															assign node15664 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node15668 = (inp[11]) ? 4'b1011 : node15669;
															assign node15669 = (inp[0]) ? node15671 : 4'b1011;
																assign node15671 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node15675 = (inp[1]) ? node15679 : node15676;
														assign node15676 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15679 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node15682 = (inp[5]) ? node15698 : node15683;
													assign node15683 = (inp[11]) ? node15687 : node15684;
														assign node15684 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node15687 = (inp[10]) ? node15693 : node15688;
															assign node15688 = (inp[1]) ? node15690 : 4'b1110;
																assign node15690 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node15693 = (inp[1]) ? node15695 : 4'b1111;
																assign node15695 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node15698 = (inp[1]) ? node15704 : node15699;
														assign node15699 = (inp[10]) ? node15701 : 4'b1011;
															assign node15701 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node15704 = (inp[10]) ? 4'b1110 : node15705;
															assign node15705 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node15709 = (inp[2]) ? node15735 : node15710;
												assign node15710 = (inp[5]) ? node15722 : node15711;
													assign node15711 = (inp[10]) ? node15713 : 4'b1111;
														assign node15713 = (inp[1]) ? node15717 : node15714;
															assign node15714 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15717 = (inp[11]) ? 4'b1110 : node15718;
																assign node15718 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node15722 = (inp[1]) ? node15730 : node15723;
														assign node15723 = (inp[11]) ? 4'b1010 : node15724;
															assign node15724 = (inp[10]) ? node15726 : 4'b1011;
																assign node15726 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node15730 = (inp[0]) ? 4'b1110 : node15731;
															assign node15731 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node15735 = (inp[1]) ? node15747 : node15736;
													assign node15736 = (inp[5]) ? node15742 : node15737;
														assign node15737 = (inp[10]) ? node15739 : 4'b1010;
															assign node15739 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node15742 = (inp[0]) ? 4'b1110 : node15743;
															assign node15743 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node15747 = (inp[10]) ? node15755 : node15748;
														assign node15748 = (inp[11]) ? 4'b1010 : node15749;
															assign node15749 = (inp[5]) ? 4'b1011 : node15750;
																assign node15750 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node15755 = (inp[0]) ? node15757 : 4'b1011;
															assign node15757 = (inp[11]) ? node15759 : 4'b1010;
																assign node15759 = (inp[5]) ? 4'b1010 : 4'b1011;
										assign node15762 = (inp[1]) ? node15826 : node15763;
											assign node15763 = (inp[10]) ? node15797 : node15764;
												assign node15764 = (inp[2]) ? node15780 : node15765;
													assign node15765 = (inp[13]) ? node15773 : node15766;
														assign node15766 = (inp[5]) ? node15770 : node15767;
															assign node15767 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node15770 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15773 = (inp[5]) ? node15775 : 4'b1110;
															assign node15775 = (inp[0]) ? node15777 : 4'b1010;
																assign node15777 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node15780 = (inp[13]) ? node15792 : node15781;
														assign node15781 = (inp[5]) ? node15787 : node15782;
															assign node15782 = (inp[0]) ? node15784 : 4'b1111;
																assign node15784 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15787 = (inp[11]) ? node15789 : 4'b1010;
																assign node15789 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node15792 = (inp[5]) ? node15794 : 4'b1011;
															assign node15794 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node15797 = (inp[2]) ? node15811 : node15798;
													assign node15798 = (inp[13]) ? node15804 : node15799;
														assign node15799 = (inp[11]) ? node15801 : 4'b1110;
															assign node15801 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node15804 = (inp[5]) ? 4'b1011 : node15805;
															assign node15805 = (inp[0]) ? 4'b1111 : node15806;
																assign node15806 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node15811 = (inp[13]) ? node15819 : node15812;
														assign node15812 = (inp[5]) ? 4'b1010 : node15813;
															assign node15813 = (inp[0]) ? node15815 : 4'b1110;
																assign node15815 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node15819 = (inp[5]) ? 4'b1110 : node15820;
															assign node15820 = (inp[11]) ? node15822 : 4'b1010;
																assign node15822 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node15826 = (inp[10]) ? node15856 : node15827;
												assign node15827 = (inp[2]) ? node15847 : node15828;
													assign node15828 = (inp[13]) ? node15840 : node15829;
														assign node15829 = (inp[5]) ? node15835 : node15830;
															assign node15830 = (inp[0]) ? node15832 : 4'b1011;
																assign node15832 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node15835 = (inp[11]) ? node15837 : 4'b1010;
																assign node15837 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node15840 = (inp[11]) ? 4'b1110 : node15841;
															assign node15841 = (inp[0]) ? 4'b1111 : node15842;
																assign node15842 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node15847 = (inp[13]) ? node15849 : 4'b1110;
														assign node15849 = (inp[11]) ? node15851 : 4'b1010;
															assign node15851 = (inp[5]) ? node15853 : 4'b1011;
																assign node15853 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node15856 = (inp[0]) ? node15876 : node15857;
													assign node15857 = (inp[5]) ? node15865 : node15858;
														assign node15858 = (inp[13]) ? node15862 : node15859;
															assign node15859 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node15862 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node15865 = (inp[2]) ? node15871 : node15866;
															assign node15866 = (inp[13]) ? node15868 : 4'b1010;
																assign node15868 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15871 = (inp[13]) ? node15873 : 4'b1111;
																assign node15873 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node15876 = (inp[2]) ? node15886 : node15877;
														assign node15877 = (inp[13]) ? node15883 : node15878;
															assign node15878 = (inp[5]) ? 4'b1011 : node15879;
																assign node15879 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node15883 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node15886 = (inp[13]) ? node15888 : 4'b1111;
															assign node15888 = (inp[5]) ? 4'b1011 : node15889;
																assign node15889 = (inp[11]) ? 4'b1010 : 4'b1011;
								assign node15893 = (inp[2]) ? node16141 : node15894;
									assign node15894 = (inp[5]) ? node16012 : node15895;
										assign node15895 = (inp[10]) ? node15947 : node15896;
											assign node15896 = (inp[9]) ? node15926 : node15897;
												assign node15897 = (inp[0]) ? node15915 : node15898;
													assign node15898 = (inp[11]) ? node15908 : node15899;
														assign node15899 = (inp[1]) ? 4'b1100 : node15900;
															assign node15900 = (inp[13]) ? node15904 : node15901;
																assign node15901 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node15904 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node15908 = (inp[13]) ? node15912 : node15909;
															assign node15909 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node15912 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node15915 = (inp[15]) ? node15919 : node15916;
														assign node15916 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node15919 = (inp[13]) ? 4'b1000 : node15920;
															assign node15920 = (inp[1]) ? node15922 : 4'b1100;
																assign node15922 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node15926 = (inp[0]) ? node15936 : node15927;
													assign node15927 = (inp[11]) ? node15931 : node15928;
														assign node15928 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node15931 = (inp[15]) ? 4'b1100 : node15932;
															assign node15932 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node15936 = (inp[15]) ? node15940 : node15937;
														assign node15937 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node15940 = (inp[13]) ? node15944 : node15941;
															assign node15941 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node15944 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node15947 = (inp[9]) ? node15983 : node15948;
												assign node15948 = (inp[0]) ? node15968 : node15949;
													assign node15949 = (inp[11]) ? node15959 : node15950;
														assign node15950 = (inp[1]) ? node15954 : node15951;
															assign node15951 = (inp[13]) ? 4'b1000 : 4'b1101;
															assign node15954 = (inp[13]) ? node15956 : 4'b1001;
																assign node15956 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node15959 = (inp[15]) ? node15963 : node15960;
															assign node15960 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node15963 = (inp[13]) ? 4'b1000 : node15964;
																assign node15964 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node15968 = (inp[15]) ? node15972 : node15969;
														assign node15969 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node15972 = (inp[13]) ? node15978 : node15973;
															assign node15973 = (inp[11]) ? 4'b1101 : node15974;
																assign node15974 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node15978 = (inp[1]) ? 4'b1001 : node15979;
																assign node15979 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node15983 = (inp[11]) ? node15997 : node15984;
													assign node15984 = (inp[1]) ? node15990 : node15985;
														assign node15985 = (inp[13]) ? 4'b1100 : node15986;
															assign node15986 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node15990 = (inp[13]) ? node15994 : node15991;
															assign node15991 = (inp[15]) ? 4'b1101 : 4'b1000;
															assign node15994 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node15997 = (inp[0]) ? node16005 : node15998;
														assign node15998 = (inp[13]) ? node16002 : node15999;
															assign node15999 = (inp[15]) ? 4'b1100 : 4'b1001;
															assign node16002 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node16005 = (inp[15]) ? node16009 : node16006;
															assign node16006 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node16009 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node16012 = (inp[13]) ? node16092 : node16013;
											assign node16013 = (inp[9]) ? node16059 : node16014;
												assign node16014 = (inp[0]) ? node16036 : node16015;
													assign node16015 = (inp[1]) ? node16027 : node16016;
														assign node16016 = (inp[15]) ? node16020 : node16017;
															assign node16017 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node16020 = (inp[11]) ? node16024 : node16021;
																assign node16021 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node16024 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node16027 = (inp[15]) ? node16033 : node16028;
															assign node16028 = (inp[11]) ? node16030 : 4'b1000;
																assign node16030 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node16033 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node16036 = (inp[10]) ? node16048 : node16037;
														assign node16037 = (inp[11]) ? node16041 : node16038;
															assign node16038 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node16041 = (inp[15]) ? node16045 : node16042;
																assign node16042 = (inp[1]) ? 4'b1001 : 4'b1100;
																assign node16045 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node16048 = (inp[15]) ? node16054 : node16049;
															assign node16049 = (inp[1]) ? 4'b1000 : node16050;
																assign node16050 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node16054 = (inp[1]) ? node16056 : 4'b1000;
																assign node16056 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node16059 = (inp[11]) ? node16079 : node16060;
													assign node16060 = (inp[10]) ? node16068 : node16061;
														assign node16061 = (inp[0]) ? node16065 : node16062;
															assign node16062 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node16065 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node16068 = (inp[1]) ? node16074 : node16069;
															assign node16069 = (inp[15]) ? 4'b1001 : node16070;
																assign node16070 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node16074 = (inp[15]) ? node16076 : 4'b1001;
																assign node16076 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node16079 = (inp[1]) ? node16085 : node16080;
														assign node16080 = (inp[15]) ? 4'b1000 : node16081;
															assign node16081 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node16085 = (inp[15]) ? 4'b1100 : node16086;
															assign node16086 = (inp[0]) ? 4'b1000 : node16087;
																assign node16087 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node16092 = (inp[1]) ? node16116 : node16093;
												assign node16093 = (inp[15]) ? node16109 : node16094;
													assign node16094 = (inp[0]) ? node16102 : node16095;
														assign node16095 = (inp[10]) ? 4'b1000 : node16096;
															assign node16096 = (inp[11]) ? 4'b1000 : node16097;
																assign node16097 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node16102 = (inp[9]) ? node16106 : node16103;
															assign node16103 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node16106 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node16109 = (inp[11]) ? node16111 : 4'b1100;
														assign node16111 = (inp[10]) ? 4'b1100 : node16112;
															assign node16112 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node16116 = (inp[15]) ? node16128 : node16117;
													assign node16117 = (inp[9]) ? node16121 : node16118;
														assign node16118 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node16121 = (inp[10]) ? node16123 : 4'b1100;
															assign node16123 = (inp[0]) ? 4'b1101 : node16124;
																assign node16124 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16128 = (inp[11]) ? node16136 : node16129;
														assign node16129 = (inp[0]) ? node16131 : 4'b1000;
															assign node16131 = (inp[10]) ? node16133 : 4'b1000;
																assign node16133 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node16136 = (inp[0]) ? 4'b1001 : node16137;
															assign node16137 = (inp[10]) ? 4'b1000 : 4'b1001;
									assign node16141 = (inp[15]) ? node16253 : node16142;
										assign node16142 = (inp[13]) ? node16204 : node16143;
											assign node16143 = (inp[1]) ? node16175 : node16144;
												assign node16144 = (inp[5]) ? node16162 : node16145;
													assign node16145 = (inp[11]) ? node16157 : node16146;
														assign node16146 = (inp[10]) ? node16152 : node16147;
															assign node16147 = (inp[9]) ? 4'b1101 : node16148;
																assign node16148 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node16152 = (inp[9]) ? 4'b1100 : node16153;
																assign node16153 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node16157 = (inp[10]) ? 4'b1101 : node16158;
															assign node16158 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node16162 = (inp[10]) ? node16168 : node16163;
														assign node16163 = (inp[9]) ? 4'b1001 : node16164;
															assign node16164 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node16168 = (inp[9]) ? 4'b1000 : node16169;
															assign node16169 = (inp[11]) ? 4'b1001 : node16170;
																assign node16170 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node16175 = (inp[11]) ? node16195 : node16176;
													assign node16176 = (inp[10]) ? node16190 : node16177;
														assign node16177 = (inp[9]) ? node16183 : node16178;
															assign node16178 = (inp[5]) ? 4'b1100 : node16179;
																assign node16179 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node16183 = (inp[0]) ? node16187 : node16184;
																assign node16184 = (inp[5]) ? 4'b1101 : 4'b1100;
																assign node16187 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node16190 = (inp[0]) ? node16192 : 4'b1101;
															assign node16192 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node16195 = (inp[10]) ? node16197 : 4'b1101;
														assign node16197 = (inp[5]) ? node16201 : node16198;
															assign node16198 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node16201 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node16204 = (inp[5]) ? node16230 : node16205;
												assign node16205 = (inp[11]) ? node16223 : node16206;
													assign node16206 = (inp[1]) ? node16214 : node16207;
														assign node16207 = (inp[9]) ? node16211 : node16208;
															assign node16208 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node16211 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node16214 = (inp[0]) ? 4'b1000 : node16215;
															assign node16215 = (inp[10]) ? node16219 : node16216;
																assign node16216 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node16219 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node16223 = (inp[1]) ? 4'b1001 : node16224;
														assign node16224 = (inp[9]) ? 4'b1001 : node16225;
															assign node16225 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node16230 = (inp[1]) ? node16248 : node16231;
													assign node16231 = (inp[10]) ? node16243 : node16232;
														assign node16232 = (inp[9]) ? node16238 : node16233;
															assign node16233 = (inp[11]) ? 4'b1100 : node16234;
																assign node16234 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node16238 = (inp[11]) ? 4'b1101 : node16239;
																assign node16239 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node16243 = (inp[9]) ? node16245 : 4'b1101;
															assign node16245 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16248 = (inp[0]) ? node16250 : 4'b1000;
														assign node16250 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node16253 = (inp[13]) ? node16331 : node16254;
											assign node16254 = (inp[5]) ? node16288 : node16255;
												assign node16255 = (inp[9]) ? node16279 : node16256;
													assign node16256 = (inp[10]) ? node16268 : node16257;
														assign node16257 = (inp[11]) ? node16263 : node16258;
															assign node16258 = (inp[1]) ? node16260 : 4'b1000;
																assign node16260 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node16263 = (inp[0]) ? 4'b1000 : node16264;
																assign node16264 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node16268 = (inp[0]) ? node16274 : node16269;
															assign node16269 = (inp[1]) ? 4'b1001 : node16270;
																assign node16270 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16274 = (inp[1]) ? node16276 : 4'b1001;
																assign node16276 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16279 = (inp[10]) ? 4'b1000 : node16280;
														assign node16280 = (inp[1]) ? 4'b1000 : node16281;
															assign node16281 = (inp[11]) ? node16283 : 4'b1001;
																assign node16283 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node16288 = (inp[1]) ? node16308 : node16289;
													assign node16289 = (inp[10]) ? node16299 : node16290;
														assign node16290 = (inp[11]) ? 4'b1101 : node16291;
															assign node16291 = (inp[0]) ? node16295 : node16292;
																assign node16292 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node16295 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node16299 = (inp[11]) ? node16305 : node16300;
															assign node16300 = (inp[0]) ? node16302 : 4'b1101;
																assign node16302 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node16305 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node16308 = (inp[0]) ? node16316 : node16309;
														assign node16309 = (inp[10]) ? node16313 : node16310;
															assign node16310 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node16313 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node16316 = (inp[9]) ? node16324 : node16317;
															assign node16317 = (inp[10]) ? node16321 : node16318;
																assign node16318 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node16321 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16324 = (inp[10]) ? node16328 : node16325;
																assign node16325 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node16328 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node16331 = (inp[1]) ? node16359 : node16332;
												assign node16332 = (inp[5]) ? node16346 : node16333;
													assign node16333 = (inp[11]) ? 4'b1101 : node16334;
														assign node16334 = (inp[0]) ? node16340 : node16335;
															assign node16335 = (inp[10]) ? node16337 : 4'b1101;
																assign node16337 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node16340 = (inp[10]) ? node16342 : 4'b1100;
																assign node16342 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node16346 = (inp[10]) ? node16354 : node16347;
														assign node16347 = (inp[11]) ? node16349 : 4'b1001;
															assign node16349 = (inp[0]) ? 4'b1001 : node16350;
																assign node16350 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node16354 = (inp[9]) ? 4'b1000 : node16355;
															assign node16355 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node16359 = (inp[5]) ? node16375 : node16360;
													assign node16360 = (inp[9]) ? node16370 : node16361;
														assign node16361 = (inp[10]) ? node16367 : node16362;
															assign node16362 = (inp[11]) ? 4'b1101 : node16363;
																assign node16363 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node16367 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node16370 = (inp[10]) ? 4'b1101 : node16371;
															assign node16371 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16375 = (inp[0]) ? node16381 : node16376;
														assign node16376 = (inp[10]) ? node16378 : 4'b1101;
															assign node16378 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node16381 = (inp[10]) ? node16383 : 4'b1100;
															assign node16383 = (inp[9]) ? node16387 : node16384;
																assign node16384 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node16387 = (inp[11]) ? 4'b1100 : 4'b1101;
							assign node16390 = (inp[4]) ? node16888 : node16391;
								assign node16391 = (inp[15]) ? node16661 : node16392;
									assign node16392 = (inp[1]) ? node16532 : node16393;
										assign node16393 = (inp[2]) ? node16467 : node16394;
											assign node16394 = (inp[10]) ? node16432 : node16395;
												assign node16395 = (inp[13]) ? node16411 : node16396;
													assign node16396 = (inp[5]) ? node16406 : node16397;
														assign node16397 = (inp[9]) ? node16403 : node16398;
															assign node16398 = (inp[11]) ? node16400 : 4'b1010;
																assign node16400 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node16403 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node16406 = (inp[0]) ? node16408 : 4'b1111;
															assign node16408 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node16411 = (inp[5]) ? node16423 : node16412;
														assign node16412 = (inp[9]) ? node16418 : node16413;
															assign node16413 = (inp[11]) ? node16415 : 4'b1110;
																assign node16415 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node16418 = (inp[0]) ? 4'b1111 : node16419;
																assign node16419 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node16423 = (inp[9]) ? node16429 : node16424;
															assign node16424 = (inp[11]) ? 4'b1011 : node16425;
																assign node16425 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node16429 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node16432 = (inp[0]) ? node16454 : node16433;
													assign node16433 = (inp[11]) ? node16443 : node16434;
														assign node16434 = (inp[9]) ? node16440 : node16435;
															assign node16435 = (inp[5]) ? 4'b1010 : node16436;
																assign node16436 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node16440 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node16443 = (inp[5]) ? node16447 : node16444;
															assign node16444 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node16447 = (inp[13]) ? node16451 : node16448;
																assign node16448 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node16451 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node16454 = (inp[9]) ? node16462 : node16455;
														assign node16455 = (inp[5]) ? node16459 : node16456;
															assign node16456 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node16459 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node16462 = (inp[11]) ? node16464 : 4'b1010;
															assign node16464 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node16467 = (inp[10]) ? node16499 : node16468;
												assign node16468 = (inp[9]) ? node16482 : node16469;
													assign node16469 = (inp[13]) ? node16477 : node16470;
														assign node16470 = (inp[5]) ? node16472 : 4'b1110;
															assign node16472 = (inp[0]) ? 4'b1010 : node16473;
																assign node16473 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16477 = (inp[5]) ? node16479 : 4'b1011;
															assign node16479 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node16482 = (inp[5]) ? node16494 : node16483;
														assign node16483 = (inp[13]) ? node16489 : node16484;
															assign node16484 = (inp[0]) ? node16486 : 4'b1111;
																assign node16486 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node16489 = (inp[0]) ? 4'b1010 : node16490;
																assign node16490 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16494 = (inp[13]) ? 4'b1111 : node16495;
															assign node16495 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node16499 = (inp[9]) ? node16517 : node16500;
													assign node16500 = (inp[5]) ? node16510 : node16501;
														assign node16501 = (inp[13]) ? node16505 : node16502;
															assign node16502 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node16505 = (inp[11]) ? node16507 : 4'b1010;
																assign node16507 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16510 = (inp[13]) ? node16512 : 4'b1011;
															assign node16512 = (inp[11]) ? node16514 : 4'b1111;
																assign node16514 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node16517 = (inp[0]) ? node16527 : node16518;
														assign node16518 = (inp[5]) ? node16522 : node16519;
															assign node16519 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node16522 = (inp[13]) ? 4'b1111 : node16523;
																assign node16523 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16527 = (inp[5]) ? 4'b1110 : node16528;
															assign node16528 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node16532 = (inp[5]) ? node16600 : node16533;
											assign node16533 = (inp[13]) ? node16571 : node16534;
												assign node16534 = (inp[2]) ? node16550 : node16535;
													assign node16535 = (inp[9]) ? node16541 : node16536;
														assign node16536 = (inp[10]) ? 4'b1011 : node16537;
															assign node16537 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16541 = (inp[11]) ? node16543 : 4'b1010;
															assign node16543 = (inp[0]) ? node16547 : node16544;
																assign node16544 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node16547 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node16550 = (inp[10]) ? node16562 : node16551;
														assign node16551 = (inp[9]) ? node16557 : node16552;
															assign node16552 = (inp[0]) ? node16554 : 4'b1110;
																assign node16554 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node16557 = (inp[0]) ? node16559 : 4'b1111;
																assign node16559 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node16562 = (inp[9]) ? node16566 : node16563;
															assign node16563 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node16566 = (inp[0]) ? node16568 : 4'b1110;
																assign node16568 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node16571 = (inp[2]) ? node16585 : node16572;
													assign node16572 = (inp[11]) ? node16576 : node16573;
														assign node16573 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node16576 = (inp[9]) ? 4'b1111 : node16577;
															assign node16577 = (inp[0]) ? node16581 : node16578;
																assign node16578 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node16581 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node16585 = (inp[10]) ? node16591 : node16586;
														assign node16586 = (inp[9]) ? node16588 : 4'b1011;
															assign node16588 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16591 = (inp[0]) ? 4'b1010 : node16592;
															assign node16592 = (inp[11]) ? node16596 : node16593;
																assign node16593 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node16596 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node16600 = (inp[9]) ? node16630 : node16601;
												assign node16601 = (inp[11]) ? node16617 : node16602;
													assign node16602 = (inp[0]) ? node16610 : node16603;
														assign node16603 = (inp[2]) ? node16607 : node16604;
															assign node16604 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node16607 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node16610 = (inp[10]) ? 4'b1010 : node16611;
															assign node16611 = (inp[2]) ? 4'b1110 : node16612;
																assign node16612 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node16617 = (inp[10]) ? node16625 : node16618;
														assign node16618 = (inp[2]) ? node16622 : node16619;
															assign node16619 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node16622 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node16625 = (inp[13]) ? 4'b1110 : node16626;
															assign node16626 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node16630 = (inp[10]) ? node16644 : node16631;
													assign node16631 = (inp[11]) ? node16639 : node16632;
														assign node16632 = (inp[2]) ? node16636 : node16633;
															assign node16633 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node16636 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16639 = (inp[0]) ? node16641 : 4'b1110;
															assign node16641 = (inp[2]) ? 4'b1111 : 4'b1010;
													assign node16644 = (inp[11]) ? node16656 : node16645;
														assign node16645 = (inp[13]) ? node16649 : node16646;
															assign node16646 = (inp[0]) ? 4'b1010 : 4'b1110;
															assign node16649 = (inp[2]) ? node16653 : node16650;
																assign node16650 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node16653 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node16656 = (inp[2]) ? 4'b1110 : node16657;
															assign node16657 = (inp[13]) ? 4'b1111 : 4'b1011;
									assign node16661 = (inp[0]) ? node16783 : node16662;
										assign node16662 = (inp[5]) ? node16730 : node16663;
											assign node16663 = (inp[10]) ? node16695 : node16664;
												assign node16664 = (inp[9]) ? node16680 : node16665;
													assign node16665 = (inp[1]) ? node16673 : node16666;
														assign node16666 = (inp[13]) ? 4'b1001 : node16667;
															assign node16667 = (inp[2]) ? node16669 : 4'b1100;
																assign node16669 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node16673 = (inp[11]) ? 4'b1101 : node16674;
															assign node16674 = (inp[2]) ? 4'b1001 : node16675;
																assign node16675 = (inp[13]) ? 4'b1100 : 4'b1001;
													assign node16680 = (inp[1]) ? node16682 : 4'b1000;
														assign node16682 = (inp[13]) ? node16688 : node16683;
															assign node16683 = (inp[2]) ? 4'b1100 : node16684;
																assign node16684 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node16688 = (inp[2]) ? node16692 : node16689;
																assign node16689 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node16692 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node16695 = (inp[13]) ? node16705 : node16696;
													assign node16696 = (inp[11]) ? 4'b1000 : node16697;
														assign node16697 = (inp[9]) ? node16701 : node16698;
															assign node16698 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node16701 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node16705 = (inp[9]) ? node16719 : node16706;
														assign node16706 = (inp[2]) ? node16712 : node16707;
															assign node16707 = (inp[1]) ? node16709 : 4'b1000;
																assign node16709 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node16712 = (inp[1]) ? node16716 : node16713;
																assign node16713 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node16716 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node16719 = (inp[2]) ? node16725 : node16720;
															assign node16720 = (inp[1]) ? node16722 : 4'b1001;
																assign node16722 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node16725 = (inp[1]) ? 4'b1000 : node16726;
																assign node16726 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node16730 = (inp[2]) ? node16750 : node16731;
												assign node16731 = (inp[13]) ? node16743 : node16732;
													assign node16732 = (inp[10]) ? 4'b1101 : node16733;
														assign node16733 = (inp[9]) ? node16737 : node16734;
															assign node16734 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node16737 = (inp[1]) ? node16739 : 4'b1100;
																assign node16739 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16743 = (inp[11]) ? 4'b1001 : node16744;
														assign node16744 = (inp[1]) ? node16746 : 4'b1000;
															assign node16746 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node16750 = (inp[13]) ? node16770 : node16751;
													assign node16751 = (inp[11]) ? node16765 : node16752;
														assign node16752 = (inp[1]) ? node16758 : node16753;
															assign node16753 = (inp[9]) ? 4'b1000 : node16754;
																assign node16754 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node16758 = (inp[10]) ? node16762 : node16759;
																assign node16759 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node16762 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node16765 = (inp[1]) ? node16767 : 4'b1001;
															assign node16767 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node16770 = (inp[10]) ? node16776 : node16771;
														assign node16771 = (inp[11]) ? node16773 : 4'b1101;
															assign node16773 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node16776 = (inp[9]) ? node16778 : 4'b1100;
															assign node16778 = (inp[1]) ? node16780 : 4'b1101;
																assign node16780 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node16783 = (inp[13]) ? node16827 : node16784;
											assign node16784 = (inp[2]) ? node16800 : node16785;
												assign node16785 = (inp[1]) ? node16795 : node16786;
													assign node16786 = (inp[9]) ? node16792 : node16787;
														assign node16787 = (inp[11]) ? 4'b1101 : node16788;
															assign node16788 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node16792 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node16795 = (inp[5]) ? 4'b1100 : node16796;
														assign node16796 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node16800 = (inp[1]) ? node16818 : node16801;
													assign node16801 = (inp[5]) ? node16811 : node16802;
														assign node16802 = (inp[11]) ? node16804 : 4'b1000;
															assign node16804 = (inp[9]) ? node16808 : node16805;
																assign node16805 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node16808 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node16811 = (inp[11]) ? 4'b1000 : node16812;
															assign node16812 = (inp[9]) ? 4'b1001 : node16813;
																assign node16813 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node16818 = (inp[5]) ? node16824 : node16819;
														assign node16819 = (inp[9]) ? node16821 : 4'b1100;
															assign node16821 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node16824 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node16827 = (inp[2]) ? node16851 : node16828;
												assign node16828 = (inp[5]) ? node16842 : node16829;
													assign node16829 = (inp[1]) ? node16833 : node16830;
														assign node16830 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node16833 = (inp[11]) ? 4'b1100 : node16834;
															assign node16834 = (inp[9]) ? node16838 : node16835;
																assign node16835 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node16838 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node16842 = (inp[11]) ? 4'b1000 : node16843;
														assign node16843 = (inp[1]) ? 4'b1001 : node16844;
															assign node16844 = (inp[9]) ? 4'b1000 : node16845;
																assign node16845 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node16851 = (inp[5]) ? node16875 : node16852;
													assign node16852 = (inp[1]) ? node16866 : node16853;
														assign node16853 = (inp[11]) ? node16859 : node16854;
															assign node16854 = (inp[10]) ? 4'b1100 : node16855;
																assign node16855 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node16859 = (inp[10]) ? node16863 : node16860;
																assign node16860 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node16863 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node16866 = (inp[11]) ? 4'b1000 : node16867;
															assign node16867 = (inp[10]) ? node16871 : node16868;
																assign node16868 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node16871 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node16875 = (inp[10]) ? node16885 : node16876;
														assign node16876 = (inp[9]) ? node16880 : node16877;
															assign node16877 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node16880 = (inp[11]) ? node16882 : 4'b1101;
																assign node16882 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node16885 = (inp[9]) ? 4'b1100 : 4'b1101;
								assign node16888 = (inp[0]) ? node17162 : node16889;
									assign node16889 = (inp[11]) ? node17015 : node16890;
										assign node16890 = (inp[10]) ? node16948 : node16891;
											assign node16891 = (inp[9]) ? node16917 : node16892;
												assign node16892 = (inp[13]) ? node16912 : node16893;
													assign node16893 = (inp[2]) ? node16903 : node16894;
														assign node16894 = (inp[1]) ? node16900 : node16895;
															assign node16895 = (inp[5]) ? node16897 : 4'b1010;
																assign node16897 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node16900 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node16903 = (inp[15]) ? node16909 : node16904;
															assign node16904 = (inp[1]) ? 4'b1111 : node16905;
																assign node16905 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node16909 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node16912 = (inp[1]) ? 4'b1110 : node16913;
														assign node16913 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node16917 = (inp[1]) ? node16937 : node16918;
													assign node16918 = (inp[15]) ? node16930 : node16919;
														assign node16919 = (inp[2]) ? node16925 : node16920;
															assign node16920 = (inp[13]) ? 4'b1011 : node16921;
																assign node16921 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node16925 = (inp[13]) ? 4'b1110 : node16926;
																assign node16926 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node16930 = (inp[13]) ? 4'b1010 : node16931;
															assign node16931 = (inp[5]) ? 4'b1011 : node16932;
																assign node16932 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node16937 = (inp[13]) ? node16945 : node16938;
														assign node16938 = (inp[2]) ? node16942 : node16939;
															assign node16939 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node16942 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node16945 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node16948 = (inp[9]) ? node16982 : node16949;
												assign node16949 = (inp[5]) ? node16963 : node16950;
													assign node16950 = (inp[15]) ? node16952 : 4'b1011;
														assign node16952 = (inp[1]) ? node16960 : node16953;
															assign node16953 = (inp[13]) ? node16957 : node16954;
																assign node16954 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node16957 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node16960 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node16963 = (inp[1]) ? node16973 : node16964;
														assign node16964 = (inp[15]) ? node16970 : node16965;
															assign node16965 = (inp[13]) ? 4'b1110 : node16966;
																assign node16966 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node16970 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node16973 = (inp[13]) ? node16979 : node16974;
															assign node16974 = (inp[2]) ? 4'b1110 : node16975;
																assign node16975 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node16979 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node16982 = (inp[13]) ? node17004 : node16983;
													assign node16983 = (inp[15]) ? node16993 : node16984;
														assign node16984 = (inp[2]) ? node16988 : node16985;
															assign node16985 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node16988 = (inp[1]) ? 4'b1111 : node16989;
																assign node16989 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node16993 = (inp[2]) ? node16999 : node16994;
															assign node16994 = (inp[1]) ? 4'b1011 : node16995;
																assign node16995 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node16999 = (inp[5]) ? node17001 : 4'b1110;
																assign node17001 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node17004 = (inp[2]) ? node17012 : node17005;
														assign node17005 = (inp[1]) ? 4'b1110 : node17006;
															assign node17006 = (inp[15]) ? 4'b1111 : node17007;
																assign node17007 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node17012 = (inp[1]) ? 4'b1010 : 4'b1011;
										assign node17015 = (inp[13]) ? node17091 : node17016;
											assign node17016 = (inp[2]) ? node17060 : node17017;
												assign node17017 = (inp[5]) ? node17045 : node17018;
													assign node17018 = (inp[1]) ? node17032 : node17019;
														assign node17019 = (inp[9]) ? node17025 : node17020;
															assign node17020 = (inp[10]) ? 4'b1010 : node17021;
																assign node17021 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node17025 = (inp[10]) ? node17029 : node17026;
																assign node17026 = (inp[15]) ? 4'b1011 : 4'b1010;
																assign node17029 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node17032 = (inp[15]) ? node17040 : node17033;
															assign node17033 = (inp[9]) ? node17037 : node17034;
																assign node17034 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node17037 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node17040 = (inp[9]) ? 4'b1011 : node17041;
																assign node17041 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node17045 = (inp[1]) ? 4'b1010 : node17046;
														assign node17046 = (inp[15]) ? node17054 : node17047;
															assign node17047 = (inp[9]) ? node17051 : node17048;
																assign node17048 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17051 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17054 = (inp[10]) ? 4'b1111 : node17055;
																assign node17055 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node17060 = (inp[1]) ? node17078 : node17061;
													assign node17061 = (inp[5]) ? node17069 : node17062;
														assign node17062 = (inp[15]) ? node17064 : 4'b1111;
															assign node17064 = (inp[9]) ? node17066 : 4'b1111;
																assign node17066 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node17069 = (inp[15]) ? node17071 : 4'b1010;
															assign node17071 = (inp[9]) ? node17075 : node17072;
																assign node17072 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node17075 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node17078 = (inp[10]) ? node17084 : node17079;
														assign node17079 = (inp[9]) ? 4'b1111 : node17080;
															assign node17080 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node17084 = (inp[9]) ? node17088 : node17085;
															assign node17085 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node17088 = (inp[15]) ? 4'b1110 : 4'b1111;
											assign node17091 = (inp[2]) ? node17123 : node17092;
												assign node17092 = (inp[5]) ? node17108 : node17093;
													assign node17093 = (inp[15]) ? node17101 : node17094;
														assign node17094 = (inp[10]) ? node17098 : node17095;
															assign node17095 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node17098 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node17101 = (inp[9]) ? node17105 : node17102;
															assign node17102 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node17105 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node17108 = (inp[1]) ? node17114 : node17109;
														assign node17109 = (inp[9]) ? node17111 : 4'b1011;
															assign node17111 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node17114 = (inp[15]) ? 4'b1111 : node17115;
															assign node17115 = (inp[9]) ? node17119 : node17116;
																assign node17116 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17119 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node17123 = (inp[1]) ? node17145 : node17124;
													assign node17124 = (inp[5]) ? node17130 : node17125;
														assign node17125 = (inp[9]) ? node17127 : 4'b1010;
															assign node17127 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node17130 = (inp[15]) ? node17138 : node17131;
															assign node17131 = (inp[9]) ? node17135 : node17132;
																assign node17132 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17135 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17138 = (inp[10]) ? node17142 : node17139;
																assign node17139 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node17142 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node17145 = (inp[5]) ? node17153 : node17146;
														assign node17146 = (inp[9]) ? node17150 : node17147;
															assign node17147 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node17150 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node17153 = (inp[15]) ? node17155 : 4'b1011;
															assign node17155 = (inp[9]) ? node17159 : node17156;
																assign node17156 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node17159 = (inp[10]) ? 4'b1011 : 4'b1010;
									assign node17162 = (inp[15]) ? node17288 : node17163;
										assign node17163 = (inp[11]) ? node17223 : node17164;
											assign node17164 = (inp[10]) ? node17194 : node17165;
												assign node17165 = (inp[9]) ? node17181 : node17166;
													assign node17166 = (inp[2]) ? node17176 : node17167;
														assign node17167 = (inp[1]) ? node17173 : node17168;
															assign node17168 = (inp[5]) ? node17170 : 4'b1010;
																assign node17170 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node17173 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node17176 = (inp[1]) ? node17178 : 4'b1110;
															assign node17178 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node17181 = (inp[5]) ? node17189 : node17182;
														assign node17182 = (inp[2]) ? node17186 : node17183;
															assign node17183 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node17186 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node17189 = (inp[13]) ? 4'b1011 : node17190;
															assign node17190 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node17194 = (inp[9]) ? node17208 : node17195;
													assign node17195 = (inp[5]) ? node17197 : 4'b1111;
														assign node17197 = (inp[2]) ? node17203 : node17198;
															assign node17198 = (inp[13]) ? 4'b1111 : node17199;
																assign node17199 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node17203 = (inp[13]) ? 4'b1011 : node17204;
																assign node17204 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node17208 = (inp[1]) ? node17216 : node17209;
														assign node17209 = (inp[2]) ? node17211 : 4'b1110;
															assign node17211 = (inp[13]) ? node17213 : 4'b1110;
																assign node17213 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node17216 = (inp[2]) ? node17220 : node17217;
															assign node17217 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node17220 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node17223 = (inp[10]) ? node17253 : node17224;
												assign node17224 = (inp[13]) ? node17236 : node17225;
													assign node17225 = (inp[9]) ? node17229 : node17226;
														assign node17226 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node17229 = (inp[2]) ? node17231 : 4'b1110;
															assign node17231 = (inp[5]) ? node17233 : 4'b1110;
																assign node17233 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node17236 = (inp[9]) ? node17246 : node17237;
														assign node17237 = (inp[2]) ? node17243 : node17238;
															assign node17238 = (inp[1]) ? 4'b1110 : node17239;
																assign node17239 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node17243 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node17246 = (inp[2]) ? node17250 : node17247;
															assign node17247 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node17250 = (inp[5]) ? 4'b1110 : 4'b1011;
												assign node17253 = (inp[9]) ? node17269 : node17254;
													assign node17254 = (inp[5]) ? node17260 : node17255;
														assign node17255 = (inp[2]) ? 4'b1011 : node17256;
															assign node17256 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node17260 = (inp[2]) ? node17262 : 4'b1111;
															assign node17262 = (inp[13]) ? node17266 : node17263;
																assign node17263 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node17266 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node17269 = (inp[13]) ? node17277 : node17270;
														assign node17270 = (inp[2]) ? 4'b1111 : node17271;
															assign node17271 = (inp[1]) ? 4'b1010 : node17272;
																assign node17272 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node17277 = (inp[2]) ? node17283 : node17278;
															assign node17278 = (inp[1]) ? 4'b1110 : node17279;
																assign node17279 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node17283 = (inp[1]) ? 4'b1010 : node17284;
																assign node17284 = (inp[5]) ? 4'b1111 : 4'b1010;
										assign node17288 = (inp[5]) ? node17352 : node17289;
											assign node17289 = (inp[2]) ? node17323 : node17290;
												assign node17290 = (inp[13]) ? node17302 : node17291;
													assign node17291 = (inp[9]) ? node17293 : 4'b1011;
														assign node17293 = (inp[1]) ? 4'b1010 : node17294;
															assign node17294 = (inp[11]) ? node17298 : node17295;
																assign node17295 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node17298 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node17302 = (inp[1]) ? node17316 : node17303;
														assign node17303 = (inp[11]) ? node17311 : node17304;
															assign node17304 = (inp[9]) ? node17308 : node17305;
																assign node17305 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node17308 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node17311 = (inp[10]) ? 4'b1110 : node17312;
																assign node17312 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node17316 = (inp[9]) ? node17320 : node17317;
															assign node17317 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17320 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node17323 = (inp[13]) ? node17339 : node17324;
													assign node17324 = (inp[1]) ? node17332 : node17325;
														assign node17325 = (inp[9]) ? node17329 : node17326;
															assign node17326 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17329 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node17332 = (inp[11]) ? node17334 : 4'b1110;
															assign node17334 = (inp[10]) ? 4'b1110 : node17335;
																assign node17335 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node17339 = (inp[10]) ? node17345 : node17340;
														assign node17340 = (inp[9]) ? node17342 : 4'b1010;
															assign node17342 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node17345 = (inp[1]) ? 4'b1011 : node17346;
															assign node17346 = (inp[9]) ? node17348 : 4'b1010;
																assign node17348 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node17352 = (inp[11]) ? node17406 : node17353;
												assign node17353 = (inp[9]) ? node17383 : node17354;
													assign node17354 = (inp[10]) ? node17368 : node17355;
														assign node17355 = (inp[13]) ? node17363 : node17356;
															assign node17356 = (inp[1]) ? node17360 : node17357;
																assign node17357 = (inp[2]) ? 4'b1010 : 4'b1110;
																assign node17360 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node17363 = (inp[1]) ? node17365 : 4'b1111;
																assign node17365 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node17368 = (inp[1]) ? node17376 : node17369;
															assign node17369 = (inp[2]) ? node17373 : node17370;
																assign node17370 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node17373 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node17376 = (inp[13]) ? node17380 : node17377;
																assign node17377 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node17380 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node17383 = (inp[2]) ? node17391 : node17384;
														assign node17384 = (inp[1]) ? node17388 : node17385;
															assign node17385 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node17388 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node17391 = (inp[13]) ? node17399 : node17392;
															assign node17392 = (inp[1]) ? node17396 : node17393;
																assign node17393 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node17396 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17399 = (inp[1]) ? node17403 : node17400;
																assign node17400 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node17403 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node17406 = (inp[1]) ? node17428 : node17407;
													assign node17407 = (inp[10]) ? node17417 : node17408;
														assign node17408 = (inp[13]) ? node17412 : node17409;
															assign node17409 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node17412 = (inp[9]) ? 4'b1010 : node17413;
																assign node17413 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node17417 = (inp[13]) ? node17423 : node17418;
															assign node17418 = (inp[9]) ? 4'b1110 : node17419;
																assign node17419 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node17423 = (inp[2]) ? node17425 : 4'b1011;
																assign node17425 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node17428 = (inp[9]) ? node17436 : node17429;
														assign node17429 = (inp[10]) ? node17433 : node17430;
															assign node17430 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node17433 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node17436 = (inp[2]) ? node17444 : node17437;
															assign node17437 = (inp[13]) ? node17441 : node17438;
																assign node17438 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node17441 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node17444 = (inp[13]) ? 4'b1011 : 4'b1111;
						assign node17447 = (inp[7]) ? node18551 : node17448;
							assign node17448 = (inp[15]) ? node18002 : node17449;
								assign node17449 = (inp[5]) ? node17729 : node17450;
									assign node17450 = (inp[4]) ? node17594 : node17451;
										assign node17451 = (inp[11]) ? node17529 : node17452;
											assign node17452 = (inp[9]) ? node17488 : node17453;
												assign node17453 = (inp[10]) ? node17471 : node17454;
													assign node17454 = (inp[2]) ? node17462 : node17455;
														assign node17455 = (inp[1]) ? node17459 : node17456;
															assign node17456 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node17459 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node17462 = (inp[1]) ? node17468 : node17463;
															assign node17463 = (inp[13]) ? 4'b1011 : node17464;
																assign node17464 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node17468 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node17471 = (inp[1]) ? node17479 : node17472;
														assign node17472 = (inp[13]) ? node17476 : node17473;
															assign node17473 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node17476 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node17479 = (inp[2]) ? node17485 : node17480;
															assign node17480 = (inp[13]) ? node17482 : 4'b1110;
																assign node17482 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node17485 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node17488 = (inp[0]) ? node17504 : node17489;
													assign node17489 = (inp[13]) ? node17501 : node17490;
														assign node17490 = (inp[10]) ? node17498 : node17491;
															assign node17491 = (inp[2]) ? node17495 : node17492;
																assign node17492 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node17495 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node17498 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node17501 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node17504 = (inp[2]) ? node17518 : node17505;
														assign node17505 = (inp[10]) ? node17511 : node17506;
															assign node17506 = (inp[13]) ? 4'b1011 : node17507;
																assign node17507 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node17511 = (inp[1]) ? node17515 : node17512;
																assign node17512 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node17515 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node17518 = (inp[13]) ? node17526 : node17519;
															assign node17519 = (inp[1]) ? node17523 : node17520;
																assign node17520 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node17523 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node17526 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node17529 = (inp[13]) ? node17563 : node17530;
												assign node17530 = (inp[2]) ? node17546 : node17531;
													assign node17531 = (inp[1]) ? 4'b1111 : node17532;
														assign node17532 = (inp[9]) ? node17538 : node17533;
															assign node17533 = (inp[10]) ? 4'b1011 : node17534;
																assign node17534 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node17538 = (inp[0]) ? node17542 : node17539;
																assign node17539 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node17542 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node17546 = (inp[1]) ? node17556 : node17547;
														assign node17547 = (inp[0]) ? node17549 : 4'b1111;
															assign node17549 = (inp[10]) ? node17553 : node17550;
																assign node17550 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node17553 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node17556 = (inp[0]) ? node17558 : 4'b1010;
															assign node17558 = (inp[9]) ? 4'b1011 : node17559;
																assign node17559 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node17563 = (inp[1]) ? node17585 : node17564;
													assign node17564 = (inp[2]) ? node17572 : node17565;
														assign node17565 = (inp[10]) ? 4'b1110 : node17566;
															assign node17566 = (inp[9]) ? node17568 : 4'b1111;
																assign node17568 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17572 = (inp[9]) ? node17578 : node17573;
															assign node17573 = (inp[0]) ? 4'b1011 : node17574;
																assign node17574 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node17578 = (inp[0]) ? node17582 : node17579;
																assign node17579 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node17582 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node17585 = (inp[2]) ? node17587 : 4'b1010;
														assign node17587 = (inp[9]) ? 4'b1110 : node17588;
															assign node17588 = (inp[0]) ? 4'b1111 : node17589;
																assign node17589 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node17594 = (inp[11]) ? node17662 : node17595;
											assign node17595 = (inp[2]) ? node17633 : node17596;
												assign node17596 = (inp[13]) ? node17614 : node17597;
													assign node17597 = (inp[1]) ? node17603 : node17598;
														assign node17598 = (inp[9]) ? node17600 : 4'b1111;
															assign node17600 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node17603 = (inp[10]) ? node17609 : node17604;
															assign node17604 = (inp[0]) ? 4'b1010 : node17605;
																assign node17605 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node17609 = (inp[0]) ? 4'b1011 : node17610;
																assign node17610 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node17614 = (inp[1]) ? node17622 : node17615;
														assign node17615 = (inp[10]) ? 4'b1010 : node17616;
															assign node17616 = (inp[9]) ? node17618 : 4'b1011;
																assign node17618 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17622 = (inp[10]) ? node17628 : node17623;
															assign node17623 = (inp[0]) ? 4'b1110 : node17624;
																assign node17624 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node17628 = (inp[9]) ? 4'b1111 : node17629;
																assign node17629 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node17633 = (inp[10]) ? node17651 : node17634;
													assign node17634 = (inp[9]) ? node17644 : node17635;
														assign node17635 = (inp[1]) ? node17639 : node17636;
															assign node17636 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node17639 = (inp[13]) ? node17641 : 4'b1111;
																assign node17641 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node17644 = (inp[0]) ? 4'b1011 : node17645;
															assign node17645 = (inp[1]) ? node17647 : 4'b1011;
																assign node17647 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node17651 = (inp[9]) ? node17657 : node17652;
														assign node17652 = (inp[1]) ? node17654 : 4'b1011;
															assign node17654 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node17657 = (inp[13]) ? node17659 : 4'b1010;
															assign node17659 = (inp[1]) ? 4'b1010 : 4'b1110;
											assign node17662 = (inp[1]) ? node17698 : node17663;
												assign node17663 = (inp[0]) ? node17683 : node17664;
													assign node17664 = (inp[2]) ? node17674 : node17665;
														assign node17665 = (inp[13]) ? 4'b1011 : node17666;
															assign node17666 = (inp[10]) ? node17670 : node17667;
																assign node17667 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node17670 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node17674 = (inp[13]) ? node17678 : node17675;
															assign node17675 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node17678 = (inp[10]) ? node17680 : 4'b1110;
																assign node17680 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node17683 = (inp[9]) ? node17691 : node17684;
														assign node17684 = (inp[10]) ? 4'b1111 : node17685;
															assign node17685 = (inp[13]) ? 4'b1110 : node17686;
																assign node17686 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node17691 = (inp[10]) ? node17693 : 4'b1111;
															assign node17693 = (inp[13]) ? node17695 : 4'b1110;
																assign node17695 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node17698 = (inp[10]) ? node17720 : node17699;
													assign node17699 = (inp[9]) ? node17711 : node17700;
														assign node17700 = (inp[0]) ? node17704 : node17701;
															assign node17701 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node17704 = (inp[13]) ? node17708 : node17705;
																assign node17705 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node17708 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node17711 = (inp[2]) ? node17715 : node17712;
															assign node17712 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node17715 = (inp[0]) ? node17717 : 4'b1111;
																assign node17717 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node17720 = (inp[9]) ? node17722 : 4'b1010;
														assign node17722 = (inp[13]) ? node17726 : node17723;
															assign node17723 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node17726 = (inp[2]) ? 4'b1011 : 4'b1111;
									assign node17729 = (inp[4]) ? node17855 : node17730;
										assign node17730 = (inp[1]) ? node17786 : node17731;
											assign node17731 = (inp[13]) ? node17761 : node17732;
												assign node17732 = (inp[2]) ? node17740 : node17733;
													assign node17733 = (inp[9]) ? node17737 : node17734;
														assign node17734 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node17737 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node17740 = (inp[0]) ? node17756 : node17741;
														assign node17741 = (inp[9]) ? node17749 : node17742;
															assign node17742 = (inp[11]) ? node17746 : node17743;
																assign node17743 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17746 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17749 = (inp[10]) ? node17753 : node17750;
																assign node17750 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node17753 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node17756 = (inp[10]) ? node17758 : 4'b1111;
															assign node17758 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node17761 = (inp[2]) ? node17769 : node17762;
													assign node17762 = (inp[10]) ? 4'b1110 : node17763;
														assign node17763 = (inp[9]) ? 4'b1111 : node17764;
															assign node17764 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node17769 = (inp[0]) ? node17777 : node17770;
														assign node17770 = (inp[9]) ? node17774 : node17771;
															assign node17771 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node17774 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node17777 = (inp[10]) ? 4'b1011 : node17778;
															assign node17778 = (inp[11]) ? node17782 : node17779;
																assign node17779 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node17782 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node17786 = (inp[9]) ? node17816 : node17787;
												assign node17787 = (inp[13]) ? node17801 : node17788;
													assign node17788 = (inp[2]) ? node17794 : node17789;
														assign node17789 = (inp[10]) ? 4'b1010 : node17790;
															assign node17790 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node17794 = (inp[11]) ? node17796 : 4'b1110;
															assign node17796 = (inp[0]) ? 4'b1111 : node17797;
																assign node17797 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node17801 = (inp[2]) ? node17813 : node17802;
														assign node17802 = (inp[10]) ? node17808 : node17803;
															assign node17803 = (inp[11]) ? 4'b1111 : node17804;
																assign node17804 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node17808 = (inp[11]) ? 4'b1110 : node17809;
																assign node17809 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17813 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node17816 = (inp[10]) ? node17836 : node17817;
													assign node17817 = (inp[2]) ? node17825 : node17818;
														assign node17818 = (inp[13]) ? 4'b1110 : node17819;
															assign node17819 = (inp[11]) ? 4'b1010 : node17820;
																assign node17820 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node17825 = (inp[13]) ? node17831 : node17826;
															assign node17826 = (inp[11]) ? node17828 : 4'b1111;
																assign node17828 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node17831 = (inp[0]) ? node17833 : 4'b1011;
																assign node17833 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node17836 = (inp[2]) ? node17844 : node17837;
														assign node17837 = (inp[13]) ? node17839 : 4'b1011;
															assign node17839 = (inp[0]) ? node17841 : 4'b1111;
																assign node17841 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node17844 = (inp[13]) ? node17850 : node17845;
															assign node17845 = (inp[0]) ? 4'b1110 : node17846;
																assign node17846 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node17850 = (inp[0]) ? node17852 : 4'b1010;
																assign node17852 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node17855 = (inp[1]) ? node17935 : node17856;
											assign node17856 = (inp[0]) ? node17898 : node17857;
												assign node17857 = (inp[9]) ? node17875 : node17858;
													assign node17858 = (inp[2]) ? node17866 : node17859;
														assign node17859 = (inp[13]) ? node17863 : node17860;
															assign node17860 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17863 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node17866 = (inp[13]) ? node17868 : 4'b1011;
															assign node17868 = (inp[11]) ? node17872 : node17869;
																assign node17869 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17872 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node17875 = (inp[13]) ? node17889 : node17876;
														assign node17876 = (inp[2]) ? node17884 : node17877;
															assign node17877 = (inp[11]) ? node17881 : node17878;
																assign node17878 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node17881 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node17884 = (inp[11]) ? node17886 : 4'b1010;
																assign node17886 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node17889 = (inp[2]) ? node17893 : node17890;
															assign node17890 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node17893 = (inp[10]) ? 4'b1111 : node17894;
																assign node17894 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node17898 = (inp[9]) ? node17920 : node17899;
													assign node17899 = (inp[10]) ? node17911 : node17900;
														assign node17900 = (inp[11]) ? node17904 : node17901;
															assign node17901 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node17904 = (inp[2]) ? node17908 : node17905;
																assign node17905 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node17908 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node17911 = (inp[2]) ? node17917 : node17912;
															assign node17912 = (inp[13]) ? node17914 : 4'b1110;
																assign node17914 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node17917 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node17920 = (inp[10]) ? node17928 : node17921;
														assign node17921 = (inp[2]) ? node17925 : node17922;
															assign node17922 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node17925 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node17928 = (inp[13]) ? node17932 : node17929;
															assign node17929 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node17932 = (inp[2]) ? 4'b1111 : 4'b1010;
											assign node17935 = (inp[11]) ? node17961 : node17936;
												assign node17936 = (inp[13]) ? node17944 : node17937;
													assign node17937 = (inp[2]) ? node17939 : 4'b1111;
														assign node17939 = (inp[9]) ? node17941 : 4'b1010;
															assign node17941 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node17944 = (inp[2]) ? node17952 : node17945;
														assign node17945 = (inp[0]) ? node17947 : 4'b1011;
															assign node17947 = (inp[10]) ? node17949 : 4'b1010;
																assign node17949 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node17952 = (inp[0]) ? node17956 : node17953;
															assign node17953 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17956 = (inp[10]) ? node17958 : 4'b1111;
																assign node17958 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node17961 = (inp[9]) ? node17985 : node17962;
													assign node17962 = (inp[13]) ? node17974 : node17963;
														assign node17963 = (inp[2]) ? node17971 : node17964;
															assign node17964 = (inp[0]) ? node17968 : node17965;
																assign node17965 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node17968 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node17971 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node17974 = (inp[2]) ? node17978 : node17975;
															assign node17975 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node17978 = (inp[10]) ? node17982 : node17979;
																assign node17979 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node17982 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node17985 = (inp[2]) ? node17995 : node17986;
														assign node17986 = (inp[13]) ? 4'b1011 : node17987;
															assign node17987 = (inp[10]) ? node17991 : node17988;
																assign node17988 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node17991 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node17995 = (inp[13]) ? node17997 : 4'b1011;
															assign node17997 = (inp[10]) ? 4'b1110 : node17998;
																assign node17998 = (inp[0]) ? 4'b1111 : 4'b1110;
								assign node18002 = (inp[4]) ? node18268 : node18003;
									assign node18003 = (inp[9]) ? node18141 : node18004;
										assign node18004 = (inp[10]) ? node18080 : node18005;
											assign node18005 = (inp[0]) ? node18043 : node18006;
												assign node18006 = (inp[2]) ? node18024 : node18007;
													assign node18007 = (inp[13]) ? node18015 : node18008;
														assign node18008 = (inp[1]) ? node18010 : 4'b1000;
															assign node18010 = (inp[5]) ? node18012 : 4'b1101;
																assign node18012 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node18015 = (inp[1]) ? node18019 : node18016;
															assign node18016 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node18019 = (inp[5]) ? 4'b1001 : node18020;
																assign node18020 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node18024 = (inp[13]) ? node18034 : node18025;
														assign node18025 = (inp[11]) ? node18029 : node18026;
															assign node18026 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node18029 = (inp[5]) ? node18031 : 4'b1000;
																assign node18031 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node18034 = (inp[5]) ? node18040 : node18035;
															assign node18035 = (inp[11]) ? 4'b1101 : node18036;
																assign node18036 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node18040 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node18043 = (inp[2]) ? node18061 : node18044;
													assign node18044 = (inp[5]) ? node18052 : node18045;
														assign node18045 = (inp[13]) ? 4'b1001 : node18046;
															assign node18046 = (inp[1]) ? node18048 : 4'b1100;
																assign node18048 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node18052 = (inp[1]) ? node18058 : node18053;
															assign node18053 = (inp[13]) ? 4'b1100 : node18054;
																assign node18054 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node18058 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node18061 = (inp[13]) ? node18071 : node18062;
														assign node18062 = (inp[1]) ? node18066 : node18063;
															assign node18063 = (inp[11]) ? 4'b1101 : 4'b1001;
															assign node18066 = (inp[5]) ? 4'b1001 : node18067;
																assign node18067 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node18071 = (inp[1]) ? node18075 : node18072;
															assign node18072 = (inp[5]) ? 4'b1001 : 4'b1100;
															assign node18075 = (inp[11]) ? node18077 : 4'b1100;
																assign node18077 = (inp[5]) ? 4'b1100 : 4'b1101;
											assign node18080 = (inp[0]) ? node18112 : node18081;
												assign node18081 = (inp[13]) ? node18097 : node18082;
													assign node18082 = (inp[2]) ? node18090 : node18083;
														assign node18083 = (inp[11]) ? 4'b1100 : node18084;
															assign node18084 = (inp[1]) ? node18086 : 4'b1101;
																assign node18086 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node18090 = (inp[5]) ? node18094 : node18091;
															assign node18091 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node18094 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node18097 = (inp[2]) ? node18107 : node18098;
														assign node18098 = (inp[5]) ? node18104 : node18099;
															assign node18099 = (inp[1]) ? node18101 : 4'b1000;
																assign node18101 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18104 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node18107 = (inp[1]) ? 4'b1100 : node18108;
															assign node18108 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node18112 = (inp[13]) ? node18130 : node18113;
													assign node18113 = (inp[2]) ? node18125 : node18114;
														assign node18114 = (inp[1]) ? node18120 : node18115;
															assign node18115 = (inp[5]) ? node18117 : 4'b1101;
																assign node18117 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18120 = (inp[11]) ? node18122 : 4'b1101;
																assign node18122 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node18125 = (inp[5]) ? node18127 : 4'b1000;
															assign node18127 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node18130 = (inp[2]) ? node18136 : node18131;
														assign node18131 = (inp[5]) ? node18133 : 4'b1000;
															assign node18133 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node18136 = (inp[5]) ? node18138 : 4'b1101;
															assign node18138 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node18141 = (inp[5]) ? node18201 : node18142;
											assign node18142 = (inp[10]) ? node18172 : node18143;
												assign node18143 = (inp[0]) ? node18159 : node18144;
													assign node18144 = (inp[2]) ? node18150 : node18145;
														assign node18145 = (inp[13]) ? node18147 : 4'b1100;
															assign node18147 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18150 = (inp[13]) ? node18154 : node18151;
															assign node18151 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node18154 = (inp[1]) ? 4'b1100 : node18155;
																assign node18155 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node18159 = (inp[1]) ? node18165 : node18160;
														assign node18160 = (inp[2]) ? node18162 : 4'b1101;
															assign node18162 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node18165 = (inp[2]) ? node18167 : 4'b1000;
															assign node18167 = (inp[13]) ? 4'b1101 : node18168;
																assign node18168 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node18172 = (inp[13]) ? node18188 : node18173;
													assign node18173 = (inp[2]) ? node18181 : node18174;
														assign node18174 = (inp[11]) ? node18176 : 4'b1100;
															assign node18176 = (inp[0]) ? node18178 : 4'b1101;
																assign node18178 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node18181 = (inp[0]) ? node18183 : 4'b1000;
															assign node18183 = (inp[11]) ? node18185 : 4'b1001;
																assign node18185 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node18188 = (inp[2]) ? node18196 : node18189;
														assign node18189 = (inp[1]) ? 4'b1001 : node18190;
															assign node18190 = (inp[0]) ? node18192 : 4'b1001;
																assign node18192 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18196 = (inp[0]) ? node18198 : 4'b1101;
															assign node18198 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node18201 = (inp[13]) ? node18241 : node18202;
												assign node18202 = (inp[11]) ? node18222 : node18203;
													assign node18203 = (inp[0]) ? node18215 : node18204;
														assign node18204 = (inp[1]) ? node18210 : node18205;
															assign node18205 = (inp[2]) ? node18207 : 4'b1001;
																assign node18207 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node18210 = (inp[2]) ? 4'b1001 : node18211;
																assign node18211 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node18215 = (inp[10]) ? node18217 : 4'b1101;
															assign node18217 = (inp[1]) ? 4'b1001 : node18218;
																assign node18218 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node18222 = (inp[0]) ? node18228 : node18223;
														assign node18223 = (inp[10]) ? 4'b1101 : node18224;
															assign node18224 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node18228 = (inp[2]) ? node18234 : node18229;
															assign node18229 = (inp[10]) ? node18231 : 4'b1101;
																assign node18231 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node18234 = (inp[1]) ? node18238 : node18235;
																assign node18235 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node18238 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node18241 = (inp[1]) ? node18253 : node18242;
													assign node18242 = (inp[2]) ? node18246 : node18243;
														assign node18243 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node18246 = (inp[10]) ? 4'b1000 : node18247;
															assign node18247 = (inp[0]) ? node18249 : 4'b1001;
																assign node18249 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node18253 = (inp[2]) ? node18259 : node18254;
														assign node18254 = (inp[11]) ? node18256 : 4'b1001;
															assign node18256 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node18259 = (inp[10]) ? node18265 : node18260;
															assign node18260 = (inp[11]) ? node18262 : 4'b1101;
																assign node18262 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node18265 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node18268 = (inp[0]) ? node18412 : node18269;
										assign node18269 = (inp[11]) ? node18347 : node18270;
											assign node18270 = (inp[2]) ? node18306 : node18271;
												assign node18271 = (inp[13]) ? node18289 : node18272;
													assign node18272 = (inp[1]) ? node18280 : node18273;
														assign node18273 = (inp[10]) ? node18275 : 4'b1010;
															assign node18275 = (inp[9]) ? node18277 : 4'b1010;
																assign node18277 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node18280 = (inp[5]) ? 4'b1010 : node18281;
															assign node18281 = (inp[10]) ? node18285 : node18282;
																assign node18282 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node18285 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node18289 = (inp[5]) ? node18299 : node18290;
														assign node18290 = (inp[1]) ? 4'b1010 : node18291;
															assign node18291 = (inp[9]) ? node18295 : node18292;
																assign node18292 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node18295 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node18299 = (inp[9]) ? node18303 : node18300;
															assign node18300 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node18303 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node18306 = (inp[13]) ? node18332 : node18307;
													assign node18307 = (inp[1]) ? node18321 : node18308;
														assign node18308 = (inp[5]) ? node18316 : node18309;
															assign node18309 = (inp[10]) ? node18313 : node18310;
																assign node18310 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node18313 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node18316 = (inp[10]) ? node18318 : 4'b1110;
																assign node18318 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node18321 = (inp[5]) ? node18327 : node18322;
															assign node18322 = (inp[9]) ? 4'b1010 : node18323;
																assign node18323 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node18327 = (inp[10]) ? 4'b1110 : node18328;
																assign node18328 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node18332 = (inp[1]) ? node18342 : node18333;
														assign node18333 = (inp[10]) ? node18335 : 4'b1011;
															assign node18335 = (inp[5]) ? node18339 : node18336;
																assign node18336 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node18339 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node18342 = (inp[5]) ? 4'b1010 : node18343;
															assign node18343 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node18347 = (inp[9]) ? node18379 : node18348;
												assign node18348 = (inp[2]) ? node18364 : node18349;
													assign node18349 = (inp[1]) ? node18353 : node18350;
														assign node18350 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node18353 = (inp[13]) ? node18359 : node18354;
															assign node18354 = (inp[5]) ? node18356 : 4'b1111;
																assign node18356 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node18359 = (inp[5]) ? 4'b1110 : node18360;
																assign node18360 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node18364 = (inp[13]) ? node18374 : node18365;
														assign node18365 = (inp[5]) ? node18371 : node18366;
															assign node18366 = (inp[1]) ? node18368 : 4'b1110;
																assign node18368 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node18371 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node18374 = (inp[10]) ? 4'b1010 : node18375;
															assign node18375 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node18379 = (inp[10]) ? node18395 : node18380;
													assign node18380 = (inp[2]) ? node18392 : node18381;
														assign node18381 = (inp[13]) ? node18389 : node18382;
															assign node18382 = (inp[5]) ? node18386 : node18383;
																assign node18383 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node18386 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node18389 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node18392 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node18395 = (inp[2]) ? node18405 : node18396;
														assign node18396 = (inp[1]) ? node18400 : node18397;
															assign node18397 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node18400 = (inp[5]) ? 4'b1111 : node18401;
																assign node18401 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node18405 = (inp[13]) ? node18409 : node18406;
															assign node18406 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node18409 = (inp[5]) ? 4'b1011 : 4'b1110;
										assign node18412 = (inp[9]) ? node18474 : node18413;
											assign node18413 = (inp[10]) ? node18445 : node18414;
												assign node18414 = (inp[1]) ? node18430 : node18415;
													assign node18415 = (inp[11]) ? node18423 : node18416;
														assign node18416 = (inp[2]) ? node18420 : node18417;
															assign node18417 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node18420 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node18423 = (inp[13]) ? node18425 : 4'b1111;
															assign node18425 = (inp[2]) ? 4'b1010 : node18426;
																assign node18426 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node18430 = (inp[5]) ? node18440 : node18431;
														assign node18431 = (inp[13]) ? node18435 : node18432;
															assign node18432 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node18435 = (inp[2]) ? 4'b1111 : node18436;
																assign node18436 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node18440 = (inp[13]) ? 4'b1010 : node18441;
															assign node18441 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node18445 = (inp[13]) ? node18459 : node18446;
													assign node18446 = (inp[5]) ? node18454 : node18447;
														assign node18447 = (inp[2]) ? node18451 : node18448;
															assign node18448 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node18451 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node18454 = (inp[2]) ? node18456 : 4'b1011;
															assign node18456 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18459 = (inp[2]) ? node18469 : node18460;
														assign node18460 = (inp[1]) ? node18466 : node18461;
															assign node18461 = (inp[11]) ? 4'b1110 : node18462;
																assign node18462 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node18466 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node18469 = (inp[5]) ? 4'b1011 : node18470;
															assign node18470 = (inp[11]) ? 4'b1110 : 4'b1011;
											assign node18474 = (inp[10]) ? node18516 : node18475;
												assign node18475 = (inp[1]) ? node18501 : node18476;
													assign node18476 = (inp[5]) ? node18490 : node18477;
														assign node18477 = (inp[11]) ? node18485 : node18478;
															assign node18478 = (inp[13]) ? node18482 : node18479;
																assign node18479 = (inp[2]) ? 4'b1111 : 4'b1010;
																assign node18482 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node18485 = (inp[13]) ? node18487 : 4'b1011;
																assign node18487 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node18490 = (inp[13]) ? node18496 : node18491;
															assign node18491 = (inp[2]) ? 4'b1110 : node18492;
																assign node18492 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node18496 = (inp[11]) ? 4'b1011 : node18497;
																assign node18497 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node18501 = (inp[13]) ? node18511 : node18502;
														assign node18502 = (inp[5]) ? node18506 : node18503;
															assign node18503 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node18506 = (inp[2]) ? node18508 : 4'b1010;
																assign node18508 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node18511 = (inp[5]) ? node18513 : 4'b1110;
															assign node18513 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node18516 = (inp[1]) ? node18538 : node18517;
													assign node18517 = (inp[5]) ? node18525 : node18518;
														assign node18518 = (inp[2]) ? 4'b1010 : node18519;
															assign node18519 = (inp[13]) ? node18521 : 4'b1010;
																assign node18521 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node18525 = (inp[11]) ? node18533 : node18526;
															assign node18526 = (inp[13]) ? node18530 : node18527;
																assign node18527 = (inp[2]) ? 4'b1111 : 4'b1010;
																assign node18530 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node18533 = (inp[13]) ? node18535 : 4'b1011;
																assign node18535 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node18538 = (inp[13]) ? node18544 : node18539;
														assign node18539 = (inp[5]) ? node18541 : 4'b1010;
															assign node18541 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18544 = (inp[11]) ? node18546 : 4'b1010;
															assign node18546 = (inp[5]) ? 4'b1010 : node18547;
																assign node18547 = (inp[2]) ? 4'b1111 : 4'b1011;
							assign node18551 = (inp[4]) ? node19107 : node18552;
								assign node18552 = (inp[15]) ? node18854 : node18553;
									assign node18553 = (inp[11]) ? node18699 : node18554;
										assign node18554 = (inp[1]) ? node18638 : node18555;
											assign node18555 = (inp[0]) ? node18599 : node18556;
												assign node18556 = (inp[5]) ? node18578 : node18557;
													assign node18557 = (inp[9]) ? node18569 : node18558;
														assign node18558 = (inp[13]) ? node18566 : node18559;
															assign node18559 = (inp[2]) ? node18563 : node18560;
																assign node18560 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node18563 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node18566 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node18569 = (inp[10]) ? node18571 : 4'b1100;
															assign node18571 = (inp[2]) ? node18575 : node18572;
																assign node18572 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node18575 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node18578 = (inp[13]) ? node18592 : node18579;
														assign node18579 = (inp[2]) ? node18587 : node18580;
															assign node18580 = (inp[10]) ? node18584 : node18581;
																assign node18581 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node18584 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node18587 = (inp[10]) ? 4'b1100 : node18588;
																assign node18588 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node18592 = (inp[2]) ? 4'b1000 : node18593;
															assign node18593 = (inp[10]) ? node18595 : 4'b1100;
																assign node18595 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node18599 = (inp[5]) ? node18615 : node18600;
													assign node18600 = (inp[13]) ? node18610 : node18601;
														assign node18601 = (inp[2]) ? node18607 : node18602;
															assign node18602 = (inp[9]) ? 4'b1101 : node18603;
																assign node18603 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node18607 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node18610 = (inp[2]) ? 4'b1100 : node18611;
															assign node18611 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node18615 = (inp[9]) ? node18625 : node18616;
														assign node18616 = (inp[2]) ? node18622 : node18617;
															assign node18617 = (inp[13]) ? 4'b1101 : node18618;
																assign node18618 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node18622 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node18625 = (inp[2]) ? node18633 : node18626;
															assign node18626 = (inp[10]) ? node18630 : node18627;
																assign node18627 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node18630 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node18633 = (inp[10]) ? node18635 : 4'b1000;
																assign node18635 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node18638 = (inp[10]) ? node18664 : node18639;
												assign node18639 = (inp[9]) ? node18649 : node18640;
													assign node18640 = (inp[5]) ? node18642 : 4'b1000;
														assign node18642 = (inp[2]) ? node18646 : node18643;
															assign node18643 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node18646 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node18649 = (inp[13]) ? node18661 : node18650;
														assign node18650 = (inp[2]) ? node18656 : node18651;
															assign node18651 = (inp[0]) ? node18653 : 4'b1100;
																assign node18653 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node18656 = (inp[5]) ? 4'b1001 : node18657;
																assign node18657 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node18661 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node18664 = (inp[9]) ? node18678 : node18665;
													assign node18665 = (inp[2]) ? node18671 : node18666;
														assign node18666 = (inp[0]) ? node18668 : 4'b1100;
															assign node18668 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node18671 = (inp[13]) ? node18673 : 4'b1001;
															assign node18673 = (inp[5]) ? 4'b1101 : node18674;
																assign node18674 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node18678 = (inp[2]) ? node18688 : node18679;
														assign node18679 = (inp[13]) ? node18685 : node18680;
															assign node18680 = (inp[0]) ? node18682 : 4'b1101;
																assign node18682 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node18685 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node18688 = (inp[13]) ? node18694 : node18689;
															assign node18689 = (inp[0]) ? node18691 : 4'b1000;
																assign node18691 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node18694 = (inp[0]) ? node18696 : 4'b1100;
																assign node18696 = (inp[5]) ? 4'b1100 : 4'b1101;
										assign node18699 = (inp[9]) ? node18773 : node18700;
											assign node18700 = (inp[0]) ? node18738 : node18701;
												assign node18701 = (inp[1]) ? node18723 : node18702;
													assign node18702 = (inp[5]) ? node18712 : node18703;
														assign node18703 = (inp[10]) ? node18707 : node18704;
															assign node18704 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node18707 = (inp[2]) ? node18709 : 4'b1001;
																assign node18709 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node18712 = (inp[13]) ? node18716 : node18713;
															assign node18713 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node18716 = (inp[2]) ? node18720 : node18717;
																assign node18717 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node18720 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node18723 = (inp[10]) ? node18731 : node18724;
														assign node18724 = (inp[13]) ? 4'b1001 : node18725;
															assign node18725 = (inp[2]) ? node18727 : 4'b1100;
																assign node18727 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node18731 = (inp[2]) ? node18735 : node18732;
															assign node18732 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node18735 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node18738 = (inp[2]) ? node18756 : node18739;
													assign node18739 = (inp[1]) ? node18751 : node18740;
														assign node18740 = (inp[5]) ? node18744 : node18741;
															assign node18741 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node18744 = (inp[10]) ? node18748 : node18745;
																assign node18745 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node18748 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node18751 = (inp[13]) ? 4'b1001 : node18752;
															assign node18752 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node18756 = (inp[13]) ? node18766 : node18757;
														assign node18757 = (inp[1]) ? node18763 : node18758;
															assign node18758 = (inp[5]) ? node18760 : 4'b1000;
																assign node18760 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node18763 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node18766 = (inp[5]) ? node18768 : 4'b1100;
															assign node18768 = (inp[1]) ? 4'b1100 : node18769;
																assign node18769 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node18773 = (inp[2]) ? node18811 : node18774;
												assign node18774 = (inp[13]) ? node18792 : node18775;
													assign node18775 = (inp[1]) ? node18787 : node18776;
														assign node18776 = (inp[5]) ? node18780 : node18777;
															assign node18777 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node18780 = (inp[10]) ? node18784 : node18781;
																assign node18781 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node18784 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node18787 = (inp[10]) ? node18789 : 4'b1100;
															assign node18789 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node18792 = (inp[1]) ? node18800 : node18793;
														assign node18793 = (inp[5]) ? node18795 : 4'b1001;
															assign node18795 = (inp[0]) ? 4'b1100 : node18796;
																assign node18796 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node18800 = (inp[10]) ? node18806 : node18801;
															assign node18801 = (inp[0]) ? node18803 : 4'b1000;
																assign node18803 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node18806 = (inp[5]) ? 4'b1001 : node18807;
																assign node18807 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node18811 = (inp[13]) ? node18829 : node18812;
													assign node18812 = (inp[5]) ? node18820 : node18813;
														assign node18813 = (inp[1]) ? node18817 : node18814;
															assign node18814 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node18817 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node18820 = (inp[1]) ? node18824 : node18821;
															assign node18821 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node18824 = (inp[10]) ? 4'b1001 : node18825;
																assign node18825 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node18829 = (inp[5]) ? node18843 : node18830;
														assign node18830 = (inp[0]) ? node18836 : node18831;
															assign node18831 = (inp[1]) ? 4'b1101 : node18832;
																assign node18832 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node18836 = (inp[1]) ? node18840 : node18837;
																assign node18837 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node18840 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node18843 = (inp[1]) ? node18849 : node18844;
															assign node18844 = (inp[0]) ? 4'b1001 : node18845;
																assign node18845 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node18849 = (inp[0]) ? node18851 : 4'b1101;
																assign node18851 = (inp[10]) ? 4'b1100 : 4'b1101;
									assign node18854 = (inp[10]) ? node18986 : node18855;
										assign node18855 = (inp[0]) ? node18925 : node18856;
											assign node18856 = (inp[5]) ? node18882 : node18857;
												assign node18857 = (inp[13]) ? node18865 : node18858;
													assign node18858 = (inp[2]) ? 4'b1110 : node18859;
														assign node18859 = (inp[9]) ? node18861 : 4'b1010;
															assign node18861 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node18865 = (inp[2]) ? node18873 : node18866;
														assign node18866 = (inp[9]) ? 4'b1110 : node18867;
															assign node18867 = (inp[1]) ? 4'b1111 : node18868;
																assign node18868 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node18873 = (inp[11]) ? 4'b1011 : node18874;
															assign node18874 = (inp[9]) ? node18878 : node18875;
																assign node18875 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node18878 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node18882 = (inp[13]) ? node18908 : node18883;
													assign node18883 = (inp[9]) ? node18893 : node18884;
														assign node18884 = (inp[11]) ? node18888 : node18885;
															assign node18885 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node18888 = (inp[2]) ? node18890 : 4'b1011;
																assign node18890 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node18893 = (inp[11]) ? node18901 : node18894;
															assign node18894 = (inp[1]) ? node18898 : node18895;
																assign node18895 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node18898 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node18901 = (inp[2]) ? node18905 : node18902;
																assign node18902 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node18905 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node18908 = (inp[9]) ? node18918 : node18909;
														assign node18909 = (inp[11]) ? node18915 : node18910;
															assign node18910 = (inp[2]) ? node18912 : 4'b1111;
																assign node18912 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node18915 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node18918 = (inp[2]) ? node18922 : node18919;
															assign node18919 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node18922 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node18925 = (inp[2]) ? node18955 : node18926;
												assign node18926 = (inp[13]) ? node18938 : node18927;
													assign node18927 = (inp[1]) ? node18933 : node18928;
														assign node18928 = (inp[5]) ? node18930 : 4'b1010;
															assign node18930 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node18933 = (inp[9]) ? node18935 : 4'b1010;
															assign node18935 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node18938 = (inp[1]) ? node18944 : node18939;
														assign node18939 = (inp[5]) ? 4'b1010 : node18940;
															assign node18940 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node18944 = (inp[9]) ? node18950 : node18945;
															assign node18945 = (inp[11]) ? 4'b1111 : node18946;
																assign node18946 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node18950 = (inp[5]) ? 4'b1110 : node18951;
																assign node18951 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node18955 = (inp[13]) ? node18975 : node18956;
													assign node18956 = (inp[9]) ? node18968 : node18957;
														assign node18957 = (inp[1]) ? node18963 : node18958;
															assign node18958 = (inp[5]) ? 4'b1011 : node18959;
																assign node18959 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node18963 = (inp[11]) ? node18965 : 4'b1111;
																assign node18965 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node18968 = (inp[5]) ? node18972 : node18969;
															assign node18969 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node18972 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node18975 = (inp[5]) ? node18981 : node18976;
														assign node18976 = (inp[9]) ? node18978 : 4'b1011;
															assign node18978 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node18981 = (inp[9]) ? node18983 : 4'b1110;
															assign node18983 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node18986 = (inp[5]) ? node19054 : node18987;
											assign node18987 = (inp[13]) ? node19027 : node18988;
												assign node18988 = (inp[2]) ? node19010 : node18989;
													assign node18989 = (inp[1]) ? node19001 : node18990;
														assign node18990 = (inp[9]) ? node18996 : node18991;
															assign node18991 = (inp[0]) ? 4'b1010 : node18992;
																assign node18992 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18996 = (inp[11]) ? node18998 : 4'b1011;
																assign node18998 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node19001 = (inp[9]) ? node19005 : node19002;
															assign node19002 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node19005 = (inp[11]) ? 4'b1010 : node19006;
																assign node19006 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node19010 = (inp[9]) ? node19020 : node19011;
														assign node19011 = (inp[11]) ? node19017 : node19012;
															assign node19012 = (inp[1]) ? 4'b1110 : node19013;
																assign node19013 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node19017 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node19020 = (inp[0]) ? node19022 : 4'b1111;
															assign node19022 = (inp[1]) ? 4'b1111 : node19023;
																assign node19023 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node19027 = (inp[2]) ? node19041 : node19028;
													assign node19028 = (inp[11]) ? node19034 : node19029;
														assign node19029 = (inp[1]) ? node19031 : 4'b1110;
															assign node19031 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node19034 = (inp[9]) ? node19038 : node19035;
															assign node19035 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node19038 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node19041 = (inp[9]) ? node19049 : node19042;
														assign node19042 = (inp[0]) ? node19044 : 4'b1011;
															assign node19044 = (inp[11]) ? node19046 : 4'b1010;
																assign node19046 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node19049 = (inp[1]) ? 4'b1010 : node19050;
															assign node19050 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node19054 = (inp[9]) ? node19080 : node19055;
												assign node19055 = (inp[13]) ? node19065 : node19056;
													assign node19056 = (inp[1]) ? 4'b1011 : node19057;
														assign node19057 = (inp[2]) ? node19061 : node19058;
															assign node19058 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node19061 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19065 = (inp[0]) ? node19071 : node19066;
														assign node19066 = (inp[11]) ? node19068 : 4'b1111;
															assign node19068 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node19071 = (inp[2]) ? node19077 : node19072;
															assign node19072 = (inp[1]) ? 4'b1110 : node19073;
																assign node19073 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19077 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node19080 = (inp[2]) ? node19094 : node19081;
													assign node19081 = (inp[11]) ? node19085 : node19082;
														assign node19082 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node19085 = (inp[13]) ? node19091 : node19086;
															assign node19086 = (inp[0]) ? 4'b1110 : node19087;
																assign node19087 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node19091 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node19094 = (inp[1]) ? node19100 : node19095;
														assign node19095 = (inp[13]) ? 4'b1111 : node19096;
															assign node19096 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node19100 = (inp[13]) ? node19102 : 4'b1110;
															assign node19102 = (inp[0]) ? 4'b1010 : node19103;
																assign node19103 = (inp[11]) ? 4'b1011 : 4'b1010;
								assign node19107 = (inp[1]) ? node19427 : node19108;
									assign node19108 = (inp[0]) ? node19256 : node19109;
										assign node19109 = (inp[10]) ? node19175 : node19110;
											assign node19110 = (inp[9]) ? node19138 : node19111;
												assign node19111 = (inp[11]) ? node19133 : node19112;
													assign node19112 = (inp[13]) ? node19120 : node19113;
														assign node19113 = (inp[15]) ? node19115 : 4'b1100;
															assign node19115 = (inp[2]) ? 4'b1001 : node19116;
																assign node19116 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node19120 = (inp[15]) ? node19126 : node19121;
															assign node19121 = (inp[5]) ? node19123 : 4'b1001;
																assign node19123 = (inp[2]) ? 4'b1100 : 4'b1001;
															assign node19126 = (inp[5]) ? node19130 : node19127;
																assign node19127 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node19130 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node19133 = (inp[13]) ? 4'b1000 : node19134;
														assign node19134 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node19138 = (inp[11]) ? node19162 : node19139;
													assign node19139 = (inp[5]) ? node19151 : node19140;
														assign node19140 = (inp[15]) ? node19148 : node19141;
															assign node19141 = (inp[2]) ? node19145 : node19142;
																assign node19142 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node19145 = (inp[13]) ? 4'b1000 : 4'b1101;
															assign node19148 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19151 = (inp[13]) ? node19157 : node19152;
															assign node19152 = (inp[2]) ? node19154 : 4'b1100;
																assign node19154 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node19157 = (inp[2]) ? 4'b1101 : node19158;
																assign node19158 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node19162 = (inp[2]) ? node19168 : node19163;
														assign node19163 = (inp[13]) ? 4'b1101 : node19164;
															assign node19164 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node19168 = (inp[5]) ? node19172 : node19169;
															assign node19169 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node19172 = (inp[13]) ? 4'b1100 : 4'b1001;
											assign node19175 = (inp[9]) ? node19211 : node19176;
												assign node19176 = (inp[11]) ? node19190 : node19177;
													assign node19177 = (inp[13]) ? node19185 : node19178;
														assign node19178 = (inp[5]) ? node19182 : node19179;
															assign node19179 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node19182 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node19185 = (inp[2]) ? node19187 : 4'b1101;
															assign node19187 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node19190 = (inp[15]) ? node19198 : node19191;
														assign node19191 = (inp[13]) ? 4'b1101 : node19192;
															assign node19192 = (inp[5]) ? 4'b1101 : node19193;
																assign node19193 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node19198 = (inp[13]) ? node19206 : node19199;
															assign node19199 = (inp[5]) ? node19203 : node19200;
																assign node19200 = (inp[2]) ? 4'b1101 : 4'b1000;
																assign node19203 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node19206 = (inp[5]) ? node19208 : 4'b1001;
																assign node19208 = (inp[2]) ? 4'b1100 : 4'b1001;
												assign node19211 = (inp[11]) ? node19229 : node19212;
													assign node19212 = (inp[2]) ? node19220 : node19213;
														assign node19213 = (inp[13]) ? node19215 : 4'b1100;
															assign node19215 = (inp[15]) ? 4'b1100 : node19216;
																assign node19216 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node19220 = (inp[13]) ? node19226 : node19221;
															assign node19221 = (inp[15]) ? 4'b1001 : node19222;
																assign node19222 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node19226 = (inp[5]) ? 4'b1100 : 4'b1001;
													assign node19229 = (inp[15]) ? node19241 : node19230;
														assign node19230 = (inp[2]) ? node19236 : node19231;
															assign node19231 = (inp[13]) ? node19233 : 4'b1100;
																assign node19233 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node19236 = (inp[13]) ? node19238 : 4'b1000;
																assign node19238 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node19241 = (inp[2]) ? node19249 : node19242;
															assign node19242 = (inp[5]) ? node19246 : node19243;
																assign node19243 = (inp[13]) ? 4'b1100 : 4'b1001;
																assign node19246 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node19249 = (inp[13]) ? node19253 : node19250;
																assign node19250 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node19253 = (inp[5]) ? 4'b1101 : 4'b1000;
										assign node19256 = (inp[10]) ? node19336 : node19257;
											assign node19257 = (inp[9]) ? node19295 : node19258;
												assign node19258 = (inp[11]) ? node19274 : node19259;
													assign node19259 = (inp[5]) ? 4'b1001 : node19260;
														assign node19260 = (inp[15]) ? node19268 : node19261;
															assign node19261 = (inp[2]) ? node19265 : node19262;
																assign node19262 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node19265 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node19268 = (inp[13]) ? node19270 : 4'b1101;
																assign node19270 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node19274 = (inp[13]) ? node19288 : node19275;
														assign node19275 = (inp[15]) ? node19281 : node19276;
															assign node19276 = (inp[2]) ? 4'b1100 : node19277;
																assign node19277 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node19281 = (inp[5]) ? node19285 : node19282;
																assign node19282 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node19285 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node19288 = (inp[15]) ? node19292 : node19289;
															assign node19289 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19292 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node19295 = (inp[11]) ? node19317 : node19296;
													assign node19296 = (inp[2]) ? node19308 : node19297;
														assign node19297 = (inp[15]) ? node19303 : node19298;
															assign node19298 = (inp[13]) ? node19300 : 4'b1000;
																assign node19300 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node19303 = (inp[13]) ? node19305 : 4'b1100;
																assign node19305 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node19308 = (inp[13]) ? node19312 : node19309;
															assign node19309 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node19312 = (inp[5]) ? node19314 : 4'b1000;
																assign node19314 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node19317 = (inp[13]) ? node19331 : node19318;
														assign node19318 = (inp[15]) ? node19326 : node19319;
															assign node19319 = (inp[2]) ? node19323 : node19320;
																assign node19320 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node19323 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19326 = (inp[2]) ? node19328 : 4'b1100;
																assign node19328 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node19331 = (inp[5]) ? node19333 : 4'b1001;
															assign node19333 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node19336 = (inp[9]) ? node19382 : node19337;
												assign node19337 = (inp[11]) ? node19361 : node19338;
													assign node19338 = (inp[15]) ? node19350 : node19339;
														assign node19339 = (inp[5]) ? node19345 : node19340;
															assign node19340 = (inp[2]) ? 4'b1000 : node19341;
																assign node19341 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node19345 = (inp[2]) ? 4'b1100 : node19346;
																assign node19346 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node19350 = (inp[5]) ? node19354 : node19351;
															assign node19351 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node19354 = (inp[2]) ? node19358 : node19355;
																assign node19355 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node19358 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node19361 = (inp[13]) ? node19373 : node19362;
														assign node19362 = (inp[15]) ? node19366 : node19363;
															assign node19363 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node19366 = (inp[5]) ? node19370 : node19367;
																assign node19367 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node19370 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node19373 = (inp[5]) ? node19379 : node19374;
															assign node19374 = (inp[15]) ? node19376 : 4'b1000;
																assign node19376 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node19379 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node19382 = (inp[11]) ? node19402 : node19383;
													assign node19383 = (inp[15]) ? node19397 : node19384;
														assign node19384 = (inp[2]) ? node19392 : node19385;
															assign node19385 = (inp[5]) ? node19389 : node19386;
																assign node19386 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node19389 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node19392 = (inp[5]) ? 4'b1001 : node19393;
																assign node19393 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node19397 = (inp[2]) ? node19399 : 4'b1000;
															assign node19399 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node19402 = (inp[5]) ? node19414 : node19403;
														assign node19403 = (inp[2]) ? node19407 : node19404;
															assign node19404 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node19407 = (inp[13]) ? node19411 : node19408;
																assign node19408 = (inp[15]) ? 4'b1101 : 4'b1100;
																assign node19411 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node19414 = (inp[15]) ? node19422 : node19415;
															assign node19415 = (inp[2]) ? node19419 : node19416;
																assign node19416 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node19419 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node19422 = (inp[13]) ? node19424 : 4'b1001;
																assign node19424 = (inp[2]) ? 4'b1100 : 4'b1000;
									assign node19427 = (inp[2]) ? node19525 : node19428;
										assign node19428 = (inp[13]) ? node19504 : node19429;
											assign node19429 = (inp[5]) ? node19459 : node19430;
												assign node19430 = (inp[10]) ? node19442 : node19431;
													assign node19431 = (inp[15]) ? node19433 : 4'b1000;
														assign node19433 = (inp[9]) ? node19437 : node19434;
															assign node19434 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node19437 = (inp[11]) ? node19439 : 4'b1000;
																assign node19439 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node19442 = (inp[0]) ? node19452 : node19443;
														assign node19443 = (inp[9]) ? 4'b1001 : node19444;
															assign node19444 = (inp[11]) ? node19448 : node19445;
																assign node19445 = (inp[15]) ? 4'b1000 : 4'b1001;
																assign node19448 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node19452 = (inp[15]) ? node19456 : node19453;
															assign node19453 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node19456 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node19459 = (inp[15]) ? node19479 : node19460;
													assign node19460 = (inp[11]) ? node19470 : node19461;
														assign node19461 = (inp[0]) ? node19463 : 4'b1001;
															assign node19463 = (inp[9]) ? node19467 : node19464;
																assign node19464 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node19467 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node19470 = (inp[0]) ? 4'b1001 : node19471;
															assign node19471 = (inp[10]) ? node19475 : node19472;
																assign node19472 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node19475 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node19479 = (inp[0]) ? node19489 : node19480;
														assign node19480 = (inp[9]) ? 4'b1001 : node19481;
															assign node19481 = (inp[10]) ? node19485 : node19482;
																assign node19482 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node19485 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19489 = (inp[11]) ? node19497 : node19490;
															assign node19490 = (inp[9]) ? node19494 : node19491;
																assign node19491 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node19494 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node19497 = (inp[10]) ? node19501 : node19498;
																assign node19498 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node19501 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node19504 = (inp[10]) ? node19516 : node19505;
												assign node19505 = (inp[9]) ? node19511 : node19506;
													assign node19506 = (inp[0]) ? 4'b1100 : node19507;
														assign node19507 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node19511 = (inp[11]) ? node19513 : 4'b1101;
														assign node19513 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node19516 = (inp[9]) ? node19522 : node19517;
													assign node19517 = (inp[0]) ? 4'b1101 : node19518;
														assign node19518 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node19522 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node19525 = (inp[13]) ? node19581 : node19526;
											assign node19526 = (inp[9]) ? node19554 : node19527;
												assign node19527 = (inp[0]) ? node19539 : node19528;
													assign node19528 = (inp[11]) ? node19534 : node19529;
														assign node19529 = (inp[10]) ? node19531 : 4'b1101;
															assign node19531 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node19534 = (inp[15]) ? node19536 : 4'b1101;
															assign node19536 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node19539 = (inp[15]) ? node19547 : node19540;
														assign node19540 = (inp[11]) ? node19544 : node19541;
															assign node19541 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node19544 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node19547 = (inp[10]) ? node19551 : node19548;
															assign node19548 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19551 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19554 = (inp[11]) ? node19574 : node19555;
													assign node19555 = (inp[10]) ? node19563 : node19556;
														assign node19556 = (inp[0]) ? node19560 : node19557;
															assign node19557 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node19560 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node19563 = (inp[5]) ? node19569 : node19564;
															assign node19564 = (inp[0]) ? 4'b1100 : node19565;
																assign node19565 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node19569 = (inp[0]) ? node19571 : 4'b1101;
																assign node19571 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node19574 = (inp[15]) ? node19578 : node19575;
														assign node19575 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node19578 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node19581 = (inp[11]) ? node19589 : node19582;
												assign node19582 = (inp[10]) ? node19586 : node19583;
													assign node19583 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node19586 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node19589 = (inp[15]) ? node19597 : node19590;
													assign node19590 = (inp[10]) ? 4'b1000 : node19591;
														assign node19591 = (inp[9]) ? node19593 : 4'b1001;
															assign node19593 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node19597 = (inp[9]) ? node19605 : node19598;
														assign node19598 = (inp[0]) ? node19602 : node19599;
															assign node19599 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node19602 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node19605 = (inp[10]) ? 4'b1001 : 4'b1000;
					assign node19608 = (inp[4]) ? node21728 : node19609;
						assign node19609 = (inp[11]) ? node20629 : node19610;
							assign node19610 = (inp[2]) ? node20164 : node19611;
								assign node19611 = (inp[13]) ? node19885 : node19612;
									assign node19612 = (inp[7]) ? node19746 : node19613;
										assign node19613 = (inp[12]) ? node19675 : node19614;
											assign node19614 = (inp[15]) ? node19640 : node19615;
												assign node19615 = (inp[1]) ? node19629 : node19616;
													assign node19616 = (inp[5]) ? node19626 : node19617;
														assign node19617 = (inp[9]) ? 4'b0011 : node19618;
															assign node19618 = (inp[10]) ? node19622 : node19619;
																assign node19619 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node19622 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node19626 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node19629 = (inp[10]) ? 4'b0110 : node19630;
														assign node19630 = (inp[0]) ? node19634 : node19631;
															assign node19631 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node19634 = (inp[5]) ? 4'b0110 : node19635;
																assign node19635 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node19640 = (inp[5]) ? node19656 : node19641;
													assign node19641 = (inp[9]) ? node19649 : node19642;
														assign node19642 = (inp[10]) ? node19644 : 4'b0001;
															assign node19644 = (inp[1]) ? node19646 : 4'b0000;
																assign node19646 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19649 = (inp[1]) ? node19651 : 4'b0000;
															assign node19651 = (inp[0]) ? 4'b0000 : node19652;
																assign node19652 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node19656 = (inp[1]) ? node19662 : node19657;
														assign node19657 = (inp[10]) ? 4'b0000 : node19658;
															assign node19658 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node19662 = (inp[9]) ? node19670 : node19663;
															assign node19663 = (inp[0]) ? node19667 : node19664;
																assign node19664 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node19667 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node19670 = (inp[10]) ? 4'b0100 : node19671;
																assign node19671 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node19675 = (inp[15]) ? node19717 : node19676;
												assign node19676 = (inp[5]) ? node19698 : node19677;
													assign node19677 = (inp[1]) ? node19689 : node19678;
														assign node19678 = (inp[10]) ? node19684 : node19679;
															assign node19679 = (inp[0]) ? 4'b0100 : node19680;
																assign node19680 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node19684 = (inp[9]) ? 4'b0101 : node19685;
																assign node19685 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node19689 = (inp[0]) ? node19691 : 4'b0000;
															assign node19691 = (inp[10]) ? node19695 : node19692;
																assign node19692 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node19695 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node19698 = (inp[10]) ? node19708 : node19699;
														assign node19699 = (inp[9]) ? node19705 : node19700;
															assign node19700 = (inp[1]) ? node19702 : 4'b0000;
																assign node19702 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node19705 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node19708 = (inp[9]) ? node19714 : node19709;
															assign node19709 = (inp[0]) ? node19711 : 4'b0001;
																assign node19711 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node19714 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node19717 = (inp[5]) ? node19735 : node19718;
													assign node19718 = (inp[1]) ? node19726 : node19719;
														assign node19719 = (inp[9]) ? node19721 : 4'b0111;
															assign node19721 = (inp[10]) ? 4'b0110 : node19722;
																assign node19722 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node19726 = (inp[0]) ? 4'b0010 : node19727;
															assign node19727 = (inp[9]) ? node19731 : node19728;
																assign node19728 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node19731 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node19735 = (inp[0]) ? node19737 : 4'b0011;
														assign node19737 = (inp[1]) ? node19743 : node19738;
															assign node19738 = (inp[10]) ? 4'b0010 : node19739;
																assign node19739 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node19743 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node19746 = (inp[1]) ? node19812 : node19747;
											assign node19747 = (inp[12]) ? node19781 : node19748;
												assign node19748 = (inp[15]) ? node19766 : node19749;
													assign node19749 = (inp[5]) ? node19759 : node19750;
														assign node19750 = (inp[10]) ? 4'b0101 : node19751;
															assign node19751 = (inp[0]) ? node19755 : node19752;
																assign node19752 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node19755 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node19759 = (inp[0]) ? 4'b0001 : node19760;
															assign node19760 = (inp[10]) ? node19762 : 4'b0000;
																assign node19762 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node19766 = (inp[5]) ? node19774 : node19767;
														assign node19767 = (inp[9]) ? node19771 : node19768;
															assign node19768 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node19771 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node19774 = (inp[9]) ? node19778 : node19775;
															assign node19775 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node19778 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node19781 = (inp[15]) ? node19793 : node19782;
													assign node19782 = (inp[0]) ? node19786 : node19783;
														assign node19783 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node19786 = (inp[5]) ? 4'b0111 : node19787;
															assign node19787 = (inp[10]) ? 4'b0111 : node19788;
																assign node19788 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node19793 = (inp[5]) ? node19809 : node19794;
														assign node19794 = (inp[9]) ? node19802 : node19795;
															assign node19795 = (inp[10]) ? node19799 : node19796;
																assign node19796 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node19799 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node19802 = (inp[0]) ? node19806 : node19803;
																assign node19803 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node19806 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node19809 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node19812 = (inp[12]) ? node19846 : node19813;
												assign node19813 = (inp[15]) ? node19827 : node19814;
													assign node19814 = (inp[5]) ? node19822 : node19815;
														assign node19815 = (inp[0]) ? node19817 : 4'b0000;
															assign node19817 = (inp[9]) ? 4'b0000 : node19818;
																assign node19818 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node19822 = (inp[9]) ? 4'b0001 : node19823;
															assign node19823 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node19827 = (inp[10]) ? node19837 : node19828;
														assign node19828 = (inp[9]) ? node19832 : node19829;
															assign node19829 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node19832 = (inp[5]) ? 4'b0111 : node19833;
																assign node19833 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node19837 = (inp[9]) ? node19841 : node19838;
															assign node19838 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node19841 = (inp[0]) ? 4'b0110 : node19842;
																assign node19842 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node19846 = (inp[15]) ? node19868 : node19847;
													assign node19847 = (inp[5]) ? node19861 : node19848;
														assign node19848 = (inp[10]) ? node19854 : node19849;
															assign node19849 = (inp[9]) ? 4'b0110 : node19850;
																assign node19850 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node19854 = (inp[9]) ? node19858 : node19855;
																assign node19855 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node19858 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node19861 = (inp[0]) ? node19863 : 4'b0010;
															assign node19863 = (inp[10]) ? 4'b0011 : node19864;
																assign node19864 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node19868 = (inp[9]) ? node19874 : node19869;
														assign node19869 = (inp[10]) ? 4'b0001 : node19870;
															assign node19870 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node19874 = (inp[10]) ? node19880 : node19875;
															assign node19875 = (inp[0]) ? 4'b0001 : node19876;
																assign node19876 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node19880 = (inp[0]) ? 4'b0000 : node19881;
																assign node19881 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node19885 = (inp[12]) ? node20017 : node19886;
										assign node19886 = (inp[5]) ? node19956 : node19887;
											assign node19887 = (inp[1]) ? node19925 : node19888;
												assign node19888 = (inp[7]) ? node19908 : node19889;
													assign node19889 = (inp[15]) ? node19897 : node19890;
														assign node19890 = (inp[9]) ? node19894 : node19891;
															assign node19891 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node19894 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node19897 = (inp[0]) ? node19903 : node19898;
															assign node19898 = (inp[10]) ? 4'b0100 : node19899;
																assign node19899 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node19903 = (inp[10]) ? node19905 : 4'b0100;
																assign node19905 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node19908 = (inp[15]) ? node19914 : node19909;
														assign node19909 = (inp[0]) ? 4'b0001 : node19910;
															assign node19910 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node19914 = (inp[9]) ? node19920 : node19915;
															assign node19915 = (inp[10]) ? node19917 : 4'b0111;
																assign node19917 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node19920 = (inp[0]) ? node19922 : 4'b0110;
																assign node19922 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node19925 = (inp[10]) ? node19935 : node19926;
													assign node19926 = (inp[0]) ? 4'b0101 : node19927;
														assign node19927 = (inp[7]) ? node19931 : node19928;
															assign node19928 = (inp[15]) ? 4'b0101 : 4'b0010;
															assign node19931 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node19935 = (inp[15]) ? node19945 : node19936;
														assign node19936 = (inp[7]) ? node19940 : node19937;
															assign node19937 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node19940 = (inp[0]) ? 4'b0100 : node19941;
																assign node19941 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node19945 = (inp[7]) ? node19949 : node19946;
															assign node19946 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node19949 = (inp[0]) ? node19953 : node19950;
																assign node19950 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node19953 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node19956 = (inp[7]) ? node19988 : node19957;
												assign node19957 = (inp[15]) ? node19971 : node19958;
													assign node19958 = (inp[9]) ? node19966 : node19959;
														assign node19959 = (inp[10]) ? 4'b0010 : node19960;
															assign node19960 = (inp[0]) ? node19962 : 4'b0011;
																assign node19962 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node19966 = (inp[1]) ? 4'b0011 : node19967;
															assign node19967 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node19971 = (inp[1]) ? node19979 : node19972;
														assign node19972 = (inp[10]) ? 4'b0101 : node19973;
															assign node19973 = (inp[0]) ? 4'b0100 : node19974;
																assign node19974 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node19979 = (inp[10]) ? node19981 : 4'b0000;
															assign node19981 = (inp[0]) ? node19985 : node19982;
																assign node19982 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node19985 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node19988 = (inp[15]) ? node20004 : node19989;
													assign node19989 = (inp[10]) ? node19997 : node19990;
														assign node19990 = (inp[1]) ? 4'b0101 : node19991;
															assign node19991 = (inp[0]) ? node19993 : 4'b0101;
																assign node19993 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node19997 = (inp[9]) ? node20001 : node19998;
															assign node19998 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node20001 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node20004 = (inp[0]) ? 4'b0011 : node20005;
														assign node20005 = (inp[1]) ? node20011 : node20006;
															assign node20006 = (inp[9]) ? node20008 : 4'b0011;
																assign node20008 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node20011 = (inp[10]) ? 4'b0010 : node20012;
																assign node20012 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node20017 = (inp[1]) ? node20087 : node20018;
											assign node20018 = (inp[5]) ? node20050 : node20019;
												assign node20019 = (inp[0]) ? node20031 : node20020;
													assign node20020 = (inp[9]) ? node20024 : node20021;
														assign node20021 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node20024 = (inp[10]) ? node20026 : 4'b0000;
															assign node20026 = (inp[7]) ? node20028 : 4'b0001;
																assign node20028 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node20031 = (inp[9]) ? node20043 : node20032;
														assign node20032 = (inp[15]) ? node20036 : node20033;
															assign node20033 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node20036 = (inp[7]) ? node20040 : node20037;
																assign node20037 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node20040 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node20043 = (inp[10]) ? node20045 : 4'b0001;
															assign node20045 = (inp[15]) ? node20047 : 4'b0000;
																assign node20047 = (inp[7]) ? 4'b0000 : 4'b0011;
												assign node20050 = (inp[15]) ? node20068 : node20051;
													assign node20051 = (inp[7]) ? node20061 : node20052;
														assign node20052 = (inp[10]) ? 4'b0101 : node20053;
															assign node20053 = (inp[0]) ? node20057 : node20054;
																assign node20054 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node20057 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node20061 = (inp[0]) ? 4'b0011 : node20062;
															assign node20062 = (inp[10]) ? node20064 : 4'b0011;
																assign node20064 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node20068 = (inp[7]) ? node20074 : node20069;
														assign node20069 = (inp[0]) ? 4'b0110 : node20070;
															assign node20070 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node20074 = (inp[9]) ? node20082 : node20075;
															assign node20075 = (inp[10]) ? node20079 : node20076;
																assign node20076 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node20079 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node20082 = (inp[10]) ? node20084 : 4'b0100;
																assign node20084 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node20087 = (inp[5]) ? node20119 : node20088;
												assign node20088 = (inp[7]) ? node20106 : node20089;
													assign node20089 = (inp[15]) ? node20099 : node20090;
														assign node20090 = (inp[9]) ? 4'b0100 : node20091;
															assign node20091 = (inp[10]) ? node20095 : node20092;
																assign node20092 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node20095 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node20099 = (inp[9]) ? node20103 : node20100;
															assign node20100 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node20103 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node20106 = (inp[15]) ? node20112 : node20107;
														assign node20107 = (inp[9]) ? node20109 : 4'b0011;
															assign node20109 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node20112 = (inp[0]) ? 4'b0101 : node20113;
															assign node20113 = (inp[10]) ? node20115 : 4'b0100;
																assign node20115 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node20119 = (inp[10]) ? node20143 : node20120;
													assign node20120 = (inp[7]) ? node20130 : node20121;
														assign node20121 = (inp[15]) ? node20125 : node20122;
															assign node20122 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node20125 = (inp[9]) ? node20127 : 4'b0111;
																assign node20127 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node20130 = (inp[15]) ? node20136 : node20131;
															assign node20131 = (inp[9]) ? 4'b0110 : node20132;
																assign node20132 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node20136 = (inp[0]) ? node20140 : node20137;
																assign node20137 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node20140 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node20143 = (inp[0]) ? node20153 : node20144;
														assign node20144 = (inp[9]) ? node20146 : 4'b0101;
															assign node20146 = (inp[15]) ? node20150 : node20147;
																assign node20147 = (inp[7]) ? 4'b0110 : 4'b0100;
																assign node20150 = (inp[7]) ? 4'b0100 : 4'b0110;
														assign node20153 = (inp[9]) ? node20159 : node20154;
															assign node20154 = (inp[15]) ? node20156 : 4'b0110;
																assign node20156 = (inp[7]) ? 4'b0100 : 4'b0110;
															assign node20159 = (inp[7]) ? 4'b0111 : node20160;
																assign node20160 = (inp[15]) ? 4'b0111 : 4'b0100;
								assign node20164 = (inp[13]) ? node20398 : node20165;
									assign node20165 = (inp[7]) ? node20287 : node20166;
										assign node20166 = (inp[12]) ? node20222 : node20167;
											assign node20167 = (inp[15]) ? node20197 : node20168;
												assign node20168 = (inp[10]) ? node20180 : node20169;
													assign node20169 = (inp[5]) ? node20173 : node20170;
														assign node20170 = (inp[0]) ? 4'b0010 : 4'b0110;
														assign node20173 = (inp[0]) ? node20175 : 4'b0010;
															assign node20175 = (inp[1]) ? 4'b0010 : node20176;
																assign node20176 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node20180 = (inp[5]) ? node20188 : node20181;
														assign node20181 = (inp[1]) ? node20183 : 4'b0111;
															assign node20183 = (inp[0]) ? 4'b0011 : node20184;
																assign node20184 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node20188 = (inp[9]) ? node20194 : node20189;
															assign node20189 = (inp[1]) ? 4'b0010 : node20190;
																assign node20190 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20194 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node20197 = (inp[1]) ? node20211 : node20198;
													assign node20198 = (inp[9]) ? node20204 : node20199;
														assign node20199 = (inp[10]) ? 4'b0101 : node20200;
															assign node20200 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node20204 = (inp[10]) ? 4'b0100 : node20205;
															assign node20205 = (inp[5]) ? node20207 : 4'b0101;
																assign node20207 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node20211 = (inp[5]) ? node20217 : node20212;
														assign node20212 = (inp[9]) ? 4'b0101 : node20213;
															assign node20213 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node20217 = (inp[10]) ? 4'b0001 : node20218;
															assign node20218 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node20222 = (inp[15]) ? node20254 : node20223;
												assign node20223 = (inp[1]) ? node20235 : node20224;
													assign node20224 = (inp[9]) ? node20230 : node20225;
														assign node20225 = (inp[0]) ? 4'b0001 : node20226;
															assign node20226 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node20230 = (inp[10]) ? node20232 : 4'b0100;
															assign node20232 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node20235 = (inp[10]) ? node20247 : node20236;
														assign node20236 = (inp[9]) ? node20242 : node20237;
															assign node20237 = (inp[5]) ? 4'b0100 : node20238;
																assign node20238 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node20242 = (inp[0]) ? node20244 : 4'b0101;
																assign node20244 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node20247 = (inp[9]) ? node20249 : 4'b0101;
															assign node20249 = (inp[0]) ? node20251 : 4'b0100;
																assign node20251 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node20254 = (inp[1]) ? node20272 : node20255;
													assign node20255 = (inp[5]) ? node20265 : node20256;
														assign node20256 = (inp[10]) ? node20258 : 4'b0010;
															assign node20258 = (inp[9]) ? node20262 : node20259;
																assign node20259 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node20262 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node20265 = (inp[0]) ? node20267 : 4'b0111;
															assign node20267 = (inp[9]) ? 4'b0110 : node20268;
																assign node20268 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node20272 = (inp[10]) ? node20278 : node20273;
														assign node20273 = (inp[9]) ? node20275 : 4'b0110;
															assign node20275 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node20278 = (inp[9]) ? node20282 : node20279;
															assign node20279 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node20282 = (inp[0]) ? 4'b0110 : node20283;
																assign node20283 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node20287 = (inp[1]) ? node20341 : node20288;
											assign node20288 = (inp[12]) ? node20314 : node20289;
												assign node20289 = (inp[15]) ? node20301 : node20290;
													assign node20290 = (inp[5]) ? node20292 : 4'b0001;
														assign node20292 = (inp[0]) ? 4'b0101 : node20293;
															assign node20293 = (inp[10]) ? node20297 : node20294;
																assign node20294 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node20297 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node20301 = (inp[5]) ? node20309 : node20302;
														assign node20302 = (inp[9]) ? node20304 : 4'b0110;
															assign node20304 = (inp[10]) ? node20306 : 4'b0110;
																assign node20306 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node20309 = (inp[10]) ? node20311 : 4'b0011;
															assign node20311 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node20314 = (inp[15]) ? node20330 : node20315;
													assign node20315 = (inp[9]) ? node20323 : node20316;
														assign node20316 = (inp[10]) ? node20320 : node20317;
															assign node20317 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node20320 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node20323 = (inp[10]) ? node20327 : node20324;
															assign node20324 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20327 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node20330 = (inp[5]) ? node20338 : node20331;
														assign node20331 = (inp[0]) ? 4'b0001 : node20332;
															assign node20332 = (inp[10]) ? 4'b0001 : node20333;
																assign node20333 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node20338 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node20341 = (inp[10]) ? node20363 : node20342;
												assign node20342 = (inp[15]) ? node20354 : node20343;
													assign node20343 = (inp[12]) ? node20349 : node20344;
														assign node20344 = (inp[0]) ? node20346 : 4'b0101;
															assign node20346 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node20349 = (inp[9]) ? node20351 : 4'b0010;
															assign node20351 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node20354 = (inp[12]) ? node20360 : node20355;
														assign node20355 = (inp[9]) ? 4'b0010 : node20356;
															assign node20356 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node20360 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node20363 = (inp[15]) ? node20383 : node20364;
													assign node20364 = (inp[12]) ? node20372 : node20365;
														assign node20365 = (inp[9]) ? 4'b0100 : node20366;
															assign node20366 = (inp[5]) ? 4'b0101 : node20367;
																assign node20367 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node20372 = (inp[5]) ? node20378 : node20373;
															assign node20373 = (inp[9]) ? 4'b0010 : node20374;
																assign node20374 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20378 = (inp[0]) ? 4'b0110 : node20379;
																assign node20379 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node20383 = (inp[12]) ? node20393 : node20384;
														assign node20384 = (inp[0]) ? 4'b0011 : node20385;
															assign node20385 = (inp[5]) ? node20389 : node20386;
																assign node20386 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node20389 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node20393 = (inp[9]) ? 4'b0101 : node20394;
															assign node20394 = (inp[5]) ? 4'b0101 : 4'b0100;
									assign node20398 = (inp[7]) ? node20518 : node20399;
										assign node20399 = (inp[12]) ? node20447 : node20400;
											assign node20400 = (inp[15]) ? node20428 : node20401;
												assign node20401 = (inp[5]) ? node20421 : node20402;
													assign node20402 = (inp[1]) ? node20410 : node20403;
														assign node20403 = (inp[10]) ? node20407 : node20404;
															assign node20404 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node20407 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node20410 = (inp[0]) ? node20416 : node20411;
															assign node20411 = (inp[9]) ? 4'b0111 : node20412;
																assign node20412 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node20416 = (inp[10]) ? 4'b0110 : node20417;
																assign node20417 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node20421 = (inp[10]) ? node20425 : node20422;
														assign node20422 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node20425 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node20428 = (inp[5]) ? node20438 : node20429;
													assign node20429 = (inp[9]) ? 4'b0001 : node20430;
														assign node20430 = (inp[1]) ? node20434 : node20431;
															assign node20431 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node20434 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node20438 = (inp[1]) ? node20440 : 4'b0001;
														assign node20440 = (inp[9]) ? node20444 : node20441;
															assign node20441 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node20444 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node20447 = (inp[15]) ? node20487 : node20448;
												assign node20448 = (inp[1]) ? node20470 : node20449;
													assign node20449 = (inp[5]) ? node20463 : node20450;
														assign node20450 = (inp[0]) ? node20458 : node20451;
															assign node20451 = (inp[9]) ? node20455 : node20452;
																assign node20452 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node20455 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node20458 = (inp[9]) ? 4'b0100 : node20459;
																assign node20459 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node20463 = (inp[10]) ? node20465 : 4'b0000;
															assign node20465 = (inp[9]) ? node20467 : 4'b0001;
																assign node20467 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node20470 = (inp[10]) ? node20476 : node20471;
														assign node20471 = (inp[9]) ? node20473 : 4'b0001;
															assign node20473 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20476 = (inp[9]) ? node20482 : node20477;
															assign node20477 = (inp[5]) ? 4'b0000 : node20478;
																assign node20478 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20482 = (inp[5]) ? 4'b0001 : node20483;
																assign node20483 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node20487 = (inp[1]) ? node20501 : node20488;
													assign node20488 = (inp[5]) ? node20496 : node20489;
														assign node20489 = (inp[10]) ? node20493 : node20490;
															assign node20490 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node20493 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node20496 = (inp[10]) ? node20498 : 4'b0010;
															assign node20498 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node20501 = (inp[5]) ? node20509 : node20502;
														assign node20502 = (inp[9]) ? node20506 : node20503;
															assign node20503 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node20506 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node20509 = (inp[0]) ? 4'b0011 : node20510;
															assign node20510 = (inp[9]) ? node20514 : node20511;
																assign node20511 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node20514 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node20518 = (inp[5]) ? node20576 : node20519;
											assign node20519 = (inp[9]) ? node20545 : node20520;
												assign node20520 = (inp[10]) ? node20530 : node20521;
													assign node20521 = (inp[15]) ? node20523 : 4'b0111;
														assign node20523 = (inp[12]) ? 4'b0001 : node20524;
															assign node20524 = (inp[1]) ? 4'b0111 : node20525;
																assign node20525 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node20530 = (inp[15]) ? node20536 : node20531;
														assign node20531 = (inp[12]) ? 4'b0110 : node20532;
															assign node20532 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node20536 = (inp[12]) ? node20542 : node20537;
															assign node20537 = (inp[1]) ? 4'b0110 : node20538;
																assign node20538 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20542 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node20545 = (inp[10]) ? node20561 : node20546;
													assign node20546 = (inp[12]) ? node20556 : node20547;
														assign node20547 = (inp[15]) ? node20553 : node20548;
															assign node20548 = (inp[0]) ? node20550 : 4'b0001;
																assign node20550 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node20553 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node20556 = (inp[15]) ? 4'b0100 : node20557;
															assign node20557 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node20561 = (inp[1]) ? node20567 : node20562;
														assign node20562 = (inp[15]) ? 4'b0101 : node20563;
															assign node20563 = (inp[12]) ? 4'b0110 : 4'b0101;
														assign node20567 = (inp[15]) ? node20573 : node20568;
															assign node20568 = (inp[12]) ? 4'b0111 : node20569;
																assign node20569 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20573 = (inp[12]) ? 4'b0001 : 4'b0111;
											assign node20576 = (inp[15]) ? node20600 : node20577;
												assign node20577 = (inp[12]) ? node20593 : node20578;
													assign node20578 = (inp[1]) ? node20588 : node20579;
														assign node20579 = (inp[0]) ? node20581 : 4'b0001;
															assign node20581 = (inp[10]) ? node20585 : node20582;
																assign node20582 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node20585 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node20588 = (inp[0]) ? 4'b0000 : node20589;
															assign node20589 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node20593 = (inp[1]) ? 4'b0010 : node20594;
														assign node20594 = (inp[10]) ? 4'b0110 : node20595;
															assign node20595 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node20600 = (inp[12]) ? node20618 : node20601;
													assign node20601 = (inp[0]) ? node20609 : node20602;
														assign node20602 = (inp[9]) ? node20604 : 4'b0111;
															assign node20604 = (inp[1]) ? node20606 : 4'b0111;
																assign node20606 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node20609 = (inp[1]) ? node20611 : 4'b0110;
															assign node20611 = (inp[9]) ? node20615 : node20612;
																assign node20612 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node20615 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node20618 = (inp[0]) ? node20624 : node20619;
														assign node20619 = (inp[10]) ? node20621 : 4'b0001;
															assign node20621 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node20624 = (inp[9]) ? 4'b0000 : node20625;
															assign node20625 = (inp[10]) ? 4'b0001 : 4'b0000;
							assign node20629 = (inp[13]) ? node21173 : node20630;
								assign node20630 = (inp[2]) ? node20916 : node20631;
									assign node20631 = (inp[1]) ? node20765 : node20632;
										assign node20632 = (inp[7]) ? node20702 : node20633;
											assign node20633 = (inp[12]) ? node20667 : node20634;
												assign node20634 = (inp[15]) ? node20650 : node20635;
													assign node20635 = (inp[5]) ? node20643 : node20636;
														assign node20636 = (inp[9]) ? node20640 : node20637;
															assign node20637 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node20640 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node20643 = (inp[0]) ? 4'b0111 : node20644;
															assign node20644 = (inp[9]) ? 4'b0110 : node20645;
																assign node20645 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node20650 = (inp[0]) ? node20656 : node20651;
														assign node20651 = (inp[9]) ? node20653 : 4'b0001;
															assign node20653 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node20656 = (inp[5]) ? node20662 : node20657;
															assign node20657 = (inp[9]) ? 4'b0000 : node20658;
																assign node20658 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node20662 = (inp[10]) ? node20664 : 4'b0001;
																assign node20664 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node20667 = (inp[5]) ? node20681 : node20668;
													assign node20668 = (inp[15]) ? node20676 : node20669;
														assign node20669 = (inp[10]) ? node20673 : node20670;
															assign node20670 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node20673 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node20676 = (inp[10]) ? node20678 : 4'b0110;
															assign node20678 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node20681 = (inp[15]) ? node20691 : node20682;
														assign node20682 = (inp[10]) ? node20684 : 4'b0000;
															assign node20684 = (inp[0]) ? node20688 : node20685;
																assign node20685 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node20688 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node20691 = (inp[10]) ? node20697 : node20692;
															assign node20692 = (inp[9]) ? 4'b0010 : node20693;
																assign node20693 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20697 = (inp[9]) ? node20699 : 4'b0011;
																assign node20699 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node20702 = (inp[12]) ? node20736 : node20703;
												assign node20703 = (inp[15]) ? node20717 : node20704;
													assign node20704 = (inp[5]) ? node20710 : node20705;
														assign node20705 = (inp[10]) ? 4'b0100 : node20706;
															assign node20706 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node20710 = (inp[9]) ? node20712 : 4'b0000;
															assign node20712 = (inp[0]) ? 4'b0001 : node20713;
																assign node20713 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node20717 = (inp[5]) ? node20727 : node20718;
														assign node20718 = (inp[10]) ? node20720 : 4'b0011;
															assign node20720 = (inp[0]) ? node20724 : node20721;
																assign node20721 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node20724 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node20727 = (inp[9]) ? 4'b0110 : node20728;
															assign node20728 = (inp[10]) ? node20732 : node20729;
																assign node20729 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node20732 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node20736 = (inp[15]) ? node20750 : node20737;
													assign node20737 = (inp[10]) ? node20743 : node20738;
														assign node20738 = (inp[9]) ? 4'b0110 : node20739;
															assign node20739 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node20743 = (inp[9]) ? node20745 : 4'b0110;
															assign node20745 = (inp[5]) ? 4'b0111 : node20746;
																assign node20746 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node20750 = (inp[5]) ? node20758 : node20751;
														assign node20751 = (inp[9]) ? node20755 : node20752;
															assign node20752 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node20755 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node20758 = (inp[0]) ? node20760 : 4'b0001;
															assign node20760 = (inp[9]) ? node20762 : 4'b0000;
																assign node20762 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node20765 = (inp[12]) ? node20851 : node20766;
											assign node20766 = (inp[5]) ? node20812 : node20767;
												assign node20767 = (inp[7]) ? node20789 : node20768;
													assign node20768 = (inp[15]) ? node20776 : node20769;
														assign node20769 = (inp[0]) ? node20771 : 4'b0110;
															assign node20771 = (inp[10]) ? 4'b0110 : node20772;
																assign node20772 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node20776 = (inp[0]) ? node20782 : node20777;
															assign node20777 = (inp[10]) ? 4'b0000 : node20778;
																assign node20778 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node20782 = (inp[9]) ? node20786 : node20783;
																assign node20783 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node20786 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node20789 = (inp[15]) ? node20805 : node20790;
														assign node20790 = (inp[0]) ? node20798 : node20791;
															assign node20791 = (inp[10]) ? node20795 : node20792;
																assign node20792 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node20795 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node20798 = (inp[10]) ? node20802 : node20799;
																assign node20799 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node20802 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node20805 = (inp[0]) ? 4'b0110 : node20806;
															assign node20806 = (inp[9]) ? node20808 : 4'b0111;
																assign node20808 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node20812 = (inp[15]) ? node20834 : node20813;
													assign node20813 = (inp[7]) ? node20825 : node20814;
														assign node20814 = (inp[10]) ? node20820 : node20815;
															assign node20815 = (inp[0]) ? node20817 : 4'b0111;
																assign node20817 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node20820 = (inp[9]) ? node20822 : 4'b0110;
																assign node20822 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node20825 = (inp[0]) ? node20827 : 4'b0000;
															assign node20827 = (inp[10]) ? node20831 : node20828;
																assign node20828 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node20831 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node20834 = (inp[7]) ? node20842 : node20835;
														assign node20835 = (inp[0]) ? node20837 : 4'b0101;
															assign node20837 = (inp[9]) ? node20839 : 4'b0100;
																assign node20839 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node20842 = (inp[9]) ? 4'b0111 : node20843;
															assign node20843 = (inp[0]) ? node20847 : node20844;
																assign node20844 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node20847 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node20851 = (inp[5]) ? node20875 : node20852;
												assign node20852 = (inp[15]) ? node20862 : node20853;
													assign node20853 = (inp[7]) ? node20857 : node20854;
														assign node20854 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node20857 = (inp[9]) ? 4'b0110 : node20858;
															assign node20858 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node20862 = (inp[7]) ? node20870 : node20863;
														assign node20863 = (inp[10]) ? node20867 : node20864;
															assign node20864 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node20867 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node20870 = (inp[0]) ? 4'b0001 : node20871;
															assign node20871 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node20875 = (inp[10]) ? node20893 : node20876;
													assign node20876 = (inp[9]) ? node20888 : node20877;
														assign node20877 = (inp[7]) ? node20881 : node20878;
															assign node20878 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node20881 = (inp[15]) ? node20885 : node20882;
																assign node20882 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node20885 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20888 = (inp[15]) ? node20890 : 4'b0000;
															assign node20890 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node20893 = (inp[15]) ? node20905 : node20894;
														assign node20894 = (inp[7]) ? node20898 : node20895;
															assign node20895 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node20898 = (inp[0]) ? node20902 : node20899;
																assign node20899 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node20902 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node20905 = (inp[7]) ? node20911 : node20906;
															assign node20906 = (inp[0]) ? 4'b0011 : node20907;
																assign node20907 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node20911 = (inp[9]) ? node20913 : 4'b0001;
																assign node20913 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node20916 = (inp[7]) ? node21050 : node20917;
										assign node20917 = (inp[15]) ? node20969 : node20918;
											assign node20918 = (inp[12]) ? node20944 : node20919;
												assign node20919 = (inp[5]) ? node20929 : node20920;
													assign node20920 = (inp[1]) ? 4'b0011 : node20921;
														assign node20921 = (inp[10]) ? node20923 : 4'b0110;
															assign node20923 = (inp[9]) ? node20925 : 4'b0111;
																assign node20925 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node20929 = (inp[0]) ? 4'b0010 : node20930;
														assign node20930 = (inp[10]) ? node20936 : node20931;
															assign node20931 = (inp[9]) ? node20933 : 4'b0010;
																assign node20933 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node20936 = (inp[9]) ? node20940 : node20937;
																assign node20937 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node20940 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node20944 = (inp[5]) ? node20956 : node20945;
													assign node20945 = (inp[1]) ? node20953 : node20946;
														assign node20946 = (inp[0]) ? node20948 : 4'b0001;
															assign node20948 = (inp[9]) ? 4'b0000 : node20949;
																assign node20949 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node20953 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node20956 = (inp[10]) ? node20962 : node20957;
														assign node20957 = (inp[9]) ? node20959 : 4'b0100;
															assign node20959 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node20962 = (inp[9]) ? node20964 : 4'b0101;
															assign node20964 = (inp[0]) ? node20966 : 4'b0100;
																assign node20966 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node20969 = (inp[12]) ? node21003 : node20970;
												assign node20970 = (inp[5]) ? node20992 : node20971;
													assign node20971 = (inp[0]) ? node20985 : node20972;
														assign node20972 = (inp[10]) ? node20978 : node20973;
															assign node20973 = (inp[9]) ? node20975 : 4'b0100;
																assign node20975 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node20978 = (inp[9]) ? node20982 : node20979;
																assign node20979 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node20982 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node20985 = (inp[9]) ? node20987 : 4'b0100;
															assign node20987 = (inp[1]) ? node20989 : 4'b0100;
																assign node20989 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node20992 = (inp[1]) ? node20998 : node20993;
														assign node20993 = (inp[9]) ? node20995 : 4'b0101;
															assign node20995 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node20998 = (inp[0]) ? node21000 : 4'b0001;
															assign node21000 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21003 = (inp[5]) ? node21025 : node21004;
													assign node21004 = (inp[1]) ? node21012 : node21005;
														assign node21005 = (inp[9]) ? node21009 : node21006;
															assign node21006 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node21009 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node21012 = (inp[0]) ? node21018 : node21013;
															assign node21013 = (inp[10]) ? 4'b0110 : node21014;
																assign node21014 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node21018 = (inp[10]) ? node21022 : node21019;
																assign node21019 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node21022 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node21025 = (inp[0]) ? node21037 : node21026;
														assign node21026 = (inp[1]) ? node21032 : node21027;
															assign node21027 = (inp[9]) ? 4'b0111 : node21028;
																assign node21028 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node21032 = (inp[9]) ? node21034 : 4'b0111;
																assign node21034 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node21037 = (inp[1]) ? node21045 : node21038;
															assign node21038 = (inp[9]) ? node21042 : node21039;
																assign node21039 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node21042 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node21045 = (inp[10]) ? 4'b0110 : node21046;
																assign node21046 = (inp[9]) ? 4'b0111 : 4'b0110;
										assign node21050 = (inp[1]) ? node21116 : node21051;
											assign node21051 = (inp[5]) ? node21087 : node21052;
												assign node21052 = (inp[12]) ? node21072 : node21053;
													assign node21053 = (inp[15]) ? node21063 : node21054;
														assign node21054 = (inp[0]) ? 4'b0000 : node21055;
															assign node21055 = (inp[9]) ? node21059 : node21056;
																assign node21056 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node21059 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node21063 = (inp[0]) ? node21065 : 4'b0111;
															assign node21065 = (inp[9]) ? node21069 : node21066;
																assign node21066 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node21069 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21072 = (inp[15]) ? node21080 : node21073;
														assign node21073 = (inp[0]) ? node21075 : 4'b0010;
															assign node21075 = (inp[10]) ? 4'b0011 : node21076;
																assign node21076 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node21080 = (inp[10]) ? node21084 : node21081;
															assign node21081 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node21084 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node21087 = (inp[12]) ? node21101 : node21088;
													assign node21088 = (inp[15]) ? node21094 : node21089;
														assign node21089 = (inp[10]) ? 4'b0100 : node21090;
															assign node21090 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node21094 = (inp[9]) ? node21096 : 4'b0010;
															assign node21096 = (inp[10]) ? 4'b0011 : node21097;
																assign node21097 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node21101 = (inp[15]) ? node21109 : node21102;
														assign node21102 = (inp[10]) ? node21106 : node21103;
															assign node21103 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node21106 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node21109 = (inp[9]) ? node21113 : node21110;
															assign node21110 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node21113 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node21116 = (inp[15]) ? node21148 : node21117;
												assign node21117 = (inp[12]) ? node21137 : node21118;
													assign node21118 = (inp[0]) ? node21124 : node21119;
														assign node21119 = (inp[5]) ? 4'b0100 : node21120;
															assign node21120 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21124 = (inp[10]) ? node21130 : node21125;
															assign node21125 = (inp[5]) ? node21127 : 4'b0101;
																assign node21127 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node21130 = (inp[9]) ? node21134 : node21131;
																assign node21131 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node21134 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node21137 = (inp[5]) ? node21143 : node21138;
														assign node21138 = (inp[0]) ? node21140 : 4'b0011;
															assign node21140 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node21143 = (inp[10]) ? 4'b0110 : node21144;
															assign node21144 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node21148 = (inp[12]) ? node21160 : node21149;
													assign node21149 = (inp[9]) ? node21151 : 4'b0010;
														assign node21151 = (inp[0]) ? node21155 : node21152;
															assign node21152 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node21155 = (inp[10]) ? node21157 : 4'b0011;
																assign node21157 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node21160 = (inp[9]) ? node21168 : node21161;
														assign node21161 = (inp[0]) ? node21165 : node21162;
															assign node21162 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node21165 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21168 = (inp[0]) ? 4'b0100 : node21169;
															assign node21169 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node21173 = (inp[2]) ? node21435 : node21174;
									assign node21174 = (inp[7]) ? node21308 : node21175;
										assign node21175 = (inp[15]) ? node21239 : node21176;
											assign node21176 = (inp[12]) ? node21206 : node21177;
												assign node21177 = (inp[1]) ? node21193 : node21178;
													assign node21178 = (inp[5]) ? node21188 : node21179;
														assign node21179 = (inp[10]) ? node21181 : 4'b0110;
															assign node21181 = (inp[0]) ? node21185 : node21182;
																assign node21182 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node21185 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node21188 = (inp[10]) ? node21190 : 4'b0010;
															assign node21190 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node21193 = (inp[9]) ? node21203 : node21194;
														assign node21194 = (inp[5]) ? node21196 : 4'b0010;
															assign node21196 = (inp[0]) ? node21200 : node21197;
																assign node21197 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node21200 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node21203 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node21206 = (inp[5]) ? node21222 : node21207;
													assign node21207 = (inp[1]) ? node21215 : node21208;
														assign node21208 = (inp[9]) ? node21212 : node21209;
															assign node21209 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node21212 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node21215 = (inp[9]) ? node21219 : node21216;
															assign node21216 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node21219 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node21222 = (inp[9]) ? node21230 : node21223;
														assign node21223 = (inp[1]) ? node21225 : 4'b0100;
															assign node21225 = (inp[0]) ? node21227 : 4'b0100;
																assign node21227 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node21230 = (inp[10]) ? node21234 : node21231;
															assign node21231 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node21234 = (inp[0]) ? node21236 : 4'b0100;
																assign node21236 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node21239 = (inp[12]) ? node21271 : node21240;
												assign node21240 = (inp[1]) ? node21256 : node21241;
													assign node21241 = (inp[9]) ? node21247 : node21242;
														assign node21242 = (inp[10]) ? 4'b0100 : node21243;
															assign node21243 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node21247 = (inp[10]) ? node21251 : node21248;
															assign node21248 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node21251 = (inp[5]) ? 4'b0101 : node21252;
																assign node21252 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node21256 = (inp[5]) ? node21264 : node21257;
														assign node21257 = (inp[10]) ? 4'b0101 : node21258;
															assign node21258 = (inp[9]) ? node21260 : 4'b0101;
																assign node21260 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node21264 = (inp[9]) ? node21268 : node21265;
															assign node21265 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node21268 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21271 = (inp[1]) ? node21287 : node21272;
													assign node21272 = (inp[5]) ? node21280 : node21273;
														assign node21273 = (inp[10]) ? node21277 : node21274;
															assign node21274 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node21277 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node21280 = (inp[10]) ? node21284 : node21281;
															assign node21281 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node21284 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node21287 = (inp[9]) ? node21299 : node21288;
														assign node21288 = (inp[10]) ? node21294 : node21289;
															assign node21289 = (inp[5]) ? 4'b0111 : node21290;
																assign node21290 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node21294 = (inp[5]) ? 4'b0110 : node21295;
																assign node21295 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node21299 = (inp[5]) ? 4'b0110 : node21300;
															assign node21300 = (inp[10]) ? node21304 : node21301;
																assign node21301 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node21304 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node21308 = (inp[1]) ? node21372 : node21309;
											assign node21309 = (inp[12]) ? node21345 : node21310;
												assign node21310 = (inp[15]) ? node21324 : node21311;
													assign node21311 = (inp[5]) ? node21319 : node21312;
														assign node21312 = (inp[9]) ? node21316 : node21313;
															assign node21313 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node21316 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node21319 = (inp[9]) ? 4'b0101 : node21320;
															assign node21320 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node21324 = (inp[5]) ? node21332 : node21325;
														assign node21325 = (inp[10]) ? node21329 : node21326;
															assign node21326 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node21329 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node21332 = (inp[9]) ? node21340 : node21333;
															assign node21333 = (inp[0]) ? node21337 : node21334;
																assign node21334 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node21337 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node21340 = (inp[10]) ? node21342 : 4'b0011;
																assign node21342 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node21345 = (inp[15]) ? node21361 : node21346;
													assign node21346 = (inp[9]) ? node21356 : node21347;
														assign node21347 = (inp[0]) ? 4'b0011 : node21348;
															assign node21348 = (inp[10]) ? node21352 : node21349;
																assign node21349 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node21352 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node21356 = (inp[0]) ? node21358 : 4'b0011;
															assign node21358 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node21361 = (inp[5]) ? node21369 : node21362;
														assign node21362 = (inp[9]) ? node21366 : node21363;
															assign node21363 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node21366 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node21369 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node21372 = (inp[12]) ? node21412 : node21373;
												assign node21373 = (inp[15]) ? node21393 : node21374;
													assign node21374 = (inp[5]) ? node21386 : node21375;
														assign node21375 = (inp[0]) ? node21381 : node21376;
															assign node21376 = (inp[10]) ? node21378 : 4'b0100;
																assign node21378 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node21381 = (inp[10]) ? 4'b0100 : node21382;
																assign node21382 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node21386 = (inp[9]) ? node21390 : node21387;
															assign node21387 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node21390 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node21393 = (inp[0]) ? node21407 : node21394;
														assign node21394 = (inp[5]) ? node21402 : node21395;
															assign node21395 = (inp[10]) ? node21399 : node21396;
																assign node21396 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node21399 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node21402 = (inp[10]) ? 4'b0010 : node21403;
																assign node21403 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node21407 = (inp[10]) ? node21409 : 4'b0011;
															assign node21409 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node21412 = (inp[15]) ? node21424 : node21413;
													assign node21413 = (inp[5]) ? node21419 : node21414;
														assign node21414 = (inp[0]) ? 4'b0011 : node21415;
															assign node21415 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node21419 = (inp[9]) ? 4'b0111 : node21420;
															assign node21420 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21424 = (inp[10]) ? node21432 : node21425;
														assign node21425 = (inp[9]) ? 4'b0100 : node21426;
															assign node21426 = (inp[0]) ? 4'b0101 : node21427;
																assign node21427 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node21432 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node21435 = (inp[12]) ? node21583 : node21436;
										assign node21436 = (inp[1]) ? node21516 : node21437;
											assign node21437 = (inp[7]) ? node21479 : node21438;
												assign node21438 = (inp[15]) ? node21462 : node21439;
													assign node21439 = (inp[5]) ? node21455 : node21440;
														assign node21440 = (inp[10]) ? node21448 : node21441;
															assign node21441 = (inp[9]) ? node21445 : node21442;
																assign node21442 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node21445 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node21448 = (inp[9]) ? node21452 : node21449;
																assign node21449 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node21452 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node21455 = (inp[10]) ? node21457 : 4'b0111;
															assign node21457 = (inp[0]) ? 4'b0110 : node21458;
																assign node21458 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node21462 = (inp[5]) ? node21472 : node21463;
														assign node21463 = (inp[0]) ? 4'b0001 : node21464;
															assign node21464 = (inp[9]) ? node21468 : node21465;
																assign node21465 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node21468 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node21472 = (inp[10]) ? node21476 : node21473;
															assign node21473 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node21476 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node21479 = (inp[15]) ? node21497 : node21480;
													assign node21480 = (inp[5]) ? node21490 : node21481;
														assign node21481 = (inp[9]) ? 4'b0101 : node21482;
															assign node21482 = (inp[0]) ? node21486 : node21483;
																assign node21483 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node21486 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21490 = (inp[9]) ? node21494 : node21491;
															assign node21491 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node21494 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node21497 = (inp[5]) ? node21507 : node21498;
														assign node21498 = (inp[0]) ? node21502 : node21499;
															assign node21499 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node21502 = (inp[9]) ? 4'b0010 : node21503;
																assign node21503 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node21507 = (inp[0]) ? 4'b0111 : node21508;
															assign node21508 = (inp[10]) ? node21512 : node21509;
																assign node21509 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node21512 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node21516 = (inp[15]) ? node21548 : node21517;
												assign node21517 = (inp[7]) ? node21535 : node21518;
													assign node21518 = (inp[9]) ? node21528 : node21519;
														assign node21519 = (inp[10]) ? node21523 : node21520;
															assign node21520 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node21523 = (inp[5]) ? 4'b0110 : node21524;
																assign node21524 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node21528 = (inp[10]) ? node21532 : node21529;
															assign node21529 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node21532 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node21535 = (inp[0]) ? node21543 : node21536;
														assign node21536 = (inp[10]) ? node21540 : node21537;
															assign node21537 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node21540 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node21543 = (inp[10]) ? node21545 : 4'b0000;
															assign node21545 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node21548 = (inp[7]) ? node21566 : node21549;
													assign node21549 = (inp[5]) ? node21557 : node21550;
														assign node21550 = (inp[10]) ? node21552 : 4'b0001;
															assign node21552 = (inp[0]) ? 4'b0000 : node21553;
																assign node21553 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node21557 = (inp[0]) ? 4'b0101 : node21558;
															assign node21558 = (inp[10]) ? node21562 : node21559;
																assign node21559 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node21562 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node21566 = (inp[10]) ? node21576 : node21567;
														assign node21567 = (inp[9]) ? node21571 : node21568;
															assign node21568 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node21571 = (inp[5]) ? 4'b0111 : node21572;
																assign node21572 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node21576 = (inp[9]) ? node21578 : 4'b0111;
															assign node21578 = (inp[0]) ? 4'b0110 : node21579;
																assign node21579 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node21583 = (inp[1]) ? node21639 : node21584;
											assign node21584 = (inp[5]) ? node21616 : node21585;
												assign node21585 = (inp[7]) ? node21601 : node21586;
													assign node21586 = (inp[15]) ? node21594 : node21587;
														assign node21587 = (inp[0]) ? node21589 : 4'b0101;
															assign node21589 = (inp[10]) ? node21591 : 4'b0100;
																assign node21591 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node21594 = (inp[0]) ? node21596 : 4'b0110;
															assign node21596 = (inp[9]) ? 4'b0110 : node21597;
																assign node21597 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21601 = (inp[15]) ? node21611 : node21602;
														assign node21602 = (inp[0]) ? node21604 : 4'b0111;
															assign node21604 = (inp[10]) ? node21608 : node21605;
																assign node21605 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node21608 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node21611 = (inp[10]) ? 4'b0101 : node21612;
															assign node21612 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node21616 = (inp[15]) ? node21626 : node21617;
													assign node21617 = (inp[7]) ? node21619 : 4'b0001;
														assign node21619 = (inp[0]) ? node21621 : 4'b0111;
															assign node21621 = (inp[10]) ? 4'b0110 : node21622;
																assign node21622 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node21626 = (inp[7]) ? node21634 : node21627;
														assign node21627 = (inp[10]) ? node21631 : node21628;
															assign node21628 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node21631 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node21634 = (inp[9]) ? 4'b0000 : node21635;
															assign node21635 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node21639 = (inp[15]) ? node21679 : node21640;
												assign node21640 = (inp[7]) ? node21658 : node21641;
													assign node21641 = (inp[9]) ? node21651 : node21642;
														assign node21642 = (inp[10]) ? node21646 : node21643;
															assign node21643 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node21646 = (inp[5]) ? node21648 : 4'b0001;
																assign node21648 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node21651 = (inp[10]) ? 4'b0000 : node21652;
															assign node21652 = (inp[0]) ? 4'b0001 : node21653;
																assign node21653 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node21658 = (inp[5]) ? node21672 : node21659;
														assign node21659 = (inp[9]) ? node21667 : node21660;
															assign node21660 = (inp[10]) ? node21664 : node21661;
																assign node21661 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node21664 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node21667 = (inp[0]) ? 4'b0110 : node21668;
																assign node21668 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node21672 = (inp[10]) ? node21676 : node21673;
															assign node21673 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node21676 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node21679 = (inp[7]) ? node21703 : node21680;
													assign node21680 = (inp[0]) ? node21694 : node21681;
														assign node21681 = (inp[5]) ? node21687 : node21682;
															assign node21682 = (inp[9]) ? node21684 : 4'b0010;
																assign node21684 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node21687 = (inp[9]) ? node21691 : node21688;
																assign node21688 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node21691 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node21694 = (inp[10]) ? node21696 : 4'b0010;
															assign node21696 = (inp[9]) ? node21700 : node21697;
																assign node21697 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node21700 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node21703 = (inp[0]) ? node21713 : node21704;
														assign node21704 = (inp[10]) ? 4'b0000 : node21705;
															assign node21705 = (inp[9]) ? node21709 : node21706;
																assign node21706 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node21709 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node21713 = (inp[5]) ? node21721 : node21714;
															assign node21714 = (inp[10]) ? node21718 : node21715;
																assign node21715 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node21718 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node21721 = (inp[9]) ? node21725 : node21722;
																assign node21722 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node21725 = (inp[10]) ? 4'b0000 : 4'b0001;
						assign node21728 = (inp[1]) ? node22834 : node21729;
							assign node21729 = (inp[9]) ? node22263 : node21730;
								assign node21730 = (inp[5]) ? node22020 : node21731;
									assign node21731 = (inp[10]) ? node21873 : node21732;
										assign node21732 = (inp[2]) ? node21798 : node21733;
											assign node21733 = (inp[13]) ? node21763 : node21734;
												assign node21734 = (inp[11]) ? node21748 : node21735;
													assign node21735 = (inp[12]) ? node21743 : node21736;
														assign node21736 = (inp[7]) ? node21738 : 4'b0100;
															assign node21738 = (inp[0]) ? node21740 : 4'b0110;
																assign node21740 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node21743 = (inp[0]) ? node21745 : 4'b0010;
															assign node21745 = (inp[7]) ? 4'b0100 : 4'b0110;
													assign node21748 = (inp[12]) ? node21754 : node21749;
														assign node21749 = (inp[7]) ? 4'b0111 : node21750;
															assign node21750 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node21754 = (inp[7]) ? 4'b0100 : node21755;
															assign node21755 = (inp[15]) ? node21759 : node21756;
																assign node21756 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node21759 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node21763 = (inp[7]) ? node21775 : node21764;
													assign node21764 = (inp[15]) ? node21770 : node21765;
														assign node21765 = (inp[0]) ? 4'b0110 : node21766;
															assign node21766 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node21770 = (inp[12]) ? node21772 : 4'b0001;
															assign node21772 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node21775 = (inp[12]) ? node21787 : node21776;
														assign node21776 = (inp[0]) ? node21782 : node21777;
															assign node21777 = (inp[15]) ? 4'b0010 : node21778;
																assign node21778 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node21782 = (inp[15]) ? node21784 : 4'b0010;
																assign node21784 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node21787 = (inp[15]) ? node21793 : node21788;
															assign node21788 = (inp[0]) ? 4'b0001 : node21789;
																assign node21789 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21793 = (inp[0]) ? node21795 : 4'b0001;
																assign node21795 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node21798 = (inp[13]) ? node21830 : node21799;
												assign node21799 = (inp[7]) ? node21819 : node21800;
													assign node21800 = (inp[15]) ? node21808 : node21801;
														assign node21801 = (inp[12]) ? 4'b0111 : node21802;
															assign node21802 = (inp[0]) ? node21804 : 4'b0101;
																assign node21804 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node21808 = (inp[12]) ? node21814 : node21809;
															assign node21809 = (inp[11]) ? 4'b0001 : node21810;
																assign node21810 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node21814 = (inp[11]) ? node21816 : 4'b0010;
																assign node21816 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node21819 = (inp[12]) ? node21827 : node21820;
														assign node21820 = (inp[15]) ? 4'b0010 : node21821;
															assign node21821 = (inp[11]) ? 4'b0011 : node21822;
																assign node21822 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node21827 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node21830 = (inp[15]) ? node21848 : node21831;
													assign node21831 = (inp[7]) ? node21841 : node21832;
														assign node21832 = (inp[12]) ? node21836 : node21833;
															assign node21833 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node21836 = (inp[0]) ? 4'b0010 : node21837;
																assign node21837 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21841 = (inp[12]) ? 4'b0101 : node21842;
															assign node21842 = (inp[0]) ? node21844 : 4'b0110;
																assign node21844 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node21848 = (inp[0]) ? node21862 : node21849;
														assign node21849 = (inp[11]) ? node21857 : node21850;
															assign node21850 = (inp[12]) ? node21854 : node21851;
																assign node21851 = (inp[7]) ? 4'b0110 : 4'b0101;
																assign node21854 = (inp[7]) ? 4'b0101 : 4'b0110;
															assign node21857 = (inp[7]) ? 4'b0111 : node21858;
																assign node21858 = (inp[12]) ? 4'b0111 : 4'b0101;
														assign node21862 = (inp[11]) ? node21868 : node21863;
															assign node21863 = (inp[7]) ? node21865 : 4'b0111;
																assign node21865 = (inp[12]) ? 4'b0100 : 4'b0111;
															assign node21868 = (inp[12]) ? 4'b0100 : node21869;
																assign node21869 = (inp[7]) ? 4'b0111 : 4'b0100;
										assign node21873 = (inp[15]) ? node21939 : node21874;
											assign node21874 = (inp[13]) ? node21910 : node21875;
												assign node21875 = (inp[12]) ? node21897 : node21876;
													assign node21876 = (inp[7]) ? node21888 : node21877;
														assign node21877 = (inp[2]) ? node21883 : node21878;
															assign node21878 = (inp[0]) ? 4'b0000 : node21879;
																assign node21879 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node21883 = (inp[0]) ? node21885 : 4'b0100;
																assign node21885 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node21888 = (inp[2]) ? node21894 : node21889;
															assign node21889 = (inp[0]) ? 4'b0110 : node21890;
																assign node21890 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node21894 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node21897 = (inp[7]) ? node21903 : node21898;
														assign node21898 = (inp[2]) ? node21900 : 4'b0011;
															assign node21900 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node21903 = (inp[2]) ? 4'b0001 : node21904;
															assign node21904 = (inp[11]) ? 4'b0101 : node21905;
																assign node21905 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node21910 = (inp[12]) ? node21926 : node21911;
													assign node21911 = (inp[7]) ? node21915 : node21912;
														assign node21912 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node21915 = (inp[2]) ? node21921 : node21916;
															assign node21916 = (inp[11]) ? 4'b0011 : node21917;
																assign node21917 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node21921 = (inp[0]) ? node21923 : 4'b0111;
																assign node21923 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node21926 = (inp[7]) ? node21936 : node21927;
														assign node21927 = (inp[2]) ? node21931 : node21928;
															assign node21928 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node21931 = (inp[0]) ? 4'b0011 : node21932;
																assign node21932 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node21936 = (inp[0]) ? 4'b0000 : 4'b0100;
											assign node21939 = (inp[0]) ? node21977 : node21940;
												assign node21940 = (inp[11]) ? node21962 : node21941;
													assign node21941 = (inp[13]) ? node21953 : node21942;
														assign node21942 = (inp[2]) ? node21948 : node21943;
															assign node21943 = (inp[7]) ? 4'b0100 : node21944;
																assign node21944 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node21948 = (inp[12]) ? 4'b0000 : node21949;
																assign node21949 = (inp[7]) ? 4'b0011 : 4'b0001;
														assign node21953 = (inp[2]) ? node21955 : 4'b0011;
															assign node21955 = (inp[12]) ? node21959 : node21956;
																assign node21956 = (inp[7]) ? 4'b0111 : 4'b0100;
																assign node21959 = (inp[7]) ? 4'b0100 : 4'b0111;
													assign node21962 = (inp[7]) ? node21968 : node21963;
														assign node21963 = (inp[12]) ? node21965 : 4'b0100;
															assign node21965 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node21968 = (inp[12]) ? node21974 : node21969;
															assign node21969 = (inp[2]) ? node21971 : 4'b0011;
																assign node21971 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node21974 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node21977 = (inp[7]) ? node21997 : node21978;
													assign node21978 = (inp[12]) ? node21988 : node21979;
														assign node21979 = (inp[2]) ? node21983 : node21980;
															assign node21980 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node21983 = (inp[13]) ? node21985 : 4'b0000;
																assign node21985 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node21988 = (inp[11]) ? node21994 : node21989;
															assign node21989 = (inp[2]) ? 4'b0110 : node21990;
																assign node21990 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node21994 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node21997 = (inp[12]) ? node22007 : node21998;
														assign node21998 = (inp[11]) ? node22004 : node21999;
															assign node21999 = (inp[13]) ? 4'b0110 : node22000;
																assign node22000 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node22004 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node22007 = (inp[11]) ? node22013 : node22008;
															assign node22008 = (inp[13]) ? 4'b0101 : node22009;
																assign node22009 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node22013 = (inp[13]) ? node22017 : node22014;
																assign node22014 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node22017 = (inp[2]) ? 4'b0101 : 4'b0001;
									assign node22020 = (inp[15]) ? node22142 : node22021;
										assign node22021 = (inp[2]) ? node22083 : node22022;
											assign node22022 = (inp[13]) ? node22052 : node22023;
												assign node22023 = (inp[7]) ? node22037 : node22024;
													assign node22024 = (inp[12]) ? node22030 : node22025;
														assign node22025 = (inp[10]) ? 4'b0001 : node22026;
															assign node22026 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node22030 = (inp[10]) ? 4'b0111 : node22031;
															assign node22031 = (inp[11]) ? 4'b0110 : node22032;
																assign node22032 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node22037 = (inp[12]) ? node22043 : node22038;
														assign node22038 = (inp[10]) ? 4'b0010 : node22039;
															assign node22039 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22043 = (inp[10]) ? node22047 : node22044;
															assign node22044 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22047 = (inp[11]) ? 4'b0001 : node22048;
																assign node22048 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node22052 = (inp[7]) ? node22068 : node22053;
													assign node22053 = (inp[12]) ? node22059 : node22054;
														assign node22054 = (inp[10]) ? node22056 : 4'b0101;
															assign node22056 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22059 = (inp[0]) ? 4'b0011 : node22060;
															assign node22060 = (inp[11]) ? node22064 : node22061;
																assign node22061 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node22064 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node22068 = (inp[12]) ? node22074 : node22069;
														assign node22069 = (inp[10]) ? node22071 : 4'b0110;
															assign node22071 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node22074 = (inp[10]) ? node22080 : node22075;
															assign node22075 = (inp[0]) ? node22077 : 4'b0101;
																assign node22077 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node22080 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node22083 = (inp[13]) ? node22111 : node22084;
												assign node22084 = (inp[7]) ? node22098 : node22085;
													assign node22085 = (inp[12]) ? node22089 : node22086;
														assign node22086 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node22089 = (inp[10]) ? node22093 : node22090;
															assign node22090 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node22093 = (inp[11]) ? 4'b0011 : node22094;
																assign node22094 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node22098 = (inp[12]) ? node22104 : node22099;
														assign node22099 = (inp[10]) ? node22101 : 4'b0111;
															assign node22101 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22104 = (inp[10]) ? node22108 : node22105;
															assign node22105 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node22108 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node22111 = (inp[12]) ? node22125 : node22112;
													assign node22112 = (inp[7]) ? node22116 : node22113;
														assign node22113 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node22116 = (inp[10]) ? node22122 : node22117;
															assign node22117 = (inp[0]) ? node22119 : 4'b0010;
																assign node22119 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22122 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node22125 = (inp[7]) ? node22137 : node22126;
														assign node22126 = (inp[10]) ? node22132 : node22127;
															assign node22127 = (inp[0]) ? node22129 : 4'b0111;
																assign node22129 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node22132 = (inp[11]) ? node22134 : 4'b0110;
																assign node22134 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22137 = (inp[11]) ? 4'b0001 : node22138;
															assign node22138 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node22142 = (inp[7]) ? node22206 : node22143;
											assign node22143 = (inp[12]) ? node22173 : node22144;
												assign node22144 = (inp[10]) ? node22160 : node22145;
													assign node22145 = (inp[0]) ? node22155 : node22146;
														assign node22146 = (inp[11]) ? 4'b0100 : node22147;
															assign node22147 = (inp[2]) ? node22151 : node22148;
																assign node22148 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node22151 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node22155 = (inp[13]) ? 4'b0000 : node22156;
															assign node22156 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node22160 = (inp[11]) ? node22166 : node22161;
														assign node22161 = (inp[13]) ? 4'b0101 : node22162;
															assign node22162 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node22166 = (inp[0]) ? 4'b0001 : node22167;
															assign node22167 = (inp[13]) ? 4'b0101 : node22168;
																assign node22168 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node22173 = (inp[13]) ? node22191 : node22174;
													assign node22174 = (inp[2]) ? node22182 : node22175;
														assign node22175 = (inp[10]) ? 4'b0010 : node22176;
															assign node22176 = (inp[11]) ? node22178 : 4'b0011;
																assign node22178 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node22182 = (inp[11]) ? 4'b0110 : node22183;
															assign node22183 = (inp[10]) ? node22187 : node22184;
																assign node22184 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node22187 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node22191 = (inp[2]) ? node22199 : node22192;
														assign node22192 = (inp[0]) ? 4'b0111 : node22193;
															assign node22193 = (inp[11]) ? 4'b0111 : node22194;
																assign node22194 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node22199 = (inp[10]) ? node22201 : 4'b0010;
															assign node22201 = (inp[11]) ? 4'b0011 : node22202;
																assign node22202 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node22206 = (inp[12]) ? node22244 : node22207;
												assign node22207 = (inp[11]) ? node22227 : node22208;
													assign node22208 = (inp[10]) ? node22218 : node22209;
														assign node22209 = (inp[0]) ? node22213 : node22210;
															assign node22210 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node22213 = (inp[13]) ? node22215 : 4'b0010;
																assign node22215 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node22218 = (inp[0]) ? node22224 : node22219;
															assign node22219 = (inp[2]) ? 4'b0011 : node22220;
																assign node22220 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node22224 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node22227 = (inp[10]) ? node22235 : node22228;
														assign node22228 = (inp[2]) ? node22232 : node22229;
															assign node22229 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node22232 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node22235 = (inp[13]) ? node22241 : node22236;
															assign node22236 = (inp[2]) ? 4'b0110 : node22237;
																assign node22237 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node22241 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node22244 = (inp[13]) ? node22256 : node22245;
													assign node22245 = (inp[2]) ? 4'b0101 : node22246;
														assign node22246 = (inp[10]) ? node22252 : node22247;
															assign node22247 = (inp[0]) ? node22249 : 4'b0001;
																assign node22249 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22252 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node22256 = (inp[2]) ? node22258 : 4'b0101;
														assign node22258 = (inp[0]) ? node22260 : 4'b0000;
															assign node22260 = (inp[10]) ? 4'b0001 : 4'b0000;
								assign node22263 = (inp[15]) ? node22529 : node22264;
									assign node22264 = (inp[5]) ? node22408 : node22265;
										assign node22265 = (inp[11]) ? node22335 : node22266;
											assign node22266 = (inp[0]) ? node22298 : node22267;
												assign node22267 = (inp[7]) ? node22287 : node22268;
													assign node22268 = (inp[12]) ? node22274 : node22269;
														assign node22269 = (inp[2]) ? 4'b0100 : node22270;
															assign node22270 = (inp[10]) ? 4'b0100 : 4'b0001;
														assign node22274 = (inp[2]) ? node22282 : node22275;
															assign node22275 = (inp[13]) ? node22279 : node22276;
																assign node22276 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node22279 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node22282 = (inp[13]) ? 4'b0010 : node22283;
																assign node22283 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node22287 = (inp[12]) ? node22295 : node22288;
														assign node22288 = (inp[2]) ? node22292 : node22289;
															assign node22289 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node22292 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node22295 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node22298 = (inp[13]) ? node22314 : node22299;
													assign node22299 = (inp[10]) ? node22307 : node22300;
														assign node22300 = (inp[12]) ? 4'b0011 : node22301;
															assign node22301 = (inp[7]) ? 4'b0110 : node22302;
																assign node22302 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node22307 = (inp[7]) ? node22311 : node22308;
															assign node22308 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node22311 = (inp[12]) ? 4'b0000 : 4'b0011;
													assign node22314 = (inp[10]) ? node22322 : node22315;
														assign node22315 = (inp[12]) ? node22317 : 4'b0011;
															assign node22317 = (inp[7]) ? node22319 : 4'b0111;
																assign node22319 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node22322 = (inp[7]) ? node22330 : node22323;
															assign node22323 = (inp[12]) ? node22327 : node22324;
																assign node22324 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node22327 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node22330 = (inp[12]) ? 4'b0101 : node22331;
																assign node22331 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node22335 = (inp[12]) ? node22371 : node22336;
												assign node22336 = (inp[7]) ? node22358 : node22337;
													assign node22337 = (inp[10]) ? node22347 : node22338;
														assign node22338 = (inp[2]) ? node22342 : node22339;
															assign node22339 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node22342 = (inp[13]) ? 4'b0001 : node22343;
																assign node22343 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22347 = (inp[13]) ? node22351 : node22348;
															assign node22348 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node22351 = (inp[0]) ? node22355 : node22352;
																assign node22352 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node22355 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node22358 = (inp[10]) ? node22362 : node22359;
														assign node22359 = (inp[0]) ? 4'b0110 : 4'b0010;
														assign node22362 = (inp[13]) ? node22366 : node22363;
															assign node22363 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node22366 = (inp[0]) ? 4'b0111 : node22367;
																assign node22367 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node22371 = (inp[7]) ? node22387 : node22372;
													assign node22372 = (inp[10]) ? node22380 : node22373;
														assign node22373 = (inp[13]) ? node22377 : node22374;
															assign node22374 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node22377 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node22380 = (inp[13]) ? node22384 : node22381;
															assign node22381 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node22384 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node22387 = (inp[0]) ? node22397 : node22388;
														assign node22388 = (inp[13]) ? node22392 : node22389;
															assign node22389 = (inp[10]) ? 4'b0000 : 4'b0101;
															assign node22392 = (inp[10]) ? 4'b0101 : node22393;
																assign node22393 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node22397 = (inp[2]) ? node22403 : node22398;
															assign node22398 = (inp[13]) ? node22400 : 4'b0100;
																assign node22400 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node22403 = (inp[13]) ? 4'b0101 : node22404;
																assign node22404 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node22408 = (inp[13]) ? node22470 : node22409;
											assign node22409 = (inp[2]) ? node22439 : node22410;
												assign node22410 = (inp[7]) ? node22424 : node22411;
													assign node22411 = (inp[12]) ? node22421 : node22412;
														assign node22412 = (inp[10]) ? node22418 : node22413;
															assign node22413 = (inp[11]) ? 4'b0001 : node22414;
																assign node22414 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node22418 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node22421 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node22424 = (inp[12]) ? node22432 : node22425;
														assign node22425 = (inp[10]) ? node22427 : 4'b0010;
															assign node22427 = (inp[0]) ? 4'b0011 : node22428;
																assign node22428 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22432 = (inp[10]) ? 4'b0000 : node22433;
															assign node22433 = (inp[0]) ? 4'b0001 : node22434;
																assign node22434 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node22439 = (inp[12]) ? node22455 : node22440;
													assign node22440 = (inp[7]) ? node22446 : node22441;
														assign node22441 = (inp[10]) ? 4'b0100 : node22442;
															assign node22442 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node22446 = (inp[10]) ? node22452 : node22447;
															assign node22447 = (inp[0]) ? node22449 : 4'b0110;
																assign node22449 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node22452 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node22455 = (inp[7]) ? node22463 : node22456;
														assign node22456 = (inp[10]) ? 4'b0010 : node22457;
															assign node22457 = (inp[0]) ? 4'b0011 : node22458;
																assign node22458 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22463 = (inp[0]) ? node22465 : 4'b0100;
															assign node22465 = (inp[11]) ? node22467 : 4'b0101;
																assign node22467 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node22470 = (inp[2]) ? node22498 : node22471;
												assign node22471 = (inp[10]) ? node22485 : node22472;
													assign node22472 = (inp[12]) ? node22478 : node22473;
														assign node22473 = (inp[7]) ? 4'b0111 : node22474;
															assign node22474 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node22478 = (inp[7]) ? node22482 : node22479;
															assign node22479 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node22482 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node22485 = (inp[7]) ? node22489 : node22486;
														assign node22486 = (inp[12]) ? 4'b0011 : 4'b0101;
														assign node22489 = (inp[12]) ? node22493 : node22490;
															assign node22490 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node22493 = (inp[11]) ? node22495 : 4'b0101;
																assign node22495 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node22498 = (inp[12]) ? node22512 : node22499;
													assign node22499 = (inp[7]) ? 4'b0011 : node22500;
														assign node22500 = (inp[10]) ? node22506 : node22501;
															assign node22501 = (inp[0]) ? node22503 : 4'b0000;
																assign node22503 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node22506 = (inp[11]) ? node22508 : 4'b0001;
																assign node22508 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node22512 = (inp[7]) ? node22522 : node22513;
														assign node22513 = (inp[11]) ? node22515 : 4'b0110;
															assign node22515 = (inp[10]) ? node22519 : node22516;
																assign node22516 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node22519 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node22522 = (inp[10]) ? 4'b0001 : node22523;
															assign node22523 = (inp[0]) ? node22525 : 4'b0000;
																assign node22525 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node22529 = (inp[11]) ? node22665 : node22530;
										assign node22530 = (inp[13]) ? node22598 : node22531;
											assign node22531 = (inp[10]) ? node22565 : node22532;
												assign node22532 = (inp[7]) ? node22552 : node22533;
													assign node22533 = (inp[12]) ? node22543 : node22534;
														assign node22534 = (inp[2]) ? node22538 : node22535;
															assign node22535 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node22538 = (inp[0]) ? 4'b0000 : node22539;
																assign node22539 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node22543 = (inp[5]) ? node22547 : node22544;
															assign node22544 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node22547 = (inp[2]) ? node22549 : 4'b0010;
																assign node22549 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node22552 = (inp[12]) ? node22562 : node22553;
														assign node22553 = (inp[2]) ? node22557 : node22554;
															assign node22554 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node22557 = (inp[5]) ? node22559 : 4'b0011;
																assign node22559 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node22562 = (inp[2]) ? 4'b0101 : 4'b0000;
												assign node22565 = (inp[12]) ? node22583 : node22566;
													assign node22566 = (inp[7]) ? node22578 : node22567;
														assign node22567 = (inp[2]) ? node22573 : node22568;
															assign node22568 = (inp[5]) ? node22570 : 4'b0101;
																assign node22570 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node22573 = (inp[0]) ? node22575 : 4'b0000;
																assign node22575 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node22578 = (inp[0]) ? node22580 : 4'b0010;
															assign node22580 = (inp[5]) ? 4'b0111 : 4'b0010;
													assign node22583 = (inp[7]) ? node22589 : node22584;
														assign node22584 = (inp[5]) ? node22586 : 4'b0110;
															assign node22586 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node22589 = (inp[2]) ? node22593 : node22590;
															assign node22590 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node22593 = (inp[5]) ? node22595 : 4'b0001;
																assign node22595 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node22598 = (inp[2]) ? node22628 : node22599;
												assign node22599 = (inp[5]) ? node22603 : node22600;
													assign node22600 = (inp[10]) ? 4'b0010 : 4'b0000;
													assign node22603 = (inp[12]) ? node22613 : node22604;
														assign node22604 = (inp[7]) ? node22606 : 4'b0001;
															assign node22606 = (inp[0]) ? node22610 : node22607;
																assign node22607 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node22610 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node22613 = (inp[7]) ? node22621 : node22614;
															assign node22614 = (inp[0]) ? node22618 : node22615;
																assign node22615 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node22618 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node22621 = (inp[0]) ? node22625 : node22622;
																assign node22622 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node22625 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node22628 = (inp[5]) ? node22644 : node22629;
													assign node22629 = (inp[10]) ? node22637 : node22630;
														assign node22630 = (inp[7]) ? node22632 : 4'b0100;
															assign node22632 = (inp[12]) ? node22634 : 4'b0111;
																assign node22634 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22637 = (inp[0]) ? node22639 : 4'b0101;
															assign node22639 = (inp[12]) ? 4'b0111 : node22640;
																assign node22640 = (inp[7]) ? 4'b0111 : 4'b0101;
													assign node22644 = (inp[10]) ? node22658 : node22645;
														assign node22645 = (inp[7]) ? node22651 : node22646;
															assign node22646 = (inp[12]) ? node22648 : 4'b0101;
																assign node22648 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node22651 = (inp[12]) ? node22655 : node22652;
																assign node22652 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node22655 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node22658 = (inp[7]) ? node22662 : node22659;
															assign node22659 = (inp[0]) ? 4'b0010 : 4'b0100;
															assign node22662 = (inp[12]) ? 4'b0000 : 4'b0010;
										assign node22665 = (inp[0]) ? node22749 : node22666;
											assign node22666 = (inp[10]) ? node22708 : node22667;
												assign node22667 = (inp[7]) ? node22685 : node22668;
													assign node22668 = (inp[12]) ? node22676 : node22669;
														assign node22669 = (inp[5]) ? node22671 : 4'b0000;
															assign node22671 = (inp[2]) ? node22673 : 4'b0001;
																assign node22673 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node22676 = (inp[13]) ? node22680 : node22677;
															assign node22677 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node22680 = (inp[5]) ? node22682 : 4'b0011;
																assign node22682 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node22685 = (inp[12]) ? node22697 : node22686;
														assign node22686 = (inp[13]) ? node22694 : node22687;
															assign node22687 = (inp[2]) ? node22691 : node22688;
																assign node22688 = (inp[5]) ? 4'b0011 : 4'b0111;
																assign node22691 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node22694 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node22697 = (inp[13]) ? node22703 : node22698;
															assign node22698 = (inp[5]) ? node22700 : 4'b0000;
																assign node22700 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node22703 = (inp[2]) ? node22705 : 4'b0101;
																assign node22705 = (inp[5]) ? 4'b0001 : 4'b0101;
												assign node22708 = (inp[2]) ? node22728 : node22709;
													assign node22709 = (inp[13]) ? node22723 : node22710;
														assign node22710 = (inp[5]) ? node22716 : node22711;
															assign node22711 = (inp[7]) ? 4'b0110 : node22712;
																assign node22712 = (inp[12]) ? 4'b0110 : 4'b0101;
															assign node22716 = (inp[12]) ? node22720 : node22717;
																assign node22717 = (inp[7]) ? 4'b0010 : 4'b0100;
																assign node22720 = (inp[7]) ? 4'b0001 : 4'b0011;
														assign node22723 = (inp[12]) ? node22725 : 4'b0111;
															assign node22725 = (inp[7]) ? 4'b0100 : 4'b0110;
													assign node22728 = (inp[5]) ? node22738 : node22729;
														assign node22729 = (inp[13]) ? 4'b0111 : node22730;
															assign node22730 = (inp[12]) ? node22734 : node22731;
																assign node22731 = (inp[7]) ? 4'b0010 : 4'b0001;
																assign node22734 = (inp[7]) ? 4'b0001 : 4'b0010;
														assign node22738 = (inp[7]) ? node22746 : node22739;
															assign node22739 = (inp[12]) ? node22743 : node22740;
																assign node22740 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node22743 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node22746 = (inp[12]) ? 4'b0000 : 4'b0011;
											assign node22749 = (inp[10]) ? node22785 : node22750;
												assign node22750 = (inp[5]) ? node22766 : node22751;
													assign node22751 = (inp[2]) ? node22763 : node22752;
														assign node22752 = (inp[13]) ? node22758 : node22753;
															assign node22753 = (inp[12]) ? 4'b0101 : node22754;
																assign node22754 = (inp[7]) ? 4'b0110 : 4'b0100;
															assign node22758 = (inp[12]) ? 4'b0010 : node22759;
																assign node22759 = (inp[7]) ? 4'b0010 : 4'b0000;
														assign node22763 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node22766 = (inp[12]) ? node22778 : node22767;
														assign node22767 = (inp[7]) ? node22773 : node22768;
															assign node22768 = (inp[13]) ? 4'b0100 : node22769;
																assign node22769 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node22773 = (inp[13]) ? 4'b0110 : node22774;
																assign node22774 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node22778 = (inp[7]) ? 4'b0101 : node22779;
															assign node22779 = (inp[13]) ? node22781 : 4'b0111;
																assign node22781 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node22785 = (inp[12]) ? node22811 : node22786;
													assign node22786 = (inp[7]) ? node22798 : node22787;
														assign node22787 = (inp[13]) ? node22791 : node22788;
															assign node22788 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node22791 = (inp[2]) ? node22795 : node22792;
																assign node22792 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node22795 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node22798 = (inp[5]) ? node22804 : node22799;
															assign node22799 = (inp[2]) ? 4'b0111 : node22800;
																assign node22800 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node22804 = (inp[2]) ? node22808 : node22805;
																assign node22805 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node22808 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node22811 = (inp[7]) ? node22825 : node22812;
														assign node22812 = (inp[5]) ? node22818 : node22813;
															assign node22813 = (inp[2]) ? 4'b0011 : node22814;
																assign node22814 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node22818 = (inp[2]) ? node22822 : node22819;
																assign node22819 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node22822 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node22825 = (inp[13]) ? 4'b0000 : node22826;
															assign node22826 = (inp[2]) ? node22830 : node22827;
																assign node22827 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node22830 = (inp[5]) ? 4'b0100 : 4'b0000;
							assign node22834 = (inp[2]) ? node23288 : node22835;
								assign node22835 = (inp[13]) ? node23087 : node22836;
									assign node22836 = (inp[7]) ? node22974 : node22837;
										assign node22837 = (inp[12]) ? node22909 : node22838;
											assign node22838 = (inp[5]) ? node22874 : node22839;
												assign node22839 = (inp[15]) ? node22845 : node22840;
													assign node22840 = (inp[11]) ? 4'b0000 : node22841;
														assign node22841 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node22845 = (inp[11]) ? node22861 : node22846;
														assign node22846 = (inp[0]) ? node22854 : node22847;
															assign node22847 = (inp[10]) ? node22851 : node22848;
																assign node22848 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node22851 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node22854 = (inp[10]) ? node22858 : node22855;
																assign node22855 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node22858 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node22861 = (inp[0]) ? node22867 : node22862;
															assign node22862 = (inp[9]) ? 4'b0100 : node22863;
																assign node22863 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node22867 = (inp[10]) ? node22871 : node22868;
																assign node22868 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node22871 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node22874 = (inp[15]) ? node22898 : node22875;
													assign node22875 = (inp[11]) ? node22889 : node22876;
														assign node22876 = (inp[10]) ? node22882 : node22877;
															assign node22877 = (inp[0]) ? node22879 : 4'b0101;
																assign node22879 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node22882 = (inp[9]) ? node22886 : node22883;
																assign node22883 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node22886 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node22889 = (inp[0]) ? node22891 : 4'b0100;
															assign node22891 = (inp[10]) ? node22895 : node22892;
																assign node22892 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node22895 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node22898 = (inp[9]) ? node22900 : 4'b0001;
														assign node22900 = (inp[10]) ? node22906 : node22901;
															assign node22901 = (inp[0]) ? 4'b0000 : node22902;
																assign node22902 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22906 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node22909 = (inp[15]) ? node22947 : node22910;
												assign node22910 = (inp[5]) ? node22928 : node22911;
													assign node22911 = (inp[10]) ? node22921 : node22912;
														assign node22912 = (inp[9]) ? node22916 : node22913;
															assign node22913 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node22916 = (inp[0]) ? node22918 : 4'b0110;
																assign node22918 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22921 = (inp[9]) ? node22925 : node22922;
															assign node22922 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node22925 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node22928 = (inp[0]) ? node22936 : node22929;
														assign node22929 = (inp[9]) ? node22933 : node22930;
															assign node22930 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node22933 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node22936 = (inp[9]) ? node22942 : node22937;
															assign node22937 = (inp[10]) ? 4'b0110 : node22938;
																assign node22938 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node22942 = (inp[11]) ? node22944 : 4'b0111;
																assign node22944 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node22947 = (inp[0]) ? node22961 : node22948;
													assign node22948 = (inp[5]) ? node22956 : node22949;
														assign node22949 = (inp[9]) ? node22953 : node22950;
															assign node22950 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node22953 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node22956 = (inp[10]) ? 4'b0011 : node22957;
															assign node22957 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node22961 = (inp[9]) ? 4'b0010 : node22962;
														assign node22962 = (inp[10]) ? node22968 : node22963;
															assign node22963 = (inp[5]) ? 4'b0011 : node22964;
																assign node22964 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22968 = (inp[11]) ? 4'b0010 : node22969;
																assign node22969 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node22974 = (inp[12]) ? node23046 : node22975;
											assign node22975 = (inp[5]) ? node23011 : node22976;
												assign node22976 = (inp[0]) ? node22990 : node22977;
													assign node22977 = (inp[15]) ? node22985 : node22978;
														assign node22978 = (inp[10]) ? node22982 : node22979;
															assign node22979 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node22982 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node22985 = (inp[10]) ? node22987 : 4'b0010;
															assign node22987 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node22990 = (inp[9]) ? node23002 : node22991;
														assign node22991 = (inp[11]) ? node22997 : node22992;
															assign node22992 = (inp[15]) ? 4'b0011 : node22993;
																assign node22993 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node22997 = (inp[15]) ? 4'b0010 : node22998;
																assign node22998 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node23002 = (inp[11]) ? 4'b0011 : node23003;
															assign node23003 = (inp[15]) ? node23007 : node23004;
																assign node23004 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node23007 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node23011 = (inp[10]) ? node23029 : node23012;
													assign node23012 = (inp[11]) ? node23020 : node23013;
														assign node23013 = (inp[9]) ? node23017 : node23014;
															assign node23014 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node23017 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node23020 = (inp[15]) ? 4'b0011 : node23021;
															assign node23021 = (inp[0]) ? node23025 : node23022;
																assign node23022 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node23025 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node23029 = (inp[9]) ? node23039 : node23030;
														assign node23030 = (inp[15]) ? node23036 : node23031;
															assign node23031 = (inp[11]) ? node23033 : 4'b0011;
																assign node23033 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node23036 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node23039 = (inp[15]) ? node23041 : 4'b0010;
															assign node23041 = (inp[0]) ? node23043 : 4'b0011;
																assign node23043 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node23046 = (inp[15]) ? node23066 : node23047;
												assign node23047 = (inp[10]) ? node23057 : node23048;
													assign node23048 = (inp[9]) ? node23052 : node23049;
														assign node23049 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23052 = (inp[0]) ? node23054 : 4'b0001;
															assign node23054 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node23057 = (inp[9]) ? node23063 : node23058;
														assign node23058 = (inp[0]) ? node23060 : 4'b0001;
															assign node23060 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node23063 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node23066 = (inp[10]) ? node23078 : node23067;
													assign node23067 = (inp[9]) ? node23073 : node23068;
														assign node23068 = (inp[11]) ? node23070 : 4'b0001;
															assign node23070 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node23073 = (inp[11]) ? node23075 : 4'b0000;
															assign node23075 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node23078 = (inp[9]) ? node23084 : node23079;
														assign node23079 = (inp[11]) ? node23081 : 4'b0000;
															assign node23081 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node23084 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node23087 = (inp[7]) ? node23221 : node23088;
										assign node23088 = (inp[12]) ? node23148 : node23089;
											assign node23089 = (inp[9]) ? node23119 : node23090;
												assign node23090 = (inp[0]) ? node23106 : node23091;
													assign node23091 = (inp[10]) ? node23099 : node23092;
														assign node23092 = (inp[11]) ? node23094 : 4'b0000;
															assign node23094 = (inp[5]) ? 4'b0101 : node23095;
																assign node23095 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node23099 = (inp[5]) ? node23103 : node23100;
															assign node23100 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node23103 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node23106 = (inp[10]) ? node23114 : node23107;
														assign node23107 = (inp[11]) ? node23111 : node23108;
															assign node23108 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node23111 = (inp[15]) ? 4'b0100 : 4'b0001;
														assign node23114 = (inp[5]) ? node23116 : 4'b0001;
															assign node23116 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node23119 = (inp[15]) ? node23135 : node23120;
													assign node23120 = (inp[5]) ? node23130 : node23121;
														assign node23121 = (inp[10]) ? node23125 : node23122;
															assign node23122 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node23125 = (inp[0]) ? 4'b0100 : node23126;
																assign node23126 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node23130 = (inp[10]) ? node23132 : 4'b0000;
															assign node23132 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node23135 = (inp[5]) ? node23143 : node23136;
														assign node23136 = (inp[10]) ? 4'b0000 : node23137;
															assign node23137 = (inp[0]) ? 4'b0001 : node23138;
																assign node23138 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node23143 = (inp[11]) ? 4'b0101 : node23144;
															assign node23144 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node23148 = (inp[15]) ? node23184 : node23149;
												assign node23149 = (inp[5]) ? node23163 : node23150;
													assign node23150 = (inp[10]) ? 4'b0011 : node23151;
														assign node23151 = (inp[9]) ? node23157 : node23152;
															assign node23152 = (inp[11]) ? node23154 : 4'b0010;
																assign node23154 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node23157 = (inp[11]) ? node23159 : 4'b0011;
																assign node23159 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node23163 = (inp[0]) ? node23171 : node23164;
														assign node23164 = (inp[10]) ? node23168 : node23165;
															assign node23165 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node23168 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node23171 = (inp[11]) ? node23179 : node23172;
															assign node23172 = (inp[9]) ? node23176 : node23173;
																assign node23173 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node23176 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node23179 = (inp[10]) ? node23181 : 4'b0011;
																assign node23181 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node23184 = (inp[5]) ? node23202 : node23185;
													assign node23185 = (inp[9]) ? node23197 : node23186;
														assign node23186 = (inp[10]) ? node23192 : node23187;
															assign node23187 = (inp[0]) ? 4'b0111 : node23188;
																assign node23188 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node23192 = (inp[11]) ? 4'b0110 : node23193;
																assign node23193 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node23197 = (inp[10]) ? 4'b0111 : node23198;
															assign node23198 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node23202 = (inp[0]) ? node23214 : node23203;
														assign node23203 = (inp[9]) ? node23209 : node23204;
															assign node23204 = (inp[10]) ? 4'b0110 : node23205;
																assign node23205 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node23209 = (inp[10]) ? 4'b0111 : node23210;
																assign node23210 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node23214 = (inp[10]) ? node23218 : node23215;
															assign node23215 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node23218 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node23221 = (inp[12]) ? node23245 : node23222;
											assign node23222 = (inp[10]) ? node23234 : node23223;
												assign node23223 = (inp[9]) ? node23229 : node23224;
													assign node23224 = (inp[11]) ? 4'b0110 : node23225;
														assign node23225 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node23229 = (inp[11]) ? 4'b0111 : node23230;
														assign node23230 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node23234 = (inp[9]) ? node23240 : node23235;
													assign node23235 = (inp[11]) ? 4'b0111 : node23236;
														assign node23236 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node23240 = (inp[11]) ? 4'b0110 : node23241;
														assign node23241 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node23245 = (inp[0]) ? node23261 : node23246;
												assign node23246 = (inp[10]) ? node23254 : node23247;
													assign node23247 = (inp[9]) ? node23251 : node23248;
														assign node23248 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node23251 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23254 = (inp[15]) ? node23256 : 4'b0100;
														assign node23256 = (inp[9]) ? node23258 : 4'b0100;
															assign node23258 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node23261 = (inp[5]) ? node23269 : node23262;
													assign node23262 = (inp[10]) ? node23266 : node23263;
														assign node23263 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node23266 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23269 = (inp[15]) ? node23283 : node23270;
														assign node23270 = (inp[11]) ? node23278 : node23271;
															assign node23271 = (inp[10]) ? node23275 : node23272;
																assign node23272 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node23275 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23278 = (inp[10]) ? node23280 : 4'b0100;
																assign node23280 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node23283 = (inp[9]) ? node23285 : 4'b0101;
															assign node23285 = (inp[10]) ? 4'b0100 : 4'b0101;
								assign node23288 = (inp[13]) ? node23548 : node23289;
									assign node23289 = (inp[7]) ? node23435 : node23290;
										assign node23290 = (inp[12]) ? node23378 : node23291;
											assign node23291 = (inp[0]) ? node23333 : node23292;
												assign node23292 = (inp[9]) ? node23318 : node23293;
													assign node23293 = (inp[10]) ? node23305 : node23294;
														assign node23294 = (inp[15]) ? node23300 : node23295;
															assign node23295 = (inp[5]) ? 4'b0000 : node23296;
																assign node23296 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node23300 = (inp[5]) ? 4'b0101 : node23301;
																assign node23301 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node23305 = (inp[15]) ? node23313 : node23306;
															assign node23306 = (inp[5]) ? node23310 : node23307;
																assign node23307 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node23310 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23313 = (inp[5]) ? 4'b0100 : node23314;
																assign node23314 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node23318 = (inp[10]) ? node23328 : node23319;
														assign node23319 = (inp[15]) ? node23325 : node23320;
															assign node23320 = (inp[5]) ? 4'b0001 : node23321;
																assign node23321 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node23325 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node23328 = (inp[5]) ? node23330 : 4'b0001;
															assign node23330 = (inp[15]) ? 4'b0101 : 4'b0001;
												assign node23333 = (inp[11]) ? node23351 : node23334;
													assign node23334 = (inp[10]) ? node23342 : node23335;
														assign node23335 = (inp[9]) ? 4'b0100 : node23336;
															assign node23336 = (inp[15]) ? node23338 : 4'b0000;
																assign node23338 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node23342 = (inp[9]) ? node23344 : 4'b0100;
															assign node23344 = (inp[15]) ? node23348 : node23345;
																assign node23345 = (inp[5]) ? 4'b0000 : 4'b0101;
																assign node23348 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node23351 = (inp[5]) ? node23367 : node23352;
														assign node23352 = (inp[15]) ? node23360 : node23353;
															assign node23353 = (inp[9]) ? node23357 : node23354;
																assign node23354 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node23357 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node23360 = (inp[9]) ? node23364 : node23361;
																assign node23361 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node23364 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23367 = (inp[15]) ? node23375 : node23368;
															assign node23368 = (inp[9]) ? node23372 : node23369;
																assign node23369 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node23372 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node23375 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node23378 = (inp[15]) ? node23402 : node23379;
												assign node23379 = (inp[10]) ? node23393 : node23380;
													assign node23380 = (inp[5]) ? node23386 : node23381;
														assign node23381 = (inp[9]) ? node23383 : 4'b0011;
															assign node23383 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node23386 = (inp[9]) ? node23388 : 4'b0010;
															assign node23388 = (inp[0]) ? node23390 : 4'b0011;
																assign node23390 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node23393 = (inp[11]) ? 4'b0010 : node23394;
														assign node23394 = (inp[5]) ? node23398 : node23395;
															assign node23395 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node23398 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node23402 = (inp[9]) ? node23416 : node23403;
													assign node23403 = (inp[5]) ? node23407 : node23404;
														assign node23404 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node23407 = (inp[0]) ? node23413 : node23408;
															assign node23408 = (inp[11]) ? 4'b0111 : node23409;
																assign node23409 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node23413 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node23416 = (inp[5]) ? node23424 : node23417;
														assign node23417 = (inp[10]) ? 4'b0111 : node23418;
															assign node23418 = (inp[0]) ? 4'b0110 : node23419;
																assign node23419 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node23424 = (inp[10]) ? node23430 : node23425;
															assign node23425 = (inp[11]) ? 4'b0111 : node23426;
																assign node23426 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node23430 = (inp[0]) ? 4'b0110 : node23431;
																assign node23431 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node23435 = (inp[12]) ? node23489 : node23436;
											assign node23436 = (inp[10]) ? node23468 : node23437;
												assign node23437 = (inp[5]) ? node23453 : node23438;
													assign node23438 = (inp[15]) ? node23448 : node23439;
														assign node23439 = (inp[9]) ? node23445 : node23440;
															assign node23440 = (inp[0]) ? 4'b0111 : node23441;
																assign node23441 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node23445 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node23448 = (inp[9]) ? 4'b0111 : node23449;
															assign node23449 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node23453 = (inp[9]) ? node23461 : node23454;
														assign node23454 = (inp[15]) ? 4'b0110 : node23455;
															assign node23455 = (inp[11]) ? 4'b0111 : node23456;
																assign node23456 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node23461 = (inp[15]) ? 4'b0111 : node23462;
															assign node23462 = (inp[0]) ? 4'b0110 : node23463;
																assign node23463 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node23468 = (inp[9]) ? node23478 : node23469;
													assign node23469 = (inp[0]) ? 4'b0110 : node23470;
														assign node23470 = (inp[15]) ? node23474 : node23471;
															assign node23471 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node23474 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node23478 = (inp[15]) ? node23484 : node23479;
														assign node23479 = (inp[11]) ? 4'b0111 : node23480;
															assign node23480 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node23484 = (inp[11]) ? 4'b0110 : node23485;
															assign node23485 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node23489 = (inp[5]) ? node23519 : node23490;
												assign node23490 = (inp[9]) ? node23508 : node23491;
													assign node23491 = (inp[11]) ? node23501 : node23492;
														assign node23492 = (inp[10]) ? 4'b0101 : node23493;
															assign node23493 = (inp[15]) ? node23497 : node23494;
																assign node23494 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node23497 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node23501 = (inp[0]) ? node23503 : 4'b0100;
															assign node23503 = (inp[15]) ? 4'b0101 : node23504;
																assign node23504 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node23508 = (inp[10]) ? 4'b0101 : node23509;
														assign node23509 = (inp[15]) ? node23513 : node23510;
															assign node23510 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node23513 = (inp[11]) ? 4'b0101 : node23514;
																assign node23514 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node23519 = (inp[10]) ? node23535 : node23520;
													assign node23520 = (inp[15]) ? node23528 : node23521;
														assign node23521 = (inp[9]) ? node23523 : 4'b0101;
															assign node23523 = (inp[11]) ? 4'b0100 : node23524;
																assign node23524 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node23528 = (inp[9]) ? node23530 : 4'b0100;
															assign node23530 = (inp[0]) ? 4'b0101 : node23531;
																assign node23531 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23535 = (inp[15]) ? node23541 : node23536;
														assign node23536 = (inp[9]) ? node23538 : 4'b0100;
															assign node23538 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node23541 = (inp[9]) ? node23543 : 4'b0101;
															assign node23543 = (inp[11]) ? 4'b0100 : node23544;
																assign node23544 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node23548 = (inp[7]) ? node23682 : node23549;
										assign node23549 = (inp[12]) ? node23607 : node23550;
											assign node23550 = (inp[9]) ? node23580 : node23551;
												assign node23551 = (inp[10]) ? node23565 : node23552;
													assign node23552 = (inp[5]) ? node23558 : node23553;
														assign node23553 = (inp[15]) ? 4'b0100 : node23554;
															assign node23554 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node23558 = (inp[15]) ? 4'b0001 : node23559;
															assign node23559 = (inp[11]) ? node23561 : 4'b0101;
																assign node23561 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node23565 = (inp[5]) ? node23573 : node23566;
														assign node23566 = (inp[15]) ? 4'b0101 : node23567;
															assign node23567 = (inp[11]) ? 4'b0001 : node23568;
																assign node23568 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23573 = (inp[15]) ? node23575 : 4'b0100;
															assign node23575 = (inp[11]) ? node23577 : 4'b0000;
																assign node23577 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node23580 = (inp[10]) ? node23596 : node23581;
													assign node23581 = (inp[11]) ? node23589 : node23582;
														assign node23582 = (inp[15]) ? node23586 : node23583;
															assign node23583 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node23586 = (inp[5]) ? 4'b0000 : 4'b0101;
														assign node23589 = (inp[15]) ? node23591 : 4'b0001;
															assign node23591 = (inp[5]) ? node23593 : 4'b0100;
																assign node23593 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node23596 = (inp[5]) ? node23604 : node23597;
														assign node23597 = (inp[15]) ? node23601 : node23598;
															assign node23598 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node23601 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node23604 = (inp[15]) ? 4'b0000 : 4'b0101;
											assign node23607 = (inp[15]) ? node23647 : node23608;
												assign node23608 = (inp[5]) ? node23632 : node23609;
													assign node23609 = (inp[0]) ? node23621 : node23610;
														assign node23610 = (inp[11]) ? node23616 : node23611;
															assign node23611 = (inp[10]) ? 4'b0110 : node23612;
																assign node23612 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node23616 = (inp[10]) ? 4'b0111 : node23617;
																assign node23617 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node23621 = (inp[11]) ? node23627 : node23622;
															assign node23622 = (inp[9]) ? node23624 : 4'b0110;
																assign node23624 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node23627 = (inp[9]) ? 4'b0110 : node23628;
																assign node23628 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node23632 = (inp[0]) ? node23640 : node23633;
														assign node23633 = (inp[10]) ? 4'b0111 : node23634;
															assign node23634 = (inp[9]) ? node23636 : 4'b0111;
																assign node23636 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node23640 = (inp[11]) ? node23642 : 4'b0111;
															assign node23642 = (inp[10]) ? 4'b0110 : node23643;
																assign node23643 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node23647 = (inp[10]) ? node23669 : node23648;
													assign node23648 = (inp[0]) ? node23664 : node23649;
														assign node23649 = (inp[9]) ? node23657 : node23650;
															assign node23650 = (inp[11]) ? node23654 : node23651;
																assign node23651 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node23654 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node23657 = (inp[5]) ? node23661 : node23658;
																assign node23658 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node23661 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node23664 = (inp[9]) ? 4'b0011 : node23665;
															assign node23665 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node23669 = (inp[9]) ? 4'b0010 : node23670;
														assign node23670 = (inp[5]) ? node23676 : node23671;
															assign node23671 = (inp[0]) ? 4'b0010 : node23672;
																assign node23672 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node23676 = (inp[0]) ? 4'b0011 : node23677;
																assign node23677 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node23682 = (inp[12]) ? node23706 : node23683;
											assign node23683 = (inp[9]) ? node23695 : node23684;
												assign node23684 = (inp[10]) ? node23690 : node23685;
													assign node23685 = (inp[0]) ? 4'b0010 : node23686;
														assign node23686 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node23690 = (inp[11]) ? 4'b0011 : node23691;
														assign node23691 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node23695 = (inp[10]) ? node23701 : node23696;
													assign node23696 = (inp[0]) ? 4'b0011 : node23697;
														assign node23697 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node23701 = (inp[0]) ? 4'b0010 : node23702;
														assign node23702 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node23706 = (inp[5]) ? node23744 : node23707;
												assign node23707 = (inp[11]) ? node23729 : node23708;
													assign node23708 = (inp[15]) ? node23714 : node23709;
														assign node23709 = (inp[9]) ? node23711 : 4'b0000;
															assign node23711 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23714 = (inp[0]) ? node23722 : node23715;
															assign node23715 = (inp[10]) ? node23719 : node23716;
																assign node23716 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node23719 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node23722 = (inp[9]) ? node23726 : node23723;
																assign node23723 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node23726 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node23729 = (inp[0]) ? node23737 : node23730;
														assign node23730 = (inp[9]) ? node23734 : node23731;
															assign node23731 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node23734 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23737 = (inp[9]) ? node23741 : node23738;
															assign node23738 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node23741 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node23744 = (inp[10]) ? node23756 : node23745;
													assign node23745 = (inp[9]) ? node23751 : node23746;
														assign node23746 = (inp[0]) ? 4'b0000 : node23747;
															assign node23747 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node23751 = (inp[0]) ? 4'b0001 : node23752;
															assign node23752 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node23756 = (inp[9]) ? node23758 : 4'b0001;
														assign node23758 = (inp[15]) ? node23760 : 4'b0000;
															assign node23760 = (inp[11]) ? 4'b0000 : 4'b0001;
				assign node23763 = (inp[7]) ? node25929 : node23764;
					assign node23764 = (inp[4]) ? node24822 : node23765;
						assign node23765 = (inp[3]) ? node24147 : node23766;
							assign node23766 = (inp[2]) ? node23948 : node23767;
								assign node23767 = (inp[9]) ? node23857 : node23768;
									assign node23768 = (inp[0]) ? node23806 : node23769;
										assign node23769 = (inp[13]) ? node23787 : node23770;
											assign node23770 = (inp[1]) ? node23774 : node23771;
												assign node23771 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node23774 = (inp[5]) ? node23782 : node23775;
													assign node23775 = (inp[12]) ? node23779 : node23776;
														assign node23776 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node23779 = (inp[15]) ? 4'b0000 : 4'b0101;
													assign node23782 = (inp[12]) ? node23784 : 4'b0101;
														assign node23784 = (inp[15]) ? 4'b0000 : 4'b0101;
											assign node23787 = (inp[12]) ? node23793 : node23788;
												assign node23788 = (inp[15]) ? node23790 : 4'b0100;
													assign node23790 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node23793 = (inp[15]) ? node23801 : node23794;
													assign node23794 = (inp[5]) ? node23798 : node23795;
														assign node23795 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node23798 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node23801 = (inp[1]) ? 4'b0101 : node23802;
														assign node23802 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node23806 = (inp[5]) ? node23832 : node23807;
											assign node23807 = (inp[12]) ? node23819 : node23808;
												assign node23808 = (inp[13]) ? node23814 : node23809;
													assign node23809 = (inp[15]) ? node23811 : 4'b0000;
														assign node23811 = (inp[1]) ? 4'b0101 : 4'b0000;
													assign node23814 = (inp[15]) ? node23816 : 4'b0100;
														assign node23816 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node23819 = (inp[13]) ? node23825 : node23820;
													assign node23820 = (inp[1]) ? node23822 : 4'b0100;
														assign node23822 = (inp[15]) ? 4'b0000 : 4'b0101;
													assign node23825 = (inp[1]) ? node23829 : node23826;
														assign node23826 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node23829 = (inp[15]) ? 4'b0101 : 4'b0000;
											assign node23832 = (inp[13]) ? node23844 : node23833;
												assign node23833 = (inp[12]) ? node23839 : node23834;
													assign node23834 = (inp[1]) ? node23836 : 4'b0001;
														assign node23836 = (inp[15]) ? 4'b0101 : 4'b0001;
													assign node23839 = (inp[1]) ? node23841 : 4'b0101;
														assign node23841 = (inp[15]) ? 4'b0001 : 4'b0100;
												assign node23844 = (inp[12]) ? node23850 : node23845;
													assign node23845 = (inp[15]) ? node23847 : 4'b0101;
														assign node23847 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node23850 = (inp[15]) ? node23854 : node23851;
														assign node23851 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node23854 = (inp[1]) ? 4'b0100 : 4'b0000;
									assign node23857 = (inp[0]) ? node23893 : node23858;
										assign node23858 = (inp[12]) ? node23872 : node23859;
											assign node23859 = (inp[13]) ? node23867 : node23860;
												assign node23860 = (inp[15]) ? node23862 : 4'b0001;
													assign node23862 = (inp[1]) ? node23864 : 4'b0001;
														assign node23864 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node23867 = (inp[15]) ? node23869 : 4'b0101;
													assign node23869 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node23872 = (inp[13]) ? node23878 : node23873;
												assign node23873 = (inp[1]) ? node23875 : 4'b0101;
													assign node23875 = (inp[15]) ? 4'b0001 : 4'b0100;
												assign node23878 = (inp[5]) ? node23886 : node23879;
													assign node23879 = (inp[15]) ? node23883 : node23880;
														assign node23880 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node23883 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node23886 = (inp[1]) ? node23890 : node23887;
														assign node23887 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node23890 = (inp[15]) ? 4'b0100 : 4'b0001;
										assign node23893 = (inp[5]) ? node23923 : node23894;
											assign node23894 = (inp[15]) ? node23906 : node23895;
												assign node23895 = (inp[12]) ? node23899 : node23896;
													assign node23896 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node23899 = (inp[13]) ? node23903 : node23900;
														assign node23900 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node23903 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node23906 = (inp[1]) ? node23914 : node23907;
													assign node23907 = (inp[12]) ? node23911 : node23908;
														assign node23908 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node23911 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node23914 = (inp[11]) ? 4'b0100 : node23915;
														assign node23915 = (inp[12]) ? node23919 : node23916;
															assign node23916 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node23919 = (inp[13]) ? 4'b0100 : 4'b0001;
											assign node23923 = (inp[12]) ? node23935 : node23924;
												assign node23924 = (inp[13]) ? node23930 : node23925;
													assign node23925 = (inp[15]) ? node23927 : 4'b0000;
														assign node23927 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node23930 = (inp[15]) ? node23932 : 4'b0100;
														assign node23932 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node23935 = (inp[13]) ? node23941 : node23936;
													assign node23936 = (inp[1]) ? node23938 : 4'b0100;
														assign node23938 = (inp[15]) ? 4'b0000 : 4'b0101;
													assign node23941 = (inp[1]) ? node23945 : node23942;
														assign node23942 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node23945 = (inp[15]) ? 4'b0101 : 4'b0001;
								assign node23948 = (inp[9]) ? node24046 : node23949;
									assign node23949 = (inp[5]) ? node23989 : node23950;
										assign node23950 = (inp[12]) ? node23964 : node23951;
											assign node23951 = (inp[13]) ? node23959 : node23952;
												assign node23952 = (inp[1]) ? node23954 : 4'b0001;
													assign node23954 = (inp[15]) ? node23956 : 4'b0001;
														assign node23956 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node23959 = (inp[15]) ? node23961 : 4'b0101;
													assign node23961 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node23964 = (inp[1]) ? node23974 : node23965;
												assign node23965 = (inp[13]) ? node23967 : 4'b0101;
													assign node23967 = (inp[15]) ? node23971 : node23968;
														assign node23968 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node23971 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node23974 = (inp[0]) ? node23982 : node23975;
													assign node23975 = (inp[13]) ? node23979 : node23976;
														assign node23976 = (inp[15]) ? 4'b0001 : 4'b0100;
														assign node23979 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node23982 = (inp[15]) ? node23986 : node23983;
														assign node23983 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node23986 = (inp[13]) ? 4'b0100 : 4'b0001;
										assign node23989 = (inp[0]) ? node24017 : node23990;
											assign node23990 = (inp[15]) ? node24002 : node23991;
												assign node23991 = (inp[12]) ? node23995 : node23992;
													assign node23992 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node23995 = (inp[13]) ? node23999 : node23996;
														assign node23996 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node23999 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node24002 = (inp[1]) ? node24010 : node24003;
													assign node24003 = (inp[13]) ? node24007 : node24004;
														assign node24004 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node24007 = (inp[12]) ? 4'b0001 : 4'b0100;
													assign node24010 = (inp[12]) ? node24014 : node24011;
														assign node24011 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node24014 = (inp[13]) ? 4'b0100 : 4'b0001;
											assign node24017 = (inp[12]) ? node24031 : node24018;
												assign node24018 = (inp[13]) ? node24024 : node24019;
													assign node24019 = (inp[1]) ? node24021 : 4'b0000;
														assign node24021 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node24024 = (inp[1]) ? node24028 : node24025;
														assign node24025 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node24028 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node24031 = (inp[13]) ? node24039 : node24032;
													assign node24032 = (inp[15]) ? node24036 : node24033;
														assign node24033 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node24036 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node24039 = (inp[15]) ? node24043 : node24040;
														assign node24040 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node24043 = (inp[1]) ? 4'b0101 : 4'b0001;
									assign node24046 = (inp[5]) ? node24082 : node24047;
										assign node24047 = (inp[12]) ? node24061 : node24048;
											assign node24048 = (inp[13]) ? node24056 : node24049;
												assign node24049 = (inp[15]) ? node24051 : 4'b0000;
													assign node24051 = (inp[1]) ? node24053 : 4'b0000;
														assign node24053 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node24056 = (inp[15]) ? node24058 : 4'b0100;
													assign node24058 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node24061 = (inp[13]) ? node24069 : node24062;
												assign node24062 = (inp[15]) ? node24066 : node24063;
													assign node24063 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node24066 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node24069 = (inp[15]) ? node24077 : node24070;
													assign node24070 = (inp[0]) ? node24074 : node24071;
														assign node24071 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node24074 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node24077 = (inp[1]) ? 4'b0101 : node24078;
														assign node24078 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node24082 = (inp[0]) ? node24120 : node24083;
											assign node24083 = (inp[15]) ? node24095 : node24084;
												assign node24084 = (inp[12]) ? node24088 : node24085;
													assign node24085 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node24088 = (inp[13]) ? node24092 : node24089;
														assign node24089 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node24092 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node24095 = (inp[13]) ? node24103 : node24096;
													assign node24096 = (inp[12]) ? node24100 : node24097;
														assign node24097 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node24100 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node24103 = (inp[10]) ? node24111 : node24104;
														assign node24104 = (inp[12]) ? node24108 : node24105;
															assign node24105 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node24108 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node24111 = (inp[11]) ? 4'b0101 : node24112;
															assign node24112 = (inp[1]) ? node24116 : node24113;
																assign node24113 = (inp[12]) ? 4'b0000 : 4'b0101;
																assign node24116 = (inp[12]) ? 4'b0101 : 4'b0000;
											assign node24120 = (inp[12]) ? node24134 : node24121;
												assign node24121 = (inp[13]) ? node24127 : node24122;
													assign node24122 = (inp[15]) ? node24124 : 4'b0001;
														assign node24124 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node24127 = (inp[1]) ? node24131 : node24128;
														assign node24128 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node24131 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node24134 = (inp[13]) ? node24140 : node24135;
													assign node24135 = (inp[15]) ? 4'b0001 : node24136;
														assign node24136 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node24140 = (inp[1]) ? node24144 : node24141;
														assign node24141 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node24144 = (inp[11]) ? 4'b0000 : 4'b0100;
							assign node24147 = (inp[0]) ? node24441 : node24148;
								assign node24148 = (inp[15]) ? node24276 : node24149;
									assign node24149 = (inp[13]) ? node24201 : node24150;
										assign node24150 = (inp[2]) ? node24170 : node24151;
											assign node24151 = (inp[9]) ? node24161 : node24152;
												assign node24152 = (inp[12]) ? node24156 : node24153;
													assign node24153 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node24156 = (inp[1]) ? node24158 : 4'b0110;
														assign node24158 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node24161 = (inp[1]) ? node24165 : node24162;
													assign node24162 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node24165 = (inp[12]) ? node24167 : 4'b0111;
														assign node24167 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node24170 = (inp[9]) ? node24192 : node24171;
												assign node24171 = (inp[5]) ? node24179 : node24172;
													assign node24172 = (inp[1]) ? node24176 : node24173;
														assign node24173 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node24176 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node24179 = (inp[11]) ? node24187 : node24180;
														assign node24180 = (inp[10]) ? node24182 : 4'b0011;
															assign node24182 = (inp[1]) ? 4'b0011 : node24183;
																assign node24183 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node24187 = (inp[1]) ? node24189 : 4'b0011;
															assign node24189 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node24192 = (inp[12]) ? node24196 : node24193;
													assign node24193 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node24196 = (inp[1]) ? node24198 : 4'b0110;
														assign node24198 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node24201 = (inp[9]) ? node24243 : node24202;
											assign node24202 = (inp[2]) ? node24222 : node24203;
												assign node24203 = (inp[11]) ? node24213 : node24204;
													assign node24204 = (inp[1]) ? node24210 : node24205;
														assign node24205 = (inp[12]) ? 4'b0011 : node24206;
															assign node24206 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24210 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node24213 = (inp[1]) ? node24219 : node24214;
														assign node24214 = (inp[12]) ? 4'b0011 : node24215;
															assign node24215 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24219 = (inp[12]) ? 4'b0110 : 4'b0011;
												assign node24222 = (inp[11]) ? node24234 : node24223;
													assign node24223 = (inp[10]) ? node24225 : 4'b0010;
														assign node24225 = (inp[5]) ? node24231 : node24226;
															assign node24226 = (inp[1]) ? 4'b0010 : node24227;
																assign node24227 = (inp[12]) ? 4'b0010 : 4'b0111;
															assign node24231 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node24234 = (inp[12]) ? node24240 : node24235;
														assign node24235 = (inp[10]) ? 4'b0010 : node24236;
															assign node24236 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node24240 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node24243 = (inp[2]) ? node24253 : node24244;
												assign node24244 = (inp[12]) ? node24250 : node24245;
													assign node24245 = (inp[1]) ? 4'b0010 : node24246;
														assign node24246 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node24250 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node24253 = (inp[5]) ? node24269 : node24254;
													assign node24254 = (inp[10]) ? node24262 : node24255;
														assign node24255 = (inp[12]) ? node24259 : node24256;
															assign node24256 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node24259 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node24262 = (inp[11]) ? node24264 : 4'b0110;
															assign node24264 = (inp[1]) ? node24266 : 4'b0011;
																assign node24266 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node24269 = (inp[1]) ? node24273 : node24270;
														assign node24270 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node24273 = (inp[12]) ? 4'b0110 : 4'b0011;
									assign node24276 = (inp[13]) ? node24340 : node24277;
										assign node24277 = (inp[12]) ? node24333 : node24278;
											assign node24278 = (inp[10]) ? node24302 : node24279;
												assign node24279 = (inp[2]) ? node24289 : node24280;
													assign node24280 = (inp[11]) ? node24282 : 4'b0010;
														assign node24282 = (inp[1]) ? node24286 : node24283;
															assign node24283 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node24286 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node24289 = (inp[11]) ? node24295 : node24290;
														assign node24290 = (inp[1]) ? 4'b0011 : node24291;
															assign node24291 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24295 = (inp[5]) ? 4'b0010 : node24296;
															assign node24296 = (inp[9]) ? node24298 : 4'b0011;
																assign node24298 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node24302 = (inp[9]) ? node24324 : node24303;
													assign node24303 = (inp[11]) ? node24317 : node24304;
														assign node24304 = (inp[5]) ? node24312 : node24305;
															assign node24305 = (inp[1]) ? node24309 : node24306;
																assign node24306 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node24309 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24312 = (inp[2]) ? node24314 : 4'b0011;
																assign node24314 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node24317 = (inp[1]) ? node24321 : node24318;
															assign node24318 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24321 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node24324 = (inp[11]) ? node24326 : 4'b0011;
														assign node24326 = (inp[2]) ? node24330 : node24327;
															assign node24327 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node24330 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node24333 = (inp[2]) ? node24337 : node24334;
												assign node24334 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node24337 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node24340 = (inp[12]) ? node24404 : node24341;
											assign node24341 = (inp[10]) ? node24367 : node24342;
												assign node24342 = (inp[1]) ? node24352 : node24343;
													assign node24343 = (inp[9]) ? node24345 : 4'b0110;
														assign node24345 = (inp[5]) ? node24349 : node24346;
															assign node24346 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node24349 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node24352 = (inp[2]) ? node24362 : node24353;
														assign node24353 = (inp[11]) ? node24355 : 4'b0111;
															assign node24355 = (inp[9]) ? node24359 : node24356;
																assign node24356 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node24359 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node24362 = (inp[5]) ? 4'b0110 : node24363;
															assign node24363 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node24367 = (inp[1]) ? node24381 : node24368;
													assign node24368 = (inp[5]) ? node24376 : node24369;
														assign node24369 = (inp[2]) ? node24373 : node24370;
															assign node24370 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node24373 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node24376 = (inp[2]) ? 4'b0111 : node24377;
															assign node24377 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node24381 = (inp[9]) ? node24397 : node24382;
														assign node24382 = (inp[11]) ? node24390 : node24383;
															assign node24383 = (inp[2]) ? node24387 : node24384;
																assign node24384 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node24387 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24390 = (inp[5]) ? node24394 : node24391;
																assign node24391 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node24394 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24397 = (inp[2]) ? node24401 : node24398;
															assign node24398 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24401 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node24404 = (inp[1]) ? node24434 : node24405;
												assign node24405 = (inp[5]) ? node24415 : node24406;
													assign node24406 = (inp[10]) ? 4'b0010 : node24407;
														assign node24407 = (inp[11]) ? 4'b0011 : node24408;
															assign node24408 = (inp[2]) ? 4'b0010 : node24409;
																assign node24409 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node24415 = (inp[10]) ? node24421 : node24416;
														assign node24416 = (inp[2]) ? node24418 : 4'b0010;
															assign node24418 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node24421 = (inp[11]) ? node24429 : node24422;
															assign node24422 = (inp[9]) ? node24426 : node24423;
																assign node24423 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node24426 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24429 = (inp[9]) ? 4'b0011 : node24430;
																assign node24430 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node24434 = (inp[2]) ? node24438 : node24435;
													assign node24435 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node24438 = (inp[9]) ? 4'b0010 : 4'b0011;
								assign node24441 = (inp[13]) ? node24647 : node24442;
									assign node24442 = (inp[12]) ? node24554 : node24443;
										assign node24443 = (inp[1]) ? node24489 : node24444;
											assign node24444 = (inp[11]) ? node24460 : node24445;
												assign node24445 = (inp[5]) ? node24453 : node24446;
													assign node24446 = (inp[2]) ? node24450 : node24447;
														assign node24447 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24450 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node24453 = (inp[2]) ? node24457 : node24454;
														assign node24454 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24457 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node24460 = (inp[15]) ? node24476 : node24461;
													assign node24461 = (inp[9]) ? node24471 : node24462;
														assign node24462 = (inp[10]) ? node24464 : 4'b0010;
															assign node24464 = (inp[5]) ? node24468 : node24465;
																assign node24465 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node24468 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24471 = (inp[5]) ? node24473 : 4'b0011;
															assign node24473 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node24476 = (inp[5]) ? node24484 : node24477;
														assign node24477 = (inp[10]) ? 4'b0010 : node24478;
															assign node24478 = (inp[2]) ? 4'b0011 : node24479;
																assign node24479 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24484 = (inp[2]) ? node24486 : 4'b0011;
															assign node24486 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node24489 = (inp[15]) ? node24529 : node24490;
												assign node24490 = (inp[2]) ? node24512 : node24491;
													assign node24491 = (inp[10]) ? node24505 : node24492;
														assign node24492 = (inp[11]) ? node24498 : node24493;
															assign node24493 = (inp[9]) ? 4'b0111 : node24494;
																assign node24494 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24498 = (inp[9]) ? node24502 : node24499;
																assign node24499 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node24502 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24505 = (inp[9]) ? node24509 : node24506;
															assign node24506 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24509 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24512 = (inp[11]) ? node24522 : node24513;
														assign node24513 = (inp[10]) ? 4'b0111 : node24514;
															assign node24514 = (inp[5]) ? node24518 : node24515;
																assign node24515 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node24518 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node24522 = (inp[9]) ? node24526 : node24523;
															assign node24523 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node24526 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node24529 = (inp[5]) ? node24543 : node24530;
													assign node24530 = (inp[10]) ? node24538 : node24531;
														assign node24531 = (inp[9]) ? node24535 : node24532;
															assign node24532 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24535 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node24538 = (inp[9]) ? 4'b0010 : node24539;
															assign node24539 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node24543 = (inp[11]) ? node24551 : node24544;
														assign node24544 = (inp[10]) ? node24546 : 4'b0011;
															assign node24546 = (inp[2]) ? 4'b0011 : node24547;
																assign node24547 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24551 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node24554 = (inp[1]) ? node24608 : node24555;
											assign node24555 = (inp[11]) ? node24585 : node24556;
												assign node24556 = (inp[9]) ? node24564 : node24557;
													assign node24557 = (inp[2]) ? node24561 : node24558;
														assign node24558 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node24561 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24564 = (inp[10]) ? node24572 : node24565;
														assign node24565 = (inp[15]) ? 4'b0111 : node24566;
															assign node24566 = (inp[2]) ? node24568 : 4'b0111;
																assign node24568 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node24572 = (inp[15]) ? node24578 : node24573;
															assign node24573 = (inp[2]) ? 4'b0111 : node24574;
																assign node24574 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node24578 = (inp[5]) ? node24582 : node24579;
																assign node24579 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node24582 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node24585 = (inp[9]) ? node24601 : node24586;
													assign node24586 = (inp[15]) ? node24594 : node24587;
														assign node24587 = (inp[5]) ? node24591 : node24588;
															assign node24588 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node24591 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node24594 = (inp[5]) ? node24598 : node24595;
															assign node24595 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node24598 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node24601 = (inp[2]) ? node24605 : node24602;
														assign node24602 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24605 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node24608 = (inp[15]) ? node24632 : node24609;
												assign node24609 = (inp[10]) ? node24617 : node24610;
													assign node24610 = (inp[2]) ? node24614 : node24611;
														assign node24611 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24614 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node24617 = (inp[5]) ? node24619 : 4'b0010;
														assign node24619 = (inp[11]) ? node24627 : node24620;
															assign node24620 = (inp[9]) ? node24624 : node24621;
																assign node24621 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node24624 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24627 = (inp[2]) ? node24629 : 4'b0010;
																assign node24629 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node24632 = (inp[5]) ? node24640 : node24633;
													assign node24633 = (inp[9]) ? node24637 : node24634;
														assign node24634 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24637 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node24640 = (inp[2]) ? node24644 : node24641;
														assign node24641 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node24644 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node24647 = (inp[12]) ? node24689 : node24648;
										assign node24648 = (inp[1]) ? node24664 : node24649;
											assign node24649 = (inp[2]) ? node24657 : node24650;
												assign node24650 = (inp[9]) ? node24654 : node24651;
													assign node24651 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node24654 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node24657 = (inp[15]) ? node24661 : node24658;
													assign node24658 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node24661 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node24664 = (inp[15]) ? node24682 : node24665;
												assign node24665 = (inp[5]) ? node24675 : node24666;
													assign node24666 = (inp[11]) ? node24668 : 4'b0010;
														assign node24668 = (inp[2]) ? node24672 : node24669;
															assign node24669 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node24672 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node24675 = (inp[2]) ? node24679 : node24676;
														assign node24676 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24679 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node24682 = (inp[2]) ? node24686 : node24683;
													assign node24683 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node24686 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node24689 = (inp[1]) ? node24751 : node24690;
											assign node24690 = (inp[15]) ? node24736 : node24691;
												assign node24691 = (inp[10]) ? node24709 : node24692;
													assign node24692 = (inp[9]) ? node24698 : node24693;
														assign node24693 = (inp[11]) ? 4'b0010 : node24694;
															assign node24694 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24698 = (inp[11]) ? node24704 : node24699;
															assign node24699 = (inp[5]) ? 4'b0010 : node24700;
																assign node24700 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24704 = (inp[2]) ? 4'b0011 : node24705;
																assign node24705 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node24709 = (inp[9]) ? node24725 : node24710;
														assign node24710 = (inp[11]) ? node24718 : node24711;
															assign node24711 = (inp[2]) ? node24715 : node24712;
																assign node24712 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node24715 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node24718 = (inp[5]) ? node24722 : node24719;
																assign node24719 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node24722 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node24725 = (inp[11]) ? node24731 : node24726;
															assign node24726 = (inp[2]) ? node24728 : 4'b0010;
																assign node24728 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node24731 = (inp[2]) ? 4'b0010 : node24732;
																assign node24732 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node24736 = (inp[9]) ? node24744 : node24737;
													assign node24737 = (inp[10]) ? 4'b0011 : node24738;
														assign node24738 = (inp[5]) ? 4'b0011 : node24739;
															assign node24739 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node24744 = (inp[2]) ? node24748 : node24745;
														assign node24745 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24748 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node24751 = (inp[15]) ? node24787 : node24752;
												assign node24752 = (inp[11]) ? node24772 : node24753;
													assign node24753 = (inp[10]) ? node24765 : node24754;
														assign node24754 = (inp[5]) ? node24760 : node24755;
															assign node24755 = (inp[9]) ? 4'b0110 : node24756;
																assign node24756 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node24760 = (inp[9]) ? 4'b0111 : node24761;
																assign node24761 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node24765 = (inp[9]) ? 4'b0111 : node24766;
															assign node24766 = (inp[5]) ? 4'b0111 : node24767;
																assign node24767 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node24772 = (inp[10]) ? 4'b0110 : node24773;
														assign node24773 = (inp[9]) ? node24779 : node24774;
															assign node24774 = (inp[5]) ? 4'b0110 : node24775;
																assign node24775 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node24779 = (inp[5]) ? node24783 : node24780;
																assign node24780 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node24783 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node24787 = (inp[5]) ? node24805 : node24788;
													assign node24788 = (inp[11]) ? node24798 : node24789;
														assign node24789 = (inp[10]) ? 4'b0011 : node24790;
															assign node24790 = (inp[9]) ? node24794 : node24791;
																assign node24791 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node24794 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24798 = (inp[10]) ? node24800 : 4'b0011;
															assign node24800 = (inp[2]) ? 4'b0010 : node24801;
																assign node24801 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node24805 = (inp[10]) ? node24815 : node24806;
														assign node24806 = (inp[11]) ? node24812 : node24807;
															assign node24807 = (inp[9]) ? node24809 : 4'b0010;
																assign node24809 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24812 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24815 = (inp[2]) ? node24819 : node24816;
															assign node24816 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node24819 = (inp[9]) ? 4'b0010 : 4'b0011;
						assign node24822 = (inp[12]) ? node25424 : node24823;
							assign node24823 = (inp[13]) ? node25075 : node24824;
								assign node24824 = (inp[15]) ? node24928 : node24825;
									assign node24825 = (inp[0]) ? node24833 : node24826;
										assign node24826 = (inp[5]) ? node24830 : node24827;
											assign node24827 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node24830 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node24833 = (inp[1]) ? node24887 : node24834;
											assign node24834 = (inp[10]) ? node24860 : node24835;
												assign node24835 = (inp[5]) ? node24853 : node24836;
													assign node24836 = (inp[11]) ? node24844 : node24837;
														assign node24837 = (inp[9]) ? node24841 : node24838;
															assign node24838 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node24841 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node24844 = (inp[2]) ? node24846 : 4'b0010;
															assign node24846 = (inp[9]) ? node24850 : node24847;
																assign node24847 = (inp[3]) ? 4'b0011 : 4'b0010;
																assign node24850 = (inp[3]) ? 4'b0010 : 4'b0011;
													assign node24853 = (inp[3]) ? node24857 : node24854;
														assign node24854 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24857 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node24860 = (inp[5]) ? node24868 : node24861;
													assign node24861 = (inp[9]) ? node24865 : node24862;
														assign node24862 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node24865 = (inp[3]) ? 4'b0010 : 4'b0011;
													assign node24868 = (inp[2]) ? node24880 : node24869;
														assign node24869 = (inp[11]) ? node24875 : node24870;
															assign node24870 = (inp[3]) ? 4'b0011 : node24871;
																assign node24871 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24875 = (inp[3]) ? node24877 : 4'b0011;
																assign node24877 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24880 = (inp[3]) ? node24884 : node24881;
															assign node24881 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24884 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node24887 = (inp[2]) ? node24905 : node24888;
												assign node24888 = (inp[10]) ? node24896 : node24889;
													assign node24889 = (inp[9]) ? node24893 : node24890;
														assign node24890 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24893 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node24896 = (inp[3]) ? 4'b0010 : node24897;
														assign node24897 = (inp[5]) ? node24901 : node24898;
															assign node24898 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node24901 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node24905 = (inp[3]) ? node24923 : node24906;
													assign node24906 = (inp[11]) ? node24916 : node24907;
														assign node24907 = (inp[10]) ? 4'b0011 : node24908;
															assign node24908 = (inp[9]) ? node24912 : node24909;
																assign node24909 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node24912 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node24916 = (inp[5]) ? node24920 : node24917;
															assign node24917 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node24920 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node24923 = (inp[5]) ? 4'b0011 : node24924;
														assign node24924 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node24928 = (inp[10]) ? node25000 : node24929;
										assign node24929 = (inp[5]) ? node24963 : node24930;
											assign node24930 = (inp[9]) ? node24950 : node24931;
												assign node24931 = (inp[3]) ? node24937 : node24932;
													assign node24932 = (inp[1]) ? node24934 : 4'b0110;
														assign node24934 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node24937 = (inp[11]) ? node24945 : node24938;
														assign node24938 = (inp[2]) ? node24940 : 4'b0111;
															assign node24940 = (inp[0]) ? node24942 : 4'b0110;
																assign node24942 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node24945 = (inp[1]) ? 4'b0111 : node24946;
															assign node24946 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node24950 = (inp[0]) ? node24956 : node24951;
													assign node24951 = (inp[1]) ? node24953 : 4'b0111;
														assign node24953 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node24956 = (inp[3]) ? node24960 : node24957;
														assign node24957 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node24960 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node24963 = (inp[9]) ? node24985 : node24964;
												assign node24964 = (inp[3]) ? node24970 : node24965;
													assign node24965 = (inp[0]) ? node24967 : 4'b0111;
														assign node24967 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node24970 = (inp[2]) ? node24978 : node24971;
														assign node24971 = (inp[0]) ? node24975 : node24972;
															assign node24972 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node24975 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node24978 = (inp[1]) ? node24982 : node24979;
															assign node24979 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node24982 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node24985 = (inp[1]) ? node24991 : node24986;
													assign node24986 = (inp[3]) ? node24988 : 4'b0110;
														assign node24988 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node24991 = (inp[2]) ? node24995 : node24992;
														assign node24992 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node24995 = (inp[0]) ? 4'b0111 : node24996;
															assign node24996 = (inp[3]) ? 4'b0111 : 4'b0110;
										assign node25000 = (inp[9]) ? node25038 : node25001;
											assign node25001 = (inp[1]) ? node25013 : node25002;
												assign node25002 = (inp[5]) ? node25008 : node25003;
													assign node25003 = (inp[0]) ? node25005 : 4'b0110;
														assign node25005 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node25008 = (inp[0]) ? node25010 : 4'b0111;
														assign node25010 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node25013 = (inp[5]) ? node25027 : node25014;
													assign node25014 = (inp[11]) ? node25022 : node25015;
														assign node25015 = (inp[0]) ? node25019 : node25016;
															assign node25016 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node25019 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node25022 = (inp[2]) ? 4'b0110 : node25023;
															assign node25023 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node25027 = (inp[2]) ? node25029 : 4'b0110;
														assign node25029 = (inp[11]) ? node25031 : 4'b0110;
															assign node25031 = (inp[3]) ? node25035 : node25032;
																assign node25032 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node25035 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node25038 = (inp[5]) ? node25064 : node25039;
												assign node25039 = (inp[1]) ? node25045 : node25040;
													assign node25040 = (inp[3]) ? node25042 : 4'b0111;
														assign node25042 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node25045 = (inp[2]) ? node25057 : node25046;
														assign node25046 = (inp[11]) ? node25052 : node25047;
															assign node25047 = (inp[0]) ? node25049 : 4'b0111;
																assign node25049 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node25052 = (inp[3]) ? node25054 : 4'b0111;
																assign node25054 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25057 = (inp[3]) ? node25061 : node25058;
															assign node25058 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node25061 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node25064 = (inp[1]) ? node25070 : node25065;
													assign node25065 = (inp[0]) ? node25067 : 4'b0110;
														assign node25067 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node25070 = (inp[0]) ? 4'b0111 : node25071;
														assign node25071 = (inp[3]) ? 4'b0111 : 4'b0110;
								assign node25075 = (inp[15]) ? node25181 : node25076;
									assign node25076 = (inp[1]) ? node25084 : node25077;
										assign node25077 = (inp[5]) ? node25081 : node25078;
											assign node25078 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node25081 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node25084 = (inp[10]) ? node25116 : node25085;
											assign node25085 = (inp[0]) ? node25109 : node25086;
												assign node25086 = (inp[9]) ? node25098 : node25087;
													assign node25087 = (inp[11]) ? node25093 : node25088;
														assign node25088 = (inp[5]) ? node25090 : 4'b0110;
															assign node25090 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node25093 = (inp[3]) ? node25095 : 4'b0110;
															assign node25095 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node25098 = (inp[2]) ? 4'b0111 : node25099;
														assign node25099 = (inp[11]) ? 4'b0111 : node25100;
															assign node25100 = (inp[3]) ? node25104 : node25101;
																assign node25101 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node25104 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node25109 = (inp[9]) ? node25113 : node25110;
													assign node25110 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node25113 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node25116 = (inp[11]) ? node25142 : node25117;
												assign node25117 = (inp[9]) ? node25131 : node25118;
													assign node25118 = (inp[5]) ? node25126 : node25119;
														assign node25119 = (inp[2]) ? 4'b0110 : node25120;
															assign node25120 = (inp[0]) ? 4'b0110 : node25121;
																assign node25121 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node25126 = (inp[3]) ? node25128 : 4'b0111;
															assign node25128 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25131 = (inp[5]) ? node25137 : node25132;
														assign node25132 = (inp[0]) ? 4'b0111 : node25133;
															assign node25133 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node25137 = (inp[0]) ? 4'b0110 : node25138;
															assign node25138 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node25142 = (inp[0]) ? node25160 : node25143;
													assign node25143 = (inp[3]) ? node25149 : node25144;
														assign node25144 = (inp[5]) ? 4'b0111 : node25145;
															assign node25145 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25149 = (inp[2]) ? node25155 : node25150;
															assign node25150 = (inp[5]) ? node25152 : 4'b0111;
																assign node25152 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25155 = (inp[5]) ? 4'b0110 : node25156;
																assign node25156 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25160 = (inp[3]) ? node25168 : node25161;
														assign node25161 = (inp[9]) ? node25165 : node25162;
															assign node25162 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25165 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25168 = (inp[2]) ? node25176 : node25169;
															assign node25169 = (inp[5]) ? node25173 : node25170;
																assign node25170 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node25173 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node25176 = (inp[5]) ? node25178 : 4'b0110;
																assign node25178 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node25181 = (inp[10]) ? node25299 : node25182;
										assign node25182 = (inp[11]) ? node25236 : node25183;
											assign node25183 = (inp[0]) ? node25215 : node25184;
												assign node25184 = (inp[2]) ? node25196 : node25185;
													assign node25185 = (inp[1]) ? node25187 : 4'b0010;
														assign node25187 = (inp[9]) ? node25189 : 4'b0010;
															assign node25189 = (inp[5]) ? node25193 : node25190;
																assign node25190 = (inp[3]) ? 4'b0010 : 4'b0011;
																assign node25193 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node25196 = (inp[9]) ? node25202 : node25197;
														assign node25197 = (inp[1]) ? 4'b0011 : node25198;
															assign node25198 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node25202 = (inp[3]) ? node25210 : node25203;
															assign node25203 = (inp[5]) ? node25207 : node25204;
																assign node25204 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node25207 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node25210 = (inp[1]) ? 4'b0010 : node25211;
																assign node25211 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25215 = (inp[2]) ? node25225 : node25216;
													assign node25216 = (inp[3]) ? node25222 : node25217;
														assign node25217 = (inp[9]) ? node25219 : 4'b0011;
															assign node25219 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node25222 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25225 = (inp[3]) ? node25229 : node25226;
														assign node25226 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25229 = (inp[1]) ? node25231 : 4'b0011;
															assign node25231 = (inp[5]) ? 4'b0010 : node25232;
																assign node25232 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node25236 = (inp[2]) ? node25272 : node25237;
												assign node25237 = (inp[1]) ? node25257 : node25238;
													assign node25238 = (inp[5]) ? node25252 : node25239;
														assign node25239 = (inp[9]) ? node25245 : node25240;
															assign node25240 = (inp[0]) ? node25242 : 4'b0010;
																assign node25242 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node25245 = (inp[3]) ? node25249 : node25246;
																assign node25246 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node25249 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25252 = (inp[9]) ? 4'b0010 : node25253;
															assign node25253 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node25257 = (inp[3]) ? node25261 : node25258;
														assign node25258 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25261 = (inp[5]) ? node25267 : node25262;
															assign node25262 = (inp[0]) ? 4'b0011 : node25263;
																assign node25263 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node25267 = (inp[9]) ? node25269 : 4'b0010;
																assign node25269 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node25272 = (inp[0]) ? node25292 : node25273;
													assign node25273 = (inp[9]) ? node25285 : node25274;
														assign node25274 = (inp[1]) ? node25280 : node25275;
															assign node25275 = (inp[5]) ? node25277 : 4'b0011;
																assign node25277 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node25280 = (inp[3]) ? 4'b0010 : node25281;
																assign node25281 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25285 = (inp[3]) ? 4'b0010 : node25286;
															assign node25286 = (inp[1]) ? 4'b0010 : node25287;
																assign node25287 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25292 = (inp[1]) ? node25294 : 4'b0010;
														assign node25294 = (inp[9]) ? node25296 : 4'b0010;
															assign node25296 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node25299 = (inp[11]) ? node25357 : node25300;
											assign node25300 = (inp[1]) ? node25328 : node25301;
												assign node25301 = (inp[0]) ? node25319 : node25302;
													assign node25302 = (inp[9]) ? node25312 : node25303;
														assign node25303 = (inp[2]) ? node25309 : node25304;
															assign node25304 = (inp[5]) ? 4'b0010 : node25305;
																assign node25305 = (inp[3]) ? 4'b0010 : 4'b0011;
															assign node25309 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node25312 = (inp[5]) ? node25316 : node25313;
															assign node25313 = (inp[3]) ? 4'b0011 : 4'b0010;
															assign node25316 = (inp[3]) ? 4'b0010 : 4'b0011;
													assign node25319 = (inp[2]) ? node25323 : node25320;
														assign node25320 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node25323 = (inp[3]) ? 4'b0010 : node25324;
															assign node25324 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node25328 = (inp[0]) ? node25342 : node25329;
													assign node25329 = (inp[5]) ? node25337 : node25330;
														assign node25330 = (inp[2]) ? node25332 : 4'b0010;
															assign node25332 = (inp[3]) ? 4'b0010 : node25333;
																assign node25333 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node25337 = (inp[9]) ? node25339 : 4'b0011;
															assign node25339 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node25342 = (inp[3]) ? node25350 : node25343;
														assign node25343 = (inp[9]) ? node25347 : node25344;
															assign node25344 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25347 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node25350 = (inp[5]) ? node25354 : node25351;
															assign node25351 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node25354 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node25357 = (inp[1]) ? node25399 : node25358;
												assign node25358 = (inp[3]) ? node25376 : node25359;
													assign node25359 = (inp[2]) ? node25367 : node25360;
														assign node25360 = (inp[9]) ? node25362 : 4'b0011;
															assign node25362 = (inp[5]) ? node25364 : 4'b0010;
																assign node25364 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25367 = (inp[9]) ? 4'b0011 : node25368;
															assign node25368 = (inp[5]) ? node25372 : node25369;
																assign node25369 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node25372 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25376 = (inp[0]) ? node25392 : node25377;
														assign node25377 = (inp[2]) ? node25385 : node25378;
															assign node25378 = (inp[9]) ? node25382 : node25379;
																assign node25379 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node25382 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node25385 = (inp[5]) ? node25389 : node25386;
																assign node25386 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node25389 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node25392 = (inp[9]) ? node25396 : node25393;
															assign node25393 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node25396 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node25399 = (inp[3]) ? node25407 : node25400;
													assign node25400 = (inp[5]) ? node25404 : node25401;
														assign node25401 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node25404 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node25407 = (inp[9]) ? node25415 : node25408;
														assign node25408 = (inp[5]) ? node25412 : node25409;
															assign node25409 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node25412 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node25415 = (inp[2]) ? node25419 : node25416;
															assign node25416 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25419 = (inp[0]) ? node25421 : 4'b0011;
																assign node25421 = (inp[5]) ? 4'b0010 : 4'b0011;
							assign node25424 = (inp[10]) ? node25730 : node25425;
								assign node25425 = (inp[13]) ? node25609 : node25426;
									assign node25426 = (inp[15]) ? node25512 : node25427;
										assign node25427 = (inp[1]) ? node25451 : node25428;
											assign node25428 = (inp[9]) ? node25440 : node25429;
												assign node25429 = (inp[5]) ? node25435 : node25430;
													assign node25430 = (inp[3]) ? 4'b0010 : node25431;
														assign node25431 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25435 = (inp[3]) ? 4'b0011 : node25436;
														assign node25436 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node25440 = (inp[5]) ? node25446 : node25441;
													assign node25441 = (inp[0]) ? node25443 : 4'b0011;
														assign node25443 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node25446 = (inp[0]) ? node25448 : 4'b0010;
														assign node25448 = (inp[3]) ? 4'b0010 : 4'b0011;
											assign node25451 = (inp[9]) ? node25483 : node25452;
												assign node25452 = (inp[11]) ? node25470 : node25453;
													assign node25453 = (inp[2]) ? node25463 : node25454;
														assign node25454 = (inp[3]) ? node25456 : 4'b0011;
															assign node25456 = (inp[5]) ? node25460 : node25457;
																assign node25457 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node25460 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25463 = (inp[3]) ? node25465 : 4'b0010;
															assign node25465 = (inp[0]) ? 4'b0010 : node25466;
																assign node25466 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25470 = (inp[2]) ? node25472 : 4'b0010;
														assign node25472 = (inp[3]) ? node25478 : node25473;
															assign node25473 = (inp[5]) ? 4'b0010 : node25474;
																assign node25474 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node25478 = (inp[0]) ? node25480 : 4'b0011;
																assign node25480 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25483 = (inp[11]) ? node25503 : node25484;
													assign node25484 = (inp[0]) ? node25492 : node25485;
														assign node25485 = (inp[3]) ? node25489 : node25486;
															assign node25486 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25489 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node25492 = (inp[2]) ? node25498 : node25493;
															assign node25493 = (inp[3]) ? 4'b0011 : node25494;
																assign node25494 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node25498 = (inp[5]) ? node25500 : 4'b0010;
																assign node25500 = (inp[3]) ? 4'b0011 : 4'b0010;
													assign node25503 = (inp[2]) ? 4'b0011 : node25504;
														assign node25504 = (inp[3]) ? node25508 : node25505;
															assign node25505 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25508 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node25512 = (inp[1]) ? node25576 : node25513;
											assign node25513 = (inp[0]) ? node25539 : node25514;
												assign node25514 = (inp[3]) ? node25532 : node25515;
													assign node25515 = (inp[2]) ? node25521 : node25516;
														assign node25516 = (inp[5]) ? node25518 : 4'b0110;
															assign node25518 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node25521 = (inp[11]) ? node25527 : node25522;
															assign node25522 = (inp[9]) ? node25524 : 4'b0110;
																assign node25524 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25527 = (inp[9]) ? 4'b0110 : node25528;
																assign node25528 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node25532 = (inp[5]) ? node25536 : node25533;
														assign node25533 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25536 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node25539 = (inp[2]) ? node25557 : node25540;
													assign node25540 = (inp[9]) ? node25548 : node25541;
														assign node25541 = (inp[3]) ? node25545 : node25542;
															assign node25542 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25545 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node25548 = (inp[11]) ? node25554 : node25549;
															assign node25549 = (inp[3]) ? 4'b0111 : node25550;
																assign node25550 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25554 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node25557 = (inp[3]) ? node25565 : node25558;
														assign node25558 = (inp[9]) ? node25562 : node25559;
															assign node25559 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25562 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node25565 = (inp[11]) ? node25571 : node25566;
															assign node25566 = (inp[5]) ? node25568 : 4'b0110;
																assign node25568 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node25571 = (inp[5]) ? 4'b0110 : node25572;
																assign node25572 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node25576 = (inp[0]) ? node25602 : node25577;
												assign node25577 = (inp[11]) ? node25593 : node25578;
													assign node25578 = (inp[2]) ? node25586 : node25579;
														assign node25579 = (inp[9]) ? node25583 : node25580;
															assign node25580 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25583 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25586 = (inp[5]) ? node25590 : node25587;
															assign node25587 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25590 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25593 = (inp[3]) ? 4'b0110 : node25594;
														assign node25594 = (inp[5]) ? node25598 : node25595;
															assign node25595 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25598 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node25602 = (inp[5]) ? node25606 : node25603;
													assign node25603 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node25606 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node25609 = (inp[15]) ? node25699 : node25610;
										assign node25610 = (inp[5]) ? node25644 : node25611;
											assign node25611 = (inp[9]) ? node25631 : node25612;
												assign node25612 = (inp[2]) ? node25622 : node25613;
													assign node25613 = (inp[0]) ? 4'b0110 : node25614;
														assign node25614 = (inp[1]) ? node25618 : node25615;
															assign node25615 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node25618 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node25622 = (inp[0]) ? 4'b0111 : node25623;
														assign node25623 = (inp[1]) ? node25627 : node25624;
															assign node25624 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node25627 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node25631 = (inp[11]) ? node25633 : 4'b0111;
													assign node25633 = (inp[3]) ? node25639 : node25634;
														assign node25634 = (inp[1]) ? 4'b0110 : node25635;
															assign node25635 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node25639 = (inp[0]) ? 4'b0111 : node25640;
															assign node25640 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node25644 = (inp[9]) ? node25676 : node25645;
												assign node25645 = (inp[3]) ? node25671 : node25646;
													assign node25646 = (inp[11]) ? node25656 : node25647;
														assign node25647 = (inp[2]) ? 4'b0110 : node25648;
															assign node25648 = (inp[1]) ? node25652 : node25649;
																assign node25649 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node25652 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25656 = (inp[2]) ? node25664 : node25657;
															assign node25657 = (inp[0]) ? node25661 : node25658;
																assign node25658 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node25661 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node25664 = (inp[0]) ? node25668 : node25665;
																assign node25665 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node25668 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node25671 = (inp[0]) ? 4'b0111 : node25672;
														assign node25672 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node25676 = (inp[0]) ? node25694 : node25677;
													assign node25677 = (inp[2]) ? node25685 : node25678;
														assign node25678 = (inp[1]) ? node25682 : node25679;
															assign node25679 = (inp[3]) ? 4'b0111 : 4'b0110;
															assign node25682 = (inp[3]) ? 4'b0110 : 4'b0111;
														assign node25685 = (inp[11]) ? 4'b0111 : node25686;
															assign node25686 = (inp[3]) ? node25690 : node25687;
																assign node25687 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node25690 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node25694 = (inp[2]) ? 4'b0110 : node25695;
														assign node25695 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node25699 = (inp[9]) ? node25715 : node25700;
											assign node25700 = (inp[5]) ? node25708 : node25701;
												assign node25701 = (inp[1]) ? node25703 : 4'b0010;
													assign node25703 = (inp[3]) ? 4'b0010 : node25704;
														assign node25704 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node25708 = (inp[1]) ? node25710 : 4'b0011;
													assign node25710 = (inp[0]) ? 4'b0011 : node25711;
														assign node25711 = (inp[3]) ? 4'b0011 : 4'b0010;
											assign node25715 = (inp[5]) ? node25723 : node25716;
												assign node25716 = (inp[1]) ? node25718 : 4'b0011;
													assign node25718 = (inp[0]) ? 4'b0011 : node25719;
														assign node25719 = (inp[3]) ? 4'b0011 : 4'b0010;
												assign node25723 = (inp[3]) ? 4'b0010 : node25724;
													assign node25724 = (inp[1]) ? node25726 : 4'b0010;
														assign node25726 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node25730 = (inp[9]) ? node25824 : node25731;
									assign node25731 = (inp[5]) ? node25775 : node25732;
										assign node25732 = (inp[15]) ? node25760 : node25733;
											assign node25733 = (inp[13]) ? node25747 : node25734;
												assign node25734 = (inp[0]) ? node25740 : node25735;
													assign node25735 = (inp[3]) ? 4'b0010 : node25736;
														assign node25736 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node25740 = (inp[1]) ? node25744 : node25741;
														assign node25741 = (inp[3]) ? 4'b0010 : 4'b0011;
														assign node25744 = (inp[3]) ? 4'b0011 : 4'b0010;
												assign node25747 = (inp[1]) ? node25755 : node25748;
													assign node25748 = (inp[0]) ? node25752 : node25749;
														assign node25749 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node25752 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node25755 = (inp[0]) ? 4'b0110 : node25756;
														assign node25756 = (inp[3]) ? 4'b0110 : 4'b0111;
											assign node25760 = (inp[13]) ? node25768 : node25761;
												assign node25761 = (inp[0]) ? node25763 : 4'b0110;
													assign node25763 = (inp[1]) ? 4'b0110 : node25764;
														assign node25764 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node25768 = (inp[1]) ? node25770 : 4'b0010;
													assign node25770 = (inp[11]) ? node25772 : 4'b0010;
														assign node25772 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node25775 = (inp[15]) ? node25809 : node25776;
											assign node25776 = (inp[13]) ? node25790 : node25777;
												assign node25777 = (inp[0]) ? node25783 : node25778;
													assign node25778 = (inp[3]) ? 4'b0011 : node25779;
														assign node25779 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node25783 = (inp[1]) ? node25787 : node25784;
														assign node25784 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node25787 = (inp[3]) ? 4'b0010 : 4'b0011;
												assign node25790 = (inp[2]) ? node25798 : node25791;
													assign node25791 = (inp[1]) ? 4'b0111 : node25792;
														assign node25792 = (inp[3]) ? node25794 : 4'b0111;
															assign node25794 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25798 = (inp[3]) ? node25804 : node25799;
														assign node25799 = (inp[0]) ? 4'b0110 : node25800;
															assign node25800 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25804 = (inp[1]) ? 4'b0111 : node25805;
															assign node25805 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node25809 = (inp[13]) ? node25817 : node25810;
												assign node25810 = (inp[0]) ? node25812 : 4'b0111;
													assign node25812 = (inp[3]) ? 4'b0111 : node25813;
														assign node25813 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node25817 = (inp[0]) ? 4'b0011 : node25818;
													assign node25818 = (inp[1]) ? node25820 : 4'b0011;
														assign node25820 = (inp[3]) ? 4'b0011 : 4'b0010;
									assign node25824 = (inp[5]) ? node25876 : node25825;
										assign node25825 = (inp[15]) ? node25861 : node25826;
											assign node25826 = (inp[13]) ? node25840 : node25827;
												assign node25827 = (inp[0]) ? node25833 : node25828;
													assign node25828 = (inp[3]) ? 4'b0011 : node25829;
														assign node25829 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25833 = (inp[1]) ? node25837 : node25834;
														assign node25834 = (inp[3]) ? 4'b0011 : 4'b0010;
														assign node25837 = (inp[3]) ? 4'b0010 : 4'b0011;
												assign node25840 = (inp[1]) ? node25856 : node25841;
													assign node25841 = (inp[2]) ? node25849 : node25842;
														assign node25842 = (inp[0]) ? node25846 : node25843;
															assign node25843 = (inp[3]) ? 4'b0110 : 4'b0111;
															assign node25846 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node25849 = (inp[3]) ? node25853 : node25850;
															assign node25850 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node25853 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25856 = (inp[3]) ? 4'b0111 : node25857;
														assign node25857 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node25861 = (inp[13]) ? node25869 : node25862;
												assign node25862 = (inp[0]) ? node25864 : 4'b0111;
													assign node25864 = (inp[1]) ? 4'b0111 : node25865;
														assign node25865 = (inp[3]) ? 4'b0111 : 4'b0110;
												assign node25869 = (inp[0]) ? 4'b0011 : node25870;
													assign node25870 = (inp[1]) ? node25872 : 4'b0011;
														assign node25872 = (inp[3]) ? 4'b0011 : 4'b0010;
										assign node25876 = (inp[3]) ? node25914 : node25877;
											assign node25877 = (inp[15]) ? node25903 : node25878;
												assign node25878 = (inp[13]) ? node25886 : node25879;
													assign node25879 = (inp[0]) ? node25883 : node25880;
														assign node25880 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node25883 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25886 = (inp[11]) ? node25898 : node25887;
														assign node25887 = (inp[2]) ? node25893 : node25888;
															assign node25888 = (inp[1]) ? 4'b0111 : node25889;
																assign node25889 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node25893 = (inp[1]) ? node25895 : 4'b0110;
																assign node25895 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node25898 = (inp[1]) ? node25900 : 4'b0111;
															assign node25900 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node25903 = (inp[13]) ? node25909 : node25904;
													assign node25904 = (inp[0]) ? node25906 : 4'b0110;
														assign node25906 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node25909 = (inp[1]) ? node25911 : 4'b0010;
														assign node25911 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node25914 = (inp[15]) ? node25926 : node25915;
												assign node25915 = (inp[13]) ? node25921 : node25916;
													assign node25916 = (inp[1]) ? node25918 : 4'b0010;
														assign node25918 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25921 = (inp[0]) ? 4'b0110 : node25922;
														assign node25922 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25926 = (inp[13]) ? 4'b0010 : 4'b0110;
					assign node25929 = (inp[4]) ? node26851 : node25930;
						assign node25930 = (inp[3]) ? node26462 : node25931;
							assign node25931 = (inp[12]) ? node26197 : node25932;
								assign node25932 = (inp[13]) ? node26080 : node25933;
									assign node25933 = (inp[1]) ? node26015 : node25934;
										assign node25934 = (inp[15]) ? node25958 : node25935;
											assign node25935 = (inp[2]) ? node25947 : node25936;
												assign node25936 = (inp[9]) ? node25942 : node25937;
													assign node25937 = (inp[0]) ? 4'b0010 : node25938;
														assign node25938 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25942 = (inp[5]) ? node25944 : 4'b0011;
														assign node25944 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node25947 = (inp[9]) ? node25953 : node25948;
													assign node25948 = (inp[5]) ? node25950 : 4'b0011;
														assign node25950 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25953 = (inp[0]) ? 4'b0010 : node25954;
														assign node25954 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node25958 = (inp[10]) ? node25982 : node25959;
												assign node25959 = (inp[2]) ? node25971 : node25960;
													assign node25960 = (inp[9]) ? node25966 : node25961;
														assign node25961 = (inp[5]) ? node25963 : 4'b0110;
															assign node25963 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node25966 = (inp[0]) ? 4'b0111 : node25967;
															assign node25967 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node25971 = (inp[9]) ? node25977 : node25972;
														assign node25972 = (inp[0]) ? 4'b0111 : node25973;
															assign node25973 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25977 = (inp[0]) ? 4'b0110 : node25978;
															assign node25978 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node25982 = (inp[5]) ? node25998 : node25983;
													assign node25983 = (inp[11]) ? node25991 : node25984;
														assign node25984 = (inp[2]) ? node25988 : node25985;
															assign node25985 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25988 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node25991 = (inp[9]) ? node25995 : node25992;
															assign node25992 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node25995 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node25998 = (inp[9]) ? node26006 : node25999;
														assign node25999 = (inp[0]) ? node26003 : node26000;
															assign node26000 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node26003 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node26006 = (inp[11]) ? node26010 : node26007;
															assign node26007 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node26010 = (inp[2]) ? node26012 : 4'b0110;
																assign node26012 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node26015 = (inp[2]) ? node26039 : node26016;
											assign node26016 = (inp[15]) ? node26028 : node26017;
												assign node26017 = (inp[9]) ? node26023 : node26018;
													assign node26018 = (inp[0]) ? 4'b0010 : node26019;
														assign node26019 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node26023 = (inp[5]) ? node26025 : 4'b0011;
														assign node26025 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node26028 = (inp[9]) ? node26034 : node26029;
													assign node26029 = (inp[0]) ? 4'b0011 : node26030;
														assign node26030 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node26034 = (inp[0]) ? 4'b0010 : node26035;
														assign node26035 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node26039 = (inp[0]) ? node26055 : node26040;
												assign node26040 = (inp[5]) ? node26048 : node26041;
													assign node26041 = (inp[9]) ? node26045 : node26042;
														assign node26042 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node26045 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node26048 = (inp[9]) ? node26052 : node26049;
														assign node26049 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node26052 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node26055 = (inp[11]) ? node26073 : node26056;
													assign node26056 = (inp[5]) ? node26066 : node26057;
														assign node26057 = (inp[10]) ? 4'b0011 : node26058;
															assign node26058 = (inp[15]) ? node26062 : node26059;
																assign node26059 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node26062 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node26066 = (inp[10]) ? node26068 : 4'b0011;
															assign node26068 = (inp[9]) ? 4'b0010 : node26069;
																assign node26069 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node26073 = (inp[15]) ? node26077 : node26074;
														assign node26074 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node26077 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node26080 = (inp[1]) ? node26150 : node26081;
										assign node26081 = (inp[15]) ? node26127 : node26082;
											assign node26082 = (inp[10]) ? node26104 : node26083;
												assign node26083 = (inp[9]) ? node26095 : node26084;
													assign node26084 = (inp[2]) ? node26090 : node26085;
														assign node26085 = (inp[0]) ? 4'b0110 : node26086;
															assign node26086 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node26090 = (inp[0]) ? 4'b0111 : node26091;
															assign node26091 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node26095 = (inp[0]) ? 4'b0111 : node26096;
														assign node26096 = (inp[11]) ? node26098 : 4'b0110;
															assign node26098 = (inp[5]) ? 4'b0111 : node26099;
																assign node26099 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node26104 = (inp[5]) ? node26112 : node26105;
													assign node26105 = (inp[9]) ? node26109 : node26106;
														assign node26106 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node26109 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node26112 = (inp[9]) ? node26120 : node26113;
														assign node26113 = (inp[11]) ? node26115 : 4'b0110;
															assign node26115 = (inp[0]) ? 4'b0111 : node26116;
																assign node26116 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node26120 = (inp[11]) ? 4'b0110 : node26121;
															assign node26121 = (inp[0]) ? node26123 : 4'b0110;
																assign node26123 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node26127 = (inp[9]) ? node26139 : node26128;
												assign node26128 = (inp[2]) ? node26134 : node26129;
													assign node26129 = (inp[0]) ? node26131 : 4'b0011;
														assign node26131 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node26134 = (inp[0]) ? node26136 : 4'b0010;
														assign node26136 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node26139 = (inp[2]) ? node26145 : node26140;
													assign node26140 = (inp[0]) ? node26142 : 4'b0010;
														assign node26142 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node26145 = (inp[0]) ? node26147 : 4'b0011;
														assign node26147 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node26150 = (inp[11]) ? node26174 : node26151;
											assign node26151 = (inp[9]) ? node26163 : node26152;
												assign node26152 = (inp[2]) ? node26158 : node26153;
													assign node26153 = (inp[0]) ? 4'b0110 : node26154;
														assign node26154 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node26158 = (inp[0]) ? 4'b0111 : node26159;
														assign node26159 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node26163 = (inp[2]) ? node26169 : node26164;
													assign node26164 = (inp[5]) ? node26166 : 4'b0111;
														assign node26166 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node26169 = (inp[5]) ? node26171 : 4'b0110;
														assign node26171 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node26174 = (inp[9]) ? node26186 : node26175;
												assign node26175 = (inp[2]) ? node26181 : node26176;
													assign node26176 = (inp[5]) ? node26178 : 4'b0110;
														assign node26178 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node26181 = (inp[5]) ? node26183 : 4'b0111;
														assign node26183 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node26186 = (inp[2]) ? node26192 : node26187;
													assign node26187 = (inp[5]) ? node26189 : 4'b0111;
														assign node26189 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node26192 = (inp[5]) ? node26194 : 4'b0110;
														assign node26194 = (inp[0]) ? 4'b0110 : 4'b0111;
								assign node26197 = (inp[13]) ? node26323 : node26198;
									assign node26198 = (inp[15]) ? node26246 : node26199;
										assign node26199 = (inp[2]) ? node26223 : node26200;
											assign node26200 = (inp[1]) ? node26212 : node26201;
												assign node26201 = (inp[9]) ? node26207 : node26202;
													assign node26202 = (inp[5]) ? 4'b0110 : node26203;
														assign node26203 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node26207 = (inp[5]) ? 4'b0111 : node26208;
														assign node26208 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node26212 = (inp[9]) ? node26218 : node26213;
													assign node26213 = (inp[0]) ? node26215 : 4'b0111;
														assign node26215 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node26218 = (inp[5]) ? 4'b0110 : node26219;
														assign node26219 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node26223 = (inp[9]) ? node26235 : node26224;
												assign node26224 = (inp[1]) ? node26230 : node26225;
													assign node26225 = (inp[0]) ? node26227 : 4'b0111;
														assign node26227 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node26230 = (inp[5]) ? 4'b0110 : node26231;
														assign node26231 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node26235 = (inp[1]) ? node26241 : node26236;
													assign node26236 = (inp[0]) ? node26238 : 4'b0110;
														assign node26238 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node26241 = (inp[5]) ? 4'b0111 : node26242;
														assign node26242 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node26246 = (inp[1]) ? node26270 : node26247;
											assign node26247 = (inp[9]) ? node26259 : node26248;
												assign node26248 = (inp[2]) ? node26254 : node26249;
													assign node26249 = (inp[5]) ? node26251 : 4'b0011;
														assign node26251 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node26254 = (inp[0]) ? 4'b0010 : node26255;
														assign node26255 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node26259 = (inp[2]) ? node26265 : node26260;
													assign node26260 = (inp[5]) ? node26262 : 4'b0010;
														assign node26262 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node26265 = (inp[0]) ? 4'b0011 : node26266;
														assign node26266 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node26270 = (inp[10]) ? node26292 : node26271;
												assign node26271 = (inp[5]) ? node26285 : node26272;
													assign node26272 = (inp[0]) ? node26280 : node26273;
														assign node26273 = (inp[9]) ? node26277 : node26274;
															assign node26274 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node26277 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node26280 = (inp[9]) ? node26282 : 4'b0110;
															assign node26282 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node26285 = (inp[2]) ? node26289 : node26286;
														assign node26286 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node26289 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node26292 = (inp[11]) ? node26316 : node26293;
													assign node26293 = (inp[5]) ? node26309 : node26294;
														assign node26294 = (inp[9]) ? node26302 : node26295;
															assign node26295 = (inp[0]) ? node26299 : node26296;
																assign node26296 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node26299 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node26302 = (inp[2]) ? node26306 : node26303;
																assign node26303 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node26306 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node26309 = (inp[2]) ? node26313 : node26310;
															assign node26310 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node26313 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node26316 = (inp[2]) ? node26318 : 4'b0110;
														assign node26318 = (inp[9]) ? node26320 : 4'b0111;
															assign node26320 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node26323 = (inp[1]) ? node26379 : node26324;
										assign node26324 = (inp[15]) ? node26348 : node26325;
											assign node26325 = (inp[9]) ? node26337 : node26326;
												assign node26326 = (inp[2]) ? node26332 : node26327;
													assign node26327 = (inp[5]) ? node26329 : 4'b0011;
														assign node26329 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node26332 = (inp[5]) ? node26334 : 4'b0010;
														assign node26334 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node26337 = (inp[2]) ? node26343 : node26338;
													assign node26338 = (inp[5]) ? node26340 : 4'b0010;
														assign node26340 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node26343 = (inp[0]) ? 4'b0011 : node26344;
														assign node26344 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node26348 = (inp[10]) ? node26366 : node26349;
												assign node26349 = (inp[0]) ? node26359 : node26350;
													assign node26350 = (inp[5]) ? 4'b0110 : node26351;
														assign node26351 = (inp[9]) ? node26355 : node26352;
															assign node26352 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node26355 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node26359 = (inp[9]) ? node26363 : node26360;
														assign node26360 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node26363 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node26366 = (inp[9]) ? node26372 : node26367;
													assign node26367 = (inp[2]) ? 4'b0111 : node26368;
														assign node26368 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node26372 = (inp[0]) ? node26376 : node26373;
														assign node26373 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node26376 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node26379 = (inp[10]) ? node26403 : node26380;
											assign node26380 = (inp[5]) ? node26388 : node26381;
												assign node26381 = (inp[2]) ? node26385 : node26382;
													assign node26382 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node26385 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node26388 = (inp[2]) ? node26396 : node26389;
													assign node26389 = (inp[9]) ? node26393 : node26390;
														assign node26390 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node26393 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node26396 = (inp[0]) ? node26400 : node26397;
														assign node26397 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node26400 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node26403 = (inp[11]) ? node26445 : node26404;
												assign node26404 = (inp[5]) ? node26422 : node26405;
													assign node26405 = (inp[15]) ? node26415 : node26406;
														assign node26406 = (inp[0]) ? node26408 : 4'b0011;
															assign node26408 = (inp[9]) ? node26412 : node26409;
																assign node26409 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node26412 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node26415 = (inp[2]) ? node26419 : node26416;
															assign node26416 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node26419 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node26422 = (inp[0]) ? node26430 : node26423;
														assign node26423 = (inp[2]) ? node26427 : node26424;
															assign node26424 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node26427 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node26430 = (inp[15]) ? node26438 : node26431;
															assign node26431 = (inp[2]) ? node26435 : node26432;
																assign node26432 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node26435 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node26438 = (inp[2]) ? node26442 : node26439;
																assign node26439 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node26442 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node26445 = (inp[2]) ? node26451 : node26446;
													assign node26446 = (inp[9]) ? node26448 : 4'b0010;
														assign node26448 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node26451 = (inp[9]) ? node26457 : node26452;
														assign node26452 = (inp[0]) ? 4'b0011 : node26453;
															assign node26453 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node26457 = (inp[0]) ? 4'b0010 : node26458;
															assign node26458 = (inp[5]) ? 4'b0011 : 4'b0010;
							assign node26462 = (inp[9]) ? node26660 : node26463;
								assign node26463 = (inp[2]) ? node26551 : node26464;
									assign node26464 = (inp[0]) ? node26518 : node26465;
										assign node26465 = (inp[5]) ? node26493 : node26466;
											assign node26466 = (inp[12]) ? node26482 : node26467;
												assign node26467 = (inp[13]) ? node26475 : node26468;
													assign node26468 = (inp[15]) ? node26472 : node26469;
														assign node26469 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node26472 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node26475 = (inp[15]) ? node26479 : node26476;
														assign node26476 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node26479 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node26482 = (inp[13]) ? node26488 : node26483;
													assign node26483 = (inp[15]) ? 4'b0101 : node26484;
														assign node26484 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node26488 = (inp[15]) ? 4'b0001 : node26489;
														assign node26489 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node26493 = (inp[13]) ? node26507 : node26494;
												assign node26494 = (inp[12]) ? node26502 : node26495;
													assign node26495 = (inp[1]) ? node26499 : node26496;
														assign node26496 = (inp[15]) ? 4'b0000 : 4'b0101;
														assign node26499 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node26502 = (inp[1]) ? 4'b0101 : node26503;
														assign node26503 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node26507 = (inp[12]) ? node26513 : node26508;
													assign node26508 = (inp[1]) ? 4'b0100 : node26509;
														assign node26509 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node26513 = (inp[15]) ? 4'b0000 : node26514;
														assign node26514 = (inp[1]) ? 4'b0000 : 4'b0101;
										assign node26518 = (inp[13]) ? node26538 : node26519;
											assign node26519 = (inp[12]) ? node26533 : node26520;
												assign node26520 = (inp[1]) ? node26526 : node26521;
													assign node26521 = (inp[15]) ? node26523 : 4'b0101;
														assign node26523 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node26526 = (inp[15]) ? node26530 : node26527;
														assign node26527 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node26530 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node26533 = (inp[15]) ? 4'b0100 : node26534;
													assign node26534 = (inp[1]) ? 4'b0101 : 4'b0000;
											assign node26538 = (inp[12]) ? node26544 : node26539;
												assign node26539 = (inp[1]) ? 4'b0100 : node26540;
													assign node26540 = (inp[15]) ? 4'b0101 : 4'b0000;
												assign node26544 = (inp[1]) ? 4'b0000 : node26545;
													assign node26545 = (inp[15]) ? 4'b0000 : node26546;
														assign node26546 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node26551 = (inp[5]) ? node26605 : node26552;
										assign node26552 = (inp[0]) ? node26578 : node26553;
											assign node26553 = (inp[12]) ? node26567 : node26554;
												assign node26554 = (inp[1]) ? node26562 : node26555;
													assign node26555 = (inp[13]) ? node26559 : node26556;
														assign node26556 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node26559 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node26562 = (inp[13]) ? 4'b0100 : node26563;
														assign node26563 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node26567 = (inp[13]) ? node26573 : node26568;
													assign node26568 = (inp[15]) ? 4'b0100 : node26569;
														assign node26569 = (inp[1]) ? 4'b0101 : 4'b0000;
													assign node26573 = (inp[1]) ? 4'b0000 : node26574;
														assign node26574 = (inp[15]) ? 4'b0000 : 4'b0100;
											assign node26578 = (inp[1]) ? node26594 : node26579;
												assign node26579 = (inp[15]) ? node26587 : node26580;
													assign node26580 = (inp[13]) ? node26584 : node26581;
														assign node26581 = (inp[12]) ? 4'b0001 : 4'b0100;
														assign node26584 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node26587 = (inp[12]) ? node26591 : node26588;
														assign node26588 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node26591 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node26594 = (inp[13]) ? node26602 : node26595;
													assign node26595 = (inp[12]) ? node26599 : node26596;
														assign node26596 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node26599 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node26602 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node26605 = (inp[13]) ? node26641 : node26606;
											assign node26606 = (inp[12]) ? node26636 : node26607;
												assign node26607 = (inp[1]) ? node26613 : node26608;
													assign node26608 = (inp[15]) ? node26610 : 4'b0100;
														assign node26610 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node26613 = (inp[11]) ? node26623 : node26614;
														assign node26614 = (inp[10]) ? 4'b0001 : node26615;
															assign node26615 = (inp[0]) ? node26619 : node26616;
																assign node26616 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node26619 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node26623 = (inp[10]) ? node26631 : node26624;
															assign node26624 = (inp[0]) ? node26628 : node26625;
																assign node26625 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node26628 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node26631 = (inp[0]) ? 4'b0000 : node26632;
																assign node26632 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node26636 = (inp[15]) ? 4'b0101 : node26637;
													assign node26637 = (inp[1]) ? 4'b0100 : 4'b0001;
											assign node26641 = (inp[1]) ? node26657 : node26642;
												assign node26642 = (inp[0]) ? node26650 : node26643;
													assign node26643 = (inp[12]) ? node26647 : node26644;
														assign node26644 = (inp[15]) ? 4'b0100 : 4'b0001;
														assign node26647 = (inp[15]) ? 4'b0001 : 4'b0100;
													assign node26650 = (inp[15]) ? node26654 : node26651;
														assign node26651 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node26654 = (inp[12]) ? 4'b0001 : 4'b0100;
												assign node26657 = (inp[12]) ? 4'b0001 : 4'b0101;
								assign node26660 = (inp[2]) ? node26756 : node26661;
									assign node26661 = (inp[0]) ? node26723 : node26662;
										assign node26662 = (inp[5]) ? node26692 : node26663;
											assign node26663 = (inp[13]) ? node26679 : node26664;
												assign node26664 = (inp[12]) ? node26672 : node26665;
													assign node26665 = (inp[15]) ? node26669 : node26666;
														assign node26666 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node26669 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node26672 = (inp[1]) ? node26676 : node26673;
														assign node26673 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node26676 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node26679 = (inp[12]) ? node26687 : node26680;
													assign node26680 = (inp[15]) ? node26684 : node26681;
														assign node26681 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node26684 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node26687 = (inp[15]) ? 4'b0000 : node26688;
														assign node26688 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node26692 = (inp[12]) ? node26712 : node26693;
												assign node26693 = (inp[15]) ? node26705 : node26694;
													assign node26694 = (inp[11]) ? node26700 : node26695;
														assign node26695 = (inp[1]) ? 4'b0001 : node26696;
															assign node26696 = (inp[13]) ? 4'b0001 : 4'b0100;
														assign node26700 = (inp[13]) ? node26702 : 4'b0001;
															assign node26702 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node26705 = (inp[13]) ? node26709 : node26706;
														assign node26706 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node26709 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node26712 = (inp[15]) ? node26720 : node26713;
													assign node26713 = (inp[13]) ? node26717 : node26714;
														assign node26714 = (inp[1]) ? 4'b0100 : 4'b0001;
														assign node26717 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node26720 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node26723 = (inp[12]) ? node26743 : node26724;
											assign node26724 = (inp[13]) ? node26738 : node26725;
												assign node26725 = (inp[15]) ? node26731 : node26726;
													assign node26726 = (inp[1]) ? node26728 : 4'b0100;
														assign node26728 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node26731 = (inp[5]) ? node26735 : node26732;
														assign node26732 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node26735 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node26738 = (inp[1]) ? 4'b0101 : node26739;
													assign node26739 = (inp[15]) ? 4'b0100 : 4'b0001;
											assign node26743 = (inp[15]) ? node26753 : node26744;
												assign node26744 = (inp[1]) ? node26750 : node26745;
													assign node26745 = (inp[13]) ? node26747 : 4'b0001;
														assign node26747 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node26750 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node26753 = (inp[13]) ? 4'b0001 : 4'b0101;
									assign node26756 = (inp[0]) ? node26812 : node26757;
										assign node26757 = (inp[5]) ? node26785 : node26758;
											assign node26758 = (inp[12]) ? node26774 : node26759;
												assign node26759 = (inp[13]) ? node26767 : node26760;
													assign node26760 = (inp[15]) ? node26764 : node26761;
														assign node26761 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node26764 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node26767 = (inp[15]) ? node26771 : node26768;
														assign node26768 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node26771 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node26774 = (inp[13]) ? node26780 : node26775;
													assign node26775 = (inp[15]) ? 4'b0101 : node26776;
														assign node26776 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node26780 = (inp[15]) ? 4'b0001 : node26781;
														assign node26781 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node26785 = (inp[13]) ? node26799 : node26786;
												assign node26786 = (inp[12]) ? node26794 : node26787;
													assign node26787 = (inp[1]) ? node26791 : node26788;
														assign node26788 = (inp[15]) ? 4'b0000 : 4'b0101;
														assign node26791 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node26794 = (inp[1]) ? 4'b0101 : node26795;
														assign node26795 = (inp[15]) ? 4'b0100 : 4'b0000;
												assign node26799 = (inp[12]) ? node26807 : node26800;
													assign node26800 = (inp[15]) ? node26804 : node26801;
														assign node26801 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node26804 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node26807 = (inp[15]) ? 4'b0000 : node26808;
														assign node26808 = (inp[1]) ? 4'b0000 : 4'b0101;
										assign node26812 = (inp[13]) ? node26838 : node26813;
											assign node26813 = (inp[12]) ? node26833 : node26814;
												assign node26814 = (inp[15]) ? node26820 : node26815;
													assign node26815 = (inp[1]) ? node26817 : 4'b0101;
														assign node26817 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node26820 = (inp[10]) ? node26826 : node26821;
														assign node26821 = (inp[5]) ? 4'b0000 : node26822;
															assign node26822 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node26826 = (inp[5]) ? node26830 : node26827;
															assign node26827 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node26830 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node26833 = (inp[15]) ? 4'b0100 : node26834;
													assign node26834 = (inp[1]) ? 4'b0101 : 4'b0000;
											assign node26838 = (inp[12]) ? node26844 : node26839;
												assign node26839 = (inp[1]) ? 4'b0100 : node26840;
													assign node26840 = (inp[15]) ? 4'b0101 : 4'b0000;
												assign node26844 = (inp[15]) ? 4'b0000 : node26845;
													assign node26845 = (inp[1]) ? 4'b0000 : node26846;
														assign node26846 = (inp[5]) ? 4'b0100 : 4'b0101;
						assign node26851 = (inp[13]) ? node27235 : node26852;
							assign node26852 = (inp[1]) ? node27056 : node26853;
								assign node26853 = (inp[3]) ? node26945 : node26854;
									assign node26854 = (inp[15]) ? node26878 : node26855;
										assign node26855 = (inp[2]) ? node26871 : node26856;
											assign node26856 = (inp[11]) ? node26864 : node26857;
												assign node26857 = (inp[12]) ? node26861 : node26858;
													assign node26858 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node26861 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node26864 = (inp[9]) ? node26868 : node26865;
													assign node26865 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node26868 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node26871 = (inp[9]) ? node26875 : node26872;
												assign node26872 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node26875 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node26878 = (inp[9]) ? node26930 : node26879;
											assign node26879 = (inp[2]) ? node26893 : node26880;
												assign node26880 = (inp[10]) ? node26886 : node26881;
													assign node26881 = (inp[0]) ? node26883 : 4'b0000;
														assign node26883 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node26886 = (inp[12]) ? node26890 : node26887;
														assign node26887 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node26890 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node26893 = (inp[5]) ? node26909 : node26894;
													assign node26894 = (inp[10]) ? node26902 : node26895;
														assign node26895 = (inp[11]) ? node26897 : 4'b0000;
															assign node26897 = (inp[0]) ? 4'b0001 : node26898;
																assign node26898 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node26902 = (inp[11]) ? 4'b0001 : node26903;
															assign node26903 = (inp[12]) ? node26905 : 4'b0001;
																assign node26905 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node26909 = (inp[10]) ? node26921 : node26910;
														assign node26910 = (inp[11]) ? node26916 : node26911;
															assign node26911 = (inp[0]) ? node26913 : 4'b0001;
																assign node26913 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node26916 = (inp[12]) ? 4'b0001 : node26917;
																assign node26917 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node26921 = (inp[11]) ? 4'b0000 : node26922;
															assign node26922 = (inp[12]) ? node26926 : node26923;
																assign node26923 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node26926 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node26930 = (inp[11]) ? node26938 : node26931;
												assign node26931 = (inp[0]) ? node26935 : node26932;
													assign node26932 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node26935 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node26938 = (inp[0]) ? node26942 : node26939;
													assign node26939 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node26942 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node26945 = (inp[5]) ? node26991 : node26946;
										assign node26946 = (inp[10]) ? node26970 : node26947;
											assign node26947 = (inp[9]) ? node26959 : node26948;
												assign node26948 = (inp[12]) ? node26954 : node26949;
													assign node26949 = (inp[0]) ? node26951 : 4'b0100;
														assign node26951 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node26954 = (inp[15]) ? 4'b0101 : node26955;
														assign node26955 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node26959 = (inp[12]) ? node26965 : node26960;
													assign node26960 = (inp[15]) ? 4'b0101 : node26961;
														assign node26961 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node26965 = (inp[15]) ? 4'b0100 : node26966;
														assign node26966 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node26970 = (inp[0]) ? node26978 : node26971;
												assign node26971 = (inp[9]) ? node26975 : node26972;
													assign node26972 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node26975 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node26978 = (inp[9]) ? node26984 : node26979;
													assign node26979 = (inp[12]) ? node26981 : 4'b0101;
														assign node26981 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node26984 = (inp[15]) ? node26988 : node26985;
														assign node26985 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node26988 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node26991 = (inp[0]) ? node26999 : node26992;
											assign node26992 = (inp[12]) ? node26996 : node26993;
												assign node26993 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node26996 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node26999 = (inp[11]) ? node27021 : node27000;
												assign node27000 = (inp[9]) ? node27006 : node27001;
													assign node27001 = (inp[15]) ? 4'b0101 : node27002;
														assign node27002 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node27006 = (inp[2]) ? node27016 : node27007;
														assign node27007 = (inp[10]) ? node27011 : node27008;
															assign node27008 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node27011 = (inp[12]) ? node27013 : 4'b0101;
																assign node27013 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node27016 = (inp[10]) ? node27018 : 4'b0100;
															assign node27018 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node27021 = (inp[12]) ? node27035 : node27022;
													assign node27022 = (inp[2]) ? node27028 : node27023;
														assign node27023 = (inp[9]) ? node27025 : 4'b0100;
															assign node27025 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27028 = (inp[9]) ? node27032 : node27029;
															assign node27029 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node27032 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node27035 = (inp[2]) ? node27043 : node27036;
														assign node27036 = (inp[15]) ? node27040 : node27037;
															assign node27037 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node27040 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node27043 = (inp[10]) ? node27049 : node27044;
															assign node27044 = (inp[9]) ? node27046 : 4'b0100;
																assign node27046 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node27049 = (inp[9]) ? node27053 : node27050;
																assign node27050 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node27053 = (inp[15]) ? 4'b0100 : 4'b0101;
								assign node27056 = (inp[12]) ? node27170 : node27057;
									assign node27057 = (inp[11]) ? node27111 : node27058;
										assign node27058 = (inp[2]) ? node27096 : node27059;
											assign node27059 = (inp[3]) ? node27075 : node27060;
												assign node27060 = (inp[0]) ? node27068 : node27061;
													assign node27061 = (inp[15]) ? node27065 : node27062;
														assign node27062 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node27065 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node27068 = (inp[9]) ? node27072 : node27069;
														assign node27069 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27072 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node27075 = (inp[10]) ? node27089 : node27076;
													assign node27076 = (inp[0]) ? node27082 : node27077;
														assign node27077 = (inp[9]) ? 4'b0100 : node27078;
															assign node27078 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27082 = (inp[15]) ? node27086 : node27083;
															assign node27083 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node27086 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node27089 = (inp[15]) ? node27093 : node27090;
														assign node27090 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node27093 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node27096 = (inp[3]) ? node27104 : node27097;
												assign node27097 = (inp[9]) ? node27101 : node27098;
													assign node27098 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node27101 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node27104 = (inp[15]) ? node27108 : node27105;
													assign node27105 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node27108 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node27111 = (inp[0]) ? node27147 : node27112;
											assign node27112 = (inp[3]) ? node27140 : node27113;
												assign node27113 = (inp[2]) ? node27121 : node27114;
													assign node27114 = (inp[15]) ? node27118 : node27115;
														assign node27115 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node27118 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node27121 = (inp[10]) ? node27131 : node27122;
														assign node27122 = (inp[5]) ? 4'b0101 : node27123;
															assign node27123 = (inp[9]) ? node27127 : node27124;
																assign node27124 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node27127 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node27131 = (inp[5]) ? node27133 : 4'b0101;
															assign node27133 = (inp[15]) ? node27137 : node27134;
																assign node27134 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node27137 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node27140 = (inp[9]) ? node27144 : node27141;
													assign node27141 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node27144 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node27147 = (inp[10]) ? node27163 : node27148;
												assign node27148 = (inp[3]) ? node27156 : node27149;
													assign node27149 = (inp[9]) ? node27153 : node27150;
														assign node27150 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27153 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node27156 = (inp[9]) ? node27160 : node27157;
														assign node27157 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27160 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node27163 = (inp[15]) ? node27167 : node27164;
													assign node27164 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node27167 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node27170 = (inp[3]) ? node27178 : node27171;
										assign node27171 = (inp[15]) ? node27175 : node27172;
											assign node27172 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node27175 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node27178 = (inp[0]) ? node27228 : node27179;
											assign node27179 = (inp[10]) ? node27203 : node27180;
												assign node27180 = (inp[11]) ? node27196 : node27181;
													assign node27181 = (inp[2]) ? node27191 : node27182;
														assign node27182 = (inp[5]) ? 4'b0101 : node27183;
															assign node27183 = (inp[15]) ? node27187 : node27184;
																assign node27184 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node27187 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node27191 = (inp[15]) ? 4'b0100 : node27192;
															assign node27192 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node27196 = (inp[9]) ? node27200 : node27197;
														assign node27197 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27200 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node27203 = (inp[11]) ? node27215 : node27204;
													assign node27204 = (inp[2]) ? node27210 : node27205;
														assign node27205 = (inp[5]) ? 4'b0101 : node27206;
															assign node27206 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node27210 = (inp[9]) ? 4'b0101 : node27211;
															assign node27211 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node27215 = (inp[2]) ? node27221 : node27216;
														assign node27216 = (inp[9]) ? 4'b0101 : node27217;
															assign node27217 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node27221 = (inp[5]) ? node27223 : 4'b0101;
															assign node27223 = (inp[9]) ? node27225 : 4'b0101;
																assign node27225 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node27228 = (inp[9]) ? node27232 : node27229;
												assign node27229 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node27232 = (inp[15]) ? 4'b0100 : 4'b0101;
							assign node27235 = (inp[1]) ? node27407 : node27236;
								assign node27236 = (inp[3]) ? node27316 : node27237;
									assign node27237 = (inp[15]) ? node27245 : node27238;
										assign node27238 = (inp[9]) ? node27242 : node27239;
											assign node27239 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node27242 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node27245 = (inp[10]) ? node27279 : node27246;
											assign node27246 = (inp[0]) ? node27272 : node27247;
												assign node27247 = (inp[5]) ? node27255 : node27248;
													assign node27248 = (inp[12]) ? node27252 : node27249;
														assign node27249 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node27252 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node27255 = (inp[11]) ? node27263 : node27256;
														assign node27256 = (inp[12]) ? node27260 : node27257;
															assign node27257 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node27260 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node27263 = (inp[2]) ? node27265 : 4'b0101;
															assign node27265 = (inp[12]) ? node27269 : node27266;
																assign node27266 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node27269 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node27272 = (inp[9]) ? node27276 : node27273;
													assign node27273 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node27276 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node27279 = (inp[9]) ? node27287 : node27280;
												assign node27280 = (inp[12]) ? node27284 : node27281;
													assign node27281 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node27284 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node27287 = (inp[2]) ? node27297 : node27288;
													assign node27288 = (inp[5]) ? 4'b0100 : node27289;
														assign node27289 = (inp[12]) ? node27293 : node27290;
															assign node27290 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node27293 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node27297 = (inp[5]) ? node27303 : node27298;
														assign node27298 = (inp[0]) ? node27300 : 4'b0100;
															assign node27300 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node27303 = (inp[11]) ? node27309 : node27304;
															assign node27304 = (inp[0]) ? 4'b0100 : node27305;
																assign node27305 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node27309 = (inp[12]) ? node27313 : node27310;
																assign node27310 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node27313 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node27316 = (inp[11]) ? node27340 : node27317;
										assign node27317 = (inp[9]) ? node27329 : node27318;
											assign node27318 = (inp[12]) ? node27324 : node27319;
												assign node27319 = (inp[0]) ? 4'b0000 : node27320;
													assign node27320 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node27324 = (inp[0]) ? 4'b0001 : node27325;
													assign node27325 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node27329 = (inp[12]) ? node27335 : node27330;
												assign node27330 = (inp[0]) ? 4'b0001 : node27331;
													assign node27331 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node27335 = (inp[0]) ? 4'b0000 : node27336;
													assign node27336 = (inp[15]) ? 4'b0000 : 4'b0001;
										assign node27340 = (inp[10]) ? node27384 : node27341;
											assign node27341 = (inp[15]) ? node27363 : node27342;
												assign node27342 = (inp[12]) ? node27350 : node27343;
													assign node27343 = (inp[0]) ? node27347 : node27344;
														assign node27344 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node27347 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node27350 = (inp[5]) ? node27358 : node27351;
														assign node27351 = (inp[0]) ? node27355 : node27352;
															assign node27352 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node27355 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node27358 = (inp[2]) ? 4'b0001 : node27359;
															assign node27359 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node27363 = (inp[2]) ? node27377 : node27364;
													assign node27364 = (inp[0]) ? node27370 : node27365;
														assign node27365 = (inp[9]) ? 4'b0001 : node27366;
															assign node27366 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node27370 = (inp[9]) ? node27374 : node27371;
															assign node27371 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node27374 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node27377 = (inp[5]) ? node27379 : 4'b0000;
														assign node27379 = (inp[9]) ? node27381 : 4'b0000;
															assign node27381 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node27384 = (inp[12]) ? node27396 : node27385;
												assign node27385 = (inp[9]) ? node27391 : node27386;
													assign node27386 = (inp[0]) ? 4'b0000 : node27387;
														assign node27387 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node27391 = (inp[15]) ? 4'b0001 : node27392;
														assign node27392 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node27396 = (inp[9]) ? node27402 : node27397;
													assign node27397 = (inp[0]) ? 4'b0001 : node27398;
														assign node27398 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node27402 = (inp[15]) ? 4'b0000 : node27403;
														assign node27403 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node27407 = (inp[9]) ? node27413 : node27408;
									assign node27408 = (inp[0]) ? 4'b0001 : node27409;
										assign node27409 = (inp[3]) ? 4'b0001 : 4'b0000;
									assign node27413 = (inp[0]) ? 4'b0000 : node27414;
										assign node27414 = (inp[3]) ? 4'b0000 : 4'b0001;
		assign node27418 = (inp[6]) ? node37778 : node27419;
			assign node27419 = (inp[3]) ? node33523 : node27420;
				assign node27420 = (inp[2]) ? node30500 : node27421;
					assign node27421 = (inp[1]) ? node28999 : node27422;
						assign node27422 = (inp[7]) ? node28188 : node27423;
							assign node27423 = (inp[14]) ? node27741 : node27424;
								assign node27424 = (inp[4]) ? node27554 : node27425;
									assign node27425 = (inp[12]) ? node27507 : node27426;
										assign node27426 = (inp[5]) ? node27472 : node27427;
											assign node27427 = (inp[11]) ? node27449 : node27428;
												assign node27428 = (inp[13]) ? node27436 : node27429;
													assign node27429 = (inp[10]) ? node27433 : node27430;
														assign node27430 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node27433 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node27436 = (inp[10]) ? node27444 : node27437;
														assign node27437 = (inp[9]) ? node27439 : 4'b1000;
															assign node27439 = (inp[15]) ? 4'b1001 : node27440;
																assign node27440 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node27444 = (inp[0]) ? node27446 : 4'b1001;
															assign node27446 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node27449 = (inp[10]) ? node27461 : node27450;
													assign node27450 = (inp[0]) ? node27456 : node27451;
														assign node27451 = (inp[15]) ? 4'b1000 : node27452;
															assign node27452 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node27456 = (inp[13]) ? node27458 : 4'b1001;
															assign node27458 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node27461 = (inp[0]) ? node27467 : node27462;
														assign node27462 = (inp[9]) ? node27464 : 4'b1001;
															assign node27464 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node27467 = (inp[13]) ? node27469 : 4'b1000;
															assign node27469 = (inp[15]) ? 4'b1000 : 4'b1001;
											assign node27472 = (inp[10]) ? node27490 : node27473;
												assign node27473 = (inp[0]) ? node27483 : node27474;
													assign node27474 = (inp[13]) ? node27476 : 4'b1000;
														assign node27476 = (inp[15]) ? node27480 : node27477;
															assign node27477 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node27480 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node27483 = (inp[13]) ? node27485 : 4'b1001;
														assign node27485 = (inp[11]) ? 4'b1001 : node27486;
															assign node27486 = (inp[15]) ? 4'b1000 : 4'b1001;
												assign node27490 = (inp[0]) ? node27498 : node27491;
													assign node27491 = (inp[13]) ? node27493 : 4'b1001;
														assign node27493 = (inp[11]) ? node27495 : 4'b1001;
															assign node27495 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node27498 = (inp[13]) ? node27500 : 4'b1000;
														assign node27500 = (inp[15]) ? node27504 : node27501;
															assign node27501 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node27504 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node27507 = (inp[15]) ? node27531 : node27508;
											assign node27508 = (inp[0]) ? node27520 : node27509;
												assign node27509 = (inp[10]) ? node27515 : node27510;
													assign node27510 = (inp[5]) ? 4'b1010 : node27511;
														assign node27511 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node27515 = (inp[13]) ? node27517 : 4'b1011;
														assign node27517 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node27520 = (inp[10]) ? node27526 : node27521;
													assign node27521 = (inp[11]) ? node27523 : 4'b1011;
														assign node27523 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node27526 = (inp[13]) ? node27528 : 4'b1010;
														assign node27528 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node27531 = (inp[10]) ? node27543 : node27532;
												assign node27532 = (inp[0]) ? node27538 : node27533;
													assign node27533 = (inp[11]) ? 4'b1010 : node27534;
														assign node27534 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node27538 = (inp[11]) ? 4'b1011 : node27539;
														assign node27539 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node27543 = (inp[0]) ? node27549 : node27544;
													assign node27544 = (inp[13]) ? node27546 : 4'b1011;
														assign node27546 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node27549 = (inp[11]) ? 4'b1010 : node27550;
														assign node27550 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node27554 = (inp[12]) ? node27650 : node27555;
										assign node27555 = (inp[15]) ? node27601 : node27556;
											assign node27556 = (inp[13]) ? node27578 : node27557;
												assign node27557 = (inp[5]) ? node27565 : node27558;
													assign node27558 = (inp[9]) ? node27560 : 4'b1010;
														assign node27560 = (inp[10]) ? node27562 : 4'b1011;
															assign node27562 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node27565 = (inp[0]) ? node27571 : node27566;
														assign node27566 = (inp[11]) ? node27568 : 4'b1011;
															assign node27568 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node27571 = (inp[10]) ? node27575 : node27572;
															assign node27572 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node27575 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node27578 = (inp[10]) ? node27590 : node27579;
													assign node27579 = (inp[5]) ? 4'b1011 : node27580;
														assign node27580 = (inp[9]) ? node27586 : node27581;
															assign node27581 = (inp[11]) ? 4'b1011 : node27582;
																assign node27582 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node27586 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node27590 = (inp[0]) ? node27596 : node27591;
														assign node27591 = (inp[5]) ? 4'b1010 : node27592;
															assign node27592 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node27596 = (inp[5]) ? 4'b1011 : node27597;
															assign node27597 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node27601 = (inp[5]) ? node27627 : node27602;
												assign node27602 = (inp[10]) ? node27616 : node27603;
													assign node27603 = (inp[9]) ? node27611 : node27604;
														assign node27604 = (inp[13]) ? node27606 : 4'b1010;
															assign node27606 = (inp[11]) ? 4'b1011 : node27607;
																assign node27607 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node27611 = (inp[0]) ? node27613 : 4'b1010;
															assign node27613 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node27616 = (inp[0]) ? node27622 : node27617;
														assign node27617 = (inp[13]) ? node27619 : 4'b1011;
															assign node27619 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node27622 = (inp[13]) ? node27624 : 4'b1010;
															assign node27624 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node27627 = (inp[9]) ? node27633 : node27628;
													assign node27628 = (inp[0]) ? node27630 : 4'b1111;
														assign node27630 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node27633 = (inp[13]) ? node27643 : node27634;
														assign node27634 = (inp[11]) ? 4'b1110 : node27635;
															assign node27635 = (inp[10]) ? node27639 : node27636;
																assign node27636 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node27639 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node27643 = (inp[0]) ? node27647 : node27644;
															assign node27644 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node27647 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node27650 = (inp[15]) ? node27686 : node27651;
											assign node27651 = (inp[5]) ? node27673 : node27652;
												assign node27652 = (inp[10]) ? node27664 : node27653;
													assign node27653 = (inp[0]) ? node27659 : node27654;
														assign node27654 = (inp[13]) ? node27656 : 4'b1100;
															assign node27656 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node27659 = (inp[11]) ? node27661 : 4'b1101;
															assign node27661 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node27664 = (inp[0]) ? node27670 : node27665;
														assign node27665 = (inp[11]) ? node27667 : 4'b1101;
															assign node27667 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node27670 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node27673 = (inp[0]) ? node27677 : node27674;
													assign node27674 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node27677 = (inp[10]) ? node27683 : node27678;
														assign node27678 = (inp[13]) ? node27680 : 4'b1000;
															assign node27680 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node27683 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node27686 = (inp[13]) ? node27706 : node27687;
												assign node27687 = (inp[5]) ? node27701 : node27688;
													assign node27688 = (inp[11]) ? node27696 : node27689;
														assign node27689 = (inp[0]) ? node27693 : node27690;
															assign node27690 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node27693 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node27696 = (inp[9]) ? node27698 : 4'b1001;
															assign node27698 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node27701 = (inp[0]) ? 4'b1001 : node27702;
														assign node27702 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node27706 = (inp[11]) ? node27714 : node27707;
													assign node27707 = (inp[0]) ? node27711 : node27708;
														assign node27708 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node27711 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node27714 = (inp[9]) ? node27728 : node27715;
														assign node27715 = (inp[5]) ? node27723 : node27716;
															assign node27716 = (inp[0]) ? node27720 : node27717;
																assign node27717 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node27720 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node27723 = (inp[0]) ? 4'b1001 : node27724;
																assign node27724 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node27728 = (inp[5]) ? node27734 : node27729;
															assign node27729 = (inp[0]) ? node27731 : 4'b1000;
																assign node27731 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node27734 = (inp[10]) ? node27738 : node27735;
																assign node27735 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node27738 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node27741 = (inp[4]) ? node27947 : node27742;
									assign node27742 = (inp[12]) ? node27856 : node27743;
										assign node27743 = (inp[15]) ? node27793 : node27744;
											assign node27744 = (inp[5]) ? node27766 : node27745;
												assign node27745 = (inp[9]) ? node27757 : node27746;
													assign node27746 = (inp[13]) ? node27754 : node27747;
														assign node27747 = (inp[10]) ? 4'b1000 : node27748;
															assign node27748 = (inp[0]) ? node27750 : 4'b1000;
																assign node27750 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node27754 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node27757 = (inp[10]) ? 4'b1001 : node27758;
														assign node27758 = (inp[0]) ? node27760 : 4'b1000;
															assign node27760 = (inp[11]) ? node27762 : 4'b1001;
																assign node27762 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node27766 = (inp[9]) ? node27780 : node27767;
													assign node27767 = (inp[10]) ? node27775 : node27768;
														assign node27768 = (inp[11]) ? node27770 : 4'b1100;
															assign node27770 = (inp[13]) ? node27772 : 4'b1101;
																assign node27772 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node27775 = (inp[0]) ? 4'b1100 : node27776;
															assign node27776 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node27780 = (inp[11]) ? node27786 : node27781;
														assign node27781 = (inp[0]) ? 4'b1101 : node27782;
															assign node27782 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node27786 = (inp[10]) ? node27790 : node27787;
															assign node27787 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node27790 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node27793 = (inp[9]) ? node27827 : node27794;
												assign node27794 = (inp[11]) ? node27816 : node27795;
													assign node27795 = (inp[13]) ? node27801 : node27796;
														assign node27796 = (inp[10]) ? 4'b1000 : node27797;
															assign node27797 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node27801 = (inp[10]) ? node27809 : node27802;
															assign node27802 = (inp[5]) ? node27806 : node27803;
																assign node27803 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node27806 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27809 = (inp[5]) ? node27813 : node27810;
																assign node27810 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node27813 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node27816 = (inp[0]) ? node27818 : 4'b1001;
														assign node27818 = (inp[5]) ? node27820 : 4'b1001;
															assign node27820 = (inp[10]) ? node27824 : node27821;
																assign node27821 = (inp[13]) ? 4'b1000 : 4'b1001;
																assign node27824 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node27827 = (inp[0]) ? node27841 : node27828;
													assign node27828 = (inp[10]) ? node27836 : node27829;
														assign node27829 = (inp[11]) ? node27831 : 4'b1000;
															assign node27831 = (inp[13]) ? 4'b1001 : node27832;
																assign node27832 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node27836 = (inp[11]) ? node27838 : 4'b1001;
															assign node27838 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node27841 = (inp[5]) ? node27851 : node27842;
														assign node27842 = (inp[10]) ? node27848 : node27843;
															assign node27843 = (inp[13]) ? 4'b1000 : node27844;
																assign node27844 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node27848 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node27851 = (inp[10]) ? 4'b1000 : node27852;
															assign node27852 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node27856 = (inp[5]) ? node27898 : node27857;
											assign node27857 = (inp[15]) ? node27877 : node27858;
												assign node27858 = (inp[10]) ? node27866 : node27859;
													assign node27859 = (inp[0]) ? node27863 : node27860;
														assign node27860 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node27863 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node27866 = (inp[0]) ? node27872 : node27867;
														assign node27867 = (inp[13]) ? 4'b1011 : node27868;
															assign node27868 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node27872 = (inp[11]) ? node27874 : 4'b1010;
															assign node27874 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node27877 = (inp[0]) ? node27889 : node27878;
													assign node27878 = (inp[10]) ? node27884 : node27879;
														assign node27879 = (inp[13]) ? 4'b1111 : node27880;
															assign node27880 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node27884 = (inp[11]) ? 4'b1110 : node27885;
															assign node27885 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node27889 = (inp[10]) ? node27893 : node27890;
														assign node27890 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node27893 = (inp[11]) ? 4'b1111 : node27894;
															assign node27894 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node27898 = (inp[11]) ? node27924 : node27899;
												assign node27899 = (inp[10]) ? node27909 : node27900;
													assign node27900 = (inp[0]) ? node27906 : node27901;
														assign node27901 = (inp[15]) ? 4'b1010 : node27902;
															assign node27902 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node27906 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node27909 = (inp[9]) ? node27915 : node27910;
														assign node27910 = (inp[0]) ? 4'b1010 : node27911;
															assign node27911 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node27915 = (inp[0]) ? node27921 : node27916;
															assign node27916 = (inp[13]) ? node27918 : 4'b1011;
																assign node27918 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node27921 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node27924 = (inp[9]) ? node27938 : node27925;
													assign node27925 = (inp[0]) ? node27933 : node27926;
														assign node27926 = (inp[13]) ? node27930 : node27927;
															assign node27927 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node27930 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node27933 = (inp[10]) ? node27935 : 4'b1011;
															assign node27935 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node27938 = (inp[0]) ? 4'b1010 : node27939;
														assign node27939 = (inp[13]) ? node27943 : node27940;
															assign node27940 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node27943 = (inp[10]) ? 4'b1010 : 4'b1011;
									assign node27947 = (inp[12]) ? node28087 : node27948;
										assign node27948 = (inp[9]) ? node28008 : node27949;
											assign node27949 = (inp[11]) ? node27987 : node27950;
												assign node27950 = (inp[10]) ? node27976 : node27951;
													assign node27951 = (inp[0]) ? node27963 : node27952;
														assign node27952 = (inp[5]) ? node27956 : node27953;
															assign node27953 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node27956 = (inp[15]) ? node27960 : node27957;
																assign node27957 = (inp[13]) ? 4'b1111 : 4'b1110;
																assign node27960 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node27963 = (inp[5]) ? node27969 : node27964;
															assign node27964 = (inp[15]) ? node27966 : 4'b1011;
																assign node27966 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node27969 = (inp[15]) ? node27973 : node27970;
																assign node27970 = (inp[13]) ? 4'b1110 : 4'b1111;
																assign node27973 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node27976 = (inp[0]) ? node27980 : node27977;
														assign node27977 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node27980 = (inp[5]) ? node27982 : 4'b1010;
															assign node27982 = (inp[15]) ? 4'b1010 : node27983;
																assign node27983 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node27987 = (inp[10]) ? node27997 : node27988;
													assign node27988 = (inp[0]) ? node27994 : node27989;
														assign node27989 = (inp[15]) ? 4'b1010 : node27990;
															assign node27990 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node27994 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node27997 = (inp[5]) ? 4'b1011 : node27998;
														assign node27998 = (inp[15]) ? node28004 : node27999;
															assign node27999 = (inp[13]) ? 4'b1011 : node28000;
																assign node28000 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28004 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node28008 = (inp[13]) ? node28052 : node28009;
												assign node28009 = (inp[15]) ? node28031 : node28010;
													assign node28010 = (inp[5]) ? node28024 : node28011;
														assign node28011 = (inp[0]) ? node28019 : node28012;
															assign node28012 = (inp[11]) ? node28016 : node28013;
																assign node28013 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node28016 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node28019 = (inp[11]) ? node28021 : 4'b1011;
																assign node28021 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node28024 = (inp[10]) ? node28028 : node28025;
															assign node28025 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node28028 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node28031 = (inp[5]) ? node28043 : node28032;
														assign node28032 = (inp[10]) ? node28038 : node28033;
															assign node28033 = (inp[11]) ? node28035 : 4'b1110;
																assign node28035 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node28038 = (inp[0]) ? 4'b1111 : node28039;
																assign node28039 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node28043 = (inp[0]) ? 4'b1010 : node28044;
															assign node28044 = (inp[11]) ? node28048 : node28045;
																assign node28045 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node28048 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node28052 = (inp[0]) ? node28068 : node28053;
													assign node28053 = (inp[11]) ? node28061 : node28054;
														assign node28054 = (inp[10]) ? 4'b1110 : node28055;
															assign node28055 = (inp[5]) ? 4'b1010 : node28056;
																assign node28056 = (inp[15]) ? 4'b1111 : 4'b1010;
														assign node28061 = (inp[5]) ? node28065 : node28062;
															assign node28062 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node28065 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node28068 = (inp[10]) ? node28076 : node28069;
														assign node28069 = (inp[15]) ? node28073 : node28070;
															assign node28070 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node28073 = (inp[5]) ? 4'b1011 : 4'b1110;
														assign node28076 = (inp[11]) ? node28082 : node28077;
															assign node28077 = (inp[15]) ? 4'b1010 : node28078;
																assign node28078 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node28082 = (inp[5]) ? node28084 : 4'b1111;
																assign node28084 = (inp[15]) ? 4'b1010 : 4'b1110;
										assign node28087 = (inp[5]) ? node28151 : node28088;
											assign node28088 = (inp[15]) ? node28120 : node28089;
												assign node28089 = (inp[9]) ? node28103 : node28090;
													assign node28090 = (inp[0]) ? 4'b1000 : node28091;
														assign node28091 = (inp[10]) ? node28097 : node28092;
															assign node28092 = (inp[13]) ? node28094 : 4'b1000;
																assign node28094 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node28097 = (inp[13]) ? node28099 : 4'b1001;
																assign node28099 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28103 = (inp[10]) ? node28111 : node28104;
														assign node28104 = (inp[0]) ? node28106 : 4'b1000;
															assign node28106 = (inp[13]) ? node28108 : 4'b1001;
																assign node28108 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node28111 = (inp[0]) ? node28117 : node28112;
															assign node28112 = (inp[11]) ? 4'b1001 : node28113;
																assign node28113 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node28117 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node28120 = (inp[11]) ? node28138 : node28121;
													assign node28121 = (inp[13]) ? node28133 : node28122;
														assign node28122 = (inp[9]) ? node28128 : node28123;
															assign node28123 = (inp[10]) ? node28125 : 4'b1101;
																assign node28125 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node28128 = (inp[0]) ? node28130 : 4'b1100;
																assign node28130 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node28133 = (inp[0]) ? node28135 : 4'b1101;
															assign node28135 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node28138 = (inp[0]) ? node28144 : node28139;
														assign node28139 = (inp[13]) ? 4'b1100 : node28140;
															assign node28140 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node28144 = (inp[10]) ? node28148 : node28145;
															assign node28145 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node28148 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node28151 = (inp[15]) ? node28173 : node28152;
												assign node28152 = (inp[0]) ? node28164 : node28153;
													assign node28153 = (inp[10]) ? node28159 : node28154;
														assign node28154 = (inp[11]) ? node28156 : 4'b1101;
															assign node28156 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node28159 = (inp[13]) ? 4'b1100 : node28160;
															assign node28160 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node28164 = (inp[10]) ? node28170 : node28165;
														assign node28165 = (inp[13]) ? 4'b1100 : node28166;
															assign node28166 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node28170 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node28173 = (inp[10]) ? node28183 : node28174;
													assign node28174 = (inp[13]) ? node28176 : 4'b1000;
														assign node28176 = (inp[11]) ? node28180 : node28177;
															assign node28177 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node28180 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node28183 = (inp[0]) ? 4'b1001 : node28184;
														assign node28184 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node28188 = (inp[14]) ? node28586 : node28189;
								assign node28189 = (inp[4]) ? node28393 : node28190;
									assign node28190 = (inp[12]) ? node28308 : node28191;
										assign node28191 = (inp[0]) ? node28235 : node28192;
											assign node28192 = (inp[13]) ? node28208 : node28193;
												assign node28193 = (inp[10]) ? node28201 : node28194;
													assign node28194 = (inp[5]) ? node28198 : node28195;
														assign node28195 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node28198 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node28201 = (inp[5]) ? node28203 : 4'b1001;
														assign node28203 = (inp[15]) ? node28205 : 4'b1100;
															assign node28205 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node28208 = (inp[15]) ? node28228 : node28209;
													assign node28209 = (inp[5]) ? node28223 : node28210;
														assign node28210 = (inp[9]) ? node28216 : node28211;
															assign node28211 = (inp[10]) ? 4'b1001 : node28212;
																assign node28212 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node28216 = (inp[11]) ? node28220 : node28217;
																assign node28217 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node28220 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node28223 = (inp[10]) ? 4'b1101 : node28224;
															assign node28224 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node28228 = (inp[10]) ? 4'b1000 : node28229;
														assign node28229 = (inp[5]) ? 4'b1001 : node28230;
															assign node28230 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node28235 = (inp[9]) ? node28271 : node28236;
												assign node28236 = (inp[11]) ? node28254 : node28237;
													assign node28237 = (inp[10]) ? node28247 : node28238;
														assign node28238 = (inp[13]) ? node28240 : 4'b1101;
															assign node28240 = (inp[5]) ? node28244 : node28241;
																assign node28241 = (inp[15]) ? 4'b1100 : 4'b1001;
																assign node28244 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node28247 = (inp[5]) ? node28251 : node28248;
															assign node28248 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node28251 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node28254 = (inp[10]) ? node28262 : node28255;
														assign node28255 = (inp[15]) ? 4'b1101 : node28256;
															assign node28256 = (inp[5]) ? node28258 : 4'b1000;
																assign node28258 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node28262 = (inp[5]) ? node28266 : node28263;
															assign node28263 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node28266 = (inp[15]) ? 4'b1000 : node28267;
																assign node28267 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node28271 = (inp[13]) ? node28287 : node28272;
													assign node28272 = (inp[15]) ? node28278 : node28273;
														assign node28273 = (inp[5]) ? node28275 : 4'b1000;
															assign node28275 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node28278 = (inp[5]) ? node28282 : node28279;
															assign node28279 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node28282 = (inp[10]) ? 4'b1000 : node28283;
																assign node28283 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28287 = (inp[10]) ? node28295 : node28288;
														assign node28288 = (inp[5]) ? 4'b1000 : node28289;
															assign node28289 = (inp[15]) ? node28291 : 4'b1001;
																assign node28291 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node28295 = (inp[15]) ? node28303 : node28296;
															assign node28296 = (inp[5]) ? node28300 : node28297;
																assign node28297 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node28300 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node28303 = (inp[5]) ? 4'b1001 : node28304;
																assign node28304 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node28308 = (inp[5]) ? node28350 : node28309;
											assign node28309 = (inp[15]) ? node28327 : node28310;
												assign node28310 = (inp[10]) ? node28320 : node28311;
													assign node28311 = (inp[0]) ? node28315 : node28312;
														assign node28312 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node28315 = (inp[11]) ? 4'b1010 : node28316;
															assign node28316 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node28320 = (inp[0]) ? node28324 : node28321;
														assign node28321 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28324 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node28327 = (inp[10]) ? node28337 : node28328;
													assign node28328 = (inp[0]) ? node28334 : node28329;
														assign node28329 = (inp[11]) ? node28331 : 4'b1110;
															assign node28331 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node28334 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node28337 = (inp[0]) ? node28345 : node28338;
														assign node28338 = (inp[9]) ? 4'b1111 : node28339;
															assign node28339 = (inp[13]) ? 4'b1111 : node28340;
																assign node28340 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node28345 = (inp[13]) ? 4'b1110 : node28346;
															assign node28346 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node28350 = (inp[15]) ? node28372 : node28351;
												assign node28351 = (inp[11]) ? node28367 : node28352;
													assign node28352 = (inp[10]) ? node28360 : node28353;
														assign node28353 = (inp[0]) ? node28357 : node28354;
															assign node28354 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node28357 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node28360 = (inp[0]) ? node28364 : node28361;
															assign node28361 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node28364 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node28367 = (inp[10]) ? node28369 : 4'b1111;
														assign node28369 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node28372 = (inp[0]) ? node28382 : node28373;
													assign node28373 = (inp[10]) ? node28377 : node28374;
														assign node28374 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28377 = (inp[9]) ? 4'b1011 : node28378;
															assign node28378 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node28382 = (inp[10]) ? node28388 : node28383;
														assign node28383 = (inp[13]) ? node28385 : 4'b1011;
															assign node28385 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node28388 = (inp[13]) ? node28390 : 4'b1010;
															assign node28390 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node28393 = (inp[12]) ? node28505 : node28394;
										assign node28394 = (inp[15]) ? node28440 : node28395;
											assign node28395 = (inp[5]) ? node28421 : node28396;
												assign node28396 = (inp[9]) ? node28410 : node28397;
													assign node28397 = (inp[13]) ? node28405 : node28398;
														assign node28398 = (inp[0]) ? node28402 : node28399;
															assign node28399 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node28402 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28405 = (inp[10]) ? 4'b1011 : node28406;
															assign node28406 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node28410 = (inp[11]) ? 4'b1010 : node28411;
														assign node28411 = (inp[13]) ? 4'b1010 : node28412;
															assign node28412 = (inp[10]) ? node28416 : node28413;
																assign node28413 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node28416 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node28421 = (inp[0]) ? node28429 : node28422;
													assign node28422 = (inp[10]) ? node28424 : 4'b1110;
														assign node28424 = (inp[13]) ? 4'b1111 : node28425;
															assign node28425 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node28429 = (inp[10]) ? node28435 : node28430;
														assign node28430 = (inp[13]) ? 4'b1111 : node28431;
															assign node28431 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node28435 = (inp[11]) ? 4'b1110 : node28436;
															assign node28436 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node28440 = (inp[9]) ? node28474 : node28441;
												assign node28441 = (inp[11]) ? node28455 : node28442;
													assign node28442 = (inp[5]) ? node28450 : node28443;
														assign node28443 = (inp[10]) ? node28447 : node28444;
															assign node28444 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28447 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node28450 = (inp[0]) ? 4'b1010 : node28451;
															assign node28451 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node28455 = (inp[5]) ? node28465 : node28456;
														assign node28456 = (inp[13]) ? 4'b1010 : node28457;
															assign node28457 = (inp[10]) ? node28461 : node28458;
																assign node28458 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node28461 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28465 = (inp[13]) ? 4'b1011 : node28466;
															assign node28466 = (inp[0]) ? node28470 : node28467;
																assign node28467 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node28470 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node28474 = (inp[10]) ? node28486 : node28475;
													assign node28475 = (inp[0]) ? node28481 : node28476;
														assign node28476 = (inp[5]) ? node28478 : 4'b1010;
															assign node28478 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28481 = (inp[11]) ? 4'b1011 : node28482;
															assign node28482 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node28486 = (inp[0]) ? node28498 : node28487;
														assign node28487 = (inp[11]) ? node28493 : node28488;
															assign node28488 = (inp[13]) ? node28490 : 4'b1011;
																assign node28490 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node28493 = (inp[5]) ? 4'b1011 : node28494;
																assign node28494 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node28498 = (inp[13]) ? 4'b1010 : node28499;
															assign node28499 = (inp[5]) ? 4'b1010 : node28500;
																assign node28500 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node28505 = (inp[15]) ? node28541 : node28506;
											assign node28506 = (inp[0]) ? node28528 : node28507;
												assign node28507 = (inp[10]) ? node28517 : node28508;
													assign node28508 = (inp[9]) ? node28514 : node28509;
														assign node28509 = (inp[5]) ? node28511 : 4'b1001;
															assign node28511 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node28514 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node28517 = (inp[9]) ? node28519 : 4'b1000;
														assign node28519 = (inp[5]) ? node28525 : node28520;
															assign node28520 = (inp[11]) ? node28522 : 4'b1000;
																assign node28522 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node28525 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node28528 = (inp[10]) ? node28530 : 4'b1000;
													assign node28530 = (inp[9]) ? 4'b1001 : node28531;
														assign node28531 = (inp[5]) ? node28537 : node28532;
															assign node28532 = (inp[13]) ? node28534 : 4'b1001;
																assign node28534 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node28537 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node28541 = (inp[5]) ? node28569 : node28542;
												assign node28542 = (inp[13]) ? node28550 : node28543;
													assign node28543 = (inp[0]) ? node28547 : node28544;
														assign node28544 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node28547 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node28550 = (inp[10]) ? node28562 : node28551;
														assign node28551 = (inp[9]) ? node28557 : node28552;
															assign node28552 = (inp[11]) ? node28554 : 4'b1100;
																assign node28554 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node28557 = (inp[11]) ? 4'b1100 : node28558;
																assign node28558 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node28562 = (inp[11]) ? node28566 : node28563;
															assign node28563 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node28566 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node28569 = (inp[13]) ? node28577 : node28570;
													assign node28570 = (inp[0]) ? node28574 : node28571;
														assign node28571 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node28574 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node28577 = (inp[10]) ? node28579 : 4'b1001;
														assign node28579 = (inp[0]) ? node28583 : node28580;
															assign node28580 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node28583 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node28586 = (inp[4]) ? node28810 : node28587;
									assign node28587 = (inp[12]) ? node28707 : node28588;
										assign node28588 = (inp[15]) ? node28656 : node28589;
											assign node28589 = (inp[9]) ? node28617 : node28590;
												assign node28590 = (inp[10]) ? node28600 : node28591;
													assign node28591 = (inp[13]) ? node28595 : node28592;
														assign node28592 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node28595 = (inp[0]) ? 4'b1001 : node28596;
															assign node28596 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node28600 = (inp[5]) ? node28608 : node28601;
														assign node28601 = (inp[13]) ? 4'b1000 : node28602;
															assign node28602 = (inp[11]) ? node28604 : 4'b1001;
																assign node28604 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node28608 = (inp[11]) ? 4'b1001 : node28609;
															assign node28609 = (inp[13]) ? node28613 : node28610;
																assign node28610 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node28613 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node28617 = (inp[5]) ? node28629 : node28618;
													assign node28618 = (inp[13]) ? 4'b1000 : node28619;
														assign node28619 = (inp[0]) ? node28621 : 4'b1000;
															assign node28621 = (inp[10]) ? node28625 : node28622;
																assign node28622 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node28625 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28629 = (inp[13]) ? node28643 : node28630;
														assign node28630 = (inp[11]) ? node28638 : node28631;
															assign node28631 = (inp[0]) ? node28635 : node28632;
																assign node28632 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node28635 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node28638 = (inp[0]) ? node28640 : 4'b1001;
																assign node28640 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node28643 = (inp[10]) ? node28649 : node28644;
															assign node28644 = (inp[11]) ? node28646 : 4'b1000;
																assign node28646 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node28649 = (inp[0]) ? node28653 : node28650;
																assign node28650 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node28653 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node28656 = (inp[5]) ? node28680 : node28657;
												assign node28657 = (inp[9]) ? node28667 : node28658;
													assign node28658 = (inp[10]) ? node28664 : node28659;
														assign node28659 = (inp[0]) ? node28661 : 4'b1000;
															assign node28661 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node28664 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node28667 = (inp[13]) ? node28675 : node28668;
														assign node28668 = (inp[0]) ? node28672 : node28669;
															assign node28669 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node28672 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node28675 = (inp[10]) ? 4'b1001 : node28676;
															assign node28676 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node28680 = (inp[13]) ? node28696 : node28681;
													assign node28681 = (inp[9]) ? node28687 : node28682;
														assign node28682 = (inp[11]) ? 4'b1101 : node28683;
															assign node28683 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node28687 = (inp[11]) ? node28689 : 4'b1100;
															assign node28689 = (inp[0]) ? node28693 : node28690;
																assign node28690 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node28693 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node28696 = (inp[10]) ? node28698 : 4'b1100;
														assign node28698 = (inp[9]) ? 4'b1100 : node28699;
															assign node28699 = (inp[11]) ? node28703 : node28700;
																assign node28700 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node28703 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node28707 = (inp[15]) ? node28767 : node28708;
											assign node28708 = (inp[5]) ? node28742 : node28709;
												assign node28709 = (inp[13]) ? node28723 : node28710;
													assign node28710 = (inp[11]) ? node28716 : node28711;
														assign node28711 = (inp[10]) ? 4'b1111 : node28712;
															assign node28712 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28716 = (inp[0]) ? node28720 : node28717;
															assign node28717 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node28720 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node28723 = (inp[10]) ? node28735 : node28724;
														assign node28724 = (inp[9]) ? node28730 : node28725;
															assign node28725 = (inp[11]) ? 4'b1110 : node28726;
																assign node28726 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node28730 = (inp[0]) ? node28732 : 4'b1110;
																assign node28732 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node28735 = (inp[9]) ? 4'b1111 : node28736;
															assign node28736 = (inp[0]) ? 4'b1110 : node28737;
																assign node28737 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node28742 = (inp[13]) ? node28760 : node28743;
													assign node28743 = (inp[0]) ? node28751 : node28744;
														assign node28744 = (inp[9]) ? node28746 : 4'b1010;
															assign node28746 = (inp[11]) ? node28748 : 4'b1011;
																assign node28748 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node28751 = (inp[9]) ? 4'b1010 : node28752;
															assign node28752 = (inp[10]) ? node28756 : node28753;
																assign node28753 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node28756 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node28760 = (inp[0]) ? node28764 : node28761;
														assign node28761 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node28764 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node28767 = (inp[10]) ? node28783 : node28768;
												assign node28768 = (inp[0]) ? node28770 : 4'b1010;
													assign node28770 = (inp[9]) ? 4'b1011 : node28771;
														assign node28771 = (inp[5]) ? node28777 : node28772;
															assign node28772 = (inp[11]) ? 4'b1011 : node28773;
																assign node28773 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node28777 = (inp[13]) ? node28779 : 4'b1011;
																assign node28779 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node28783 = (inp[0]) ? node28799 : node28784;
													assign node28784 = (inp[9]) ? node28792 : node28785;
														assign node28785 = (inp[5]) ? node28789 : node28786;
															assign node28786 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node28789 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node28792 = (inp[11]) ? node28794 : 4'b1011;
															assign node28794 = (inp[13]) ? node28796 : 4'b1011;
																assign node28796 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node28799 = (inp[5]) ? node28805 : node28800;
														assign node28800 = (inp[11]) ? 4'b1010 : node28801;
															assign node28801 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node28805 = (inp[11]) ? node28807 : 4'b1010;
															assign node28807 = (inp[13]) ? 4'b1011 : 4'b1010;
									assign node28810 = (inp[12]) ? node28912 : node28811;
										assign node28811 = (inp[5]) ? node28849 : node28812;
											assign node28812 = (inp[0]) ? node28834 : node28813;
												assign node28813 = (inp[10]) ? node28821 : node28814;
													assign node28814 = (inp[11]) ? node28816 : 4'b1010;
														assign node28816 = (inp[13]) ? 4'b1011 : node28817;
															assign node28817 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node28821 = (inp[11]) ? node28823 : 4'b1011;
														assign node28823 = (inp[9]) ? node28829 : node28824;
															assign node28824 = (inp[15]) ? 4'b1011 : node28825;
																assign node28825 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node28829 = (inp[13]) ? node28831 : 4'b1011;
																assign node28831 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node28834 = (inp[10]) ? node28842 : node28835;
													assign node28835 = (inp[11]) ? node28837 : 4'b1011;
														assign node28837 = (inp[15]) ? node28839 : 4'b1010;
															assign node28839 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node28842 = (inp[11]) ? node28844 : 4'b1010;
														assign node28844 = (inp[13]) ? node28846 : 4'b1011;
															assign node28846 = (inp[15]) ? 4'b1011 : 4'b1010;
											assign node28849 = (inp[9]) ? node28887 : node28850;
												assign node28850 = (inp[11]) ? node28864 : node28851;
													assign node28851 = (inp[15]) ? node28857 : node28852;
														assign node28852 = (inp[10]) ? 4'b1011 : node28853;
															assign node28853 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28857 = (inp[0]) ? node28861 : node28858;
															assign node28858 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node28861 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node28864 = (inp[10]) ? node28880 : node28865;
														assign node28865 = (inp[13]) ? node28873 : node28866;
															assign node28866 = (inp[0]) ? node28870 : node28867;
																assign node28867 = (inp[15]) ? 4'b1010 : 4'b1011;
																assign node28870 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node28873 = (inp[15]) ? node28877 : node28874;
																assign node28874 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node28877 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node28880 = (inp[13]) ? node28882 : 4'b1010;
															assign node28882 = (inp[0]) ? node28884 : 4'b1010;
																assign node28884 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node28887 = (inp[11]) ? node28895 : node28888;
													assign node28888 = (inp[10]) ? node28892 : node28889;
														assign node28889 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28892 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node28895 = (inp[13]) ? node28897 : 4'b1011;
														assign node28897 = (inp[15]) ? node28905 : node28898;
															assign node28898 = (inp[10]) ? node28902 : node28899;
																assign node28899 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node28902 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node28905 = (inp[10]) ? node28909 : node28906;
																assign node28906 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node28909 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node28912 = (inp[15]) ? node28956 : node28913;
											assign node28913 = (inp[9]) ? node28941 : node28914;
												assign node28914 = (inp[5]) ? node28930 : node28915;
													assign node28915 = (inp[0]) ? node28925 : node28916;
														assign node28916 = (inp[10]) ? node28922 : node28917;
															assign node28917 = (inp[11]) ? node28919 : 4'b1001;
																assign node28919 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node28922 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node28925 = (inp[10]) ? 4'b1001 : node28926;
															assign node28926 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node28930 = (inp[13]) ? node28932 : 4'b1001;
														assign node28932 = (inp[11]) ? node28934 : 4'b1001;
															assign node28934 = (inp[0]) ? node28938 : node28935;
																assign node28935 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node28938 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node28941 = (inp[10]) ? node28953 : node28942;
													assign node28942 = (inp[0]) ? node28948 : node28943;
														assign node28943 = (inp[13]) ? 4'b1001 : node28944;
															assign node28944 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node28948 = (inp[13]) ? 4'b1000 : node28949;
															assign node28949 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28953 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node28956 = (inp[5]) ? node28980 : node28957;
												assign node28957 = (inp[0]) ? node28969 : node28958;
													assign node28958 = (inp[9]) ? node28960 : 4'b1000;
														assign node28960 = (inp[11]) ? node28962 : 4'b1000;
															assign node28962 = (inp[13]) ? node28966 : node28963;
																assign node28963 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node28966 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node28969 = (inp[10]) ? node28975 : node28970;
														assign node28970 = (inp[11]) ? node28972 : 4'b1000;
															assign node28972 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node28975 = (inp[11]) ? node28977 : 4'b1001;
															assign node28977 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node28980 = (inp[0]) ? node28992 : node28981;
													assign node28981 = (inp[10]) ? node28987 : node28982;
														assign node28982 = (inp[11]) ? node28984 : 4'b1001;
															assign node28984 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node28987 = (inp[11]) ? node28989 : 4'b1000;
															assign node28989 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node28992 = (inp[10]) ? node28996 : node28993;
														assign node28993 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node28996 = (inp[11]) ? 4'b1000 : 4'b1001;
						assign node28999 = (inp[15]) ? node29687 : node29000;
							assign node29000 = (inp[5]) ? node29314 : node29001;
								assign node29001 = (inp[12]) ? node29105 : node29002;
									assign node29002 = (inp[4]) ? node29052 : node29003;
										assign node29003 = (inp[0]) ? node29033 : node29004;
											assign node29004 = (inp[10]) ? node29024 : node29005;
												assign node29005 = (inp[11]) ? node29007 : 4'b1100;
													assign node29007 = (inp[7]) ? node29015 : node29008;
														assign node29008 = (inp[13]) ? node29012 : node29009;
															assign node29009 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node29012 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node29015 = (inp[9]) ? 4'b1100 : node29016;
															assign node29016 = (inp[13]) ? node29020 : node29017;
																assign node29017 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node29020 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node29024 = (inp[11]) ? node29026 : 4'b1101;
													assign node29026 = (inp[14]) ? node29030 : node29027;
														assign node29027 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node29030 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node29033 = (inp[10]) ? node29043 : node29034;
												assign node29034 = (inp[11]) ? node29036 : 4'b1101;
													assign node29036 = (inp[13]) ? node29040 : node29037;
														assign node29037 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node29040 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node29043 = (inp[11]) ? node29045 : 4'b1100;
													assign node29045 = (inp[13]) ? node29049 : node29046;
														assign node29046 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node29049 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node29052 = (inp[10]) ? node29084 : node29053;
											assign node29053 = (inp[0]) ? node29069 : node29054;
												assign node29054 = (inp[11]) ? node29056 : 4'b1110;
													assign node29056 = (inp[7]) ? node29062 : node29057;
														assign node29057 = (inp[14]) ? node29059 : 4'b1111;
															assign node29059 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node29062 = (inp[13]) ? node29066 : node29063;
															assign node29063 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node29066 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node29069 = (inp[11]) ? node29071 : 4'b1111;
													assign node29071 = (inp[9]) ? node29079 : node29072;
														assign node29072 = (inp[7]) ? 4'b1111 : node29073;
															assign node29073 = (inp[14]) ? node29075 : 4'b1111;
																assign node29075 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node29079 = (inp[13]) ? node29081 : 4'b1111;
															assign node29081 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node29084 = (inp[0]) ? node29092 : node29085;
												assign node29085 = (inp[11]) ? node29087 : 4'b1111;
													assign node29087 = (inp[14]) ? 4'b1110 : node29088;
														assign node29088 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node29092 = (inp[11]) ? node29094 : 4'b1110;
													assign node29094 = (inp[9]) ? node29102 : node29095;
														assign node29095 = (inp[14]) ? node29099 : node29096;
															assign node29096 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node29099 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node29102 = (inp[14]) ? 4'b1111 : 4'b1110;
									assign node29105 = (inp[4]) ? node29197 : node29106;
										assign node29106 = (inp[14]) ? node29156 : node29107;
											assign node29107 = (inp[10]) ? node29121 : node29108;
												assign node29108 = (inp[0]) ? node29116 : node29109;
													assign node29109 = (inp[7]) ? node29111 : 4'b1111;
														assign node29111 = (inp[13]) ? 4'b1110 : node29112;
															assign node29112 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node29116 = (inp[13]) ? node29118 : 4'b1110;
														assign node29118 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node29121 = (inp[9]) ? node29143 : node29122;
													assign node29122 = (inp[13]) ? node29132 : node29123;
														assign node29123 = (inp[7]) ? node29125 : 4'b1111;
															assign node29125 = (inp[0]) ? node29129 : node29126;
																assign node29126 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node29129 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29132 = (inp[0]) ? node29138 : node29133;
															assign node29133 = (inp[11]) ? 4'b1111 : node29134;
																assign node29134 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node29138 = (inp[7]) ? 4'b1110 : node29139;
																assign node29139 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node29143 = (inp[11]) ? node29149 : node29144;
														assign node29144 = (inp[0]) ? 4'b1111 : node29145;
															assign node29145 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node29149 = (inp[13]) ? 4'b1111 : node29150;
															assign node29150 = (inp[7]) ? node29152 : 4'b1110;
																assign node29152 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node29156 = (inp[7]) ? node29180 : node29157;
												assign node29157 = (inp[10]) ? node29169 : node29158;
													assign node29158 = (inp[0]) ? node29164 : node29159;
														assign node29159 = (inp[13]) ? 4'b1111 : node29160;
															assign node29160 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29164 = (inp[11]) ? node29166 : 4'b1110;
															assign node29166 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node29169 = (inp[0]) ? node29175 : node29170;
														assign node29170 = (inp[11]) ? node29172 : 4'b1110;
															assign node29172 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node29175 = (inp[11]) ? node29177 : 4'b1111;
															assign node29177 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node29180 = (inp[0]) ? node29186 : node29181;
													assign node29181 = (inp[10]) ? 4'b1011 : node29182;
														assign node29182 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node29186 = (inp[10]) ? node29192 : node29187;
														assign node29187 = (inp[11]) ? node29189 : 4'b1011;
															assign node29189 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node29192 = (inp[11]) ? node29194 : 4'b1010;
															assign node29194 = (inp[13]) ? 4'b1010 : 4'b1011;
										assign node29197 = (inp[14]) ? node29265 : node29198;
											assign node29198 = (inp[7]) ? node29236 : node29199;
												assign node29199 = (inp[9]) ? node29219 : node29200;
													assign node29200 = (inp[11]) ? node29212 : node29201;
														assign node29201 = (inp[10]) ? node29207 : node29202;
															assign node29202 = (inp[0]) ? 4'b1000 : node29203;
																assign node29203 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node29207 = (inp[0]) ? 4'b1001 : node29208;
																assign node29208 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node29212 = (inp[10]) ? node29216 : node29213;
															assign node29213 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29216 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node29219 = (inp[10]) ? node29225 : node29220;
														assign node29220 = (inp[13]) ? node29222 : 4'b1000;
															assign node29222 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node29225 = (inp[0]) ? node29231 : node29226;
															assign node29226 = (inp[13]) ? 4'b1001 : node29227;
																assign node29227 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node29231 = (inp[11]) ? 4'b1000 : node29232;
																assign node29232 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node29236 = (inp[13]) ? node29252 : node29237;
													assign node29237 = (inp[9]) ? node29245 : node29238;
														assign node29238 = (inp[10]) ? node29242 : node29239;
															assign node29239 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29242 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node29245 = (inp[0]) ? node29249 : node29246;
															assign node29246 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node29249 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node29252 = (inp[11]) ? node29254 : 4'b1100;
														assign node29254 = (inp[9]) ? node29260 : node29255;
															assign node29255 = (inp[10]) ? 4'b1100 : node29256;
																assign node29256 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node29260 = (inp[10]) ? node29262 : 4'b1100;
																assign node29262 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node29265 = (inp[10]) ? node29293 : node29266;
												assign node29266 = (inp[11]) ? node29282 : node29267;
													assign node29267 = (inp[13]) ? 4'b1100 : node29268;
														assign node29268 = (inp[9]) ? node29276 : node29269;
															assign node29269 = (inp[7]) ? node29273 : node29270;
																assign node29270 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node29273 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29276 = (inp[0]) ? 4'b1100 : node29277;
																assign node29277 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node29282 = (inp[13]) ? node29286 : node29283;
														assign node29283 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node29286 = (inp[0]) ? node29290 : node29287;
															assign node29287 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node29290 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node29293 = (inp[13]) ? node29303 : node29294;
													assign node29294 = (inp[0]) ? node29298 : node29295;
														assign node29295 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node29298 = (inp[7]) ? node29300 : 4'b1101;
															assign node29300 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node29303 = (inp[0]) ? node29309 : node29304;
														assign node29304 = (inp[11]) ? node29306 : 4'b1101;
															assign node29306 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node29309 = (inp[7]) ? 4'b1100 : node29310;
															assign node29310 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node29314 = (inp[12]) ? node29480 : node29315;
									assign node29315 = (inp[4]) ? node29405 : node29316;
										assign node29316 = (inp[10]) ? node29360 : node29317;
											assign node29317 = (inp[0]) ? node29337 : node29318;
												assign node29318 = (inp[7]) ? node29330 : node29319;
													assign node29319 = (inp[14]) ? node29325 : node29320;
														assign node29320 = (inp[11]) ? node29322 : 4'b1100;
															assign node29322 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node29325 = (inp[13]) ? node29327 : 4'b1000;
															assign node29327 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node29330 = (inp[14]) ? 4'b1101 : node29331;
														assign node29331 = (inp[13]) ? 4'b1000 : node29332;
															assign node29332 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node29337 = (inp[7]) ? node29349 : node29338;
													assign node29338 = (inp[14]) ? node29344 : node29339;
														assign node29339 = (inp[11]) ? node29341 : 4'b1101;
															assign node29341 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node29344 = (inp[13]) ? node29346 : 4'b1001;
															assign node29346 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node29349 = (inp[14]) ? node29355 : node29350;
														assign node29350 = (inp[13]) ? 4'b1001 : node29351;
															assign node29351 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29355 = (inp[13]) ? node29357 : 4'b1100;
															assign node29357 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node29360 = (inp[0]) ? node29384 : node29361;
												assign node29361 = (inp[14]) ? node29373 : node29362;
													assign node29362 = (inp[7]) ? node29368 : node29363;
														assign node29363 = (inp[13]) ? node29365 : 4'b1101;
															assign node29365 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29368 = (inp[13]) ? 4'b1001 : node29369;
															assign node29369 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node29373 = (inp[7]) ? node29379 : node29374;
														assign node29374 = (inp[13]) ? node29376 : 4'b1001;
															assign node29376 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29379 = (inp[13]) ? node29381 : 4'b1100;
															assign node29381 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node29384 = (inp[7]) ? node29396 : node29385;
													assign node29385 = (inp[14]) ? node29391 : node29386;
														assign node29386 = (inp[13]) ? node29388 : 4'b1100;
															assign node29388 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node29391 = (inp[11]) ? 4'b1000 : node29392;
															assign node29392 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node29396 = (inp[14]) ? node29400 : node29397;
														assign node29397 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node29400 = (inp[13]) ? node29402 : 4'b1101;
															assign node29402 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node29405 = (inp[10]) ? node29443 : node29406;
											assign node29406 = (inp[0]) ? node29430 : node29407;
												assign node29407 = (inp[7]) ? node29419 : node29408;
													assign node29408 = (inp[14]) ? node29414 : node29409;
														assign node29409 = (inp[11]) ? 4'b1111 : node29410;
															assign node29410 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node29414 = (inp[13]) ? 4'b1011 : node29415;
															assign node29415 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node29419 = (inp[14]) ? node29425 : node29420;
														assign node29420 = (inp[13]) ? node29422 : 4'b1010;
															assign node29422 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node29425 = (inp[13]) ? 4'b1110 : node29426;
															assign node29426 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node29430 = (inp[7]) ? node29434 : node29431;
													assign node29431 = (inp[14]) ? 4'b1010 : 4'b1110;
													assign node29434 = (inp[14]) ? node29440 : node29435;
														assign node29435 = (inp[11]) ? node29437 : 4'b1011;
															assign node29437 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node29440 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node29443 = (inp[13]) ? node29467 : node29444;
												assign node29444 = (inp[14]) ? node29456 : node29445;
													assign node29445 = (inp[7]) ? node29453 : node29446;
														assign node29446 = (inp[11]) ? node29450 : node29447;
															assign node29447 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node29450 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29453 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node29456 = (inp[7]) ? node29458 : 4'b1011;
														assign node29458 = (inp[9]) ? node29462 : node29459;
															assign node29459 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node29462 = (inp[0]) ? node29464 : 4'b1111;
																assign node29464 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node29467 = (inp[7]) ? node29475 : node29468;
													assign node29468 = (inp[14]) ? node29472 : node29469;
														assign node29469 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29472 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node29475 = (inp[14]) ? node29477 : 4'b1010;
														assign node29477 = (inp[0]) ? 4'b1110 : 4'b1111;
									assign node29480 = (inp[4]) ? node29574 : node29481;
										assign node29481 = (inp[7]) ? node29517 : node29482;
											assign node29482 = (inp[0]) ? node29500 : node29483;
												assign node29483 = (inp[10]) ? node29491 : node29484;
													assign node29484 = (inp[14]) ? 4'b1111 : node29485;
														assign node29485 = (inp[11]) ? node29487 : 4'b1111;
															assign node29487 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node29491 = (inp[13]) ? node29493 : 4'b1110;
														assign node29493 = (inp[9]) ? 4'b1110 : node29494;
															assign node29494 = (inp[11]) ? 4'b1111 : node29495;
																assign node29495 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node29500 = (inp[10]) ? node29508 : node29501;
													assign node29501 = (inp[13]) ? node29503 : 4'b1110;
														assign node29503 = (inp[14]) ? node29505 : 4'b1111;
															assign node29505 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node29508 = (inp[13]) ? node29510 : 4'b1111;
														assign node29510 = (inp[14]) ? node29514 : node29511;
															assign node29511 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29514 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node29517 = (inp[14]) ? node29545 : node29518;
												assign node29518 = (inp[11]) ? node29524 : node29519;
													assign node29519 = (inp[10]) ? node29521 : 4'b1010;
														assign node29521 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node29524 = (inp[9]) ? node29534 : node29525;
														assign node29525 = (inp[0]) ? 4'b1011 : node29526;
															assign node29526 = (inp[13]) ? node29530 : node29527;
																assign node29527 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node29530 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29534 = (inp[0]) ? node29540 : node29535;
															assign node29535 = (inp[13]) ? node29537 : 4'b1011;
																assign node29537 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node29540 = (inp[10]) ? 4'b1010 : node29541;
																assign node29541 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node29545 = (inp[13]) ? node29567 : node29546;
													assign node29546 = (inp[10]) ? node29552 : node29547;
														assign node29547 = (inp[11]) ? node29549 : 4'b1110;
															assign node29549 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29552 = (inp[9]) ? node29560 : node29553;
															assign node29553 = (inp[11]) ? node29557 : node29554;
																assign node29554 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node29557 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node29560 = (inp[0]) ? node29564 : node29561;
																assign node29561 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node29564 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node29567 = (inp[10]) ? node29571 : node29568;
														assign node29568 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29571 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node29574 = (inp[7]) ? node29620 : node29575;
											assign node29575 = (inp[14]) ? node29601 : node29576;
												assign node29576 = (inp[9]) ? node29586 : node29577;
													assign node29577 = (inp[13]) ? 4'b1100 : node29578;
														assign node29578 = (inp[10]) ? node29582 : node29579;
															assign node29579 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29582 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node29586 = (inp[13]) ? node29594 : node29587;
														assign node29587 = (inp[10]) ? node29591 : node29588;
															assign node29588 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29591 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node29594 = (inp[10]) ? 4'b1101 : node29595;
															assign node29595 = (inp[0]) ? node29597 : 4'b1101;
																assign node29597 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node29601 = (inp[9]) ? node29615 : node29602;
													assign node29602 = (inp[0]) ? node29608 : node29603;
														assign node29603 = (inp[10]) ? 4'b1001 : node29604;
															assign node29604 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node29608 = (inp[10]) ? node29610 : 4'b1001;
															assign node29610 = (inp[11]) ? 4'b1000 : node29611;
																assign node29611 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node29615 = (inp[11]) ? node29617 : 4'b1000;
														assign node29617 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node29620 = (inp[9]) ? node29650 : node29621;
												assign node29621 = (inp[11]) ? node29635 : node29622;
													assign node29622 = (inp[0]) ? node29630 : node29623;
														assign node29623 = (inp[10]) ? 4'b1101 : node29624;
															assign node29624 = (inp[13]) ? 4'b1100 : node29625;
																assign node29625 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node29630 = (inp[14]) ? node29632 : 4'b1100;
															assign node29632 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node29635 = (inp[10]) ? node29639 : node29636;
														assign node29636 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node29639 = (inp[0]) ? node29645 : node29640;
															assign node29640 = (inp[13]) ? 4'b1101 : node29641;
																assign node29641 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node29645 = (inp[13]) ? 4'b1100 : node29646;
																assign node29646 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node29650 = (inp[11]) ? node29660 : node29651;
													assign node29651 = (inp[0]) ? node29655 : node29652;
														assign node29652 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node29655 = (inp[10]) ? node29657 : 4'b1101;
															assign node29657 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node29660 = (inp[14]) ? node29674 : node29661;
														assign node29661 = (inp[13]) ? node29667 : node29662;
															assign node29662 = (inp[0]) ? 4'b1100 : node29663;
																assign node29663 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node29667 = (inp[10]) ? node29671 : node29668;
																assign node29668 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node29671 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node29674 = (inp[13]) ? node29682 : node29675;
															assign node29675 = (inp[10]) ? node29679 : node29676;
																assign node29676 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node29679 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29682 = (inp[0]) ? node29684 : 4'b1101;
																assign node29684 = (inp[10]) ? 4'b1100 : 4'b1101;
							assign node29687 = (inp[5]) ? node30113 : node29688;
								assign node29688 = (inp[12]) ? node29924 : node29689;
									assign node29689 = (inp[4]) ? node29809 : node29690;
										assign node29690 = (inp[7]) ? node29770 : node29691;
											assign node29691 = (inp[9]) ? node29739 : node29692;
												assign node29692 = (inp[11]) ? node29720 : node29693;
													assign node29693 = (inp[14]) ? node29705 : node29694;
														assign node29694 = (inp[13]) ? node29700 : node29695;
															assign node29695 = (inp[10]) ? 4'b1100 : node29696;
																assign node29696 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29700 = (inp[0]) ? 4'b1100 : node29701;
																assign node29701 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node29705 = (inp[13]) ? node29713 : node29706;
															assign node29706 = (inp[0]) ? node29710 : node29707;
																assign node29707 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node29710 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node29713 = (inp[10]) ? node29717 : node29714;
																assign node29714 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node29717 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node29720 = (inp[14]) ? node29728 : node29721;
														assign node29721 = (inp[10]) ? node29723 : 4'b1101;
															assign node29723 = (inp[13]) ? 4'b1100 : node29724;
																assign node29724 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node29728 = (inp[10]) ? node29734 : node29729;
															assign node29729 = (inp[13]) ? 4'b1100 : node29730;
																assign node29730 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29734 = (inp[13]) ? 4'b1101 : node29735;
																assign node29735 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node29739 = (inp[13]) ? node29755 : node29740;
													assign node29740 = (inp[10]) ? node29746 : node29741;
														assign node29741 = (inp[11]) ? 4'b1100 : node29742;
															assign node29742 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node29746 = (inp[0]) ? node29752 : node29747;
															assign node29747 = (inp[14]) ? 4'b1101 : node29748;
																assign node29748 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node29752 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node29755 = (inp[14]) ? node29761 : node29756;
														assign node29756 = (inp[0]) ? node29758 : 4'b1101;
															assign node29758 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node29761 = (inp[11]) ? 4'b1101 : node29762;
															assign node29762 = (inp[0]) ? node29766 : node29763;
																assign node29763 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node29766 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node29770 = (inp[14]) ? node29792 : node29771;
												assign node29771 = (inp[0]) ? node29781 : node29772;
													assign node29772 = (inp[10]) ? node29778 : node29773;
														assign node29773 = (inp[11]) ? 4'b1001 : node29774;
															assign node29774 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node29778 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node29781 = (inp[11]) ? node29789 : node29782;
														assign node29782 = (inp[10]) ? node29786 : node29783;
															assign node29783 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node29786 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node29789 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node29792 = (inp[10]) ? node29802 : node29793;
													assign node29793 = (inp[0]) ? node29799 : node29794;
														assign node29794 = (inp[13]) ? 4'b1100 : node29795;
															assign node29795 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29799 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node29802 = (inp[0]) ? 4'b1100 : node29803;
														assign node29803 = (inp[11]) ? 4'b1101 : node29804;
															assign node29804 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node29809 = (inp[14]) ? node29875 : node29810;
											assign node29810 = (inp[9]) ? node29842 : node29811;
												assign node29811 = (inp[13]) ? node29831 : node29812;
													assign node29812 = (inp[7]) ? node29826 : node29813;
														assign node29813 = (inp[0]) ? node29821 : node29814;
															assign node29814 = (inp[10]) ? node29818 : node29815;
																assign node29815 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node29818 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29821 = (inp[10]) ? node29823 : 4'b1111;
																assign node29823 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node29826 = (inp[0]) ? node29828 : 4'b1110;
															assign node29828 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node29831 = (inp[10]) ? node29833 : 4'b1111;
														assign node29833 = (inp[0]) ? node29839 : node29834;
															assign node29834 = (inp[11]) ? node29836 : 4'b1111;
																assign node29836 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node29839 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node29842 = (inp[0]) ? node29856 : node29843;
													assign node29843 = (inp[7]) ? node29845 : 4'b1110;
														assign node29845 = (inp[10]) ? node29851 : node29846;
															assign node29846 = (inp[13]) ? node29848 : 4'b1111;
																assign node29848 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29851 = (inp[13]) ? node29853 : 4'b1110;
																assign node29853 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node29856 = (inp[11]) ? node29864 : node29857;
														assign node29857 = (inp[10]) ? 4'b1110 : node29858;
															assign node29858 = (inp[13]) ? 4'b1111 : node29859;
																assign node29859 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node29864 = (inp[10]) ? node29870 : node29865;
															assign node29865 = (inp[7]) ? 4'b1110 : node29866;
																assign node29866 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node29870 = (inp[13]) ? node29872 : 4'b1111;
																assign node29872 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node29875 = (inp[7]) ? node29895 : node29876;
												assign node29876 = (inp[0]) ? node29884 : node29877;
													assign node29877 = (inp[10]) ? node29879 : 4'b1010;
														assign node29879 = (inp[13]) ? 4'b1011 : node29880;
															assign node29880 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node29884 = (inp[10]) ? node29890 : node29885;
														assign node29885 = (inp[13]) ? 4'b1011 : node29886;
															assign node29886 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node29890 = (inp[11]) ? 4'b1010 : node29891;
															assign node29891 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node29895 = (inp[9]) ? node29911 : node29896;
													assign node29896 = (inp[13]) ? node29902 : node29897;
														assign node29897 = (inp[11]) ? 4'b1111 : node29898;
															assign node29898 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29902 = (inp[11]) ? node29904 : 4'b1110;
															assign node29904 = (inp[0]) ? node29908 : node29905;
																assign node29905 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node29908 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node29911 = (inp[13]) ? 4'b1111 : node29912;
														assign node29912 = (inp[10]) ? node29918 : node29913;
															assign node29913 = (inp[11]) ? 4'b1110 : node29914;
																assign node29914 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node29918 = (inp[11]) ? node29920 : 4'b1111;
																assign node29920 = (inp[0]) ? 4'b1110 : 4'b1111;
									assign node29924 = (inp[4]) ? node30012 : node29925;
										assign node29925 = (inp[13]) ? node29975 : node29926;
											assign node29926 = (inp[0]) ? node29950 : node29927;
												assign node29927 = (inp[10]) ? node29937 : node29928;
													assign node29928 = (inp[14]) ? node29934 : node29929;
														assign node29929 = (inp[7]) ? 4'b1011 : node29930;
															assign node29930 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29934 = (inp[7]) ? 4'b1110 : 4'b1010;
													assign node29937 = (inp[14]) ? node29945 : node29938;
														assign node29938 = (inp[7]) ? node29942 : node29939;
															assign node29939 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29942 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node29945 = (inp[7]) ? 4'b1111 : node29946;
															assign node29946 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node29950 = (inp[10]) ? node29964 : node29951;
													assign node29951 = (inp[9]) ? node29955 : node29952;
														assign node29952 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node29955 = (inp[14]) ? node29959 : node29956;
															assign node29956 = (inp[7]) ? 4'b1010 : 4'b1110;
															assign node29959 = (inp[7]) ? 4'b1111 : node29960;
																assign node29960 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node29964 = (inp[14]) ? node29972 : node29965;
														assign node29965 = (inp[7]) ? node29969 : node29966;
															assign node29966 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29969 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node29972 = (inp[7]) ? 4'b1110 : 4'b1010;
											assign node29975 = (inp[0]) ? node29995 : node29976;
												assign node29976 = (inp[7]) ? node29984 : node29977;
													assign node29977 = (inp[14]) ? node29981 : node29978;
														assign node29978 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node29981 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node29984 = (inp[14]) ? node29988 : node29985;
														assign node29985 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29988 = (inp[10]) ? node29992 : node29989;
															assign node29989 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29992 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node29995 = (inp[7]) ? node30003 : node29996;
													assign node29996 = (inp[14]) ? node30000 : node29997;
														assign node29997 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node30000 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node30003 = (inp[14]) ? node30007 : node30004;
														assign node30004 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node30007 = (inp[11]) ? 4'b1111 : node30008;
															assign node30008 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node30012 = (inp[13]) ? node30058 : node30013;
											assign node30013 = (inp[10]) ? node30037 : node30014;
												assign node30014 = (inp[11]) ? node30026 : node30015;
													assign node30015 = (inp[0]) ? node30021 : node30016;
														assign node30016 = (inp[7]) ? node30018 : 4'b1100;
															assign node30018 = (inp[14]) ? 4'b1101 : 4'b1001;
														assign node30021 = (inp[9]) ? node30023 : 4'b1100;
															assign node30023 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node30026 = (inp[14]) ? node30034 : node30027;
														assign node30027 = (inp[7]) ? node30031 : node30028;
															assign node30028 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30031 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node30034 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node30037 = (inp[0]) ? node30045 : node30038;
													assign node30038 = (inp[14]) ? node30040 : 4'b1000;
														assign node30040 = (inp[7]) ? node30042 : 4'b1001;
															assign node30042 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30045 = (inp[11]) ? node30053 : node30046;
														assign node30046 = (inp[7]) ? node30050 : node30047;
															assign node30047 = (inp[14]) ? 4'b1000 : 4'b1100;
															assign node30050 = (inp[14]) ? 4'b1101 : 4'b1001;
														assign node30053 = (inp[7]) ? 4'b1100 : node30054;
															assign node30054 = (inp[14]) ? 4'b1000 : 4'b1100;
											assign node30058 = (inp[7]) ? node30092 : node30059;
												assign node30059 = (inp[14]) ? node30077 : node30060;
													assign node30060 = (inp[11]) ? node30062 : 4'b1101;
														assign node30062 = (inp[9]) ? node30070 : node30063;
															assign node30063 = (inp[0]) ? node30067 : node30064;
																assign node30064 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node30067 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node30070 = (inp[10]) ? node30074 : node30071;
																assign node30071 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node30074 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30077 = (inp[10]) ? node30087 : node30078;
														assign node30078 = (inp[9]) ? 4'b1000 : node30079;
															assign node30079 = (inp[0]) ? node30083 : node30080;
																assign node30080 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node30083 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30087 = (inp[9]) ? 4'b1001 : node30088;
															assign node30088 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node30092 = (inp[14]) ? node30106 : node30093;
													assign node30093 = (inp[9]) ? node30099 : node30094;
														assign node30094 = (inp[10]) ? node30096 : 4'b1001;
															assign node30096 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node30099 = (inp[0]) ? node30101 : 4'b1000;
															assign node30101 = (inp[11]) ? node30103 : 4'b1000;
																assign node30103 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node30106 = (inp[0]) ? node30110 : node30107;
														assign node30107 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node30110 = (inp[10]) ? 4'b1100 : 4'b1101;
								assign node30113 = (inp[12]) ? node30309 : node30114;
									assign node30114 = (inp[4]) ? node30192 : node30115;
										assign node30115 = (inp[14]) ? node30151 : node30116;
											assign node30116 = (inp[0]) ? node30134 : node30117;
												assign node30117 = (inp[10]) ? node30125 : node30118;
													assign node30118 = (inp[9]) ? node30120 : 4'b1100;
														assign node30120 = (inp[13]) ? 4'b1101 : node30121;
															assign node30121 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30125 = (inp[9]) ? 4'b1101 : node30126;
														assign node30126 = (inp[13]) ? node30128 : 4'b1101;
															assign node30128 = (inp[11]) ? 4'b1101 : node30129;
																assign node30129 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node30134 = (inp[10]) ? node30146 : node30135;
													assign node30135 = (inp[11]) ? node30141 : node30136;
														assign node30136 = (inp[13]) ? node30138 : 4'b1101;
															assign node30138 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node30141 = (inp[7]) ? 4'b1101 : node30142;
															assign node30142 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node30146 = (inp[11]) ? node30148 : 4'b1100;
														assign node30148 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node30151 = (inp[7]) ? node30173 : node30152;
												assign node30152 = (inp[10]) ? node30162 : node30153;
													assign node30153 = (inp[11]) ? node30159 : node30154;
														assign node30154 = (inp[13]) ? 4'b1101 : node30155;
															assign node30155 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30159 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node30162 = (inp[13]) ? 4'b1100 : node30163;
														assign node30163 = (inp[9]) ? node30165 : 4'b1100;
															assign node30165 = (inp[0]) ? node30169 : node30166;
																assign node30166 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node30169 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node30173 = (inp[0]) ? node30185 : node30174;
													assign node30174 = (inp[10]) ? node30180 : node30175;
														assign node30175 = (inp[11]) ? node30177 : 4'b1000;
															assign node30177 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node30180 = (inp[11]) ? node30182 : 4'b1001;
															assign node30182 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node30185 = (inp[10]) ? 4'b1000 : node30186;
														assign node30186 = (inp[11]) ? node30188 : 4'b1001;
															assign node30188 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node30192 = (inp[14]) ? node30256 : node30193;
											assign node30193 = (inp[7]) ? node30227 : node30194;
												assign node30194 = (inp[13]) ? node30212 : node30195;
													assign node30195 = (inp[11]) ? node30207 : node30196;
														assign node30196 = (inp[9]) ? node30202 : node30197;
															assign node30197 = (inp[0]) ? node30199 : 4'b1011;
																assign node30199 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node30202 = (inp[0]) ? node30204 : 4'b1010;
																assign node30204 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node30207 = (inp[10]) ? 4'b1010 : node30208;
															assign node30208 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node30212 = (inp[11]) ? node30224 : node30213;
														assign node30213 = (inp[9]) ? node30219 : node30214;
															assign node30214 = (inp[10]) ? node30216 : 4'b1010;
																assign node30216 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node30219 = (inp[10]) ? node30221 : 4'b1011;
																assign node30221 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30224 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node30227 = (inp[11]) ? node30235 : node30228;
													assign node30228 = (inp[10]) ? node30232 : node30229;
														assign node30229 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node30232 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node30235 = (inp[9]) ? node30249 : node30236;
														assign node30236 = (inp[0]) ? node30242 : node30237;
															assign node30237 = (inp[13]) ? node30239 : 4'b1110;
																assign node30239 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node30242 = (inp[13]) ? node30246 : node30243;
																assign node30243 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node30246 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node30249 = (inp[13]) ? 4'b1110 : node30250;
															assign node30250 = (inp[10]) ? node30252 : 4'b1110;
																assign node30252 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node30256 = (inp[9]) ? node30282 : node30257;
												assign node30257 = (inp[10]) ? node30267 : node30258;
													assign node30258 = (inp[0]) ? node30264 : node30259;
														assign node30259 = (inp[7]) ? 4'b1110 : node30260;
															assign node30260 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node30264 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node30267 = (inp[13]) ? node30273 : node30268;
														assign node30268 = (inp[0]) ? node30270 : 4'b1110;
															assign node30270 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node30273 = (inp[0]) ? node30277 : node30274;
															assign node30274 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node30277 = (inp[7]) ? 4'b1110 : node30278;
																assign node30278 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node30282 = (inp[13]) ? node30298 : node30283;
													assign node30283 = (inp[10]) ? node30289 : node30284;
														assign node30284 = (inp[0]) ? 4'b1110 : node30285;
															assign node30285 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node30289 = (inp[7]) ? node30293 : node30290;
															assign node30290 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node30293 = (inp[0]) ? node30295 : 4'b1111;
																assign node30295 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node30298 = (inp[0]) ? node30300 : 4'b1111;
														assign node30300 = (inp[10]) ? node30304 : node30301;
															assign node30301 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node30304 = (inp[7]) ? 4'b1110 : node30305;
																assign node30305 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node30309 = (inp[4]) ? node30417 : node30310;
										assign node30310 = (inp[7]) ? node30370 : node30311;
											assign node30311 = (inp[13]) ? node30351 : node30312;
												assign node30312 = (inp[14]) ? node30326 : node30313;
													assign node30313 = (inp[0]) ? node30321 : node30314;
														assign node30314 = (inp[11]) ? node30318 : node30315;
															assign node30315 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node30318 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node30321 = (inp[11]) ? 4'b1110 : node30322;
															assign node30322 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node30326 = (inp[10]) ? node30336 : node30327;
														assign node30327 = (inp[9]) ? node30333 : node30328;
															assign node30328 = (inp[0]) ? 4'b1111 : node30329;
																assign node30329 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node30333 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30336 = (inp[9]) ? node30344 : node30337;
															assign node30337 = (inp[11]) ? node30341 : node30338;
																assign node30338 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30341 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node30344 = (inp[11]) ? node30348 : node30345;
																assign node30345 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30348 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node30351 = (inp[14]) ? node30359 : node30352;
													assign node30352 = (inp[0]) ? node30356 : node30353;
														assign node30353 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node30356 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node30359 = (inp[11]) ? node30361 : 4'b1110;
														assign node30361 = (inp[9]) ? 4'b1110 : node30362;
															assign node30362 = (inp[10]) ? node30366 : node30363;
																assign node30363 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30366 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node30370 = (inp[10]) ? node30398 : node30371;
												assign node30371 = (inp[0]) ? node30381 : node30372;
													assign node30372 = (inp[13]) ? 4'b1111 : node30373;
														assign node30373 = (inp[14]) ? node30377 : node30374;
															assign node30374 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node30377 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node30381 = (inp[13]) ? 4'b1110 : node30382;
														assign node30382 = (inp[9]) ? node30390 : node30383;
															assign node30383 = (inp[11]) ? node30387 : node30384;
																assign node30384 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node30387 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node30390 = (inp[11]) ? node30394 : node30391;
																assign node30391 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node30394 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node30398 = (inp[0]) ? node30408 : node30399;
													assign node30399 = (inp[13]) ? 4'b1110 : node30400;
														assign node30400 = (inp[11]) ? node30404 : node30401;
															assign node30401 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node30404 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node30408 = (inp[13]) ? 4'b1111 : node30409;
														assign node30409 = (inp[11]) ? node30413 : node30410;
															assign node30410 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node30413 = (inp[14]) ? 4'b1111 : 4'b1110;
										assign node30417 = (inp[14]) ? node30477 : node30418;
											assign node30418 = (inp[13]) ? node30440 : node30419;
												assign node30419 = (inp[10]) ? node30421 : 4'b1101;
													assign node30421 = (inp[9]) ? node30427 : node30422;
														assign node30422 = (inp[11]) ? node30424 : 4'b1101;
															assign node30424 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node30427 = (inp[7]) ? node30433 : node30428;
															assign node30428 = (inp[0]) ? node30430 : 4'b1101;
																assign node30430 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node30433 = (inp[11]) ? node30437 : node30434;
																assign node30434 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node30437 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node30440 = (inp[7]) ? node30466 : node30441;
													assign node30441 = (inp[9]) ? node30453 : node30442;
														assign node30442 = (inp[11]) ? node30448 : node30443;
															assign node30443 = (inp[10]) ? 4'b1100 : node30444;
																assign node30444 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30448 = (inp[10]) ? node30450 : 4'b1100;
																assign node30450 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30453 = (inp[11]) ? node30459 : node30454;
															assign node30454 = (inp[10]) ? 4'b1101 : node30455;
																assign node30455 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30459 = (inp[0]) ? node30463 : node30460;
																assign node30460 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node30463 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node30466 = (inp[11]) ? node30472 : node30467;
														assign node30467 = (inp[0]) ? node30469 : 4'b1100;
															assign node30469 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30472 = (inp[10]) ? 4'b1101 : node30473;
															assign node30473 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node30477 = (inp[10]) ? node30489 : node30478;
												assign node30478 = (inp[0]) ? node30484 : node30479;
													assign node30479 = (inp[13]) ? 4'b1100 : node30480;
														assign node30480 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node30484 = (inp[13]) ? 4'b1101 : node30485;
														assign node30485 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node30489 = (inp[0]) ? node30495 : node30490;
													assign node30490 = (inp[13]) ? 4'b1101 : node30491;
														assign node30491 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30495 = (inp[11]) ? 4'b1100 : node30496;
														assign node30496 = (inp[13]) ? 4'b1100 : 4'b1101;
					assign node30500 = (inp[1]) ? node32064 : node30501;
						assign node30501 = (inp[14]) ? node31269 : node30502;
							assign node30502 = (inp[7]) ? node30896 : node30503;
								assign node30503 = (inp[4]) ? node30677 : node30504;
									assign node30504 = (inp[12]) ? node30606 : node30505;
										assign node30505 = (inp[9]) ? node30553 : node30506;
											assign node30506 = (inp[13]) ? node30528 : node30507;
												assign node30507 = (inp[11]) ? node30515 : node30508;
													assign node30508 = (inp[0]) ? node30512 : node30509;
														assign node30509 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node30512 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node30515 = (inp[15]) ? node30521 : node30516;
														assign node30516 = (inp[0]) ? node30518 : 4'b1100;
															assign node30518 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node30521 = (inp[0]) ? node30525 : node30522;
															assign node30522 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node30525 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node30528 = (inp[10]) ? node30538 : node30529;
													assign node30529 = (inp[0]) ? node30531 : 4'b1101;
														assign node30531 = (inp[11]) ? node30535 : node30532;
															assign node30532 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node30535 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node30538 = (inp[15]) ? node30546 : node30539;
														assign node30539 = (inp[11]) ? node30543 : node30540;
															assign node30540 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node30543 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node30546 = (inp[11]) ? node30550 : node30547;
															assign node30547 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30550 = (inp[5]) ? 4'b1100 : 4'b1101;
											assign node30553 = (inp[15]) ? node30581 : node30554;
												assign node30554 = (inp[13]) ? node30568 : node30555;
													assign node30555 = (inp[5]) ? 4'b1100 : node30556;
														assign node30556 = (inp[11]) ? node30562 : node30557;
															assign node30557 = (inp[0]) ? node30559 : 4'b1100;
																assign node30559 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node30562 = (inp[10]) ? node30564 : 4'b1100;
																assign node30564 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30568 = (inp[11]) ? node30576 : node30569;
														assign node30569 = (inp[10]) ? node30573 : node30570;
															assign node30570 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30573 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30576 = (inp[10]) ? 4'b1100 : node30577;
															assign node30577 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node30581 = (inp[10]) ? node30593 : node30582;
													assign node30582 = (inp[0]) ? node30588 : node30583;
														assign node30583 = (inp[11]) ? 4'b1100 : node30584;
															assign node30584 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node30588 = (inp[13]) ? node30590 : 4'b1101;
															assign node30590 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node30593 = (inp[0]) ? node30599 : node30594;
														assign node30594 = (inp[13]) ? node30596 : 4'b1101;
															assign node30596 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30599 = (inp[5]) ? node30601 : 4'b1101;
															assign node30601 = (inp[11]) ? 4'b1100 : node30602;
																assign node30602 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node30606 = (inp[5]) ? node30644 : node30607;
											assign node30607 = (inp[10]) ? node30627 : node30608;
												assign node30608 = (inp[0]) ? node30618 : node30609;
													assign node30609 = (inp[13]) ? node30611 : 4'b1110;
														assign node30611 = (inp[15]) ? node30615 : node30612;
															assign node30612 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node30615 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node30618 = (inp[13]) ? node30620 : 4'b1111;
														assign node30620 = (inp[15]) ? node30624 : node30621;
															assign node30621 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node30624 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node30627 = (inp[0]) ? node30637 : node30628;
													assign node30628 = (inp[13]) ? node30630 : 4'b1111;
														assign node30630 = (inp[11]) ? node30634 : node30631;
															assign node30631 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node30634 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node30637 = (inp[13]) ? node30639 : 4'b1110;
														assign node30639 = (inp[9]) ? node30641 : 4'b1111;
															assign node30641 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node30644 = (inp[0]) ? node30662 : node30645;
												assign node30645 = (inp[10]) ? node30655 : node30646;
													assign node30646 = (inp[13]) ? node30648 : 4'b1110;
														assign node30648 = (inp[9]) ? 4'b1110 : node30649;
															assign node30649 = (inp[11]) ? node30651 : 4'b1111;
																assign node30651 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node30655 = (inp[13]) ? node30657 : 4'b1111;
														assign node30657 = (inp[9]) ? 4'b1110 : node30658;
															assign node30658 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node30662 = (inp[10]) ? node30668 : node30663;
													assign node30663 = (inp[13]) ? node30665 : 4'b1111;
														assign node30665 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node30668 = (inp[13]) ? node30670 : 4'b1110;
														assign node30670 = (inp[11]) ? node30674 : node30671;
															assign node30671 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node30674 = (inp[15]) ? 4'b1110 : 4'b1111;
									assign node30677 = (inp[12]) ? node30769 : node30678;
										assign node30678 = (inp[15]) ? node30722 : node30679;
											assign node30679 = (inp[10]) ? node30703 : node30680;
												assign node30680 = (inp[5]) ? node30692 : node30681;
													assign node30681 = (inp[9]) ? 4'b1111 : node30682;
														assign node30682 = (inp[11]) ? node30686 : node30683;
															assign node30683 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node30686 = (inp[13]) ? node30688 : 4'b1110;
																assign node30688 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node30692 = (inp[0]) ? node30698 : node30693;
														assign node30693 = (inp[13]) ? 4'b1110 : node30694;
															assign node30694 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30698 = (inp[11]) ? 4'b1111 : node30699;
															assign node30699 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node30703 = (inp[13]) ? node30715 : node30704;
													assign node30704 = (inp[0]) ? node30710 : node30705;
														assign node30705 = (inp[11]) ? node30707 : 4'b1110;
															assign node30707 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node30710 = (inp[11]) ? node30712 : 4'b1111;
															assign node30712 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node30715 = (inp[0]) ? 4'b1110 : node30716;
														assign node30716 = (inp[5]) ? 4'b1111 : node30717;
															assign node30717 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node30722 = (inp[5]) ? node30744 : node30723;
												assign node30723 = (inp[0]) ? node30733 : node30724;
													assign node30724 = (inp[11]) ? node30730 : node30725;
														assign node30725 = (inp[10]) ? 4'b1111 : node30726;
															assign node30726 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node30730 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node30733 = (inp[10]) ? node30739 : node30734;
														assign node30734 = (inp[13]) ? node30736 : 4'b1110;
															assign node30736 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30739 = (inp[13]) ? node30741 : 4'b1111;
															assign node30741 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node30744 = (inp[11]) ? node30758 : node30745;
													assign node30745 = (inp[9]) ? 4'b1011 : node30746;
														assign node30746 = (inp[0]) ? node30752 : node30747;
															assign node30747 = (inp[10]) ? node30749 : 4'b1011;
																assign node30749 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node30752 = (inp[13]) ? node30754 : 4'b1010;
																assign node30754 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node30758 = (inp[13]) ? node30764 : node30759;
														assign node30759 = (inp[10]) ? 4'b1010 : node30760;
															assign node30760 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30764 = (inp[10]) ? node30766 : 4'b1010;
															assign node30766 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node30769 = (inp[5]) ? node30823 : node30770;
											assign node30770 = (inp[15]) ? node30800 : node30771;
												assign node30771 = (inp[9]) ? node30781 : node30772;
													assign node30772 = (inp[13]) ? 4'b1001 : node30773;
														assign node30773 = (inp[10]) ? node30777 : node30774;
															assign node30774 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30777 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node30781 = (inp[0]) ? node30791 : node30782;
														assign node30782 = (inp[10]) ? node30786 : node30783;
															assign node30783 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node30786 = (inp[13]) ? 4'b1001 : node30787;
																assign node30787 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node30791 = (inp[10]) ? node30797 : node30792;
															assign node30792 = (inp[13]) ? 4'b1001 : node30793;
																assign node30793 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30797 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node30800 = (inp[11]) ? node30808 : node30801;
													assign node30801 = (inp[0]) ? node30805 : node30802;
														assign node30802 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node30805 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node30808 = (inp[10]) ? node30816 : node30809;
														assign node30809 = (inp[0]) ? node30813 : node30810;
															assign node30810 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node30813 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node30816 = (inp[0]) ? node30820 : node30817;
															assign node30817 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node30820 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node30823 = (inp[13]) ? node30851 : node30824;
												assign node30824 = (inp[15]) ? node30842 : node30825;
													assign node30825 = (inp[9]) ? node30833 : node30826;
														assign node30826 = (inp[0]) ? node30830 : node30827;
															assign node30827 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node30830 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node30833 = (inp[11]) ? node30835 : 4'b1101;
															assign node30835 = (inp[10]) ? node30839 : node30836;
																assign node30836 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node30839 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30842 = (inp[11]) ? 4'b1101 : node30843;
														assign node30843 = (inp[0]) ? node30847 : node30844;
															assign node30844 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node30847 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node30851 = (inp[9]) ? node30871 : node30852;
													assign node30852 = (inp[11]) ? node30862 : node30853;
														assign node30853 = (inp[15]) ? node30855 : 4'b1100;
															assign node30855 = (inp[0]) ? node30859 : node30856;
																assign node30856 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30859 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node30862 = (inp[15]) ? 4'b1101 : node30863;
															assign node30863 = (inp[0]) ? node30867 : node30864;
																assign node30864 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30867 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node30871 = (inp[15]) ? node30881 : node30872;
														assign node30872 = (inp[11]) ? node30874 : 4'b1101;
															assign node30874 = (inp[0]) ? node30878 : node30875;
																assign node30875 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30878 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node30881 = (inp[11]) ? node30889 : node30882;
															assign node30882 = (inp[0]) ? node30886 : node30883;
																assign node30883 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30886 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node30889 = (inp[10]) ? node30893 : node30890;
																assign node30890 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node30893 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node30896 = (inp[4]) ? node31084 : node30897;
									assign node30897 = (inp[12]) ? node30997 : node30898;
										assign node30898 = (inp[15]) ? node30956 : node30899;
											assign node30899 = (inp[5]) ? node30931 : node30900;
												assign node30900 = (inp[9]) ? node30916 : node30901;
													assign node30901 = (inp[0]) ? node30907 : node30902;
														assign node30902 = (inp[10]) ? node30904 : 4'b1100;
															assign node30904 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node30907 = (inp[10]) ? node30913 : node30908;
															assign node30908 = (inp[11]) ? node30910 : 4'b1101;
																assign node30910 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node30913 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30916 = (inp[11]) ? node30922 : node30917;
														assign node30917 = (inp[10]) ? 4'b1101 : node30918;
															assign node30918 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node30922 = (inp[13]) ? node30924 : 4'b1100;
															assign node30924 = (inp[0]) ? node30928 : node30925;
																assign node30925 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node30928 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node30931 = (inp[9]) ? node30941 : node30932;
													assign node30932 = (inp[10]) ? node30938 : node30933;
														assign node30933 = (inp[13]) ? node30935 : 4'b1000;
															assign node30935 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node30938 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node30941 = (inp[0]) ? node30949 : node30942;
														assign node30942 = (inp[10]) ? node30944 : 4'b1000;
															assign node30944 = (inp[13]) ? 4'b1001 : node30945;
																assign node30945 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node30949 = (inp[10]) ? node30951 : 4'b1001;
															assign node30951 = (inp[11]) ? 4'b1000 : node30952;
																assign node30952 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node30956 = (inp[5]) ? node30980 : node30957;
												assign node30957 = (inp[0]) ? node30969 : node30958;
													assign node30958 = (inp[10]) ? node30964 : node30959;
														assign node30959 = (inp[11]) ? node30961 : 4'b1000;
															assign node30961 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node30964 = (inp[11]) ? node30966 : 4'b1001;
															assign node30966 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node30969 = (inp[10]) ? node30975 : node30970;
														assign node30970 = (inp[13]) ? 4'b1001 : node30971;
															assign node30971 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30975 = (inp[13]) ? 4'b1000 : node30976;
															assign node30976 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node30980 = (inp[0]) ? node30986 : node30981;
													assign node30981 = (inp[10]) ? node30983 : 4'b1101;
														assign node30983 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node30986 = (inp[13]) ? node30994 : node30987;
														assign node30987 = (inp[11]) ? node30991 : node30988;
															assign node30988 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node30991 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node30994 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node30997 = (inp[15]) ? node31037 : node30998;
											assign node30998 = (inp[5]) ? node31020 : node30999;
												assign node30999 = (inp[0]) ? node31011 : node31000;
													assign node31000 = (inp[10]) ? node31006 : node31001;
														assign node31001 = (inp[13]) ? 4'b1111 : node31002;
															assign node31002 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node31006 = (inp[11]) ? 4'b1110 : node31007;
															assign node31007 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31011 = (inp[10]) ? node31015 : node31012;
														assign node31012 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node31015 = (inp[11]) ? 4'b1111 : node31016;
															assign node31016 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node31020 = (inp[10]) ? node31032 : node31021;
													assign node31021 = (inp[0]) ? node31027 : node31022;
														assign node31022 = (inp[13]) ? node31024 : 4'b1010;
															assign node31024 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node31027 = (inp[13]) ? node31029 : 4'b1011;
															assign node31029 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node31032 = (inp[0]) ? node31034 : 4'b1011;
														assign node31034 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node31037 = (inp[5]) ? node31067 : node31038;
												assign node31038 = (inp[11]) ? node31054 : node31039;
													assign node31039 = (inp[13]) ? 4'b1011 : node31040;
														assign node31040 = (inp[9]) ? node31048 : node31041;
															assign node31041 = (inp[0]) ? node31045 : node31042;
																assign node31042 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node31045 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31048 = (inp[10]) ? node31050 : 4'b1011;
																assign node31050 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node31054 = (inp[9]) ? node31060 : node31055;
														assign node31055 = (inp[0]) ? 4'b1010 : node31056;
															assign node31056 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31060 = (inp[10]) ? node31064 : node31061;
															assign node31061 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31064 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node31067 = (inp[11]) ? node31077 : node31068;
													assign node31068 = (inp[0]) ? 4'b1110 : node31069;
														assign node31069 = (inp[13]) ? node31073 : node31070;
															assign node31070 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31073 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node31077 = (inp[10]) ? node31081 : node31078;
														assign node31078 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31081 = (inp[0]) ? 4'b1110 : 4'b1111;
									assign node31084 = (inp[12]) ? node31190 : node31085;
										assign node31085 = (inp[15]) ? node31147 : node31086;
											assign node31086 = (inp[5]) ? node31104 : node31087;
												assign node31087 = (inp[11]) ? node31095 : node31088;
													assign node31088 = (inp[0]) ? node31092 : node31089;
														assign node31089 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31092 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31095 = (inp[0]) ? node31097 : 4'b1110;
														assign node31097 = (inp[9]) ? node31099 : 4'b1110;
															assign node31099 = (inp[10]) ? 4'b1111 : node31100;
																assign node31100 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node31104 = (inp[9]) ? node31132 : node31105;
													assign node31105 = (inp[13]) ? node31119 : node31106;
														assign node31106 = (inp[11]) ? node31112 : node31107;
															assign node31107 = (inp[10]) ? 4'b1010 : node31108;
																assign node31108 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node31112 = (inp[10]) ? node31116 : node31113;
																assign node31113 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node31116 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31119 = (inp[11]) ? node31127 : node31120;
															assign node31120 = (inp[10]) ? node31124 : node31121;
																assign node31121 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node31124 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node31127 = (inp[10]) ? node31129 : 4'b1011;
																assign node31129 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node31132 = (inp[11]) ? node31138 : node31133;
														assign node31133 = (inp[0]) ? 4'b1010 : node31134;
															assign node31134 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31138 = (inp[13]) ? 4'b1010 : node31139;
															assign node31139 = (inp[0]) ? node31143 : node31140;
																assign node31140 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node31143 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node31147 = (inp[10]) ? node31171 : node31148;
												assign node31148 = (inp[0]) ? node31160 : node31149;
													assign node31149 = (inp[5]) ? node31155 : node31150;
														assign node31150 = (inp[11]) ? node31152 : 4'b1111;
															assign node31152 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node31155 = (inp[11]) ? 4'b1111 : node31156;
															assign node31156 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31160 = (inp[11]) ? node31166 : node31161;
														assign node31161 = (inp[5]) ? node31163 : 4'b1110;
															assign node31163 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node31166 = (inp[5]) ? 4'b1110 : node31167;
															assign node31167 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node31171 = (inp[0]) ? node31177 : node31172;
													assign node31172 = (inp[5]) ? node31174 : 4'b1110;
														assign node31174 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node31177 = (inp[9]) ? node31179 : 4'b1111;
														assign node31179 = (inp[5]) ? node31185 : node31180;
															assign node31180 = (inp[11]) ? node31182 : 4'b1111;
																assign node31182 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31185 = (inp[13]) ? node31187 : 4'b1111;
																assign node31187 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node31190 = (inp[5]) ? node31234 : node31191;
											assign node31191 = (inp[15]) ? node31213 : node31192;
												assign node31192 = (inp[10]) ? node31202 : node31193;
													assign node31193 = (inp[0]) ? node31197 : node31194;
														assign node31194 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node31197 = (inp[13]) ? node31199 : 4'b1101;
															assign node31199 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node31202 = (inp[0]) ? node31208 : node31203;
														assign node31203 = (inp[11]) ? node31205 : 4'b1101;
															assign node31205 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node31208 = (inp[13]) ? node31210 : 4'b1100;
															assign node31210 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node31213 = (inp[10]) ? node31223 : node31214;
													assign node31214 = (inp[0]) ? node31218 : node31215;
														assign node31215 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node31218 = (inp[13]) ? 4'b1001 : node31219;
															assign node31219 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node31223 = (inp[0]) ? node31229 : node31224;
														assign node31224 = (inp[11]) ? node31226 : 4'b1001;
															assign node31226 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node31229 = (inp[11]) ? node31231 : 4'b1000;
															assign node31231 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node31234 = (inp[10]) ? node31252 : node31235;
												assign node31235 = (inp[0]) ? node31243 : node31236;
													assign node31236 = (inp[11]) ? 4'b1100 : node31237;
														assign node31237 = (inp[13]) ? 4'b1101 : node31238;
															assign node31238 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node31243 = (inp[11]) ? 4'b1101 : node31244;
														assign node31244 = (inp[13]) ? node31248 : node31245;
															assign node31245 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node31248 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node31252 = (inp[0]) ? node31260 : node31253;
													assign node31253 = (inp[11]) ? 4'b1101 : node31254;
														assign node31254 = (inp[13]) ? 4'b1100 : node31255;
															assign node31255 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node31260 = (inp[11]) ? 4'b1100 : node31261;
														assign node31261 = (inp[15]) ? node31265 : node31262;
															assign node31262 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node31265 = (inp[13]) ? 4'b1101 : 4'b1100;
							assign node31269 = (inp[7]) ? node31705 : node31270;
								assign node31270 = (inp[4]) ? node31462 : node31271;
									assign node31271 = (inp[12]) ? node31375 : node31272;
										assign node31272 = (inp[5]) ? node31328 : node31273;
											assign node31273 = (inp[15]) ? node31297 : node31274;
												assign node31274 = (inp[10]) ? node31286 : node31275;
													assign node31275 = (inp[0]) ? node31281 : node31276;
														assign node31276 = (inp[13]) ? node31278 : 4'b1100;
															assign node31278 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node31281 = (inp[11]) ? 4'b1101 : node31282;
															assign node31282 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node31286 = (inp[0]) ? node31292 : node31287;
														assign node31287 = (inp[13]) ? node31289 : 4'b1101;
															assign node31289 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node31292 = (inp[13]) ? node31294 : 4'b1100;
															assign node31294 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node31297 = (inp[9]) ? node31315 : node31298;
													assign node31298 = (inp[0]) ? node31306 : node31299;
														assign node31299 = (inp[10]) ? node31301 : 4'b1100;
															assign node31301 = (inp[11]) ? node31303 : 4'b1101;
																assign node31303 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node31306 = (inp[10]) ? node31312 : node31307;
															assign node31307 = (inp[11]) ? node31309 : 4'b1101;
																assign node31309 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node31312 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node31315 = (inp[10]) ? node31321 : node31316;
														assign node31316 = (inp[0]) ? 4'b1101 : node31317;
															assign node31317 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node31321 = (inp[0]) ? node31323 : 4'b1101;
															assign node31323 = (inp[13]) ? node31325 : 4'b1100;
																assign node31325 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node31328 = (inp[15]) ? node31354 : node31329;
												assign node31329 = (inp[11]) ? node31345 : node31330;
													assign node31330 = (inp[13]) ? node31338 : node31331;
														assign node31331 = (inp[0]) ? node31335 : node31332;
															assign node31332 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31335 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node31338 = (inp[0]) ? node31342 : node31339;
															assign node31339 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31342 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node31345 = (inp[13]) ? 4'b1001 : node31346;
														assign node31346 = (inp[9]) ? node31350 : node31347;
															assign node31347 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node31350 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node31354 = (inp[9]) ? node31370 : node31355;
													assign node31355 = (inp[0]) ? node31361 : node31356;
														assign node31356 = (inp[10]) ? node31358 : 4'b1100;
															assign node31358 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node31361 = (inp[11]) ? node31367 : node31362;
															assign node31362 = (inp[10]) ? node31364 : 4'b1100;
																assign node31364 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node31367 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node31370 = (inp[0]) ? node31372 : 4'b1100;
														assign node31372 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node31375 = (inp[15]) ? node31425 : node31376;
											assign node31376 = (inp[5]) ? node31394 : node31377;
												assign node31377 = (inp[0]) ? node31389 : node31378;
													assign node31378 = (inp[10]) ? node31384 : node31379;
														assign node31379 = (inp[13]) ? node31381 : 4'b1110;
															assign node31381 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node31384 = (inp[13]) ? node31386 : 4'b1111;
															assign node31386 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node31389 = (inp[10]) ? 4'b1110 : node31390;
														assign node31390 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node31394 = (inp[9]) ? node31412 : node31395;
													assign node31395 = (inp[13]) ? node31405 : node31396;
														assign node31396 = (inp[11]) ? node31398 : 4'b1110;
															assign node31398 = (inp[0]) ? node31402 : node31399;
																assign node31399 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node31402 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31405 = (inp[11]) ? 4'b1110 : node31406;
															assign node31406 = (inp[10]) ? 4'b1110 : node31407;
																assign node31407 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node31412 = (inp[0]) ? node31422 : node31413;
														assign node31413 = (inp[10]) ? node31417 : node31414;
															assign node31414 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31417 = (inp[13]) ? 4'b1110 : node31418;
																assign node31418 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node31422 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node31425 = (inp[5]) ? node31439 : node31426;
												assign node31426 = (inp[0]) ? node31432 : node31427;
													assign node31427 = (inp[10]) ? node31429 : 4'b1010;
														assign node31429 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node31432 = (inp[10]) ? node31434 : 4'b1011;
														assign node31434 = (inp[13]) ? 4'b1010 : node31435;
															assign node31435 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node31439 = (inp[13]) ? node31455 : node31440;
													assign node31440 = (inp[9]) ? node31446 : node31441;
														assign node31441 = (inp[0]) ? 4'b1111 : node31442;
															assign node31442 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31446 = (inp[0]) ? 4'b1110 : node31447;
															assign node31447 = (inp[10]) ? node31451 : node31448;
																assign node31448 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node31451 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node31455 = (inp[10]) ? node31459 : node31456;
														assign node31456 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31459 = (inp[0]) ? 4'b1110 : 4'b1111;
									assign node31462 = (inp[12]) ? node31554 : node31463;
										assign node31463 = (inp[0]) ? node31507 : node31464;
											assign node31464 = (inp[15]) ? node31484 : node31465;
												assign node31465 = (inp[5]) ? node31477 : node31466;
													assign node31466 = (inp[10]) ? node31472 : node31467;
														assign node31467 = (inp[13]) ? node31469 : 4'b1111;
															assign node31469 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node31472 = (inp[11]) ? 4'b1110 : node31473;
															assign node31473 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node31477 = (inp[10]) ? 4'b1011 : node31478;
														assign node31478 = (inp[13]) ? node31480 : 4'b1010;
															assign node31480 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node31484 = (inp[5]) ? node31496 : node31485;
													assign node31485 = (inp[10]) ? node31491 : node31486;
														assign node31486 = (inp[13]) ? 4'b1011 : node31487;
															assign node31487 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node31491 = (inp[11]) ? 4'b1010 : node31492;
															assign node31492 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node31496 = (inp[10]) ? node31502 : node31497;
														assign node31497 = (inp[11]) ? node31499 : 4'b1110;
															assign node31499 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node31502 = (inp[13]) ? node31504 : 4'b1111;
															assign node31504 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node31507 = (inp[11]) ? node31535 : node31508;
												assign node31508 = (inp[10]) ? node31526 : node31509;
													assign node31509 = (inp[13]) ? node31515 : node31510;
														assign node31510 = (inp[5]) ? node31512 : 4'b1011;
															assign node31512 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node31515 = (inp[9]) ? node31521 : node31516;
															assign node31516 = (inp[15]) ? node31518 : 4'b1111;
																assign node31518 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node31521 = (inp[15]) ? 4'b1010 : node31522;
																assign node31522 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node31526 = (inp[15]) ? 4'b1110 : node31527;
														assign node31527 = (inp[5]) ? node31531 : node31528;
															assign node31528 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node31531 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node31535 = (inp[10]) ? node31545 : node31536;
													assign node31536 = (inp[5]) ? node31540 : node31537;
														assign node31537 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node31540 = (inp[15]) ? node31542 : 4'b1011;
															assign node31542 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31545 = (inp[5]) ? node31549 : node31546;
														assign node31546 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node31549 = (inp[15]) ? node31551 : 4'b1010;
															assign node31551 = (inp[13]) ? 4'b1111 : 4'b1110;
										assign node31554 = (inp[13]) ? node31634 : node31555;
											assign node31555 = (inp[9]) ? node31591 : node31556;
												assign node31556 = (inp[10]) ? node31576 : node31557;
													assign node31557 = (inp[15]) ? node31571 : node31558;
														assign node31558 = (inp[5]) ? node31564 : node31559;
															assign node31559 = (inp[0]) ? 4'b1100 : node31560;
																assign node31560 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node31564 = (inp[11]) ? node31568 : node31565;
																assign node31565 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node31568 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node31571 = (inp[5]) ? 4'b1101 : node31572;
															assign node31572 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node31576 = (inp[5]) ? node31582 : node31577;
														assign node31577 = (inp[15]) ? node31579 : 4'b1101;
															assign node31579 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node31582 = (inp[15]) ? node31586 : node31583;
															assign node31583 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node31586 = (inp[0]) ? 4'b1101 : node31587;
																assign node31587 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node31591 = (inp[11]) ? node31615 : node31592;
													assign node31592 = (inp[10]) ? node31604 : node31593;
														assign node31593 = (inp[5]) ? node31599 : node31594;
															assign node31594 = (inp[0]) ? node31596 : 4'b1100;
																assign node31596 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node31599 = (inp[15]) ? node31601 : 4'b1001;
																assign node31601 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31604 = (inp[0]) ? node31612 : node31605;
															assign node31605 = (inp[5]) ? node31609 : node31606;
																assign node31606 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node31609 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node31612 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node31615 = (inp[0]) ? node31627 : node31616;
														assign node31616 = (inp[5]) ? node31622 : node31617;
															assign node31617 = (inp[15]) ? 4'b1001 : node31618;
																assign node31618 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node31622 = (inp[10]) ? 4'b1101 : node31623;
																assign node31623 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node31627 = (inp[15]) ? node31631 : node31628;
															assign node31628 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node31631 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node31634 = (inp[11]) ? node31678 : node31635;
												assign node31635 = (inp[9]) ? node31663 : node31636;
													assign node31636 = (inp[10]) ? node31648 : node31637;
														assign node31637 = (inp[5]) ? node31643 : node31638;
															assign node31638 = (inp[0]) ? node31640 : 4'b1000;
																assign node31640 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node31643 = (inp[15]) ? 4'b1100 : node31644;
																assign node31644 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node31648 = (inp[0]) ? node31656 : node31649;
															assign node31649 = (inp[5]) ? node31653 : node31650;
																assign node31650 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node31653 = (inp[15]) ? 4'b1101 : 4'b1000;
															assign node31656 = (inp[5]) ? node31660 : node31657;
																assign node31657 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node31660 = (inp[15]) ? 4'b1100 : 4'b1001;
													assign node31663 = (inp[0]) ? node31665 : 4'b1100;
														assign node31665 = (inp[10]) ? node31673 : node31666;
															assign node31666 = (inp[15]) ? node31670 : node31667;
																assign node31667 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node31670 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node31673 = (inp[5]) ? node31675 : 4'b1100;
																assign node31675 = (inp[15]) ? 4'b1100 : 4'b1001;
												assign node31678 = (inp[15]) ? node31690 : node31679;
													assign node31679 = (inp[5]) ? node31687 : node31680;
														assign node31680 = (inp[10]) ? node31684 : node31681;
															assign node31681 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node31684 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31687 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node31690 = (inp[5]) ? node31696 : node31691;
														assign node31691 = (inp[10]) ? node31693 : 4'b1000;
															assign node31693 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node31696 = (inp[9]) ? 4'b1100 : node31697;
															assign node31697 = (inp[0]) ? node31701 : node31698;
																assign node31698 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node31701 = (inp[10]) ? 4'b1100 : 4'b1101;
								assign node31705 = (inp[4]) ? node31905 : node31706;
									assign node31706 = (inp[12]) ? node31818 : node31707;
										assign node31707 = (inp[5]) ? node31755 : node31708;
											assign node31708 = (inp[0]) ? node31738 : node31709;
												assign node31709 = (inp[10]) ? node31721 : node31710;
													assign node31710 = (inp[11]) ? 4'b1100 : node31711;
														assign node31711 = (inp[9]) ? 4'b1100 : node31712;
															assign node31712 = (inp[15]) ? node31716 : node31713;
																assign node31713 = (inp[13]) ? 4'b1101 : 4'b1100;
																assign node31716 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node31721 = (inp[11]) ? 4'b1101 : node31722;
														assign node31722 = (inp[9]) ? node31730 : node31723;
															assign node31723 = (inp[15]) ? node31727 : node31724;
																assign node31724 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node31727 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node31730 = (inp[15]) ? node31734 : node31731;
																assign node31731 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node31734 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node31738 = (inp[10]) ? node31748 : node31739;
													assign node31739 = (inp[11]) ? 4'b1101 : node31740;
														assign node31740 = (inp[13]) ? node31744 : node31741;
															assign node31741 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node31744 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node31748 = (inp[11]) ? 4'b1100 : node31749;
														assign node31749 = (inp[13]) ? node31751 : 4'b1101;
															assign node31751 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node31755 = (inp[15]) ? node31787 : node31756;
												assign node31756 = (inp[11]) ? node31774 : node31757;
													assign node31757 = (inp[13]) ? node31767 : node31758;
														assign node31758 = (inp[9]) ? 4'b1100 : node31759;
															assign node31759 = (inp[0]) ? node31763 : node31760;
																assign node31760 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node31763 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node31767 = (inp[0]) ? node31771 : node31768;
															assign node31768 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node31771 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node31774 = (inp[0]) ? node31782 : node31775;
														assign node31775 = (inp[13]) ? node31779 : node31776;
															assign node31776 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node31779 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node31782 = (inp[13]) ? 4'b1101 : node31783;
															assign node31783 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node31787 = (inp[9]) ? node31807 : node31788;
													assign node31788 = (inp[10]) ? node31796 : node31789;
														assign node31789 = (inp[11]) ? node31791 : 4'b1000;
															assign node31791 = (inp[13]) ? 4'b1001 : node31792;
																assign node31792 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node31796 = (inp[0]) ? node31802 : node31797;
															assign node31797 = (inp[11]) ? node31799 : 4'b1001;
																assign node31799 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node31802 = (inp[13]) ? node31804 : 4'b1000;
																assign node31804 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node31807 = (inp[13]) ? node31815 : node31808;
														assign node31808 = (inp[0]) ? node31812 : node31809;
															assign node31809 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node31812 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node31815 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node31818 = (inp[15]) ? node31860 : node31819;
											assign node31819 = (inp[5]) ? node31837 : node31820;
												assign node31820 = (inp[10]) ? node31828 : node31821;
													assign node31821 = (inp[0]) ? node31823 : 4'b1011;
														assign node31823 = (inp[13]) ? node31825 : 4'b1010;
															assign node31825 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node31828 = (inp[0]) ? node31834 : node31829;
														assign node31829 = (inp[11]) ? 4'b1010 : node31830;
															assign node31830 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node31834 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node31837 = (inp[9]) ? node31851 : node31838;
													assign node31838 = (inp[0]) ? node31844 : node31839;
														assign node31839 = (inp[10]) ? 4'b1111 : node31840;
															assign node31840 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node31844 = (inp[11]) ? node31848 : node31845;
															assign node31845 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31848 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node31851 = (inp[0]) ? 4'b1110 : node31852;
														assign node31852 = (inp[10]) ? node31854 : 4'b1110;
															assign node31854 = (inp[11]) ? 4'b1111 : node31855;
																assign node31855 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node31860 = (inp[13]) ? node31888 : node31861;
												assign node31861 = (inp[5]) ? node31869 : node31862;
													assign node31862 = (inp[0]) ? node31866 : node31863;
														assign node31863 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31866 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31869 = (inp[9]) ? node31875 : node31870;
														assign node31870 = (inp[11]) ? node31872 : 4'b1111;
															assign node31872 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31875 = (inp[11]) ? node31883 : node31876;
															assign node31876 = (inp[0]) ? node31880 : node31877;
																assign node31877 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node31880 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31883 = (inp[10]) ? node31885 : 4'b1111;
																assign node31885 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node31888 = (inp[0]) ? node31900 : node31889;
													assign node31889 = (inp[10]) ? node31895 : node31890;
														assign node31890 = (inp[5]) ? 4'b1110 : node31891;
															assign node31891 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node31895 = (inp[5]) ? 4'b1111 : node31896;
															assign node31896 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node31900 = (inp[10]) ? 4'b1110 : node31901;
														assign node31901 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node31905 = (inp[12]) ? node32009 : node31906;
										assign node31906 = (inp[5]) ? node31962 : node31907;
											assign node31907 = (inp[9]) ? node31931 : node31908;
												assign node31908 = (inp[13]) ? node31918 : node31909;
													assign node31909 = (inp[15]) ? 4'b1111 : node31910;
														assign node31910 = (inp[11]) ? 4'b1110 : node31911;
															assign node31911 = (inp[10]) ? node31913 : 4'b1111;
																assign node31913 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node31918 = (inp[11]) ? node31926 : node31919;
														assign node31919 = (inp[15]) ? node31921 : 4'b1110;
															assign node31921 = (inp[0]) ? 4'b1111 : node31922;
																assign node31922 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node31926 = (inp[10]) ? node31928 : 4'b1110;
															assign node31928 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node31931 = (inp[13]) ? node31947 : node31932;
													assign node31932 = (inp[15]) ? node31940 : node31933;
														assign node31933 = (inp[10]) ? node31937 : node31934;
															assign node31934 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node31937 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31940 = (inp[10]) ? 4'b1110 : node31941;
															assign node31941 = (inp[11]) ? node31943 : 4'b1110;
																assign node31943 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node31947 = (inp[10]) ? node31953 : node31948;
														assign node31948 = (inp[0]) ? 4'b1110 : node31949;
															assign node31949 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node31953 = (inp[15]) ? node31959 : node31954;
															assign node31954 = (inp[11]) ? 4'b1110 : node31955;
																assign node31955 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node31959 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node31962 = (inp[11]) ? node31994 : node31963;
												assign node31963 = (inp[15]) ? node31979 : node31964;
													assign node31964 = (inp[0]) ? node31972 : node31965;
														assign node31965 = (inp[13]) ? node31969 : node31966;
															assign node31966 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31969 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node31972 = (inp[10]) ? node31976 : node31973;
															assign node31973 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31976 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node31979 = (inp[0]) ? node31987 : node31980;
														assign node31980 = (inp[10]) ? node31984 : node31981;
															assign node31981 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node31984 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node31987 = (inp[13]) ? node31991 : node31988;
															assign node31988 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node31991 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node31994 = (inp[13]) ? node32002 : node31995;
													assign node31995 = (inp[10]) ? node31999 : node31996;
														assign node31996 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31999 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node32002 = (inp[0]) ? node32006 : node32003;
														assign node32003 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node32006 = (inp[10]) ? 4'b1111 : 4'b1110;
										assign node32009 = (inp[10]) ? node32041 : node32010;
											assign node32010 = (inp[0]) ? node32032 : node32011;
												assign node32011 = (inp[11]) ? 4'b1100 : node32012;
													assign node32012 = (inp[9]) ? node32026 : node32013;
														assign node32013 = (inp[5]) ? node32021 : node32014;
															assign node32014 = (inp[15]) ? node32018 : node32015;
																assign node32015 = (inp[13]) ? 4'b1101 : 4'b1100;
																assign node32018 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node32021 = (inp[15]) ? 4'b1101 : node32022;
																assign node32022 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node32026 = (inp[15]) ? node32028 : 4'b1100;
															assign node32028 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node32032 = (inp[11]) ? 4'b1101 : node32033;
													assign node32033 = (inp[13]) ? node32037 : node32034;
														assign node32034 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node32037 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node32041 = (inp[0]) ? node32055 : node32042;
												assign node32042 = (inp[11]) ? 4'b1101 : node32043;
													assign node32043 = (inp[9]) ? node32049 : node32044;
														assign node32044 = (inp[13]) ? 4'b1100 : node32045;
															assign node32045 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node32049 = (inp[13]) ? node32051 : 4'b1101;
															assign node32051 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node32055 = (inp[11]) ? 4'b1100 : node32056;
													assign node32056 = (inp[13]) ? node32060 : node32057;
														assign node32057 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node32060 = (inp[15]) ? 4'b1100 : 4'b1101;
						assign node32064 = (inp[4]) ? node32848 : node32065;
							assign node32065 = (inp[12]) ? node32463 : node32066;
								assign node32066 = (inp[7]) ? node32248 : node32067;
									assign node32067 = (inp[5]) ? node32155 : node32068;
										assign node32068 = (inp[0]) ? node32120 : node32069;
											assign node32069 = (inp[10]) ? node32095 : node32070;
												assign node32070 = (inp[15]) ? node32084 : node32071;
													assign node32071 = (inp[13]) ? 4'b1001 : node32072;
														assign node32072 = (inp[9]) ? node32078 : node32073;
															assign node32073 = (inp[14]) ? 4'b1000 : node32074;
																assign node32074 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node32078 = (inp[14]) ? node32080 : 4'b1000;
																assign node32080 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node32084 = (inp[13]) ? node32086 : 4'b1001;
														assign node32086 = (inp[9]) ? node32090 : node32087;
															assign node32087 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node32090 = (inp[14]) ? node32092 : 4'b1001;
																assign node32092 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node32095 = (inp[11]) ? node32103 : node32096;
													assign node32096 = (inp[14]) ? 4'b1000 : node32097;
														assign node32097 = (inp[13]) ? 4'b1000 : node32098;
															assign node32098 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node32103 = (inp[14]) ? node32105 : 4'b1000;
														assign node32105 = (inp[9]) ? node32113 : node32106;
															assign node32106 = (inp[15]) ? node32110 : node32107;
																assign node32107 = (inp[13]) ? 4'b1000 : 4'b1001;
																assign node32110 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node32113 = (inp[15]) ? node32117 : node32114;
																assign node32114 = (inp[13]) ? 4'b1000 : 4'b1001;
																assign node32117 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node32120 = (inp[10]) ? node32138 : node32121;
												assign node32121 = (inp[11]) ? node32131 : node32122;
													assign node32122 = (inp[14]) ? 4'b1000 : node32123;
														assign node32123 = (inp[9]) ? node32125 : 4'b1000;
															assign node32125 = (inp[13]) ? 4'b1001 : node32126;
																assign node32126 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node32131 = (inp[14]) ? node32133 : 4'b1000;
														assign node32133 = (inp[15]) ? node32135 : 4'b1001;
															assign node32135 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node32138 = (inp[14]) ? node32148 : node32139;
													assign node32139 = (inp[11]) ? 4'b1001 : node32140;
														assign node32140 = (inp[15]) ? node32144 : node32141;
															assign node32141 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node32144 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node32148 = (inp[11]) ? node32150 : 4'b1001;
														assign node32150 = (inp[9]) ? 4'b1001 : node32151;
															assign node32151 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node32155 = (inp[14]) ? node32199 : node32156;
											assign node32156 = (inp[10]) ? node32174 : node32157;
												assign node32157 = (inp[0]) ? node32165 : node32158;
													assign node32158 = (inp[15]) ? node32160 : 4'b1001;
														assign node32160 = (inp[13]) ? node32162 : 4'b1001;
															assign node32162 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node32165 = (inp[11]) ? 4'b1000 : node32166;
														assign node32166 = (inp[13]) ? node32170 : node32167;
															assign node32167 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node32170 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node32174 = (inp[0]) ? node32192 : node32175;
													assign node32175 = (inp[11]) ? 4'b1000 : node32176;
														assign node32176 = (inp[9]) ? node32184 : node32177;
															assign node32177 = (inp[15]) ? node32181 : node32178;
																assign node32178 = (inp[13]) ? 4'b1000 : 4'b1001;
																assign node32181 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node32184 = (inp[13]) ? node32188 : node32185;
																assign node32185 = (inp[15]) ? 4'b1000 : 4'b1001;
																assign node32188 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node32192 = (inp[11]) ? 4'b1001 : node32193;
														assign node32193 = (inp[15]) ? node32195 : 4'b1001;
															assign node32195 = (inp[13]) ? 4'b1000 : 4'b1001;
											assign node32199 = (inp[15]) ? node32225 : node32200;
												assign node32200 = (inp[9]) ? node32210 : node32201;
													assign node32201 = (inp[10]) ? 4'b1100 : node32202;
														assign node32202 = (inp[0]) ? node32204 : 4'b1100;
															assign node32204 = (inp[13]) ? 4'b1100 : node32205;
																assign node32205 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node32210 = (inp[11]) ? node32220 : node32211;
														assign node32211 = (inp[13]) ? 4'b1101 : node32212;
															assign node32212 = (inp[10]) ? node32216 : node32213;
																assign node32213 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node32216 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node32220 = (inp[0]) ? 4'b1100 : node32221;
															assign node32221 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node32225 = (inp[11]) ? node32235 : node32226;
													assign node32226 = (inp[9]) ? 4'b1000 : node32227;
														assign node32227 = (inp[0]) ? 4'b1000 : node32228;
															assign node32228 = (inp[10]) ? 4'b1001 : node32229;
																assign node32229 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node32235 = (inp[9]) ? node32241 : node32236;
														assign node32236 = (inp[0]) ? 4'b1001 : node32237;
															assign node32237 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node32241 = (inp[10]) ? node32245 : node32242;
															assign node32242 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node32245 = (inp[0]) ? 4'b1001 : 4'b1000;
									assign node32248 = (inp[15]) ? node32358 : node32249;
										assign node32249 = (inp[5]) ? node32307 : node32250;
											assign node32250 = (inp[13]) ? node32300 : node32251;
												assign node32251 = (inp[9]) ? node32275 : node32252;
													assign node32252 = (inp[14]) ? node32262 : node32253;
														assign node32253 = (inp[10]) ? 4'b1001 : node32254;
															assign node32254 = (inp[0]) ? node32258 : node32255;
																assign node32255 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node32258 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node32262 = (inp[11]) ? node32268 : node32263;
															assign node32263 = (inp[0]) ? 4'b1001 : node32264;
																assign node32264 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node32268 = (inp[10]) ? node32272 : node32269;
																assign node32269 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node32272 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node32275 = (inp[11]) ? node32291 : node32276;
														assign node32276 = (inp[0]) ? node32284 : node32277;
															assign node32277 = (inp[14]) ? node32281 : node32278;
																assign node32278 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node32281 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node32284 = (inp[14]) ? node32288 : node32285;
																assign node32285 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node32288 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node32291 = (inp[14]) ? node32293 : 4'b1000;
															assign node32293 = (inp[10]) ? node32297 : node32294;
																assign node32294 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node32297 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node32300 = (inp[0]) ? node32304 : node32301;
													assign node32301 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node32304 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node32307 = (inp[14]) ? node32325 : node32308;
												assign node32308 = (inp[9]) ? node32314 : node32309;
													assign node32309 = (inp[11]) ? 4'b1100 : node32310;
														assign node32310 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node32314 = (inp[11]) ? node32320 : node32315;
														assign node32315 = (inp[0]) ? 4'b1100 : node32316;
															assign node32316 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node32320 = (inp[0]) ? 4'b1101 : node32321;
															assign node32321 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node32325 = (inp[13]) ? node32345 : node32326;
													assign node32326 = (inp[11]) ? node32332 : node32327;
														assign node32327 = (inp[0]) ? 4'b1001 : node32328;
															assign node32328 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node32332 = (inp[9]) ? node32340 : node32333;
															assign node32333 = (inp[0]) ? node32337 : node32334;
																assign node32334 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node32337 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node32340 = (inp[0]) ? node32342 : 4'b1001;
																assign node32342 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node32345 = (inp[0]) ? node32353 : node32346;
														assign node32346 = (inp[11]) ? node32350 : node32347;
															assign node32347 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node32350 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node32353 = (inp[9]) ? node32355 : 4'b1000;
															assign node32355 = (inp[10]) ? 4'b1000 : 4'b1001;
										assign node32358 = (inp[11]) ? node32412 : node32359;
											assign node32359 = (inp[0]) ? node32387 : node32360;
												assign node32360 = (inp[10]) ? node32374 : node32361;
													assign node32361 = (inp[5]) ? node32369 : node32362;
														assign node32362 = (inp[14]) ? node32366 : node32363;
															assign node32363 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node32366 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node32369 = (inp[14]) ? node32371 : 4'b1000;
															assign node32371 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node32374 = (inp[5]) ? node32382 : node32375;
														assign node32375 = (inp[14]) ? node32379 : node32376;
															assign node32376 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node32379 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node32382 = (inp[14]) ? node32384 : 4'b1001;
															assign node32384 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node32387 = (inp[10]) ? node32401 : node32388;
													assign node32388 = (inp[5]) ? node32396 : node32389;
														assign node32389 = (inp[14]) ? node32393 : node32390;
															assign node32390 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node32393 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node32396 = (inp[14]) ? node32398 : 4'b1001;
															assign node32398 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node32401 = (inp[5]) ? node32407 : node32402;
														assign node32402 = (inp[14]) ? node32404 : 4'b1101;
															assign node32404 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node32407 = (inp[14]) ? node32409 : 4'b1000;
															assign node32409 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node32412 = (inp[14]) ? node32446 : node32413;
												assign node32413 = (inp[5]) ? node32427 : node32414;
													assign node32414 = (inp[9]) ? 4'b1100 : node32415;
														assign node32415 = (inp[13]) ? node32421 : node32416;
															assign node32416 = (inp[0]) ? 4'b1100 : node32417;
																assign node32417 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node32421 = (inp[10]) ? node32423 : 4'b1100;
																assign node32423 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node32427 = (inp[9]) ? node32437 : node32428;
														assign node32428 = (inp[0]) ? node32430 : 4'b1001;
															assign node32430 = (inp[13]) ? node32434 : node32431;
																assign node32431 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node32434 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node32437 = (inp[0]) ? node32439 : 4'b1000;
															assign node32439 = (inp[10]) ? node32443 : node32440;
																assign node32440 = (inp[13]) ? 4'b1001 : 4'b1000;
																assign node32443 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node32446 = (inp[5]) ? node32456 : node32447;
													assign node32447 = (inp[13]) ? 4'b1000 : node32448;
														assign node32448 = (inp[10]) ? node32452 : node32449;
															assign node32449 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node32452 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node32456 = (inp[0]) ? node32460 : node32457;
														assign node32457 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node32460 = (inp[10]) ? 4'b1100 : 4'b1101;
								assign node32463 = (inp[7]) ? node32639 : node32464;
									assign node32464 = (inp[14]) ? node32542 : node32465;
										assign node32465 = (inp[11]) ? node32513 : node32466;
											assign node32466 = (inp[0]) ? node32498 : node32467;
												assign node32467 = (inp[15]) ? node32475 : node32468;
													assign node32468 = (inp[13]) ? node32472 : node32469;
														assign node32469 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node32472 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node32475 = (inp[5]) ? node32485 : node32476;
														assign node32476 = (inp[9]) ? node32478 : 4'b1011;
															assign node32478 = (inp[10]) ? node32482 : node32479;
																assign node32479 = (inp[13]) ? 4'b1011 : 4'b1010;
																assign node32482 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node32485 = (inp[9]) ? node32491 : node32486;
															assign node32486 = (inp[10]) ? node32488 : 4'b1010;
																assign node32488 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node32491 = (inp[10]) ? node32495 : node32492;
																assign node32492 = (inp[13]) ? 4'b1011 : 4'b1010;
																assign node32495 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node32498 = (inp[15]) ? 4'b1010 : node32499;
													assign node32499 = (inp[5]) ? node32505 : node32500;
														assign node32500 = (inp[9]) ? 4'b1010 : node32501;
															assign node32501 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node32505 = (inp[10]) ? node32509 : node32506;
															assign node32506 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node32509 = (inp[13]) ? 4'b1010 : 4'b1011;
											assign node32513 = (inp[15]) ? node32535 : node32514;
												assign node32514 = (inp[13]) ? node32522 : node32515;
													assign node32515 = (inp[0]) ? node32519 : node32516;
														assign node32516 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node32519 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node32522 = (inp[9]) ? node32528 : node32523;
														assign node32523 = (inp[0]) ? 4'b1010 : node32524;
															assign node32524 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node32528 = (inp[10]) ? node32532 : node32529;
															assign node32529 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node32532 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node32535 = (inp[0]) ? node32539 : node32536;
													assign node32536 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node32539 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node32542 = (inp[15]) ? node32586 : node32543;
											assign node32543 = (inp[13]) ? node32567 : node32544;
												assign node32544 = (inp[11]) ? node32552 : node32545;
													assign node32545 = (inp[10]) ? node32549 : node32546;
														assign node32546 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node32549 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node32552 = (inp[0]) ? node32558 : node32553;
														assign node32553 = (inp[9]) ? node32555 : 4'b1010;
															assign node32555 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node32558 = (inp[9]) ? 4'b1010 : node32559;
															assign node32559 = (inp[10]) ? node32563 : node32560;
																assign node32560 = (inp[5]) ? 4'b1011 : 4'b1010;
																assign node32563 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node32567 = (inp[0]) ? node32575 : node32568;
													assign node32568 = (inp[10]) ? 4'b1011 : node32569;
														assign node32569 = (inp[11]) ? 4'b1010 : node32570;
															assign node32570 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node32575 = (inp[10]) ? node32581 : node32576;
														assign node32576 = (inp[11]) ? 4'b1011 : node32577;
															assign node32577 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node32581 = (inp[5]) ? node32583 : 4'b1010;
															assign node32583 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node32586 = (inp[5]) ? node32608 : node32587;
												assign node32587 = (inp[10]) ? node32599 : node32588;
													assign node32588 = (inp[0]) ? node32594 : node32589;
														assign node32589 = (inp[13]) ? node32591 : 4'b1110;
															assign node32591 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node32594 = (inp[9]) ? node32596 : 4'b1111;
															assign node32596 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node32599 = (inp[0]) ? node32605 : node32600;
														assign node32600 = (inp[13]) ? node32602 : 4'b1111;
															assign node32602 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node32605 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node32608 = (inp[9]) ? node32622 : node32609;
													assign node32609 = (inp[13]) ? node32617 : node32610;
														assign node32610 = (inp[0]) ? 4'b1010 : node32611;
															assign node32611 = (inp[10]) ? node32613 : 4'b1010;
																assign node32613 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32617 = (inp[0]) ? node32619 : 4'b1010;
															assign node32619 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node32622 = (inp[10]) ? node32634 : node32623;
														assign node32623 = (inp[0]) ? node32629 : node32624;
															assign node32624 = (inp[11]) ? 4'b1010 : node32625;
																assign node32625 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node32629 = (inp[13]) ? 4'b1011 : node32630;
																assign node32630 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32634 = (inp[0]) ? node32636 : 4'b1011;
															assign node32636 = (inp[13]) ? 4'b1010 : 4'b1011;
									assign node32639 = (inp[15]) ? node32755 : node32640;
										assign node32640 = (inp[5]) ? node32694 : node32641;
											assign node32641 = (inp[14]) ? node32665 : node32642;
												assign node32642 = (inp[10]) ? node32654 : node32643;
													assign node32643 = (inp[0]) ? node32649 : node32644;
														assign node32644 = (inp[13]) ? node32646 : 4'b1010;
															assign node32646 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32649 = (inp[13]) ? node32651 : 4'b1011;
															assign node32651 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node32654 = (inp[0]) ? node32660 : node32655;
														assign node32655 = (inp[13]) ? node32657 : 4'b1011;
															assign node32657 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32660 = (inp[13]) ? node32662 : 4'b1010;
															assign node32662 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node32665 = (inp[11]) ? node32687 : node32666;
													assign node32666 = (inp[9]) ? node32672 : node32667;
														assign node32667 = (inp[10]) ? 4'b1111 : node32668;
															assign node32668 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node32672 = (inp[10]) ? node32680 : node32673;
															assign node32673 = (inp[13]) ? node32677 : node32674;
																assign node32674 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node32677 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32680 = (inp[0]) ? node32684 : node32681;
																assign node32681 = (inp[13]) ? 4'b1110 : 4'b1111;
																assign node32684 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node32687 = (inp[10]) ? node32691 : node32688;
														assign node32688 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32691 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node32694 = (inp[14]) ? node32724 : node32695;
												assign node32695 = (inp[9]) ? node32707 : node32696;
													assign node32696 = (inp[0]) ? node32702 : node32697;
														assign node32697 = (inp[10]) ? node32699 : 4'b1111;
															assign node32699 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node32702 = (inp[10]) ? 4'b1111 : node32703;
															assign node32703 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node32707 = (inp[13]) ? node32715 : node32708;
														assign node32708 = (inp[10]) ? node32712 : node32709;
															assign node32709 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32712 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32715 = (inp[0]) ? 4'b1110 : node32716;
															assign node32716 = (inp[11]) ? node32720 : node32717;
																assign node32717 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node32720 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node32724 = (inp[9]) ? node32740 : node32725;
													assign node32725 = (inp[10]) ? node32735 : node32726;
														assign node32726 = (inp[0]) ? node32732 : node32727;
															assign node32727 = (inp[11]) ? node32729 : 4'b1010;
																assign node32729 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node32732 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32735 = (inp[0]) ? 4'b1010 : node32736;
															assign node32736 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node32740 = (inp[13]) ? node32748 : node32741;
														assign node32741 = (inp[0]) ? 4'b1011 : node32742;
															assign node32742 = (inp[10]) ? node32744 : 4'b1011;
																assign node32744 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32748 = (inp[11]) ? 4'b1010 : node32749;
															assign node32749 = (inp[10]) ? node32751 : 4'b1011;
																assign node32751 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node32755 = (inp[14]) ? node32799 : node32756;
											assign node32756 = (inp[5]) ? node32778 : node32757;
												assign node32757 = (inp[13]) ? node32771 : node32758;
													assign node32758 = (inp[10]) ? node32766 : node32759;
														assign node32759 = (inp[0]) ? node32763 : node32760;
															assign node32760 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node32763 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node32766 = (inp[11]) ? 4'b1111 : node32767;
															assign node32767 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node32771 = (inp[0]) ? node32775 : node32772;
														assign node32772 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node32775 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node32778 = (inp[13]) ? node32786 : node32779;
													assign node32779 = (inp[0]) ? node32783 : node32780;
														assign node32780 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node32783 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node32786 = (inp[10]) ? node32794 : node32787;
														assign node32787 = (inp[9]) ? node32791 : node32788;
															assign node32788 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node32791 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32794 = (inp[9]) ? 4'b1010 : node32795;
															assign node32795 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node32799 = (inp[10]) ? node32823 : node32800;
												assign node32800 = (inp[13]) ? node32812 : node32801;
													assign node32801 = (inp[0]) ? node32807 : node32802;
														assign node32802 = (inp[11]) ? node32804 : 4'b1011;
															assign node32804 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node32807 = (inp[11]) ? node32809 : 4'b1010;
															assign node32809 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node32812 = (inp[0]) ? node32818 : node32813;
														assign node32813 = (inp[11]) ? 4'b1010 : node32814;
															assign node32814 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node32818 = (inp[11]) ? 4'b1011 : node32819;
															assign node32819 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node32823 = (inp[9]) ? node32837 : node32824;
													assign node32824 = (inp[13]) ? node32830 : node32825;
														assign node32825 = (inp[5]) ? node32827 : 4'b1011;
															assign node32827 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node32830 = (inp[0]) ? node32834 : node32831;
															assign node32831 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node32834 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node32837 = (inp[13]) ? node32841 : node32838;
														assign node32838 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node32841 = (inp[0]) ? node32843 : 4'b1011;
															assign node32843 = (inp[5]) ? 4'b1010 : node32844;
																assign node32844 = (inp[11]) ? 4'b1010 : 4'b1011;
							assign node32848 = (inp[12]) ? node33186 : node32849;
								assign node32849 = (inp[7]) ? node33031 : node32850;
									assign node32850 = (inp[5]) ? node32950 : node32851;
										assign node32851 = (inp[14]) ? node32891 : node32852;
											assign node32852 = (inp[0]) ? node32876 : node32853;
												assign node32853 = (inp[10]) ? node32861 : node32854;
													assign node32854 = (inp[11]) ? 4'b1010 : node32855;
														assign node32855 = (inp[13]) ? node32857 : 4'b1010;
															assign node32857 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node32861 = (inp[11]) ? 4'b1011 : node32862;
														assign node32862 = (inp[9]) ? node32868 : node32863;
															assign node32863 = (inp[13]) ? 4'b1011 : node32864;
																assign node32864 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node32868 = (inp[15]) ? node32872 : node32869;
																assign node32869 = (inp[13]) ? 4'b1011 : 4'b1010;
																assign node32872 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node32876 = (inp[10]) ? node32884 : node32877;
													assign node32877 = (inp[11]) ? 4'b1011 : node32878;
														assign node32878 = (inp[13]) ? node32880 : 4'b1011;
															assign node32880 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node32884 = (inp[11]) ? 4'b1010 : node32885;
														assign node32885 = (inp[15]) ? 4'b1010 : node32886;
															assign node32886 = (inp[13]) ? 4'b1010 : 4'b1011;
											assign node32891 = (inp[15]) ? node32927 : node32892;
												assign node32892 = (inp[11]) ? node32912 : node32893;
													assign node32893 = (inp[9]) ? node32903 : node32894;
														assign node32894 = (inp[13]) ? 4'b1010 : node32895;
															assign node32895 = (inp[0]) ? node32899 : node32896;
																assign node32896 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node32899 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node32903 = (inp[13]) ? node32907 : node32904;
															assign node32904 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node32907 = (inp[0]) ? node32909 : 4'b1011;
																assign node32909 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node32912 = (inp[0]) ? node32920 : node32913;
														assign node32913 = (inp[9]) ? node32915 : 4'b1011;
															assign node32915 = (inp[10]) ? node32917 : 4'b1011;
																assign node32917 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node32920 = (inp[10]) ? node32924 : node32921;
															assign node32921 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node32924 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node32927 = (inp[10]) ? node32939 : node32928;
													assign node32928 = (inp[13]) ? node32932 : node32929;
														assign node32929 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32932 = (inp[9]) ? node32934 : 4'b1110;
															assign node32934 = (inp[11]) ? node32936 : 4'b1111;
																assign node32936 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node32939 = (inp[0]) ? node32945 : node32940;
														assign node32940 = (inp[11]) ? node32942 : 4'b1111;
															assign node32942 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node32945 = (inp[13]) ? node32947 : 4'b1110;
															assign node32947 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node32950 = (inp[0]) ? node32990 : node32951;
											assign node32951 = (inp[10]) ? node32973 : node32952;
												assign node32952 = (inp[14]) ? node32964 : node32953;
													assign node32953 = (inp[15]) ? node32959 : node32954;
														assign node32954 = (inp[11]) ? node32956 : 4'b1010;
															assign node32956 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node32959 = (inp[11]) ? node32961 : 4'b1110;
															assign node32961 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node32964 = (inp[15]) ? node32970 : node32965;
														assign node32965 = (inp[11]) ? 4'b1110 : node32966;
															assign node32966 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node32970 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node32973 = (inp[14]) ? node32985 : node32974;
													assign node32974 = (inp[15]) ? node32980 : node32975;
														assign node32975 = (inp[13]) ? node32977 : 4'b1011;
															assign node32977 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32980 = (inp[13]) ? 4'b1111 : node32981;
															assign node32981 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node32985 = (inp[15]) ? 4'b1010 : node32986;
														assign node32986 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node32990 = (inp[10]) ? node33012 : node32991;
												assign node32991 = (inp[15]) ? node33003 : node32992;
													assign node32992 = (inp[14]) ? node32998 : node32993;
														assign node32993 = (inp[11]) ? node32995 : 4'b1011;
															assign node32995 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node32998 = (inp[13]) ? node33000 : 4'b1111;
															assign node33000 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node33003 = (inp[14]) ? node33009 : node33004;
														assign node33004 = (inp[11]) ? node33006 : 4'b1111;
															assign node33006 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node33009 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node33012 = (inp[15]) ? node33024 : node33013;
													assign node33013 = (inp[14]) ? node33019 : node33014;
														assign node33014 = (inp[11]) ? node33016 : 4'b1010;
															assign node33016 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node33019 = (inp[11]) ? 4'b1110 : node33020;
															assign node33020 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node33024 = (inp[14]) ? 4'b1011 : node33025;
														assign node33025 = (inp[11]) ? node33027 : 4'b1110;
															assign node33027 = (inp[13]) ? 4'b1110 : 4'b1111;
									assign node33031 = (inp[5]) ? node33109 : node33032;
										assign node33032 = (inp[13]) ? node33102 : node33033;
											assign node33033 = (inp[14]) ? node33055 : node33034;
												assign node33034 = (inp[10]) ? node33048 : node33035;
													assign node33035 = (inp[15]) ? node33041 : node33036;
														assign node33036 = (inp[9]) ? 4'b1011 : node33037;
															assign node33037 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node33041 = (inp[0]) ? node33045 : node33042;
															assign node33042 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node33045 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node33048 = (inp[0]) ? node33050 : 4'b1011;
														assign node33050 = (inp[15]) ? 4'b1011 : node33051;
															assign node33051 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node33055 = (inp[9]) ? node33073 : node33056;
													assign node33056 = (inp[10]) ? node33064 : node33057;
														assign node33057 = (inp[15]) ? node33061 : node33058;
															assign node33058 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33061 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33064 = (inp[11]) ? 4'b1011 : node33065;
															assign node33065 = (inp[15]) ? node33069 : node33066;
																assign node33066 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node33069 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node33073 = (inp[10]) ? node33089 : node33074;
														assign node33074 = (inp[11]) ? node33082 : node33075;
															assign node33075 = (inp[15]) ? node33079 : node33076;
																assign node33076 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node33079 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33082 = (inp[0]) ? node33086 : node33083;
																assign node33083 = (inp[15]) ? 4'b1010 : 4'b1011;
																assign node33086 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node33089 = (inp[15]) ? node33095 : node33090;
															assign node33090 = (inp[11]) ? node33092 : 4'b1010;
																assign node33092 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node33095 = (inp[0]) ? node33099 : node33096;
																assign node33096 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node33099 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node33102 = (inp[0]) ? node33106 : node33103;
												assign node33103 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node33106 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node33109 = (inp[14]) ? node33147 : node33110;
											assign node33110 = (inp[15]) ? node33128 : node33111;
												assign node33111 = (inp[10]) ? node33117 : node33112;
													assign node33112 = (inp[0]) ? node33114 : 4'b1111;
														assign node33114 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node33117 = (inp[0]) ? node33123 : node33118;
														assign node33118 = (inp[9]) ? 4'b1110 : node33119;
															assign node33119 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node33123 = (inp[13]) ? node33125 : 4'b1111;
															assign node33125 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node33128 = (inp[13]) ? node33136 : node33129;
													assign node33129 = (inp[10]) ? node33133 : node33130;
														assign node33130 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33133 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node33136 = (inp[0]) ? node33142 : node33137;
														assign node33137 = (inp[10]) ? 4'b1011 : node33138;
															assign node33138 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node33142 = (inp[11]) ? node33144 : 4'b1010;
															assign node33144 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node33147 = (inp[10]) ? node33169 : node33148;
												assign node33148 = (inp[0]) ? node33162 : node33149;
													assign node33149 = (inp[13]) ? 4'b1010 : node33150;
														assign node33150 = (inp[9]) ? node33156 : node33151;
															assign node33151 = (inp[11]) ? node33153 : 4'b1011;
																assign node33153 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node33156 = (inp[15]) ? 4'b1011 : node33157;
																assign node33157 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node33162 = (inp[13]) ? 4'b1011 : node33163;
														assign node33163 = (inp[9]) ? 4'b1011 : node33164;
															assign node33164 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node33169 = (inp[0]) ? node33177 : node33170;
													assign node33170 = (inp[13]) ? 4'b1011 : node33171;
														assign node33171 = (inp[15]) ? node33173 : 4'b1010;
															assign node33173 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node33177 = (inp[13]) ? 4'b1010 : node33178;
														assign node33178 = (inp[11]) ? node33182 : node33179;
															assign node33179 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node33182 = (inp[15]) ? 4'b1010 : 4'b1011;
								assign node33186 = (inp[7]) ? node33388 : node33187;
									assign node33187 = (inp[5]) ? node33275 : node33188;
										assign node33188 = (inp[14]) ? node33236 : node33189;
											assign node33189 = (inp[15]) ? node33217 : node33190;
												assign node33190 = (inp[13]) ? node33204 : node33191;
													assign node33191 = (inp[11]) ? node33199 : node33192;
														assign node33192 = (inp[0]) ? node33196 : node33193;
															assign node33193 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node33196 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node33199 = (inp[0]) ? node33201 : 4'b1101;
															assign node33201 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node33204 = (inp[9]) ? node33210 : node33205;
														assign node33205 = (inp[10]) ? 4'b1100 : node33206;
															assign node33206 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33210 = (inp[0]) ? node33214 : node33211;
															assign node33211 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node33214 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node33217 = (inp[9]) ? node33229 : node33218;
													assign node33218 = (inp[0]) ? 4'b1000 : node33219;
														assign node33219 = (inp[13]) ? 4'b1001 : node33220;
															assign node33220 = (inp[11]) ? node33224 : node33221;
																assign node33221 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node33224 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node33229 = (inp[0]) ? 4'b1001 : node33230;
														assign node33230 = (inp[10]) ? 4'b1001 : node33231;
															assign node33231 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node33236 = (inp[15]) ? node33256 : node33237;
												assign node33237 = (inp[0]) ? node33249 : node33238;
													assign node33238 = (inp[10]) ? node33244 : node33239;
														assign node33239 = (inp[11]) ? 4'b1001 : node33240;
															assign node33240 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node33244 = (inp[11]) ? 4'b1000 : node33245;
															assign node33245 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node33249 = (inp[10]) ? 4'b1001 : node33250;
														assign node33250 = (inp[13]) ? node33252 : 4'b1000;
															assign node33252 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node33256 = (inp[0]) ? node33266 : node33257;
													assign node33257 = (inp[13]) ? node33263 : node33258;
														assign node33258 = (inp[10]) ? node33260 : 4'b1100;
															assign node33260 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node33263 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node33266 = (inp[10]) ? node33272 : node33267;
														assign node33267 = (inp[11]) ? 4'b1100 : node33268;
															assign node33268 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node33272 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node33275 = (inp[14]) ? node33337 : node33276;
											assign node33276 = (inp[9]) ? node33308 : node33277;
												assign node33277 = (inp[11]) ? node33301 : node33278;
													assign node33278 = (inp[0]) ? node33292 : node33279;
														assign node33279 = (inp[10]) ? node33287 : node33280;
															assign node33280 = (inp[13]) ? node33284 : node33281;
																assign node33281 = (inp[15]) ? 4'b1000 : 4'b1001;
																assign node33284 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node33287 = (inp[13]) ? 4'b1000 : node33288;
																assign node33288 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node33292 = (inp[13]) ? 4'b1001 : node33293;
															assign node33293 = (inp[10]) ? node33297 : node33294;
																assign node33294 = (inp[15]) ? 4'b1001 : 4'b1000;
																assign node33297 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node33301 = (inp[10]) ? node33305 : node33302;
														assign node33302 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33305 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node33308 = (inp[10]) ? node33322 : node33309;
													assign node33309 = (inp[11]) ? 4'b1001 : node33310;
														assign node33310 = (inp[0]) ? node33316 : node33311;
															assign node33311 = (inp[13]) ? node33313 : 4'b1000;
																assign node33313 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node33316 = (inp[15]) ? node33318 : 4'b1001;
																assign node33318 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node33322 = (inp[0]) ? node33328 : node33323;
														assign node33323 = (inp[15]) ? 4'b1001 : node33324;
															assign node33324 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node33328 = (inp[11]) ? 4'b1000 : node33329;
															assign node33329 = (inp[13]) ? node33333 : node33330;
																assign node33330 = (inp[15]) ? 4'b1000 : 4'b1001;
																assign node33333 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node33337 = (inp[15]) ? node33361 : node33338;
												assign node33338 = (inp[10]) ? node33350 : node33339;
													assign node33339 = (inp[0]) ? node33345 : node33340;
														assign node33340 = (inp[13]) ? 4'b1100 : node33341;
															assign node33341 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node33345 = (inp[13]) ? 4'b1101 : node33346;
															assign node33346 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node33350 = (inp[0]) ? node33356 : node33351;
														assign node33351 = (inp[11]) ? node33353 : 4'b1101;
															assign node33353 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node33356 = (inp[13]) ? 4'b1100 : node33357;
															assign node33357 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node33361 = (inp[13]) ? node33377 : node33362;
													assign node33362 = (inp[10]) ? node33370 : node33363;
														assign node33363 = (inp[11]) ? node33367 : node33364;
															assign node33364 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node33367 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33370 = (inp[0]) ? node33374 : node33371;
															assign node33371 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node33374 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node33377 = (inp[9]) ? node33383 : node33378;
														assign node33378 = (inp[0]) ? node33380 : 4'b1001;
															assign node33380 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node33383 = (inp[0]) ? 4'b1001 : node33384;
															assign node33384 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node33388 = (inp[14]) ? node33462 : node33389;
										assign node33389 = (inp[5]) ? node33427 : node33390;
											assign node33390 = (inp[15]) ? node33412 : node33391;
												assign node33391 = (inp[0]) ? node33401 : node33392;
													assign node33392 = (inp[10]) ? node33396 : node33393;
														assign node33393 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node33396 = (inp[11]) ? 4'b1001 : node33397;
															assign node33397 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node33401 = (inp[10]) ? node33407 : node33402;
														assign node33402 = (inp[11]) ? 4'b1001 : node33403;
															assign node33403 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node33407 = (inp[13]) ? 4'b1000 : node33408;
															assign node33408 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node33412 = (inp[10]) ? node33420 : node33413;
													assign node33413 = (inp[0]) ? node33417 : node33414;
														assign node33414 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node33417 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node33420 = (inp[0]) ? 4'b1100 : node33421;
														assign node33421 = (inp[13]) ? node33423 : 4'b1101;
															assign node33423 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node33427 = (inp[0]) ? node33445 : node33428;
												assign node33428 = (inp[10]) ? node33436 : node33429;
													assign node33429 = (inp[11]) ? node33431 : 4'b1001;
														assign node33431 = (inp[15]) ? 4'b1000 : node33432;
															assign node33432 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node33436 = (inp[11]) ? 4'b1001 : node33437;
														assign node33437 = (inp[9]) ? node33439 : 4'b1000;
															assign node33439 = (inp[15]) ? node33441 : 4'b1000;
																assign node33441 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node33445 = (inp[10]) ? node33453 : node33446;
													assign node33446 = (inp[13]) ? node33450 : node33447;
														assign node33447 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node33450 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node33453 = (inp[15]) ? node33457 : node33454;
														assign node33454 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node33457 = (inp[11]) ? 4'b1000 : node33458;
															assign node33458 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node33462 = (inp[13]) ? node33516 : node33463;
											assign node33463 = (inp[10]) ? node33501 : node33464;
												assign node33464 = (inp[0]) ? node33490 : node33465;
													assign node33465 = (inp[5]) ? node33475 : node33466;
														assign node33466 = (inp[9]) ? node33470 : node33467;
															assign node33467 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node33470 = (inp[11]) ? 4'b1000 : node33471;
																assign node33471 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node33475 = (inp[9]) ? node33483 : node33476;
															assign node33476 = (inp[15]) ? node33480 : node33477;
																assign node33477 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node33480 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node33483 = (inp[15]) ? node33487 : node33484;
																assign node33484 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node33487 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node33490 = (inp[9]) ? node33496 : node33491;
														assign node33491 = (inp[11]) ? 4'b1000 : node33492;
															assign node33492 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node33496 = (inp[11]) ? 4'b1001 : node33497;
															assign node33497 = (inp[15]) ? 4'b1000 : 4'b1001;
												assign node33501 = (inp[15]) ? node33509 : node33502;
													assign node33502 = (inp[0]) ? node33506 : node33503;
														assign node33503 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node33506 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node33509 = (inp[11]) ? node33513 : node33510;
														assign node33510 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node33513 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node33516 = (inp[10]) ? node33520 : node33517;
												assign node33517 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node33520 = (inp[0]) ? 4'b1000 : 4'b1001;
				assign node33523 = (inp[12]) ? node35821 : node33524;
					assign node33524 = (inp[15]) ? node34490 : node33525;
						assign node33525 = (inp[14]) ? node34081 : node33526;
							assign node33526 = (inp[5]) ? node33830 : node33527;
								assign node33527 = (inp[11]) ? node33589 : node33528;
									assign node33528 = (inp[13]) ? node33560 : node33529;
										assign node33529 = (inp[10]) ? node33545 : node33530;
											assign node33530 = (inp[2]) ? node33534 : node33531;
												assign node33531 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node33534 = (inp[7]) ? node33538 : node33535;
													assign node33535 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node33538 = (inp[4]) ? node33542 : node33539;
														assign node33539 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node33542 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node33545 = (inp[2]) ? node33549 : node33546;
												assign node33546 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node33549 = (inp[7]) ? node33553 : node33550;
													assign node33550 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node33553 = (inp[4]) ? node33557 : node33554;
														assign node33554 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node33557 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node33560 = (inp[10]) ? node33574 : node33561;
											assign node33561 = (inp[2]) ? node33565 : node33562;
												assign node33562 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node33565 = (inp[7]) ? node33569 : node33566;
													assign node33566 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node33569 = (inp[4]) ? 4'b0001 : node33570;
														assign node33570 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node33574 = (inp[2]) ? node33578 : node33575;
												assign node33575 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node33578 = (inp[7]) ? node33582 : node33579;
													assign node33579 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node33582 = (inp[4]) ? node33586 : node33583;
														assign node33583 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node33586 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node33589 = (inp[7]) ? node33717 : node33590;
										assign node33590 = (inp[2]) ? node33648 : node33591;
											assign node33591 = (inp[10]) ? node33619 : node33592;
												assign node33592 = (inp[4]) ? node33598 : node33593;
													assign node33593 = (inp[1]) ? node33595 : 4'b0000;
														assign node33595 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node33598 = (inp[0]) ? node33614 : node33599;
														assign node33599 = (inp[9]) ? node33607 : node33600;
															assign node33600 = (inp[1]) ? node33604 : node33601;
																assign node33601 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node33604 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33607 = (inp[1]) ? node33611 : node33608;
																assign node33608 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node33611 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node33614 = (inp[13]) ? node33616 : 4'b0000;
															assign node33616 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node33619 = (inp[9]) ? node33635 : node33620;
													assign node33620 = (inp[0]) ? node33628 : node33621;
														assign node33621 = (inp[4]) ? 4'b0000 : node33622;
															assign node33622 = (inp[1]) ? 4'b0000 : node33623;
																assign node33623 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node33628 = (inp[1]) ? node33632 : node33629;
															assign node33629 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33632 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node33635 = (inp[4]) ? node33643 : node33636;
														assign node33636 = (inp[1]) ? node33640 : node33637;
															assign node33637 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node33640 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node33643 = (inp[1]) ? node33645 : 4'b0001;
															assign node33645 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node33648 = (inp[0]) ? node33680 : node33649;
												assign node33649 = (inp[9]) ? node33661 : node33650;
													assign node33650 = (inp[10]) ? node33656 : node33651;
														assign node33651 = (inp[4]) ? node33653 : 4'b0100;
															assign node33653 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node33656 = (inp[4]) ? node33658 : 4'b0101;
															assign node33658 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node33661 = (inp[1]) ? node33671 : node33662;
														assign node33662 = (inp[10]) ? 4'b0100 : node33663;
															assign node33663 = (inp[4]) ? node33667 : node33664;
																assign node33664 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node33667 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node33671 = (inp[4]) ? node33673 : 4'b0101;
															assign node33673 = (inp[10]) ? node33677 : node33674;
																assign node33674 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node33677 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node33680 = (inp[10]) ? node33702 : node33681;
													assign node33681 = (inp[9]) ? node33693 : node33682;
														assign node33682 = (inp[1]) ? node33688 : node33683;
															assign node33683 = (inp[13]) ? node33685 : 4'b0101;
																assign node33685 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node33688 = (inp[4]) ? node33690 : 4'b0100;
																assign node33690 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node33693 = (inp[1]) ? node33695 : 4'b0100;
															assign node33695 = (inp[13]) ? node33699 : node33696;
																assign node33696 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node33699 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node33702 = (inp[13]) ? node33710 : node33703;
														assign node33703 = (inp[4]) ? node33707 : node33704;
															assign node33704 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node33707 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node33710 = (inp[9]) ? node33712 : 4'b0100;
															assign node33712 = (inp[1]) ? node33714 : 4'b0100;
																assign node33714 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node33717 = (inp[2]) ? node33765 : node33718;
											assign node33718 = (inp[10]) ? node33750 : node33719;
												assign node33719 = (inp[9]) ? node33743 : node33720;
													assign node33720 = (inp[0]) ? node33736 : node33721;
														assign node33721 = (inp[4]) ? node33729 : node33722;
															assign node33722 = (inp[1]) ? node33726 : node33723;
																assign node33723 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node33726 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node33729 = (inp[1]) ? node33733 : node33730;
																assign node33730 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node33733 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node33736 = (inp[1]) ? node33740 : node33737;
															assign node33737 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node33740 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node33743 = (inp[13]) ? node33747 : node33744;
														assign node33744 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node33747 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node33750 = (inp[9]) ? node33758 : node33751;
													assign node33751 = (inp[13]) ? node33755 : node33752;
														assign node33752 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node33755 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node33758 = (inp[13]) ? node33762 : node33759;
														assign node33759 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node33762 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node33765 = (inp[9]) ? node33795 : node33766;
												assign node33766 = (inp[10]) ? node33782 : node33767;
													assign node33767 = (inp[1]) ? 4'b0000 : node33768;
														assign node33768 = (inp[0]) ? node33774 : node33769;
															assign node33769 = (inp[4]) ? node33771 : 4'b0000;
																assign node33771 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node33774 = (inp[4]) ? node33778 : node33775;
																assign node33775 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node33778 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node33782 = (inp[1]) ? node33790 : node33783;
														assign node33783 = (inp[0]) ? node33785 : 4'b0000;
															assign node33785 = (inp[13]) ? node33787 : 4'b0000;
																assign node33787 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node33790 = (inp[4]) ? 4'b0001 : node33791;
															assign node33791 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node33795 = (inp[1]) ? node33817 : node33796;
													assign node33796 = (inp[0]) ? node33812 : node33797;
														assign node33797 = (inp[4]) ? node33805 : node33798;
															assign node33798 = (inp[10]) ? node33802 : node33799;
																assign node33799 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node33802 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node33805 = (inp[13]) ? node33809 : node33806;
																assign node33806 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node33809 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node33812 = (inp[13]) ? 4'b0001 : node33813;
															assign node33813 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node33817 = (inp[13]) ? node33825 : node33818;
														assign node33818 = (inp[10]) ? node33822 : node33819;
															assign node33819 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node33822 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node33825 = (inp[10]) ? 4'b0000 : node33826;
															assign node33826 = (inp[4]) ? 4'b0001 : 4'b0000;
								assign node33830 = (inp[11]) ? node33916 : node33831;
									assign node33831 = (inp[10]) ? node33877 : node33832;
										assign node33832 = (inp[13]) ? node33852 : node33833;
											assign node33833 = (inp[7]) ? node33843 : node33834;
												assign node33834 = (inp[4]) ? node33838 : node33835;
													assign node33835 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node33838 = (inp[2]) ? 4'b0000 : node33839;
														assign node33839 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node33843 = (inp[2]) ? node33847 : node33844;
													assign node33844 = (inp[4]) ? 4'b0000 : 4'b0101;
													assign node33847 = (inp[4]) ? 4'b0101 : node33848;
														assign node33848 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node33852 = (inp[7]) ? node33862 : node33853;
												assign node33853 = (inp[4]) ? node33857 : node33854;
													assign node33854 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node33857 = (inp[2]) ? 4'b0001 : node33858;
														assign node33858 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node33862 = (inp[1]) ? node33870 : node33863;
													assign node33863 = (inp[2]) ? node33867 : node33864;
														assign node33864 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node33867 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node33870 = (inp[2]) ? node33874 : node33871;
														assign node33871 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node33874 = (inp[4]) ? 4'b0100 : 4'b0001;
										assign node33877 = (inp[13]) ? node33897 : node33878;
											assign node33878 = (inp[7]) ? node33888 : node33879;
												assign node33879 = (inp[2]) ? node33885 : node33880;
													assign node33880 = (inp[4]) ? node33882 : 4'b0001;
														assign node33882 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node33885 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node33888 = (inp[4]) ? node33894 : node33889;
													assign node33889 = (inp[2]) ? node33891 : 4'b0100;
														assign node33891 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node33894 = (inp[2]) ? 4'b0100 : 4'b0001;
											assign node33897 = (inp[7]) ? node33907 : node33898;
												assign node33898 = (inp[2]) ? node33904 : node33899;
													assign node33899 = (inp[4]) ? node33901 : 4'b0000;
														assign node33901 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node33904 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node33907 = (inp[4]) ? node33913 : node33908;
													assign node33908 = (inp[2]) ? node33910 : 4'b0101;
														assign node33910 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node33913 = (inp[2]) ? 4'b0101 : 4'b0000;
									assign node33916 = (inp[10]) ? node33996 : node33917;
										assign node33917 = (inp[13]) ? node33955 : node33918;
											assign node33918 = (inp[1]) ? node33940 : node33919;
												assign node33919 = (inp[7]) ? node33933 : node33920;
													assign node33920 = (inp[9]) ? node33926 : node33921;
														assign node33921 = (inp[4]) ? 4'b0000 : node33922;
															assign node33922 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node33926 = (inp[4]) ? node33930 : node33927;
															assign node33927 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node33930 = (inp[2]) ? 4'b0000 : 4'b0101;
													assign node33933 = (inp[4]) ? node33937 : node33934;
														assign node33934 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node33937 = (inp[2]) ? 4'b0101 : 4'b0000;
												assign node33940 = (inp[7]) ? node33948 : node33941;
													assign node33941 = (inp[2]) ? node33945 : node33942;
														assign node33942 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node33945 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node33948 = (inp[4]) ? node33952 : node33949;
														assign node33949 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node33952 = (inp[2]) ? 4'b0100 : 4'b0001;
											assign node33955 = (inp[1]) ? node33981 : node33956;
												assign node33956 = (inp[0]) ? node33972 : node33957;
													assign node33957 = (inp[4]) ? node33965 : node33958;
														assign node33958 = (inp[2]) ? node33962 : node33959;
															assign node33959 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node33962 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node33965 = (inp[2]) ? node33969 : node33966;
															assign node33966 = (inp[7]) ? 4'b0001 : 4'b0100;
															assign node33969 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node33972 = (inp[4]) ? 4'b0001 : node33973;
														assign node33973 = (inp[2]) ? node33977 : node33974;
															assign node33974 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node33977 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node33981 = (inp[7]) ? node33989 : node33982;
													assign node33982 = (inp[4]) ? node33986 : node33983;
														assign node33983 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node33986 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node33989 = (inp[4]) ? node33993 : node33990;
														assign node33990 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node33993 = (inp[2]) ? 4'b0101 : 4'b0000;
										assign node33996 = (inp[13]) ? node34026 : node33997;
											assign node33997 = (inp[4]) ? node34013 : node33998;
												assign node33998 = (inp[1]) ? node34006 : node33999;
													assign node33999 = (inp[7]) ? node34003 : node34000;
														assign node34000 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node34003 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node34006 = (inp[7]) ? node34010 : node34007;
														assign node34007 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node34010 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node34013 = (inp[2]) ? node34019 : node34014;
													assign node34014 = (inp[7]) ? node34016 : 4'b0100;
														assign node34016 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node34019 = (inp[7]) ? node34023 : node34020;
														assign node34020 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node34023 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node34026 = (inp[4]) ? node34056 : node34027;
												assign node34027 = (inp[9]) ? node34041 : node34028;
													assign node34028 = (inp[2]) ? node34036 : node34029;
														assign node34029 = (inp[7]) ? node34033 : node34030;
															assign node34030 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node34033 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node34036 = (inp[7]) ? 4'b0000 : node34037;
															assign node34037 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node34041 = (inp[0]) ? node34049 : node34042;
														assign node34042 = (inp[7]) ? node34046 : node34043;
															assign node34043 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node34046 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node34049 = (inp[1]) ? node34053 : node34050;
															assign node34050 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node34053 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node34056 = (inp[9]) ? node34066 : node34057;
													assign node34057 = (inp[2]) ? node34059 : 4'b0101;
														assign node34059 = (inp[7]) ? node34063 : node34060;
															assign node34060 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node34063 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node34066 = (inp[1]) ? node34074 : node34067;
														assign node34067 = (inp[7]) ? node34071 : node34068;
															assign node34068 = (inp[2]) ? 4'b0000 : 4'b0101;
															assign node34071 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node34074 = (inp[2]) ? node34078 : node34075;
															assign node34075 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node34078 = (inp[7]) ? 4'b0100 : 4'b0001;
							assign node34081 = (inp[13]) ? node34277 : node34082;
								assign node34082 = (inp[10]) ? node34182 : node34083;
									assign node34083 = (inp[1]) ? node34151 : node34084;
										assign node34084 = (inp[11]) ? node34126 : node34085;
											assign node34085 = (inp[5]) ? node34095 : node34086;
												assign node34086 = (inp[2]) ? node34090 : node34087;
													assign node34087 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node34090 = (inp[7]) ? node34092 : 4'b0111;
														assign node34092 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node34095 = (inp[0]) ? node34105 : node34096;
													assign node34096 = (inp[9]) ? 4'b0011 : node34097;
														assign node34097 = (inp[7]) ? 4'b0010 : node34098;
															assign node34098 = (inp[4]) ? 4'b0011 : node34099;
																assign node34099 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node34105 = (inp[4]) ? node34119 : node34106;
														assign node34106 = (inp[9]) ? node34114 : node34107;
															assign node34107 = (inp[2]) ? node34111 : node34108;
																assign node34108 = (inp[7]) ? 4'b0011 : 4'b0110;
																assign node34111 = (inp[7]) ? 4'b0110 : 4'b0011;
															assign node34114 = (inp[7]) ? node34116 : 4'b0011;
																assign node34116 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node34119 = (inp[7]) ? node34123 : node34120;
															assign node34120 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node34123 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node34126 = (inp[2]) ? node34138 : node34127;
												assign node34127 = (inp[7]) ? node34133 : node34128;
													assign node34128 = (inp[5]) ? node34130 : 4'b0011;
														assign node34130 = (inp[4]) ? 4'b0010 : 4'b0111;
													assign node34133 = (inp[5]) ? node34135 : 4'b0111;
														assign node34135 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node34138 = (inp[7]) ? node34146 : node34139;
													assign node34139 = (inp[4]) ? node34143 : node34140;
														assign node34140 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node34143 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node34146 = (inp[4]) ? 4'b0011 : node34147;
														assign node34147 = (inp[5]) ? 4'b0111 : 4'b0010;
										assign node34151 = (inp[2]) ? node34165 : node34152;
											assign node34152 = (inp[7]) ? node34158 : node34153;
												assign node34153 = (inp[5]) ? node34155 : 4'b0010;
													assign node34155 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node34158 = (inp[4]) ? 4'b0110 : node34159;
													assign node34159 = (inp[5]) ? node34161 : 4'b0110;
														assign node34161 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node34165 = (inp[7]) ? node34177 : node34166;
												assign node34166 = (inp[11]) ? node34172 : node34167;
													assign node34167 = (inp[4]) ? node34169 : 4'b0111;
														assign node34169 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node34172 = (inp[5]) ? 4'b0110 : node34173;
														assign node34173 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node34177 = (inp[4]) ? 4'b0010 : node34178;
													assign node34178 = (inp[5]) ? 4'b0110 : 4'b0011;
									assign node34182 = (inp[1]) ? node34238 : node34183;
										assign node34183 = (inp[11]) ? node34209 : node34184;
											assign node34184 = (inp[5]) ? node34196 : node34185;
												assign node34185 = (inp[2]) ? node34189 : node34186;
													assign node34186 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node34189 = (inp[7]) ? node34193 : node34190;
														assign node34190 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node34193 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node34196 = (inp[7]) ? node34202 : node34197;
													assign node34197 = (inp[4]) ? 4'b0010 : node34198;
														assign node34198 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node34202 = (inp[2]) ? node34206 : node34203;
														assign node34203 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node34206 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node34209 = (inp[7]) ? node34225 : node34210;
												assign node34210 = (inp[2]) ? node34218 : node34211;
													assign node34211 = (inp[4]) ? node34215 : node34212;
														assign node34212 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node34215 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node34218 = (inp[5]) ? node34222 : node34219;
														assign node34219 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node34222 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node34225 = (inp[2]) ? node34231 : node34226;
													assign node34226 = (inp[4]) ? 4'b0110 : node34227;
														assign node34227 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node34231 = (inp[5]) ? node34235 : node34232;
														assign node34232 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node34235 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node34238 = (inp[2]) ? node34252 : node34239;
											assign node34239 = (inp[7]) ? node34245 : node34240;
												assign node34240 = (inp[5]) ? node34242 : 4'b0011;
													assign node34242 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node34245 = (inp[5]) ? node34247 : 4'b0111;
													assign node34247 = (inp[4]) ? 4'b0111 : node34248;
														assign node34248 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node34252 = (inp[7]) ? node34270 : node34253;
												assign node34253 = (inp[4]) ? node34259 : node34254;
													assign node34254 = (inp[5]) ? 4'b0010 : node34255;
														assign node34255 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node34259 = (inp[0]) ? node34267 : node34260;
														assign node34260 = (inp[5]) ? node34264 : node34261;
															assign node34261 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node34264 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node34267 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node34270 = (inp[5]) ? node34274 : node34271;
													assign node34271 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node34274 = (inp[4]) ? 4'b0011 : 4'b0111;
								assign node34277 = (inp[10]) ? node34381 : node34278;
									assign node34278 = (inp[1]) ? node34334 : node34279;
										assign node34279 = (inp[11]) ? node34307 : node34280;
											assign node34280 = (inp[2]) ? node34292 : node34281;
												assign node34281 = (inp[7]) ? node34287 : node34282;
													assign node34282 = (inp[5]) ? node34284 : 4'b0011;
														assign node34284 = (inp[4]) ? 4'b0010 : 4'b0111;
													assign node34287 = (inp[4]) ? 4'b0111 : node34288;
														assign node34288 = (inp[5]) ? 4'b0010 : 4'b0111;
												assign node34292 = (inp[7]) ? node34300 : node34293;
													assign node34293 = (inp[4]) ? node34297 : node34294;
														assign node34294 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node34297 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node34300 = (inp[5]) ? node34304 : node34301;
														assign node34301 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node34304 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node34307 = (inp[7]) ? node34323 : node34308;
												assign node34308 = (inp[2]) ? node34316 : node34309;
													assign node34309 = (inp[4]) ? node34313 : node34310;
														assign node34310 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node34313 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node34316 = (inp[5]) ? node34320 : node34317;
														assign node34317 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node34320 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node34323 = (inp[2]) ? node34329 : node34324;
													assign node34324 = (inp[5]) ? node34326 : 4'b0110;
														assign node34326 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node34329 = (inp[4]) ? 4'b0010 : node34330;
														assign node34330 = (inp[5]) ? 4'b0110 : 4'b0011;
										assign node34334 = (inp[7]) ? node34368 : node34335;
											assign node34335 = (inp[2]) ? node34341 : node34336;
												assign node34336 = (inp[5]) ? node34338 : 4'b0011;
													assign node34338 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node34341 = (inp[4]) ? node34347 : node34342;
													assign node34342 = (inp[5]) ? 4'b0010 : node34343;
														assign node34343 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node34347 = (inp[9]) ? node34353 : node34348;
														assign node34348 = (inp[5]) ? node34350 : 4'b0111;
															assign node34350 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node34353 = (inp[0]) ? node34361 : node34354;
															assign node34354 = (inp[5]) ? node34358 : node34355;
																assign node34355 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node34358 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node34361 = (inp[11]) ? node34365 : node34362;
																assign node34362 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node34365 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node34368 = (inp[2]) ? node34376 : node34369;
												assign node34369 = (inp[4]) ? 4'b0111 : node34370;
													assign node34370 = (inp[5]) ? node34372 : 4'b0111;
														assign node34372 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node34376 = (inp[4]) ? 4'b0011 : node34377;
													assign node34377 = (inp[5]) ? 4'b0111 : 4'b0010;
									assign node34381 = (inp[1]) ? node34445 : node34382;
										assign node34382 = (inp[11]) ? node34420 : node34383;
											assign node34383 = (inp[2]) ? node34405 : node34384;
												assign node34384 = (inp[5]) ? node34388 : node34385;
													assign node34385 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node34388 = (inp[9]) ? node34398 : node34389;
														assign node34389 = (inp[0]) ? node34393 : node34390;
															assign node34390 = (inp[7]) ? 4'b0110 : 4'b0011;
															assign node34393 = (inp[4]) ? 4'b0011 : node34394;
																assign node34394 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node34398 = (inp[0]) ? 4'b0110 : node34399;
															assign node34399 = (inp[4]) ? 4'b0011 : node34400;
																assign node34400 = (inp[7]) ? 4'b0011 : 4'b0110;
												assign node34405 = (inp[7]) ? node34413 : node34406;
													assign node34406 = (inp[5]) ? node34410 : node34407;
														assign node34407 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node34410 = (inp[4]) ? 4'b0110 : 4'b0011;
													assign node34413 = (inp[5]) ? node34417 : node34414;
														assign node34414 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node34417 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node34420 = (inp[7]) ? node34434 : node34421;
												assign node34421 = (inp[2]) ? node34429 : node34422;
													assign node34422 = (inp[4]) ? node34426 : node34423;
														assign node34423 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node34426 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node34429 = (inp[5]) ? 4'b0010 : node34430;
														assign node34430 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node34434 = (inp[2]) ? node34440 : node34435;
													assign node34435 = (inp[5]) ? node34437 : 4'b0111;
														assign node34437 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node34440 = (inp[4]) ? 4'b0011 : node34441;
														assign node34441 = (inp[5]) ? 4'b0111 : 4'b0010;
										assign node34445 = (inp[2]) ? node34463 : node34446;
											assign node34446 = (inp[5]) ? node34450 : node34447;
												assign node34447 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node34450 = (inp[11]) ? node34458 : node34451;
													assign node34451 = (inp[7]) ? node34455 : node34452;
														assign node34452 = (inp[4]) ? 4'b0011 : 4'b0110;
														assign node34455 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node34458 = (inp[7]) ? 4'b0011 : node34459;
														assign node34459 = (inp[4]) ? 4'b0011 : 4'b0110;
											assign node34463 = (inp[7]) ? node34483 : node34464;
												assign node34464 = (inp[11]) ? node34472 : node34465;
													assign node34465 = (inp[4]) ? node34469 : node34466;
														assign node34466 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node34469 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node34472 = (inp[9]) ? 4'b0110 : node34473;
														assign node34473 = (inp[0]) ? node34477 : node34474;
															assign node34474 = (inp[4]) ? 4'b0110 : 4'b0011;
															assign node34477 = (inp[4]) ? node34479 : 4'b0110;
																assign node34479 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node34483 = (inp[5]) ? node34487 : node34484;
													assign node34484 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node34487 = (inp[4]) ? 4'b0010 : 4'b0110;
						assign node34490 = (inp[5]) ? node35128 : node34491;
							assign node34491 = (inp[13]) ? node34927 : node34492;
								assign node34492 = (inp[9]) ? node34752 : node34493;
									assign node34493 = (inp[7]) ? node34615 : node34494;
										assign node34494 = (inp[1]) ? node34542 : node34495;
											assign node34495 = (inp[10]) ? node34515 : node34496;
												assign node34496 = (inp[14]) ? node34506 : node34497;
													assign node34497 = (inp[2]) ? node34501 : node34498;
														assign node34498 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node34501 = (inp[4]) ? node34503 : 4'b0110;
															assign node34503 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node34506 = (inp[11]) ? node34508 : 4'b0010;
														assign node34508 = (inp[2]) ? node34512 : node34509;
															assign node34509 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34512 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node34515 = (inp[14]) ? node34529 : node34516;
													assign node34516 = (inp[11]) ? node34522 : node34517;
														assign node34517 = (inp[2]) ? 4'b0010 : node34518;
															assign node34518 = (inp[0]) ? 4'b0011 : 4'b0111;
														assign node34522 = (inp[2]) ? node34526 : node34523;
															assign node34523 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34526 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node34529 = (inp[11]) ? node34537 : node34530;
														assign node34530 = (inp[2]) ? node34534 : node34531;
															assign node34531 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34534 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node34537 = (inp[2]) ? 4'b0010 : node34538;
															assign node34538 = (inp[0]) ? 4'b0110 : 4'b0010;
											assign node34542 = (inp[10]) ? node34580 : node34543;
												assign node34543 = (inp[11]) ? node34565 : node34544;
													assign node34544 = (inp[14]) ? node34552 : node34545;
														assign node34545 = (inp[0]) ? 4'b0010 : node34546;
															assign node34546 = (inp[2]) ? 4'b0111 : node34547;
																assign node34547 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34552 = (inp[0]) ? node34560 : node34553;
															assign node34553 = (inp[2]) ? node34557 : node34554;
																assign node34554 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node34557 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node34560 = (inp[4]) ? 4'b0111 : node34561;
																assign node34561 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node34565 = (inp[14]) ? node34573 : node34566;
														assign node34566 = (inp[2]) ? node34570 : node34567;
															assign node34567 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34570 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node34573 = (inp[2]) ? node34577 : node34574;
															assign node34574 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node34577 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node34580 = (inp[0]) ? node34598 : node34581;
													assign node34581 = (inp[14]) ? node34589 : node34582;
														assign node34582 = (inp[2]) ? node34586 : node34583;
															assign node34583 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node34586 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node34589 = (inp[4]) ? node34593 : node34590;
															assign node34590 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node34593 = (inp[11]) ? node34595 : 4'b0110;
																assign node34595 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node34598 = (inp[2]) ? node34606 : node34599;
														assign node34599 = (inp[4]) ? 4'b0110 : node34600;
															assign node34600 = (inp[11]) ? node34602 : 4'b0010;
																assign node34602 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node34606 = (inp[4]) ? node34608 : 4'b0110;
															assign node34608 = (inp[14]) ? node34612 : node34609;
																assign node34609 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node34612 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node34615 = (inp[11]) ? node34685 : node34616;
											assign node34616 = (inp[0]) ? node34652 : node34617;
												assign node34617 = (inp[1]) ? node34635 : node34618;
													assign node34618 = (inp[10]) ? node34632 : node34619;
														assign node34619 = (inp[14]) ? node34627 : node34620;
															assign node34620 = (inp[4]) ? node34624 : node34621;
																assign node34621 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node34624 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node34627 = (inp[2]) ? 4'b0111 : node34628;
																assign node34628 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node34632 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node34635 = (inp[10]) ? node34645 : node34636;
														assign node34636 = (inp[2]) ? node34640 : node34637;
															assign node34637 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34640 = (inp[4]) ? 4'b0011 : node34641;
																assign node34641 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node34645 = (inp[4]) ? node34649 : node34646;
															assign node34646 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node34649 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node34652 = (inp[2]) ? node34668 : node34653;
													assign node34653 = (inp[4]) ? node34661 : node34654;
														assign node34654 = (inp[1]) ? node34658 : node34655;
															assign node34655 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node34658 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node34661 = (inp[10]) ? node34665 : node34662;
															assign node34662 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node34665 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node34668 = (inp[4]) ? node34672 : node34669;
														assign node34669 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node34672 = (inp[14]) ? node34680 : node34673;
															assign node34673 = (inp[1]) ? node34677 : node34674;
																assign node34674 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node34677 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node34680 = (inp[10]) ? node34682 : 4'b0010;
																assign node34682 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node34685 = (inp[1]) ? node34715 : node34686;
												assign node34686 = (inp[10]) ? node34706 : node34687;
													assign node34687 = (inp[14]) ? node34693 : node34688;
														assign node34688 = (inp[2]) ? 4'b0111 : node34689;
															assign node34689 = (inp[0]) ? 4'b0011 : 4'b0111;
														assign node34693 = (inp[0]) ? node34699 : node34694;
															assign node34694 = (inp[4]) ? node34696 : 4'b0110;
																assign node34696 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node34699 = (inp[2]) ? node34703 : node34700;
																assign node34700 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node34703 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node34706 = (inp[14]) ? node34708 : 4'b0110;
														assign node34708 = (inp[4]) ? node34712 : node34709;
															assign node34709 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node34712 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node34715 = (inp[0]) ? node34733 : node34716;
													assign node34716 = (inp[2]) ? node34726 : node34717;
														assign node34717 = (inp[4]) ? 4'b0110 : node34718;
															assign node34718 = (inp[10]) ? node34722 : node34719;
																assign node34719 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node34722 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node34726 = (inp[4]) ? node34730 : node34727;
															assign node34727 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node34730 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node34733 = (inp[2]) ? node34743 : node34734;
														assign node34734 = (inp[4]) ? node34736 : 4'b0011;
															assign node34736 = (inp[14]) ? node34740 : node34737;
																assign node34737 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node34740 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node34743 = (inp[4]) ? node34749 : node34744;
															assign node34744 = (inp[10]) ? node34746 : 4'b0110;
																assign node34746 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node34749 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node34752 = (inp[1]) ? node34838 : node34753;
										assign node34753 = (inp[10]) ? node34799 : node34754;
											assign node34754 = (inp[11]) ? node34774 : node34755;
												assign node34755 = (inp[14]) ? node34767 : node34756;
													assign node34756 = (inp[0]) ? 4'b0010 : node34757;
														assign node34757 = (inp[2]) ? node34761 : node34758;
															assign node34758 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node34761 = (inp[7]) ? node34763 : 4'b0011;
																assign node34763 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node34767 = (inp[4]) ? node34771 : node34768;
														assign node34768 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node34771 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node34774 = (inp[14]) ? node34790 : node34775;
													assign node34775 = (inp[7]) ? node34781 : node34776;
														assign node34776 = (inp[2]) ? 4'b0010 : node34777;
															assign node34777 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node34781 = (inp[0]) ? node34787 : node34782;
															assign node34782 = (inp[2]) ? 4'b0111 : node34783;
																assign node34783 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34787 = (inp[4]) ? 4'b0010 : 4'b0111;
													assign node34790 = (inp[4]) ? node34794 : node34791;
														assign node34791 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node34794 = (inp[2]) ? 4'b0011 : node34795;
															assign node34795 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node34799 = (inp[11]) ? node34815 : node34800;
												assign node34800 = (inp[2]) ? node34804 : node34801;
													assign node34801 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node34804 = (inp[4]) ? node34810 : node34805;
														assign node34805 = (inp[7]) ? node34807 : 4'b0111;
															assign node34807 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node34810 = (inp[14]) ? 4'b0011 : node34811;
															assign node34811 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node34815 = (inp[2]) ? node34827 : node34816;
													assign node34816 = (inp[4]) ? node34824 : node34817;
														assign node34817 = (inp[14]) ? node34821 : node34818;
															assign node34818 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node34821 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node34824 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node34827 = (inp[4]) ? node34833 : node34828;
														assign node34828 = (inp[7]) ? node34830 : 4'b0111;
															assign node34830 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node34833 = (inp[14]) ? node34835 : 4'b0011;
															assign node34835 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node34838 = (inp[10]) ? node34888 : node34839;
											assign node34839 = (inp[11]) ? node34859 : node34840;
												assign node34840 = (inp[7]) ? node34850 : node34841;
													assign node34841 = (inp[2]) ? node34845 : node34842;
														assign node34842 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node34845 = (inp[4]) ? node34847 : 4'b0111;
															assign node34847 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node34850 = (inp[14]) ? node34852 : 4'b0011;
														assign node34852 = (inp[2]) ? node34856 : node34853;
															assign node34853 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node34856 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node34859 = (inp[14]) ? node34873 : node34860;
													assign node34860 = (inp[7]) ? node34866 : node34861;
														assign node34861 = (inp[4]) ? 4'b0111 : node34862;
															assign node34862 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node34866 = (inp[4]) ? node34870 : node34867;
															assign node34867 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node34870 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node34873 = (inp[7]) ? node34879 : node34874;
														assign node34874 = (inp[4]) ? 4'b0010 : node34875;
															assign node34875 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node34879 = (inp[0]) ? node34881 : 4'b0011;
															assign node34881 = (inp[2]) ? node34885 : node34882;
																assign node34882 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node34885 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node34888 = (inp[11]) ? node34900 : node34889;
												assign node34889 = (inp[2]) ? node34893 : node34890;
													assign node34890 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node34893 = (inp[4]) ? node34895 : 4'b0110;
														assign node34895 = (inp[14]) ? 4'b0010 : node34896;
															assign node34896 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node34900 = (inp[2]) ? node34916 : node34901;
													assign node34901 = (inp[4]) ? node34909 : node34902;
														assign node34902 = (inp[14]) ? node34906 : node34903;
															assign node34903 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node34906 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node34909 = (inp[14]) ? node34913 : node34910;
															assign node34910 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node34913 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node34916 = (inp[4]) ? node34922 : node34917;
														assign node34917 = (inp[7]) ? node34919 : 4'b0110;
															assign node34919 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node34922 = (inp[14]) ? node34924 : 4'b0010;
															assign node34924 = (inp[7]) ? 4'b0010 : 4'b0011;
								assign node34927 = (inp[1]) ? node35031 : node34928;
									assign node34928 = (inp[10]) ? node34982 : node34929;
										assign node34929 = (inp[11]) ? node34945 : node34930;
											assign node34930 = (inp[2]) ? node34934 : node34931;
												assign node34931 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node34934 = (inp[4]) ? node34940 : node34935;
													assign node34935 = (inp[14]) ? node34937 : 4'b0110;
														assign node34937 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node34940 = (inp[7]) ? 4'b0010 : node34941;
														assign node34941 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node34945 = (inp[2]) ? node34971 : node34946;
												assign node34946 = (inp[4]) ? node34956 : node34947;
													assign node34947 = (inp[9]) ? 4'b0010 : node34948;
														assign node34948 = (inp[14]) ? node34952 : node34949;
															assign node34949 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node34952 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node34956 = (inp[0]) ? node34964 : node34957;
														assign node34957 = (inp[7]) ? node34961 : node34958;
															assign node34958 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node34961 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node34964 = (inp[7]) ? node34968 : node34965;
															assign node34965 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node34968 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node34971 = (inp[4]) ? node34977 : node34972;
													assign node34972 = (inp[14]) ? 4'b0110 : node34973;
														assign node34973 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node34977 = (inp[14]) ? node34979 : 4'b0010;
														assign node34979 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node34982 = (inp[11]) ? node34998 : node34983;
											assign node34983 = (inp[2]) ? node34987 : node34984;
												assign node34984 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node34987 = (inp[4]) ? node34993 : node34988;
													assign node34988 = (inp[14]) ? node34990 : 4'b0111;
														assign node34990 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node34993 = (inp[7]) ? 4'b0011 : node34994;
														assign node34994 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node34998 = (inp[2]) ? node35020 : node34999;
												assign node34999 = (inp[4]) ? node35007 : node35000;
													assign node35000 = (inp[7]) ? node35004 : node35001;
														assign node35001 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node35004 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node35007 = (inp[9]) ? node35013 : node35008;
														assign node35008 = (inp[7]) ? node35010 : 4'b0111;
															assign node35010 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35013 = (inp[0]) ? node35015 : 4'b0110;
															assign node35015 = (inp[7]) ? 4'b0111 : node35016;
																assign node35016 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node35020 = (inp[4]) ? node35026 : node35021;
													assign node35021 = (inp[14]) ? 4'b0111 : node35022;
														assign node35022 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node35026 = (inp[7]) ? 4'b0011 : node35027;
														assign node35027 = (inp[14]) ? 4'b0010 : 4'b0011;
									assign node35031 = (inp[10]) ? node35079 : node35032;
										assign node35032 = (inp[11]) ? node35048 : node35033;
											assign node35033 = (inp[2]) ? node35037 : node35034;
												assign node35034 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node35037 = (inp[4]) ? node35043 : node35038;
													assign node35038 = (inp[14]) ? node35040 : 4'b0111;
														assign node35040 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node35043 = (inp[7]) ? 4'b0011 : node35044;
														assign node35044 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node35048 = (inp[2]) ? node35068 : node35049;
												assign node35049 = (inp[4]) ? node35061 : node35050;
													assign node35050 = (inp[9]) ? node35052 : 4'b0010;
														assign node35052 = (inp[0]) ? node35054 : 4'b0011;
															assign node35054 = (inp[14]) ? node35058 : node35055;
																assign node35055 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node35058 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node35061 = (inp[14]) ? node35065 : node35062;
														assign node35062 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node35065 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node35068 = (inp[4]) ? node35074 : node35069;
													assign node35069 = (inp[14]) ? 4'b0111 : node35070;
														assign node35070 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node35074 = (inp[7]) ? 4'b0011 : node35075;
														assign node35075 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node35079 = (inp[11]) ? node35095 : node35080;
											assign node35080 = (inp[2]) ? node35084 : node35081;
												assign node35081 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node35084 = (inp[4]) ? node35090 : node35085;
													assign node35085 = (inp[14]) ? node35087 : 4'b0110;
														assign node35087 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node35090 = (inp[7]) ? 4'b0010 : node35091;
														assign node35091 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node35095 = (inp[2]) ? node35117 : node35096;
												assign node35096 = (inp[4]) ? node35110 : node35097;
													assign node35097 = (inp[0]) ? node35105 : node35098;
														assign node35098 = (inp[14]) ? node35102 : node35099;
															assign node35099 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node35102 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node35105 = (inp[14]) ? node35107 : 4'b0011;
															assign node35107 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node35110 = (inp[7]) ? node35114 : node35111;
														assign node35111 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35114 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node35117 = (inp[4]) ? node35123 : node35118;
													assign node35118 = (inp[7]) ? node35120 : 4'b0110;
														assign node35120 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node35123 = (inp[7]) ? 4'b0010 : node35124;
														assign node35124 = (inp[14]) ? 4'b0011 : 4'b0010;
							assign node35128 = (inp[0]) ? node35476 : node35129;
								assign node35129 = (inp[7]) ? node35309 : node35130;
									assign node35130 = (inp[9]) ? node35218 : node35131;
										assign node35131 = (inp[1]) ? node35177 : node35132;
											assign node35132 = (inp[10]) ? node35150 : node35133;
												assign node35133 = (inp[11]) ? node35143 : node35134;
													assign node35134 = (inp[14]) ? node35136 : 4'b0110;
														assign node35136 = (inp[2]) ? node35140 : node35137;
															assign node35137 = (inp[4]) ? 4'b0111 : 4'b0010;
															assign node35140 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node35143 = (inp[4]) ? node35147 : node35144;
														assign node35144 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node35147 = (inp[2]) ? 4'b0010 : 4'b0111;
												assign node35150 = (inp[11]) ? node35164 : node35151;
													assign node35151 = (inp[14]) ? node35159 : node35152;
														assign node35152 = (inp[13]) ? node35154 : 4'b0011;
															assign node35154 = (inp[2]) ? node35156 : 4'b0111;
																assign node35156 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35159 = (inp[2]) ? node35161 : 4'b0011;
															assign node35161 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node35164 = (inp[14]) ? node35172 : node35165;
														assign node35165 = (inp[2]) ? node35169 : node35166;
															assign node35166 = (inp[4]) ? 4'b0110 : 4'b0011;
															assign node35169 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35172 = (inp[2]) ? 4'b0111 : node35173;
															assign node35173 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node35177 = (inp[10]) ? node35193 : node35178;
												assign node35178 = (inp[4]) ? node35182 : node35179;
													assign node35179 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node35182 = (inp[2]) ? node35188 : node35183;
														assign node35183 = (inp[14]) ? 4'b0110 : node35184;
															assign node35184 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node35188 = (inp[11]) ? 4'b0011 : node35189;
															assign node35189 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node35193 = (inp[11]) ? node35207 : node35194;
													assign node35194 = (inp[14]) ? node35200 : node35195;
														assign node35195 = (inp[4]) ? 4'b0010 : node35196;
															assign node35196 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node35200 = (inp[2]) ? node35204 : node35201;
															assign node35201 = (inp[4]) ? 4'b0111 : 4'b0010;
															assign node35204 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node35207 = (inp[13]) ? node35211 : node35208;
														assign node35208 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node35211 = (inp[2]) ? node35215 : node35212;
															assign node35212 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node35215 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node35218 = (inp[2]) ? node35264 : node35219;
											assign node35219 = (inp[4]) ? node35235 : node35220;
												assign node35220 = (inp[14]) ? node35228 : node35221;
													assign node35221 = (inp[10]) ? node35225 : node35222;
														assign node35222 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node35225 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node35228 = (inp[10]) ? node35232 : node35229;
														assign node35229 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node35232 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node35235 = (inp[11]) ? node35245 : node35236;
													assign node35236 = (inp[13]) ? 4'b0111 : node35237;
														assign node35237 = (inp[10]) ? node35239 : 4'b0110;
															assign node35239 = (inp[14]) ? node35241 : 4'b0111;
																assign node35241 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node35245 = (inp[13]) ? node35259 : node35246;
														assign node35246 = (inp[1]) ? node35252 : node35247;
															assign node35247 = (inp[10]) ? node35249 : 4'b0111;
																assign node35249 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35252 = (inp[14]) ? node35256 : node35253;
																assign node35253 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node35256 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node35259 = (inp[14]) ? 4'b0110 : node35260;
															assign node35260 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node35264 = (inp[4]) ? node35286 : node35265;
												assign node35265 = (inp[11]) ? node35281 : node35266;
													assign node35266 = (inp[1]) ? node35272 : node35267;
														assign node35267 = (inp[13]) ? node35269 : 4'b0110;
															assign node35269 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35272 = (inp[13]) ? node35274 : 4'b0111;
															assign node35274 = (inp[10]) ? node35278 : node35275;
																assign node35275 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35278 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node35281 = (inp[1]) ? 4'b0110 : node35282;
														assign node35282 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node35286 = (inp[10]) ? node35298 : node35287;
													assign node35287 = (inp[1]) ? node35293 : node35288;
														assign node35288 = (inp[14]) ? node35290 : 4'b0010;
															assign node35290 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node35293 = (inp[11]) ? 4'b0011 : node35294;
															assign node35294 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node35298 = (inp[1]) ? node35304 : node35299;
														assign node35299 = (inp[14]) ? node35301 : 4'b0011;
															assign node35301 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node35304 = (inp[11]) ? 4'b0010 : node35305;
															assign node35305 = (inp[14]) ? 4'b0011 : 4'b0010;
									assign node35309 = (inp[11]) ? node35431 : node35310;
										assign node35310 = (inp[13]) ? node35368 : node35311;
											assign node35311 = (inp[1]) ? node35337 : node35312;
												assign node35312 = (inp[14]) ? node35328 : node35313;
													assign node35313 = (inp[10]) ? node35321 : node35314;
														assign node35314 = (inp[2]) ? node35318 : node35315;
															assign node35315 = (inp[4]) ? 4'b0110 : 4'b0011;
															assign node35318 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35321 = (inp[4]) ? node35325 : node35322;
															assign node35322 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node35325 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node35328 = (inp[10]) ? 4'b0011 : node35329;
														assign node35329 = (inp[2]) ? node35333 : node35330;
															assign node35330 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node35333 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node35337 = (inp[2]) ? node35347 : node35338;
													assign node35338 = (inp[4]) ? node35344 : node35339;
														assign node35339 = (inp[10]) ? 4'b0011 : node35340;
															assign node35340 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node35344 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node35347 = (inp[4]) ? node35355 : node35348;
														assign node35348 = (inp[10]) ? node35352 : node35349;
															assign node35349 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35352 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node35355 = (inp[9]) ? node35361 : node35356;
															assign node35356 = (inp[10]) ? node35358 : 4'b0010;
																assign node35358 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node35361 = (inp[10]) ? node35365 : node35362;
																assign node35362 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node35365 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node35368 = (inp[1]) ? node35404 : node35369;
												assign node35369 = (inp[10]) ? node35389 : node35370;
													assign node35370 = (inp[14]) ? node35380 : node35371;
														assign node35371 = (inp[9]) ? node35373 : 4'b0011;
															assign node35373 = (inp[2]) ? node35377 : node35374;
																assign node35374 = (inp[4]) ? 4'b0110 : 4'b0011;
																assign node35377 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35380 = (inp[9]) ? node35382 : 4'b0010;
															assign node35382 = (inp[2]) ? node35386 : node35383;
																assign node35383 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node35386 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node35389 = (inp[14]) ? node35397 : node35390;
														assign node35390 = (inp[2]) ? node35394 : node35391;
															assign node35391 = (inp[4]) ? 4'b0111 : 4'b0010;
															assign node35394 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node35397 = (inp[4]) ? node35401 : node35398;
															assign node35398 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node35401 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node35404 = (inp[14]) ? node35416 : node35405;
													assign node35405 = (inp[10]) ? node35411 : node35406;
														assign node35406 = (inp[4]) ? 4'b0010 : node35407;
															assign node35407 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node35411 = (inp[4]) ? node35413 : 4'b0011;
															assign node35413 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node35416 = (inp[10]) ? node35424 : node35417;
														assign node35417 = (inp[2]) ? node35421 : node35418;
															assign node35418 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node35421 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35424 = (inp[4]) ? node35428 : node35425;
															assign node35425 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node35428 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node35431 = (inp[1]) ? node35457 : node35432;
											assign node35432 = (inp[10]) ? node35448 : node35433;
												assign node35433 = (inp[14]) ? node35441 : node35434;
													assign node35434 = (inp[2]) ? node35438 : node35435;
														assign node35435 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node35438 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node35441 = (inp[2]) ? node35445 : node35442;
														assign node35442 = (inp[4]) ? 4'b0110 : 4'b0011;
														assign node35445 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node35448 = (inp[2]) ? node35454 : node35449;
													assign node35449 = (inp[4]) ? 4'b0111 : node35450;
														assign node35450 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node35454 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node35457 = (inp[10]) ? node35467 : node35458;
												assign node35458 = (inp[4]) ? node35464 : node35459;
													assign node35459 = (inp[2]) ? 4'b0111 : node35460;
														assign node35460 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node35464 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node35467 = (inp[2]) ? node35473 : node35468;
													assign node35468 = (inp[4]) ? 4'b0110 : node35469;
														assign node35469 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node35473 = (inp[4]) ? 4'b0010 : 4'b0110;
								assign node35476 = (inp[4]) ? node35656 : node35477;
									assign node35477 = (inp[2]) ? node35593 : node35478;
										assign node35478 = (inp[11]) ? node35538 : node35479;
											assign node35479 = (inp[14]) ? node35503 : node35480;
												assign node35480 = (inp[9]) ? node35490 : node35481;
													assign node35481 = (inp[10]) ? node35483 : 4'b0011;
														assign node35483 = (inp[7]) ? node35487 : node35484;
															assign node35484 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node35487 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node35490 = (inp[1]) ? node35498 : node35491;
														assign node35491 = (inp[7]) ? node35495 : node35492;
															assign node35492 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node35495 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node35498 = (inp[10]) ? 4'b0010 : node35499;
															assign node35499 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node35503 = (inp[9]) ? node35525 : node35504;
													assign node35504 = (inp[13]) ? node35512 : node35505;
														assign node35505 = (inp[1]) ? node35509 : node35506;
															assign node35506 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node35509 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node35512 = (inp[7]) ? node35520 : node35513;
															assign node35513 = (inp[1]) ? node35517 : node35514;
																assign node35514 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node35517 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node35520 = (inp[1]) ? 4'b0010 : node35521;
																assign node35521 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node35525 = (inp[7]) ? node35533 : node35526;
														assign node35526 = (inp[10]) ? node35530 : node35527;
															assign node35527 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node35530 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node35533 = (inp[13]) ? node35535 : 4'b0011;
															assign node35535 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node35538 = (inp[13]) ? node35562 : node35539;
												assign node35539 = (inp[7]) ? node35547 : node35540;
													assign node35540 = (inp[10]) ? node35544 : node35541;
														assign node35541 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node35544 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node35547 = (inp[9]) ? node35555 : node35548;
														assign node35548 = (inp[1]) ? 4'b0011 : node35549;
															assign node35549 = (inp[10]) ? node35551 : 4'b0010;
																assign node35551 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node35555 = (inp[1]) ? 4'b0010 : node35556;
															assign node35556 = (inp[14]) ? node35558 : 4'b0011;
																assign node35558 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node35562 = (inp[9]) ? node35578 : node35563;
													assign node35563 = (inp[1]) ? node35573 : node35564;
														assign node35564 = (inp[10]) ? node35570 : node35565;
															assign node35565 = (inp[7]) ? node35567 : 4'b0010;
																assign node35567 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node35570 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node35573 = (inp[14]) ? 4'b0010 : node35574;
															assign node35574 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node35578 = (inp[10]) ? node35584 : node35579;
														assign node35579 = (inp[1]) ? 4'b0011 : node35580;
															assign node35580 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node35584 = (inp[1]) ? node35588 : node35585;
															assign node35585 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node35588 = (inp[7]) ? node35590 : 4'b0010;
																assign node35590 = (inp[14]) ? 4'b0011 : 4'b0010;
										assign node35593 = (inp[11]) ? node35641 : node35594;
											assign node35594 = (inp[9]) ? node35622 : node35595;
												assign node35595 = (inp[14]) ? node35609 : node35596;
													assign node35596 = (inp[1]) ? node35604 : node35597;
														assign node35597 = (inp[7]) ? node35601 : node35598;
															assign node35598 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node35601 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node35604 = (inp[10]) ? 4'b0110 : node35605;
															assign node35605 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node35609 = (inp[1]) ? node35615 : node35610;
														assign node35610 = (inp[7]) ? node35612 : 4'b0111;
															assign node35612 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node35615 = (inp[13]) ? 4'b0110 : node35616;
															assign node35616 = (inp[10]) ? 4'b0111 : node35617;
																assign node35617 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node35622 = (inp[7]) ? node35628 : node35623;
													assign node35623 = (inp[14]) ? node35625 : 4'b0110;
														assign node35625 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node35628 = (inp[1]) ? node35634 : node35629;
														assign node35629 = (inp[14]) ? 4'b0110 : node35630;
															assign node35630 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node35634 = (inp[10]) ? node35638 : node35635;
															assign node35635 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35638 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node35641 = (inp[13]) ? node35649 : node35642;
												assign node35642 = (inp[10]) ? node35646 : node35643;
													assign node35643 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node35646 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node35649 = (inp[10]) ? node35653 : node35650;
													assign node35650 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node35653 = (inp[1]) ? 4'b0110 : 4'b0111;
									assign node35656 = (inp[2]) ? node35720 : node35657;
										assign node35657 = (inp[1]) ? node35701 : node35658;
											assign node35658 = (inp[10]) ? node35670 : node35659;
												assign node35659 = (inp[7]) ? 4'b0110 : node35660;
													assign node35660 = (inp[13]) ? node35662 : 4'b0110;
														assign node35662 = (inp[11]) ? node35666 : node35663;
															assign node35663 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35666 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node35670 = (inp[7]) ? 4'b0111 : node35671;
													assign node35671 = (inp[9]) ? node35687 : node35672;
														assign node35672 = (inp[13]) ? node35680 : node35673;
															assign node35673 = (inp[11]) ? node35677 : node35674;
																assign node35674 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35677 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35680 = (inp[11]) ? node35684 : node35681;
																assign node35681 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35684 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35687 = (inp[13]) ? node35693 : node35688;
															assign node35688 = (inp[11]) ? node35690 : 4'b0110;
																assign node35690 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node35693 = (inp[11]) ? node35697 : node35694;
																assign node35694 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node35697 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node35701 = (inp[10]) ? node35711 : node35702;
												assign node35702 = (inp[7]) ? 4'b0111 : node35703;
													assign node35703 = (inp[14]) ? node35707 : node35704;
														assign node35704 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node35707 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node35711 = (inp[7]) ? 4'b0110 : node35712;
													assign node35712 = (inp[14]) ? node35716 : node35713;
														assign node35713 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node35716 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node35720 = (inp[9]) ? node35770 : node35721;
											assign node35721 = (inp[13]) ? node35739 : node35722;
												assign node35722 = (inp[11]) ? node35732 : node35723;
													assign node35723 = (inp[10]) ? node35725 : 4'b0010;
														assign node35725 = (inp[1]) ? node35727 : 4'b0011;
															assign node35727 = (inp[7]) ? node35729 : 4'b0010;
																assign node35729 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node35732 = (inp[1]) ? node35736 : node35733;
														assign node35733 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node35736 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node35739 = (inp[7]) ? node35755 : node35740;
													assign node35740 = (inp[1]) ? node35748 : node35741;
														assign node35741 = (inp[10]) ? node35743 : 4'b0010;
															assign node35743 = (inp[11]) ? 4'b0011 : node35744;
																assign node35744 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node35748 = (inp[10]) ? 4'b0010 : node35749;
															assign node35749 = (inp[14]) ? node35751 : 4'b0011;
																assign node35751 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node35755 = (inp[14]) ? node35763 : node35756;
														assign node35756 = (inp[1]) ? 4'b0010 : node35757;
															assign node35757 = (inp[10]) ? node35759 : 4'b0011;
																assign node35759 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node35763 = (inp[11]) ? node35765 : 4'b0011;
															assign node35765 = (inp[1]) ? 4'b0011 : node35766;
																assign node35766 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node35770 = (inp[7]) ? node35800 : node35771;
												assign node35771 = (inp[13]) ? node35785 : node35772;
													assign node35772 = (inp[1]) ? node35778 : node35773;
														assign node35773 = (inp[10]) ? node35775 : 4'b0010;
															assign node35775 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node35778 = (inp[10]) ? node35780 : 4'b0011;
															assign node35780 = (inp[14]) ? node35782 : 4'b0010;
																assign node35782 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node35785 = (inp[14]) ? node35791 : node35786;
														assign node35786 = (inp[10]) ? node35788 : 4'b0010;
															assign node35788 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node35791 = (inp[11]) ? node35793 : 4'b0010;
															assign node35793 = (inp[1]) ? node35797 : node35794;
																assign node35794 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node35797 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node35800 = (inp[10]) ? node35812 : node35801;
													assign node35801 = (inp[1]) ? node35807 : node35802;
														assign node35802 = (inp[11]) ? 4'b0010 : node35803;
															assign node35803 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node35807 = (inp[11]) ? 4'b0011 : node35808;
															assign node35808 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node35812 = (inp[1]) ? node35816 : node35813;
														assign node35813 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node35816 = (inp[11]) ? 4'b0010 : node35817;
															assign node35817 = (inp[14]) ? 4'b0010 : 4'b0011;
					assign node35821 = (inp[15]) ? node36951 : node35822;
						assign node35822 = (inp[14]) ? node36228 : node35823;
							assign node35823 = (inp[13]) ? node36023 : node35824;
								assign node35824 = (inp[10]) ? node35928 : node35825;
									assign node35825 = (inp[11]) ? node35893 : node35826;
										assign node35826 = (inp[1]) ? node35868 : node35827;
											assign node35827 = (inp[7]) ? node35853 : node35828;
												assign node35828 = (inp[4]) ? node35832 : node35829;
													assign node35829 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node35832 = (inp[0]) ? node35840 : node35833;
														assign node35833 = (inp[2]) ? node35837 : node35834;
															assign node35834 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node35837 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node35840 = (inp[9]) ? node35848 : node35841;
															assign node35841 = (inp[2]) ? node35845 : node35842;
																assign node35842 = (inp[5]) ? 4'b0011 : 4'b0110;
																assign node35845 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node35848 = (inp[2]) ? 4'b0110 : node35849;
																assign node35849 = (inp[5]) ? 4'b0011 : 4'b0110;
												assign node35853 = (inp[2]) ? node35861 : node35854;
													assign node35854 = (inp[4]) ? node35858 : node35855;
														assign node35855 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node35858 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node35861 = (inp[4]) ? node35865 : node35862;
														assign node35862 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node35865 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node35868 = (inp[7]) ? node35880 : node35869;
												assign node35869 = (inp[2]) ? node35875 : node35870;
													assign node35870 = (inp[4]) ? node35872 : 4'b0011;
														assign node35872 = (inp[5]) ? 4'b0010 : 4'b0111;
													assign node35875 = (inp[4]) ? node35877 : 4'b0111;
														assign node35877 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node35880 = (inp[2]) ? node35888 : node35881;
													assign node35881 = (inp[5]) ? node35885 : node35882;
														assign node35882 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node35885 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node35888 = (inp[5]) ? 4'b0011 : node35889;
														assign node35889 = (inp[4]) ? 4'b0111 : 4'b0010;
										assign node35893 = (inp[2]) ? node35915 : node35894;
											assign node35894 = (inp[7]) ? node35902 : node35895;
												assign node35895 = (inp[5]) ? node35899 : node35896;
													assign node35896 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node35899 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node35902 = (inp[4]) ? node35910 : node35903;
													assign node35903 = (inp[1]) ? node35907 : node35904;
														assign node35904 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node35907 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node35910 = (inp[5]) ? node35912 : 4'b0011;
														assign node35912 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node35915 = (inp[7]) ? node35923 : node35916;
												assign node35916 = (inp[5]) ? 4'b0110 : node35917;
													assign node35917 = (inp[4]) ? node35919 : 4'b0110;
														assign node35919 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node35923 = (inp[5]) ? 4'b0010 : node35924;
													assign node35924 = (inp[4]) ? 4'b0110 : 4'b0011;
									assign node35928 = (inp[11]) ? node35982 : node35929;
										assign node35929 = (inp[1]) ? node35957 : node35930;
											assign node35930 = (inp[7]) ? node35944 : node35931;
												assign node35931 = (inp[2]) ? node35939 : node35932;
													assign node35932 = (inp[5]) ? node35936 : node35933;
														assign node35933 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node35936 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node35939 = (inp[5]) ? 4'b0111 : node35940;
														assign node35940 = (inp[4]) ? 4'b0010 : 4'b0111;
												assign node35944 = (inp[2]) ? node35952 : node35945;
													assign node35945 = (inp[5]) ? node35949 : node35946;
														assign node35946 = (inp[4]) ? 4'b0010 : 4'b0111;
														assign node35949 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node35952 = (inp[5]) ? 4'b0011 : node35953;
														assign node35953 = (inp[4]) ? 4'b0111 : 4'b0010;
											assign node35957 = (inp[7]) ? node35969 : node35958;
												assign node35958 = (inp[2]) ? node35964 : node35959;
													assign node35959 = (inp[4]) ? node35961 : 4'b0010;
														assign node35961 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node35964 = (inp[5]) ? 4'b0110 : node35965;
														assign node35965 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node35969 = (inp[2]) ? node35977 : node35970;
													assign node35970 = (inp[5]) ? node35974 : node35971;
														assign node35971 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node35974 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node35977 = (inp[5]) ? 4'b0010 : node35978;
														assign node35978 = (inp[4]) ? 4'b0110 : 4'b0011;
										assign node35982 = (inp[2]) ? node36008 : node35983;
											assign node35983 = (inp[4]) ? node35991 : node35984;
												assign node35984 = (inp[7]) ? node35986 : 4'b0011;
													assign node35986 = (inp[1]) ? 4'b0111 : node35987;
														assign node35987 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node35991 = (inp[1]) ? node35999 : node35992;
													assign node35992 = (inp[5]) ? node35996 : node35993;
														assign node35993 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node35996 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node35999 = (inp[9]) ? node36001 : 4'b0111;
														assign node36001 = (inp[7]) ? node36005 : node36002;
															assign node36002 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node36005 = (inp[5]) ? 4'b0111 : 4'b0010;
											assign node36008 = (inp[7]) ? node36016 : node36009;
												assign node36009 = (inp[5]) ? 4'b0111 : node36010;
													assign node36010 = (inp[4]) ? node36012 : 4'b0111;
														assign node36012 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node36016 = (inp[4]) ? node36020 : node36017;
													assign node36017 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node36020 = (inp[5]) ? 4'b0011 : 4'b0111;
								assign node36023 = (inp[10]) ? node36131 : node36024;
									assign node36024 = (inp[11]) ? node36088 : node36025;
										assign node36025 = (inp[1]) ? node36063 : node36026;
											assign node36026 = (inp[5]) ? node36052 : node36027;
												assign node36027 = (inp[0]) ? node36033 : node36028;
													assign node36028 = (inp[4]) ? 4'b0010 : node36029;
														assign node36029 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node36033 = (inp[9]) ? node36043 : node36034;
														assign node36034 = (inp[2]) ? node36036 : 4'b0010;
															assign node36036 = (inp[7]) ? node36040 : node36037;
																assign node36037 = (inp[4]) ? 4'b0010 : 4'b0111;
																assign node36040 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node36043 = (inp[2]) ? 4'b0111 : node36044;
															assign node36044 = (inp[4]) ? node36048 : node36045;
																assign node36045 = (inp[7]) ? 4'b0111 : 4'b0011;
																assign node36048 = (inp[7]) ? 4'b0010 : 4'b0111;
												assign node36052 = (inp[2]) ? node36060 : node36053;
													assign node36053 = (inp[7]) ? node36057 : node36054;
														assign node36054 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node36057 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node36060 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node36063 = (inp[2]) ? node36077 : node36064;
												assign node36064 = (inp[7]) ? node36070 : node36065;
													assign node36065 = (inp[0]) ? 4'b0011 : node36066;
														assign node36066 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node36070 = (inp[4]) ? node36074 : node36071;
														assign node36071 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node36074 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node36077 = (inp[7]) ? node36083 : node36078;
													assign node36078 = (inp[5]) ? 4'b0110 : node36079;
														assign node36079 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node36083 = (inp[5]) ? 4'b0010 : node36084;
														assign node36084 = (inp[4]) ? 4'b0110 : 4'b0011;
										assign node36088 = (inp[7]) ? node36102 : node36089;
											assign node36089 = (inp[2]) ? node36095 : node36090;
												assign node36090 = (inp[4]) ? node36092 : 4'b0011;
													assign node36092 = (inp[5]) ? 4'b0010 : 4'b0111;
												assign node36095 = (inp[4]) ? node36097 : 4'b0111;
													assign node36097 = (inp[5]) ? 4'b0111 : node36098;
														assign node36098 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node36102 = (inp[2]) ? node36126 : node36103;
												assign node36103 = (inp[5]) ? node36109 : node36104;
													assign node36104 = (inp[4]) ? 4'b0010 : node36105;
														assign node36105 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node36109 = (inp[0]) ? node36119 : node36110;
														assign node36110 = (inp[9]) ? node36112 : 4'b0111;
															assign node36112 = (inp[1]) ? node36116 : node36113;
																assign node36113 = (inp[4]) ? 4'b0110 : 4'b0111;
																assign node36116 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node36119 = (inp[1]) ? node36123 : node36120;
															assign node36120 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node36123 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node36126 = (inp[5]) ? 4'b0011 : node36127;
													assign node36127 = (inp[4]) ? 4'b0111 : 4'b0010;
									assign node36131 = (inp[11]) ? node36195 : node36132;
										assign node36132 = (inp[1]) ? node36166 : node36133;
											assign node36133 = (inp[4]) ? node36145 : node36134;
												assign node36134 = (inp[7]) ? node36138 : node36135;
													assign node36135 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node36138 = (inp[2]) ? node36142 : node36139;
														assign node36139 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node36142 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node36145 = (inp[5]) ? node36159 : node36146;
													assign node36146 = (inp[0]) ? node36152 : node36147;
														assign node36147 = (inp[2]) ? 4'b0011 : node36148;
															assign node36148 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node36152 = (inp[7]) ? node36156 : node36153;
															assign node36153 = (inp[2]) ? 4'b0011 : 4'b0110;
															assign node36156 = (inp[2]) ? 4'b0110 : 4'b0011;
													assign node36159 = (inp[7]) ? node36163 : node36160;
														assign node36160 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node36163 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node36166 = (inp[2]) ? node36182 : node36167;
												assign node36167 = (inp[7]) ? node36175 : node36168;
													assign node36168 = (inp[5]) ? node36172 : node36169;
														assign node36169 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node36172 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node36175 = (inp[5]) ? node36179 : node36176;
														assign node36176 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node36179 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node36182 = (inp[7]) ? node36188 : node36183;
													assign node36183 = (inp[4]) ? node36185 : 4'b0111;
														assign node36185 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node36188 = (inp[4]) ? node36192 : node36189;
														assign node36189 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node36192 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node36195 = (inp[2]) ? node36215 : node36196;
											assign node36196 = (inp[7]) ? node36202 : node36197;
												assign node36197 = (inp[4]) ? node36199 : 4'b0010;
													assign node36199 = (inp[5]) ? 4'b0011 : 4'b0110;
												assign node36202 = (inp[5]) ? node36208 : node36203;
													assign node36203 = (inp[4]) ? 4'b0011 : node36204;
														assign node36204 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node36208 = (inp[1]) ? node36212 : node36209;
														assign node36209 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node36212 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node36215 = (inp[7]) ? node36223 : node36216;
												assign node36216 = (inp[4]) ? node36218 : 4'b0110;
													assign node36218 = (inp[5]) ? 4'b0110 : node36219;
														assign node36219 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node36223 = (inp[5]) ? 4'b0010 : node36224;
													assign node36224 = (inp[4]) ? 4'b0110 : 4'b0011;
							assign node36228 = (inp[2]) ? node36654 : node36229;
								assign node36229 = (inp[7]) ? node36433 : node36230;
									assign node36230 = (inp[5]) ? node36300 : node36231;
										assign node36231 = (inp[4]) ? node36257 : node36232;
											assign node36232 = (inp[10]) ? node36246 : node36233;
												assign node36233 = (inp[13]) ? node36241 : node36234;
													assign node36234 = (inp[0]) ? node36236 : 4'b0101;
														assign node36236 = (inp[1]) ? 4'b0101 : node36237;
															assign node36237 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node36241 = (inp[11]) ? 4'b0100 : node36242;
														assign node36242 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node36246 = (inp[13]) ? node36252 : node36247;
													assign node36247 = (inp[11]) ? 4'b0100 : node36248;
														assign node36248 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node36252 = (inp[1]) ? 4'b0101 : node36253;
														assign node36253 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node36257 = (inp[1]) ? node36265 : node36258;
												assign node36258 = (inp[10]) ? node36262 : node36259;
													assign node36259 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node36262 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node36265 = (inp[0]) ? node36283 : node36266;
													assign node36266 = (inp[13]) ? node36272 : node36267;
														assign node36267 = (inp[9]) ? 4'b0001 : node36268;
															assign node36268 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node36272 = (inp[9]) ? node36278 : node36273;
															assign node36273 = (inp[11]) ? 4'b0001 : node36274;
																assign node36274 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node36278 = (inp[11]) ? 4'b0000 : node36279;
																assign node36279 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node36283 = (inp[10]) ? node36291 : node36284;
														assign node36284 = (inp[13]) ? node36288 : node36285;
															assign node36285 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node36288 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node36291 = (inp[9]) ? node36293 : 4'b0001;
															assign node36293 = (inp[13]) ? node36297 : node36294;
																assign node36294 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node36297 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node36300 = (inp[9]) ? node36368 : node36301;
											assign node36301 = (inp[10]) ? node36333 : node36302;
												assign node36302 = (inp[0]) ? node36322 : node36303;
													assign node36303 = (inp[4]) ? node36313 : node36304;
														assign node36304 = (inp[13]) ? node36310 : node36305;
															assign node36305 = (inp[11]) ? node36307 : 4'b0000;
																assign node36307 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node36310 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node36313 = (inp[13]) ? node36319 : node36314;
															assign node36314 = (inp[11]) ? node36316 : 4'b0001;
																assign node36316 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node36319 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node36322 = (inp[4]) ? node36324 : 4'b0001;
														assign node36324 = (inp[11]) ? node36328 : node36325;
															assign node36325 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node36328 = (inp[13]) ? 4'b0001 : node36329;
																assign node36329 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node36333 = (inp[1]) ? node36353 : node36334;
													assign node36334 = (inp[0]) ? node36348 : node36335;
														assign node36335 = (inp[11]) ? node36343 : node36336;
															assign node36336 = (inp[13]) ? node36340 : node36337;
																assign node36337 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node36340 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node36343 = (inp[4]) ? node36345 : 4'b0000;
																assign node36345 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36348 = (inp[4]) ? 4'b0000 : node36349;
															assign node36349 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node36353 = (inp[4]) ? node36361 : node36354;
														assign node36354 = (inp[11]) ? node36358 : node36355;
															assign node36355 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node36358 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36361 = (inp[0]) ? node36365 : node36362;
															assign node36362 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node36365 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node36368 = (inp[0]) ? node36406 : node36369;
												assign node36369 = (inp[11]) ? node36391 : node36370;
													assign node36370 = (inp[1]) ? node36384 : node36371;
														assign node36371 = (inp[4]) ? node36377 : node36372;
															assign node36372 = (inp[13]) ? 4'b0001 : node36373;
																assign node36373 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node36377 = (inp[10]) ? node36381 : node36378;
																assign node36378 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node36381 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36384 = (inp[10]) ? 4'b0000 : node36385;
															assign node36385 = (inp[13]) ? 4'b0000 : node36386;
																assign node36386 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node36391 = (inp[1]) ? node36393 : 4'b0000;
														assign node36393 = (inp[10]) ? node36399 : node36394;
															assign node36394 = (inp[4]) ? 4'b0000 : node36395;
																assign node36395 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node36399 = (inp[13]) ? node36403 : node36400;
																assign node36400 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node36403 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node36406 = (inp[11]) ? node36414 : node36407;
													assign node36407 = (inp[10]) ? 4'b0000 : node36408;
														assign node36408 = (inp[4]) ? node36410 : 4'b0001;
															assign node36410 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node36414 = (inp[13]) ? node36428 : node36415;
														assign node36415 = (inp[10]) ? node36421 : node36416;
															assign node36416 = (inp[4]) ? node36418 : 4'b0000;
																assign node36418 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node36421 = (inp[1]) ? node36425 : node36422;
																assign node36422 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node36425 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node36428 = (inp[4]) ? 4'b0001 : node36429;
															assign node36429 = (inp[10]) ? 4'b0001 : 4'b0000;
									assign node36433 = (inp[5]) ? node36535 : node36434;
										assign node36434 = (inp[4]) ? node36492 : node36435;
											assign node36435 = (inp[1]) ? node36475 : node36436;
												assign node36436 = (inp[11]) ? node36462 : node36437;
													assign node36437 = (inp[9]) ? node36451 : node36438;
														assign node36438 = (inp[0]) ? node36444 : node36439;
															assign node36439 = (inp[10]) ? node36441 : 4'b0001;
																assign node36441 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node36444 = (inp[10]) ? node36448 : node36445;
																assign node36445 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node36448 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36451 = (inp[0]) ? node36457 : node36452;
															assign node36452 = (inp[10]) ? node36454 : 4'b0000;
																assign node36454 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node36457 = (inp[13]) ? node36459 : 4'b0001;
																assign node36459 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node36462 = (inp[0]) ? node36470 : node36463;
														assign node36463 = (inp[9]) ? 4'b0000 : node36464;
															assign node36464 = (inp[13]) ? node36466 : 4'b0000;
																assign node36466 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node36470 = (inp[13]) ? 4'b0000 : node36471;
															assign node36471 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node36475 = (inp[9]) ? 4'b0001 : node36476;
													assign node36476 = (inp[0]) ? node36484 : node36477;
														assign node36477 = (inp[11]) ? node36479 : 4'b0001;
															assign node36479 = (inp[10]) ? 4'b0000 : node36480;
																assign node36480 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36484 = (inp[13]) ? node36488 : node36485;
															assign node36485 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node36488 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node36492 = (inp[0]) ? node36516 : node36493;
												assign node36493 = (inp[11]) ? node36505 : node36494;
													assign node36494 = (inp[13]) ? 4'b0101 : node36495;
														assign node36495 = (inp[9]) ? node36501 : node36496;
															assign node36496 = (inp[10]) ? node36498 : 4'b0100;
																assign node36498 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node36501 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node36505 = (inp[1]) ? node36511 : node36506;
														assign node36506 = (inp[10]) ? 4'b0100 : node36507;
															assign node36507 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node36511 = (inp[10]) ? node36513 : 4'b0100;
															assign node36513 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node36516 = (inp[10]) ? node36528 : node36517;
													assign node36517 = (inp[1]) ? 4'b0101 : node36518;
														assign node36518 = (inp[9]) ? node36520 : 4'b0101;
															assign node36520 = (inp[11]) ? node36524 : node36521;
																assign node36521 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node36524 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node36528 = (inp[13]) ? 4'b0100 : node36529;
														assign node36529 = (inp[11]) ? 4'b0101 : node36530;
															assign node36530 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node36535 = (inp[9]) ? node36611 : node36536;
											assign node36536 = (inp[13]) ? node36568 : node36537;
												assign node36537 = (inp[1]) ? node36561 : node36538;
													assign node36538 = (inp[0]) ? node36552 : node36539;
														assign node36539 = (inp[11]) ? node36545 : node36540;
															assign node36540 = (inp[10]) ? node36542 : 4'b0100;
																assign node36542 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node36545 = (inp[4]) ? node36549 : node36546;
																assign node36546 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node36549 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node36552 = (inp[11]) ? node36554 : 4'b0101;
															assign node36554 = (inp[10]) ? node36558 : node36555;
																assign node36555 = (inp[4]) ? 4'b0100 : 4'b0101;
																assign node36558 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node36561 = (inp[4]) ? node36565 : node36562;
														assign node36562 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node36565 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node36568 = (inp[11]) ? node36596 : node36569;
													assign node36569 = (inp[0]) ? node36583 : node36570;
														assign node36570 = (inp[10]) ? node36576 : node36571;
															assign node36571 = (inp[1]) ? node36573 : 4'b0101;
																assign node36573 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node36576 = (inp[4]) ? node36580 : node36577;
																assign node36577 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node36580 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node36583 = (inp[1]) ? node36591 : node36584;
															assign node36584 = (inp[4]) ? node36588 : node36585;
																assign node36585 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node36588 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node36591 = (inp[10]) ? node36593 : 4'b0100;
																assign node36593 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node36596 = (inp[0]) ? node36604 : node36597;
														assign node36597 = (inp[10]) ? node36601 : node36598;
															assign node36598 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node36601 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node36604 = (inp[4]) ? node36608 : node36605;
															assign node36605 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node36608 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node36611 = (inp[10]) ? node36635 : node36612;
												assign node36612 = (inp[1]) ? node36630 : node36613;
													assign node36613 = (inp[0]) ? node36621 : node36614;
														assign node36614 = (inp[13]) ? 4'b0101 : node36615;
															assign node36615 = (inp[11]) ? 4'b0100 : node36616;
																assign node36616 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node36621 = (inp[4]) ? 4'b0100 : node36622;
															assign node36622 = (inp[11]) ? node36626 : node36623;
																assign node36623 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node36626 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node36630 = (inp[4]) ? node36632 : 4'b0100;
														assign node36632 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node36635 = (inp[13]) ? node36647 : node36636;
													assign node36636 = (inp[4]) ? node36642 : node36637;
														assign node36637 = (inp[1]) ? 4'b0100 : node36638;
															assign node36638 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node36642 = (inp[11]) ? 4'b0101 : node36643;
															assign node36643 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node36647 = (inp[4]) ? 4'b0100 : node36648;
														assign node36648 = (inp[1]) ? 4'b0101 : node36649;
															assign node36649 = (inp[11]) ? 4'b0101 : 4'b0100;
								assign node36654 = (inp[7]) ? node36790 : node36655;
									assign node36655 = (inp[4]) ? node36737 : node36656;
										assign node36656 = (inp[5]) ? node36700 : node36657;
											assign node36657 = (inp[11]) ? node36687 : node36658;
												assign node36658 = (inp[9]) ? node36670 : node36659;
													assign node36659 = (inp[1]) ? node36665 : node36660;
														assign node36660 = (inp[10]) ? node36662 : 4'b0000;
															assign node36662 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node36665 = (inp[13]) ? node36667 : 4'b0001;
															assign node36667 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node36670 = (inp[13]) ? node36676 : node36671;
														assign node36671 = (inp[1]) ? 4'b0000 : node36672;
															assign node36672 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node36676 = (inp[0]) ? node36682 : node36677;
															assign node36677 = (inp[1]) ? node36679 : 4'b0000;
																assign node36679 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node36682 = (inp[10]) ? 4'b0001 : node36683;
																assign node36683 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node36687 = (inp[9]) ? node36695 : node36688;
													assign node36688 = (inp[13]) ? node36692 : node36689;
														assign node36689 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node36692 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node36695 = (inp[10]) ? 4'b0001 : node36696;
														assign node36696 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node36700 = (inp[1]) ? node36730 : node36701;
												assign node36701 = (inp[9]) ? node36709 : node36702;
													assign node36702 = (inp[10]) ? 4'b0101 : node36703;
														assign node36703 = (inp[11]) ? 4'b0101 : node36704;
															assign node36704 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node36709 = (inp[0]) ? node36717 : node36710;
														assign node36710 = (inp[13]) ? node36712 : 4'b0101;
															assign node36712 = (inp[11]) ? node36714 : 4'b0101;
																assign node36714 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node36717 = (inp[10]) ? node36723 : node36718;
															assign node36718 = (inp[11]) ? 4'b0100 : node36719;
																assign node36719 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node36723 = (inp[13]) ? node36727 : node36724;
																assign node36724 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node36727 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node36730 = (inp[10]) ? node36734 : node36731;
													assign node36731 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node36734 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node36737 = (inp[13]) ? node36767 : node36738;
											assign node36738 = (inp[1]) ? node36760 : node36739;
												assign node36739 = (inp[11]) ? node36753 : node36740;
													assign node36740 = (inp[9]) ? node36748 : node36741;
														assign node36741 = (inp[10]) ? node36745 : node36742;
															assign node36742 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node36745 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node36748 = (inp[0]) ? 4'b0100 : node36749;
															assign node36749 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node36753 = (inp[5]) ? node36757 : node36754;
														assign node36754 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node36757 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node36760 = (inp[5]) ? node36764 : node36761;
													assign node36761 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node36764 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node36767 = (inp[5]) ? node36779 : node36768;
												assign node36768 = (inp[10]) ? node36774 : node36769;
													assign node36769 = (inp[11]) ? 4'b0100 : node36770;
														assign node36770 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node36774 = (inp[11]) ? 4'b0101 : node36775;
														assign node36775 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node36779 = (inp[10]) ? node36785 : node36780;
													assign node36780 = (inp[11]) ? 4'b0101 : node36781;
														assign node36781 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node36785 = (inp[1]) ? 4'b0100 : node36786;
														assign node36786 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node36790 = (inp[4]) ? node36838 : node36791;
										assign node36791 = (inp[5]) ? node36815 : node36792;
											assign node36792 = (inp[1]) ? node36800 : node36793;
												assign node36793 = (inp[10]) ? node36797 : node36794;
													assign node36794 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node36797 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node36800 = (inp[11]) ? node36808 : node36801;
													assign node36801 = (inp[10]) ? node36805 : node36802;
														assign node36802 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node36805 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node36808 = (inp[13]) ? node36812 : node36809;
														assign node36809 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node36812 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node36815 = (inp[13]) ? node36827 : node36816;
												assign node36816 = (inp[10]) ? node36822 : node36817;
													assign node36817 = (inp[11]) ? 4'b0000 : node36818;
														assign node36818 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node36822 = (inp[11]) ? 4'b0001 : node36823;
														assign node36823 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node36827 = (inp[10]) ? node36833 : node36828;
													assign node36828 = (inp[11]) ? 4'b0001 : node36829;
														assign node36829 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node36833 = (inp[1]) ? 4'b0000 : node36834;
														assign node36834 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node36838 = (inp[9]) ? node36910 : node36839;
											assign node36839 = (inp[0]) ? node36875 : node36840;
												assign node36840 = (inp[11]) ? node36862 : node36841;
													assign node36841 = (inp[5]) ? node36851 : node36842;
														assign node36842 = (inp[1]) ? node36844 : 4'b0000;
															assign node36844 = (inp[10]) ? node36848 : node36845;
																assign node36845 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node36848 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node36851 = (inp[1]) ? node36857 : node36852;
															assign node36852 = (inp[13]) ? 4'b0001 : node36853;
																assign node36853 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node36857 = (inp[13]) ? 4'b0000 : node36858;
																assign node36858 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node36862 = (inp[1]) ? node36870 : node36863;
														assign node36863 = (inp[10]) ? node36867 : node36864;
															assign node36864 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node36867 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node36870 = (inp[10]) ? 4'b0001 : node36871;
															assign node36871 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node36875 = (inp[11]) ? node36903 : node36876;
													assign node36876 = (inp[5]) ? node36890 : node36877;
														assign node36877 = (inp[13]) ? node36885 : node36878;
															assign node36878 = (inp[10]) ? node36882 : node36879;
																assign node36879 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node36882 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node36885 = (inp[10]) ? node36887 : 4'b0001;
																assign node36887 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node36890 = (inp[1]) ? node36896 : node36891;
															assign node36891 = (inp[10]) ? 4'b0000 : node36892;
																assign node36892 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node36896 = (inp[13]) ? node36900 : node36897;
																assign node36897 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node36900 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node36903 = (inp[13]) ? node36907 : node36904;
														assign node36904 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node36907 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node36910 = (inp[5]) ? node36932 : node36911;
												assign node36911 = (inp[11]) ? node36925 : node36912;
													assign node36912 = (inp[13]) ? node36920 : node36913;
														assign node36913 = (inp[10]) ? node36917 : node36914;
															assign node36914 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node36917 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node36920 = (inp[10]) ? node36922 : 4'b0001;
															assign node36922 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node36925 = (inp[13]) ? node36929 : node36926;
														assign node36926 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node36929 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node36932 = (inp[13]) ? node36940 : node36933;
													assign node36933 = (inp[10]) ? 4'b0001 : node36934;
														assign node36934 = (inp[11]) ? 4'b0000 : node36935;
															assign node36935 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node36940 = (inp[10]) ? node36946 : node36941;
														assign node36941 = (inp[1]) ? 4'b0001 : node36942;
															assign node36942 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node36946 = (inp[1]) ? 4'b0000 : node36947;
															assign node36947 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node36951 = (inp[2]) ? node37497 : node36952;
							assign node36952 = (inp[14]) ? node37196 : node36953;
								assign node36953 = (inp[5]) ? node37121 : node36954;
									assign node36954 = (inp[9]) ? node37038 : node36955;
										assign node36955 = (inp[1]) ? node36995 : node36956;
											assign node36956 = (inp[13]) ? node36978 : node36957;
												assign node36957 = (inp[11]) ? node36965 : node36958;
													assign node36958 = (inp[10]) ? node36962 : node36959;
														assign node36959 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node36962 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node36965 = (inp[10]) ? node36973 : node36966;
														assign node36966 = (inp[4]) ? node36970 : node36967;
															assign node36967 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node36970 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node36973 = (inp[7]) ? node36975 : 4'b0000;
															assign node36975 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node36978 = (inp[10]) ? node36988 : node36979;
													assign node36979 = (inp[7]) ? node36985 : node36980;
														assign node36980 = (inp[4]) ? node36982 : 4'b0000;
															assign node36982 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node36985 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node36988 = (inp[7]) ? node36990 : 4'b0001;
														assign node36990 = (inp[11]) ? node36992 : 4'b0000;
															assign node36992 = (inp[4]) ? 4'b0001 : 4'b0000;
											assign node36995 = (inp[13]) ? node37017 : node36996;
												assign node36996 = (inp[10]) ? node37008 : node36997;
													assign node36997 = (inp[7]) ? node37003 : node36998;
														assign node36998 = (inp[11]) ? node37000 : 4'b0000;
															assign node37000 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node37003 = (inp[11]) ? node37005 : 4'b0001;
															assign node37005 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node37008 = (inp[11]) ? node37010 : 4'b0000;
														assign node37010 = (inp[7]) ? node37014 : node37011;
															assign node37011 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node37014 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node37017 = (inp[7]) ? node37027 : node37018;
													assign node37018 = (inp[10]) ? node37022 : node37019;
														assign node37019 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node37022 = (inp[11]) ? node37024 : 4'b0001;
															assign node37024 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node37027 = (inp[10]) ? node37033 : node37028;
														assign node37028 = (inp[4]) ? node37030 : 4'b0001;
															assign node37030 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node37033 = (inp[4]) ? node37035 : 4'b0000;
															assign node37035 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node37038 = (inp[11]) ? node37062 : node37039;
											assign node37039 = (inp[13]) ? node37055 : node37040;
												assign node37040 = (inp[4]) ? node37048 : node37041;
													assign node37041 = (inp[7]) ? node37045 : node37042;
														assign node37042 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node37045 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node37048 = (inp[10]) ? node37052 : node37049;
														assign node37049 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37052 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node37055 = (inp[7]) ? node37059 : node37056;
													assign node37056 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node37059 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node37062 = (inp[1]) ? node37104 : node37063;
												assign node37063 = (inp[13]) ? node37085 : node37064;
													assign node37064 = (inp[0]) ? node37074 : node37065;
														assign node37065 = (inp[10]) ? node37067 : 4'b0001;
															assign node37067 = (inp[4]) ? node37071 : node37068;
																assign node37068 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node37071 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37074 = (inp[10]) ? node37080 : node37075;
															assign node37075 = (inp[4]) ? node37077 : 4'b0000;
																assign node37077 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node37080 = (inp[7]) ? 4'b0001 : node37081;
																assign node37081 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node37085 = (inp[10]) ? node37091 : node37086;
														assign node37086 = (inp[4]) ? 4'b0000 : node37087;
															assign node37087 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37091 = (inp[0]) ? node37099 : node37092;
															assign node37092 = (inp[4]) ? node37096 : node37093;
																assign node37093 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node37096 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37099 = (inp[4]) ? 4'b0001 : node37100;
																assign node37100 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node37104 = (inp[10]) ? node37114 : node37105;
													assign node37105 = (inp[13]) ? 4'b0001 : node37106;
														assign node37106 = (inp[4]) ? node37110 : node37107;
															assign node37107 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37110 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node37114 = (inp[4]) ? node37118 : node37115;
														assign node37115 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node37118 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node37121 = (inp[11]) ? node37165 : node37122;
										assign node37122 = (inp[13]) ? node37158 : node37123;
											assign node37123 = (inp[7]) ? node37131 : node37124;
												assign node37124 = (inp[4]) ? node37128 : node37125;
													assign node37125 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node37128 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node37131 = (inp[1]) ? node37139 : node37132;
													assign node37132 = (inp[4]) ? node37136 : node37133;
														assign node37133 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37136 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node37139 = (inp[9]) ? node37149 : node37140;
														assign node37140 = (inp[0]) ? node37142 : 4'b0100;
															assign node37142 = (inp[4]) ? node37146 : node37143;
																assign node37143 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node37146 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node37149 = (inp[0]) ? node37151 : 4'b0101;
															assign node37151 = (inp[4]) ? node37155 : node37152;
																assign node37152 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node37155 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node37158 = (inp[4]) ? node37162 : node37159;
												assign node37159 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node37162 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node37165 = (inp[9]) ? node37173 : node37166;
											assign node37166 = (inp[4]) ? node37170 : node37167;
												assign node37167 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node37170 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node37173 = (inp[1]) ? node37189 : node37174;
												assign node37174 = (inp[13]) ? node37182 : node37175;
													assign node37175 = (inp[4]) ? node37179 : node37176;
														assign node37176 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37179 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node37182 = (inp[4]) ? node37186 : node37183;
														assign node37183 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37186 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node37189 = (inp[10]) ? node37193 : node37190;
													assign node37190 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node37193 = (inp[4]) ? 4'b0100 : 4'b0101;
								assign node37196 = (inp[5]) ? node37338 : node37197;
									assign node37197 = (inp[1]) ? node37245 : node37198;
										assign node37198 = (inp[13]) ? node37222 : node37199;
											assign node37199 = (inp[7]) ? node37211 : node37200;
												assign node37200 = (inp[10]) ? node37206 : node37201;
													assign node37201 = (inp[4]) ? 4'b0100 : node37202;
														assign node37202 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node37206 = (inp[11]) ? node37208 : 4'b0101;
														assign node37208 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node37211 = (inp[10]) ? node37217 : node37212;
													assign node37212 = (inp[4]) ? 4'b0101 : node37213;
														assign node37213 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node37217 = (inp[11]) ? node37219 : 4'b0100;
														assign node37219 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node37222 = (inp[7]) ? node37234 : node37223;
												assign node37223 = (inp[10]) ? node37229 : node37224;
													assign node37224 = (inp[4]) ? 4'b0100 : node37225;
														assign node37225 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node37229 = (inp[4]) ? 4'b0101 : node37230;
														assign node37230 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node37234 = (inp[10]) ? node37240 : node37235;
													assign node37235 = (inp[4]) ? 4'b0101 : node37236;
														assign node37236 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node37240 = (inp[11]) ? node37242 : 4'b0100;
														assign node37242 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node37245 = (inp[0]) ? node37301 : node37246;
											assign node37246 = (inp[9]) ? node37282 : node37247;
												assign node37247 = (inp[11]) ? node37269 : node37248;
													assign node37248 = (inp[4]) ? node37262 : node37249;
														assign node37249 = (inp[13]) ? node37255 : node37250;
															assign node37250 = (inp[7]) ? 4'b0100 : node37251;
																assign node37251 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node37255 = (inp[10]) ? node37259 : node37256;
																assign node37256 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node37259 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node37262 = (inp[7]) ? node37266 : node37263;
															assign node37263 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node37266 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node37269 = (inp[4]) ? node37277 : node37270;
														assign node37270 = (inp[10]) ? node37274 : node37271;
															assign node37271 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node37274 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node37277 = (inp[10]) ? node37279 : 4'b0100;
															assign node37279 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node37282 = (inp[7]) ? node37292 : node37283;
													assign node37283 = (inp[10]) ? node37289 : node37284;
														assign node37284 = (inp[11]) ? node37286 : 4'b0100;
															assign node37286 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node37289 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node37292 = (inp[4]) ? 4'b0100 : node37293;
														assign node37293 = (inp[10]) ? node37297 : node37294;
															assign node37294 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node37297 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node37301 = (inp[4]) ? node37331 : node37302;
												assign node37302 = (inp[9]) ? node37316 : node37303;
													assign node37303 = (inp[7]) ? node37311 : node37304;
														assign node37304 = (inp[10]) ? node37308 : node37305;
															assign node37305 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node37308 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node37311 = (inp[10]) ? 4'b0100 : node37312;
															assign node37312 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node37316 = (inp[10]) ? node37324 : node37317;
														assign node37317 = (inp[11]) ? node37321 : node37318;
															assign node37318 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node37321 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node37324 = (inp[11]) ? node37328 : node37325;
															assign node37325 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node37328 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node37331 = (inp[7]) ? node37335 : node37332;
													assign node37332 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node37335 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node37338 = (inp[13]) ? node37404 : node37339;
										assign node37339 = (inp[0]) ? node37397 : node37340;
											assign node37340 = (inp[7]) ? node37362 : node37341;
												assign node37341 = (inp[11]) ? node37349 : node37342;
													assign node37342 = (inp[10]) ? node37346 : node37343;
														assign node37343 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node37346 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node37349 = (inp[1]) ? node37355 : node37350;
														assign node37350 = (inp[10]) ? node37352 : 4'b0101;
															assign node37352 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node37355 = (inp[10]) ? node37359 : node37356;
															assign node37356 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node37359 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node37362 = (inp[9]) ? node37390 : node37363;
													assign node37363 = (inp[1]) ? node37377 : node37364;
														assign node37364 = (inp[11]) ? node37372 : node37365;
															assign node37365 = (inp[10]) ? node37369 : node37366;
																assign node37366 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node37369 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node37372 = (inp[4]) ? 4'b0100 : node37373;
																assign node37373 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37377 = (inp[11]) ? node37385 : node37378;
															assign node37378 = (inp[10]) ? node37382 : node37379;
																assign node37379 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node37382 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node37385 = (inp[4]) ? 4'b0101 : node37386;
																assign node37386 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node37390 = (inp[4]) ? node37394 : node37391;
														assign node37391 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37394 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node37397 = (inp[4]) ? node37401 : node37398;
												assign node37398 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node37401 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node37404 = (inp[0]) ? node37440 : node37405;
											assign node37405 = (inp[9]) ? node37413 : node37406;
												assign node37406 = (inp[10]) ? node37410 : node37407;
													assign node37407 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node37410 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node37413 = (inp[1]) ? node37431 : node37414;
													assign node37414 = (inp[7]) ? node37424 : node37415;
														assign node37415 = (inp[11]) ? node37417 : 4'b0100;
															assign node37417 = (inp[10]) ? node37421 : node37418;
																assign node37418 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node37421 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node37424 = (inp[10]) ? node37428 : node37425;
															assign node37425 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node37428 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node37431 = (inp[7]) ? 4'b0100 : node37432;
														assign node37432 = (inp[4]) ? node37436 : node37433;
															assign node37433 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node37436 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node37440 = (inp[7]) ? node37460 : node37441;
												assign node37441 = (inp[1]) ? node37453 : node37442;
													assign node37442 = (inp[9]) ? node37444 : 4'b0101;
														assign node37444 = (inp[11]) ? node37448 : node37445;
															assign node37445 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node37448 = (inp[10]) ? 4'b0101 : node37449;
																assign node37449 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node37453 = (inp[4]) ? node37457 : node37454;
														assign node37454 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node37457 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node37460 = (inp[11]) ? node37484 : node37461;
													assign node37461 = (inp[1]) ? node37477 : node37462;
														assign node37462 = (inp[9]) ? node37470 : node37463;
															assign node37463 = (inp[4]) ? node37467 : node37464;
																assign node37464 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node37467 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node37470 = (inp[10]) ? node37474 : node37471;
																assign node37471 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node37474 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node37477 = (inp[10]) ? node37481 : node37478;
															assign node37478 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node37481 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node37484 = (inp[9]) ? node37492 : node37485;
														assign node37485 = (inp[4]) ? node37489 : node37486;
															assign node37486 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node37489 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node37492 = (inp[10]) ? node37494 : 4'b0101;
															assign node37494 = (inp[4]) ? 4'b0100 : 4'b0101;
							assign node37497 = (inp[5]) ? node37767 : node37498;
								assign node37498 = (inp[14]) ? node37634 : node37499;
									assign node37499 = (inp[4]) ? node37515 : node37500;
										assign node37500 = (inp[1]) ? node37508 : node37501;
											assign node37501 = (inp[7]) ? node37505 : node37502;
												assign node37502 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node37505 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node37508 = (inp[7]) ? node37512 : node37509;
												assign node37509 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node37512 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node37515 = (inp[1]) ? node37573 : node37516;
											assign node37516 = (inp[9]) ? node37542 : node37517;
												assign node37517 = (inp[11]) ? node37523 : node37518;
													assign node37518 = (inp[7]) ? 4'b0100 : node37519;
														assign node37519 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node37523 = (inp[13]) ? node37531 : node37524;
														assign node37524 = (inp[7]) ? node37528 : node37525;
															assign node37525 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37528 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node37531 = (inp[0]) ? node37537 : node37532;
															assign node37532 = (inp[7]) ? 4'b0100 : node37533;
																assign node37533 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node37537 = (inp[7]) ? node37539 : 4'b0100;
																assign node37539 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node37542 = (inp[10]) ? node37550 : node37543;
													assign node37543 = (inp[7]) ? node37547 : node37544;
														assign node37544 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node37547 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node37550 = (inp[13]) ? node37566 : node37551;
														assign node37551 = (inp[0]) ? node37559 : node37552;
															assign node37552 = (inp[7]) ? node37556 : node37553;
																assign node37553 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node37556 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node37559 = (inp[7]) ? node37563 : node37560;
																assign node37560 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node37563 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node37566 = (inp[7]) ? node37570 : node37567;
															assign node37567 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node37570 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node37573 = (inp[10]) ? node37611 : node37574;
												assign node37574 = (inp[13]) ? node37588 : node37575;
													assign node37575 = (inp[9]) ? node37583 : node37576;
														assign node37576 = (inp[11]) ? node37580 : node37577;
															assign node37577 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node37580 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node37583 = (inp[0]) ? node37585 : 4'b0101;
															assign node37585 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node37588 = (inp[9]) ? node37596 : node37589;
														assign node37589 = (inp[11]) ? node37593 : node37590;
															assign node37590 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node37593 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node37596 = (inp[0]) ? node37604 : node37597;
															assign node37597 = (inp[11]) ? node37601 : node37598;
																assign node37598 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node37601 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node37604 = (inp[7]) ? node37608 : node37605;
																assign node37605 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node37608 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node37611 = (inp[0]) ? node37625 : node37612;
													assign node37612 = (inp[13]) ? node37620 : node37613;
														assign node37613 = (inp[7]) ? node37617 : node37614;
															assign node37614 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node37617 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node37620 = (inp[11]) ? 4'b0101 : node37621;
															assign node37621 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node37625 = (inp[13]) ? node37627 : 4'b0101;
														assign node37627 = (inp[9]) ? node37629 : 4'b0101;
															assign node37629 = (inp[7]) ? node37631 : 4'b0100;
																assign node37631 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node37634 = (inp[1]) ? node37700 : node37635;
										assign node37635 = (inp[11]) ? node37673 : node37636;
											assign node37636 = (inp[9]) ? node37660 : node37637;
												assign node37637 = (inp[4]) ? node37653 : node37638;
													assign node37638 = (inp[0]) ? node37646 : node37639;
														assign node37639 = (inp[13]) ? 4'b0000 : node37640;
															assign node37640 = (inp[10]) ? node37642 : 4'b0000;
																assign node37642 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37646 = (inp[7]) ? node37650 : node37647;
															assign node37647 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node37650 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node37653 = (inp[7]) ? node37657 : node37654;
														assign node37654 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node37657 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node37660 = (inp[4]) ? node37666 : node37661;
													assign node37661 = (inp[7]) ? 4'b0001 : node37662;
														assign node37662 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node37666 = (inp[10]) ? node37670 : node37667;
														assign node37667 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37670 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node37673 = (inp[4]) ? node37681 : node37674;
												assign node37674 = (inp[7]) ? node37678 : node37675;
													assign node37675 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node37678 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node37681 = (inp[0]) ? node37695 : node37682;
													assign node37682 = (inp[13]) ? node37688 : node37683;
														assign node37683 = (inp[10]) ? 4'b0001 : node37684;
															assign node37684 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node37688 = (inp[10]) ? node37692 : node37689;
															assign node37689 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37692 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node37695 = (inp[10]) ? node37697 : 4'b0001;
														assign node37697 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node37700 = (inp[4]) ? node37724 : node37701;
											assign node37701 = (inp[7]) ? node37709 : node37702;
												assign node37702 = (inp[10]) ? node37706 : node37703;
													assign node37703 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node37706 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node37709 = (inp[13]) ? node37717 : node37710;
													assign node37710 = (inp[10]) ? node37714 : node37711;
														assign node37711 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node37714 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node37717 = (inp[10]) ? node37721 : node37718;
														assign node37718 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node37721 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node37724 = (inp[0]) ? node37746 : node37725;
												assign node37725 = (inp[11]) ? node37733 : node37726;
													assign node37726 = (inp[7]) ? node37730 : node37727;
														assign node37727 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node37730 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node37733 = (inp[9]) ? node37741 : node37734;
														assign node37734 = (inp[10]) ? node37738 : node37735;
															assign node37735 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37738 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node37741 = (inp[7]) ? 4'b0000 : node37742;
															assign node37742 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node37746 = (inp[11]) ? node37754 : node37747;
													assign node37747 = (inp[10]) ? node37751 : node37748;
														assign node37748 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node37751 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node37754 = (inp[9]) ? node37762 : node37755;
														assign node37755 = (inp[13]) ? 4'b0000 : node37756;
															assign node37756 = (inp[7]) ? node37758 : 4'b0001;
																assign node37758 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node37762 = (inp[13]) ? 4'b0001 : node37763;
															assign node37763 = (inp[10]) ? 4'b0001 : 4'b0000;
								assign node37767 = (inp[10]) ? node37773 : node37768;
									assign node37768 = (inp[11]) ? 4'b0001 : node37769;
										assign node37769 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node37773 = (inp[11]) ? 4'b0000 : node37774;
										assign node37774 = (inp[14]) ? 4'b0000 : 4'b0001;
			assign node37778 = (inp[3]) ? node41592 : node37779;
				assign node37779 = (inp[4]) ? node39957 : node37780;
					assign node37780 = (inp[15]) ? node39202 : node37781;
						assign node37781 = (inp[14]) ? node38561 : node37782;
							assign node37782 = (inp[10]) ? node38174 : node37783;
								assign node37783 = (inp[1]) ? node37967 : node37784;
									assign node37784 = (inp[5]) ? node37850 : node37785;
										assign node37785 = (inp[12]) ? node37809 : node37786;
											assign node37786 = (inp[13]) ? node37794 : node37787;
												assign node37787 = (inp[0]) ? node37791 : node37788;
													assign node37788 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node37791 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node37794 = (inp[2]) ? node37802 : node37795;
													assign node37795 = (inp[0]) ? node37799 : node37796;
														assign node37796 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node37799 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node37802 = (inp[0]) ? node37806 : node37803;
														assign node37803 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node37806 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node37809 = (inp[7]) ? node37823 : node37810;
												assign node37810 = (inp[11]) ? node37816 : node37811;
													assign node37811 = (inp[0]) ? 4'b0001 : node37812;
														assign node37812 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node37816 = (inp[0]) ? node37818 : 4'b0001;
														assign node37818 = (inp[2]) ? node37820 : 4'b0000;
															assign node37820 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node37823 = (inp[11]) ? node37839 : node37824;
													assign node37824 = (inp[9]) ? node37830 : node37825;
														assign node37825 = (inp[2]) ? 4'b0100 : node37826;
															assign node37826 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node37830 = (inp[0]) ? node37836 : node37831;
															assign node37831 = (inp[13]) ? 4'b0101 : node37832;
																assign node37832 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node37836 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node37839 = (inp[0]) ? node37845 : node37840;
														assign node37840 = (inp[13]) ? 4'b0100 : node37841;
															assign node37841 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node37845 = (inp[2]) ? 4'b0101 : node37846;
															assign node37846 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node37850 = (inp[7]) ? node37896 : node37851;
											assign node37851 = (inp[9]) ? node37873 : node37852;
												assign node37852 = (inp[11]) ? node37862 : node37853;
													assign node37853 = (inp[2]) ? node37855 : 4'b0100;
														assign node37855 = (inp[13]) ? node37859 : node37856;
															assign node37856 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37859 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node37862 = (inp[0]) ? node37868 : node37863;
														assign node37863 = (inp[2]) ? node37865 : 4'b0101;
															assign node37865 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node37868 = (inp[13]) ? node37870 : 4'b0100;
															assign node37870 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node37873 = (inp[0]) ? node37885 : node37874;
													assign node37874 = (inp[11]) ? node37880 : node37875;
														assign node37875 = (inp[2]) ? node37877 : 4'b0100;
															assign node37877 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node37880 = (inp[2]) ? node37882 : 4'b0101;
															assign node37882 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node37885 = (inp[11]) ? node37891 : node37886;
														assign node37886 = (inp[2]) ? node37888 : 4'b0101;
															assign node37888 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node37891 = (inp[2]) ? node37893 : 4'b0100;
															assign node37893 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node37896 = (inp[12]) ? node37936 : node37897;
												assign node37897 = (inp[2]) ? node37913 : node37898;
													assign node37898 = (inp[13]) ? node37908 : node37899;
														assign node37899 = (inp[9]) ? node37905 : node37900;
															assign node37900 = (inp[11]) ? 4'b0100 : node37901;
																assign node37901 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node37905 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node37908 = (inp[11]) ? 4'b0101 : node37909;
															assign node37909 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node37913 = (inp[13]) ? node37927 : node37914;
														assign node37914 = (inp[9]) ? node37922 : node37915;
															assign node37915 = (inp[11]) ? node37919 : node37916;
																assign node37916 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node37919 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37922 = (inp[11]) ? 4'b0100 : node37923;
																assign node37923 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node37927 = (inp[9]) ? node37929 : 4'b0100;
															assign node37929 = (inp[11]) ? node37933 : node37930;
																assign node37930 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node37933 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node37936 = (inp[13]) ? node37954 : node37937;
													assign node37937 = (inp[9]) ? node37939 : 4'b0001;
														assign node37939 = (inp[2]) ? node37947 : node37940;
															assign node37940 = (inp[0]) ? node37944 : node37941;
																assign node37941 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node37944 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node37947 = (inp[0]) ? node37951 : node37948;
																assign node37948 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node37951 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node37954 = (inp[2]) ? node37960 : node37955;
														assign node37955 = (inp[11]) ? node37957 : 4'b0000;
															assign node37957 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node37960 = (inp[11]) ? node37964 : node37961;
															assign node37961 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node37964 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node37967 = (inp[5]) ? node38073 : node37968;
										assign node37968 = (inp[7]) ? node38036 : node37969;
											assign node37969 = (inp[13]) ? node38005 : node37970;
												assign node37970 = (inp[2]) ? node37990 : node37971;
													assign node37971 = (inp[11]) ? node37981 : node37972;
														assign node37972 = (inp[9]) ? node37974 : 4'b0101;
															assign node37974 = (inp[0]) ? node37978 : node37975;
																assign node37975 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node37978 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node37981 = (inp[9]) ? 4'b0101 : node37982;
															assign node37982 = (inp[0]) ? node37986 : node37983;
																assign node37983 = (inp[12]) ? 4'b0100 : 4'b0101;
																assign node37986 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node37990 = (inp[11]) ? node37998 : node37991;
														assign node37991 = (inp[0]) ? node37995 : node37992;
															assign node37992 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node37995 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node37998 = (inp[0]) ? node38002 : node37999;
															assign node37999 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node38002 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node38005 = (inp[11]) ? node38021 : node38006;
													assign node38006 = (inp[2]) ? node38014 : node38007;
														assign node38007 = (inp[0]) ? node38011 : node38008;
															assign node38008 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node38011 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node38014 = (inp[12]) ? node38018 : node38015;
															assign node38015 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38018 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node38021 = (inp[2]) ? node38029 : node38022;
														assign node38022 = (inp[12]) ? node38026 : node38023;
															assign node38023 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38026 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38029 = (inp[12]) ? node38033 : node38030;
															assign node38030 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38033 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node38036 = (inp[12]) ? node38056 : node38037;
												assign node38037 = (inp[0]) ? node38047 : node38038;
													assign node38038 = (inp[11]) ? node38044 : node38039;
														assign node38039 = (inp[2]) ? node38041 : 4'b0100;
															assign node38041 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node38044 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node38047 = (inp[11]) ? node38053 : node38048;
														assign node38048 = (inp[13]) ? node38050 : 4'b0101;
															assign node38050 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node38053 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node38056 = (inp[11]) ? node38066 : node38057;
													assign node38057 = (inp[0]) ? node38063 : node38058;
														assign node38058 = (inp[13]) ? node38060 : 4'b0000;
															assign node38060 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node38063 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node38066 = (inp[0]) ? node38068 : 4'b0001;
														assign node38068 = (inp[2]) ? node38070 : 4'b0000;
															assign node38070 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node38073 = (inp[7]) ? node38129 : node38074;
											assign node38074 = (inp[11]) ? node38102 : node38075;
												assign node38075 = (inp[2]) ? node38087 : node38076;
													assign node38076 = (inp[0]) ? 4'b0001 : node38077;
														assign node38077 = (inp[9]) ? node38079 : 4'b0001;
															assign node38079 = (inp[13]) ? node38083 : node38080;
																assign node38080 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node38083 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node38087 = (inp[13]) ? node38095 : node38088;
														assign node38088 = (inp[0]) ? node38092 : node38089;
															assign node38089 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node38092 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node38095 = (inp[0]) ? node38099 : node38096;
															assign node38096 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node38099 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node38102 = (inp[2]) ? node38120 : node38103;
													assign node38103 = (inp[0]) ? node38111 : node38104;
														assign node38104 = (inp[13]) ? node38108 : node38105;
															assign node38105 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node38108 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node38111 = (inp[9]) ? node38113 : 4'b0001;
															assign node38113 = (inp[13]) ? node38117 : node38114;
																assign node38114 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node38117 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node38120 = (inp[13]) ? node38122 : 4'b0000;
														assign node38122 = (inp[0]) ? node38126 : node38123;
															assign node38123 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node38126 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node38129 = (inp[12]) ? node38155 : node38130;
												assign node38130 = (inp[13]) ? node38148 : node38131;
													assign node38131 = (inp[0]) ? node38139 : node38132;
														assign node38132 = (inp[9]) ? node38134 : 4'b0000;
															assign node38134 = (inp[2]) ? node38136 : 4'b0001;
																assign node38136 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node38139 = (inp[9]) ? node38141 : 4'b0001;
															assign node38141 = (inp[2]) ? node38145 : node38142;
																assign node38142 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node38145 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node38148 = (inp[11]) ? node38152 : node38149;
														assign node38149 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node38152 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node38155 = (inp[11]) ? node38163 : node38156;
													assign node38156 = (inp[0]) ? 4'b0100 : node38157;
														assign node38157 = (inp[13]) ? node38159 : 4'b0101;
															assign node38159 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node38163 = (inp[0]) ? node38169 : node38164;
														assign node38164 = (inp[13]) ? node38166 : 4'b0100;
															assign node38166 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node38169 = (inp[13]) ? node38171 : 4'b0101;
															assign node38171 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node38174 = (inp[5]) ? node38372 : node38175;
									assign node38175 = (inp[1]) ? node38251 : node38176;
										assign node38176 = (inp[12]) ? node38198 : node38177;
											assign node38177 = (inp[0]) ? node38187 : node38178;
												assign node38178 = (inp[11]) ? node38184 : node38179;
													assign node38179 = (inp[13]) ? node38181 : 4'b0000;
														assign node38181 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node38184 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node38187 = (inp[11]) ? node38193 : node38188;
													assign node38188 = (inp[2]) ? node38190 : 4'b0001;
														assign node38190 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node38193 = (inp[2]) ? node38195 : 4'b0000;
														assign node38195 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node38198 = (inp[7]) ? node38222 : node38199;
												assign node38199 = (inp[13]) ? node38207 : node38200;
													assign node38200 = (inp[11]) ? node38204 : node38201;
														assign node38201 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node38204 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node38207 = (inp[9]) ? node38215 : node38208;
														assign node38208 = (inp[2]) ? node38210 : 4'b0000;
															assign node38210 = (inp[11]) ? node38212 : 4'b0000;
																assign node38212 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node38215 = (inp[0]) ? 4'b0000 : node38216;
															assign node38216 = (inp[2]) ? node38218 : 4'b0001;
																assign node38218 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node38222 = (inp[13]) ? node38244 : node38223;
													assign node38223 = (inp[9]) ? node38237 : node38224;
														assign node38224 = (inp[0]) ? node38230 : node38225;
															assign node38225 = (inp[11]) ? node38227 : 4'b0100;
																assign node38227 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node38230 = (inp[11]) ? node38234 : node38231;
																assign node38231 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node38234 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node38237 = (inp[0]) ? node38239 : 4'b0100;
															assign node38239 = (inp[11]) ? node38241 : 4'b0100;
																assign node38241 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node38244 = (inp[0]) ? node38248 : node38245;
														assign node38245 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node38248 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node38251 = (inp[7]) ? node38321 : node38252;
											assign node38252 = (inp[12]) ? node38286 : node38253;
												assign node38253 = (inp[9]) ? node38277 : node38254;
													assign node38254 = (inp[0]) ? node38266 : node38255;
														assign node38255 = (inp[11]) ? node38261 : node38256;
															assign node38256 = (inp[2]) ? node38258 : 4'b0100;
																assign node38258 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node38261 = (inp[2]) ? node38263 : 4'b0101;
																assign node38263 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node38266 = (inp[11]) ? node38272 : node38267;
															assign node38267 = (inp[13]) ? node38269 : 4'b0101;
																assign node38269 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node38272 = (inp[13]) ? node38274 : 4'b0100;
																assign node38274 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node38277 = (inp[11]) ? node38281 : node38278;
														assign node38278 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38281 = (inp[0]) ? 4'b0100 : node38282;
															assign node38282 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node38286 = (inp[9]) ? node38306 : node38287;
													assign node38287 = (inp[2]) ? node38301 : node38288;
														assign node38288 = (inp[13]) ? node38294 : node38289;
															assign node38289 = (inp[11]) ? node38291 : 4'b0100;
																assign node38291 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38294 = (inp[11]) ? node38298 : node38295;
																assign node38295 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node38298 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38301 = (inp[11]) ? 4'b0100 : node38302;
															assign node38302 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node38306 = (inp[11]) ? node38314 : node38307;
														assign node38307 = (inp[0]) ? 4'b0100 : node38308;
															assign node38308 = (inp[13]) ? node38310 : 4'b0101;
																assign node38310 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node38314 = (inp[0]) ? node38318 : node38315;
															assign node38315 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node38318 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node38321 = (inp[12]) ? node38351 : node38322;
												assign node38322 = (inp[9]) ? node38336 : node38323;
													assign node38323 = (inp[2]) ? node38325 : 4'b0101;
														assign node38325 = (inp[0]) ? node38331 : node38326;
															assign node38326 = (inp[11]) ? node38328 : 4'b0101;
																assign node38328 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node38331 = (inp[11]) ? node38333 : 4'b0100;
																assign node38333 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node38336 = (inp[13]) ? node38344 : node38337;
														assign node38337 = (inp[11]) ? node38341 : node38338;
															assign node38338 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38341 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node38344 = (inp[11]) ? node38346 : 4'b0100;
															assign node38346 = (inp[0]) ? node38348 : 4'b0100;
																assign node38348 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node38351 = (inp[2]) ? node38359 : node38352;
													assign node38352 = (inp[0]) ? node38356 : node38353;
														assign node38353 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node38356 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node38359 = (inp[11]) ? node38365 : node38360;
														assign node38360 = (inp[0]) ? 4'b0000 : node38361;
															assign node38361 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node38365 = (inp[13]) ? node38369 : node38366;
															assign node38366 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node38369 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node38372 = (inp[1]) ? node38454 : node38373;
										assign node38373 = (inp[7]) ? node38397 : node38374;
											assign node38374 = (inp[0]) ? node38386 : node38375;
												assign node38375 = (inp[11]) ? node38381 : node38376;
													assign node38376 = (inp[13]) ? node38378 : 4'b0100;
														assign node38378 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node38381 = (inp[2]) ? node38383 : 4'b0101;
														assign node38383 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node38386 = (inp[11]) ? node38392 : node38387;
													assign node38387 = (inp[2]) ? node38389 : 4'b0101;
														assign node38389 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node38392 = (inp[13]) ? node38394 : 4'b0100;
														assign node38394 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node38397 = (inp[12]) ? node38433 : node38398;
												assign node38398 = (inp[9]) ? node38418 : node38399;
													assign node38399 = (inp[13]) ? node38407 : node38400;
														assign node38400 = (inp[2]) ? 4'b0100 : node38401;
															assign node38401 = (inp[0]) ? 4'b0101 : node38402;
																assign node38402 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node38407 = (inp[2]) ? node38413 : node38408;
															assign node38408 = (inp[11]) ? node38410 : 4'b0100;
																assign node38410 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node38413 = (inp[11]) ? node38415 : 4'b0101;
																assign node38415 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node38418 = (inp[2]) ? node38426 : node38419;
														assign node38419 = (inp[13]) ? node38421 : 4'b0100;
															assign node38421 = (inp[0]) ? node38423 : 4'b0101;
																assign node38423 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node38426 = (inp[13]) ? node38428 : 4'b0101;
															assign node38428 = (inp[0]) ? 4'b0101 : node38429;
																assign node38429 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node38433 = (inp[0]) ? node38445 : node38434;
													assign node38434 = (inp[11]) ? node38440 : node38435;
														assign node38435 = (inp[13]) ? node38437 : 4'b0000;
															assign node38437 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node38440 = (inp[2]) ? node38442 : 4'b0001;
															assign node38442 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node38445 = (inp[11]) ? node38451 : node38446;
														assign node38446 = (inp[2]) ? node38448 : 4'b0001;
															assign node38448 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node38451 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node38454 = (inp[7]) ? node38516 : node38455;
											assign node38455 = (inp[0]) ? node38489 : node38456;
												assign node38456 = (inp[9]) ? node38472 : node38457;
													assign node38457 = (inp[11]) ? node38463 : node38458;
														assign node38458 = (inp[12]) ? 4'b0000 : node38459;
															assign node38459 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node38463 = (inp[13]) ? node38469 : node38464;
															assign node38464 = (inp[2]) ? 4'b0001 : node38465;
																assign node38465 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node38469 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node38472 = (inp[11]) ? node38482 : node38473;
														assign node38473 = (inp[12]) ? node38479 : node38474;
															assign node38474 = (inp[2]) ? 4'b0001 : node38475;
																assign node38475 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node38479 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node38482 = (inp[12]) ? node38484 : 4'b0000;
															assign node38484 = (inp[2]) ? 4'b0001 : node38485;
																assign node38485 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node38489 = (inp[13]) ? node38505 : node38490;
													assign node38490 = (inp[11]) ? node38498 : node38491;
														assign node38491 = (inp[2]) ? node38495 : node38492;
															assign node38492 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node38495 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node38498 = (inp[12]) ? node38502 : node38499;
															assign node38499 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node38502 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node38505 = (inp[2]) ? node38509 : node38506;
														assign node38506 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node38509 = (inp[12]) ? node38513 : node38510;
															assign node38510 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node38513 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node38516 = (inp[12]) ? node38532 : node38517;
												assign node38517 = (inp[0]) ? node38525 : node38518;
													assign node38518 = (inp[11]) ? node38520 : 4'b0000;
														assign node38520 = (inp[13]) ? 4'b0001 : node38521;
															assign node38521 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node38525 = (inp[11]) ? node38527 : 4'b0001;
														assign node38527 = (inp[13]) ? 4'b0000 : node38528;
															assign node38528 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node38532 = (inp[13]) ? node38548 : node38533;
													assign node38533 = (inp[2]) ? node38537 : node38534;
														assign node38534 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node38537 = (inp[9]) ? node38543 : node38538;
															assign node38538 = (inp[0]) ? 4'b0101 : node38539;
																assign node38539 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node38543 = (inp[0]) ? 4'b0100 : node38544;
																assign node38544 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node38548 = (inp[11]) ? node38556 : node38549;
														assign node38549 = (inp[2]) ? node38553 : node38550;
															assign node38550 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node38553 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node38556 = (inp[2]) ? node38558 : 4'b0100;
															assign node38558 = (inp[0]) ? 4'b0100 : 4'b0101;
							assign node38561 = (inp[9]) ? node38927 : node38562;
								assign node38562 = (inp[11]) ? node38720 : node38563;
									assign node38563 = (inp[2]) ? node38629 : node38564;
										assign node38564 = (inp[0]) ? node38604 : node38565;
											assign node38565 = (inp[5]) ? node38577 : node38566;
												assign node38566 = (inp[12]) ? node38570 : node38567;
													assign node38567 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node38570 = (inp[1]) ? node38572 : 4'b0110;
														assign node38572 = (inp[7]) ? 4'b0010 : node38573;
															assign node38573 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node38577 = (inp[7]) ? node38589 : node38578;
													assign node38578 = (inp[13]) ? node38584 : node38579;
														assign node38579 = (inp[1]) ? 4'b0110 : node38580;
															assign node38580 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38584 = (inp[12]) ? node38586 : 4'b0111;
															assign node38586 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node38589 = (inp[13]) ? node38595 : node38590;
														assign node38590 = (inp[1]) ? node38592 : 4'b0011;
															assign node38592 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node38595 = (inp[10]) ? node38599 : node38596;
															assign node38596 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node38599 = (inp[12]) ? 4'b0010 : node38600;
																assign node38600 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node38604 = (inp[1]) ? node38618 : node38605;
												assign node38605 = (inp[12]) ? node38609 : node38606;
													assign node38606 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node38609 = (inp[13]) ? node38611 : 4'b0111;
														assign node38611 = (inp[5]) ? node38615 : node38612;
															assign node38612 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node38615 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node38618 = (inp[12]) ? 4'b0011 : node38619;
													assign node38619 = (inp[10]) ? 4'b0111 : node38620;
														assign node38620 = (inp[13]) ? node38622 : 4'b0110;
															assign node38622 = (inp[5]) ? node38624 : 4'b0111;
																assign node38624 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node38629 = (inp[0]) ? node38679 : node38630;
											assign node38630 = (inp[5]) ? node38646 : node38631;
												assign node38631 = (inp[12]) ? node38635 : node38632;
													assign node38632 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node38635 = (inp[1]) ? node38641 : node38636;
														assign node38636 = (inp[13]) ? node38638 : 4'b0111;
															assign node38638 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node38641 = (inp[13]) ? 4'b0011 : node38642;
															assign node38642 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node38646 = (inp[12]) ? node38668 : node38647;
													assign node38647 = (inp[1]) ? node38655 : node38648;
														assign node38648 = (inp[10]) ? node38650 : 4'b0011;
															assign node38650 = (inp[13]) ? 4'b0010 : node38651;
																assign node38651 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node38655 = (inp[10]) ? node38663 : node38656;
															assign node38656 = (inp[13]) ? node38660 : node38657;
																assign node38657 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node38660 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node38663 = (inp[13]) ? 4'b0110 : node38664;
																assign node38664 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node38668 = (inp[1]) ? node38674 : node38669;
														assign node38669 = (inp[13]) ? node38671 : 4'b0111;
															assign node38671 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38674 = (inp[7]) ? node38676 : 4'b0011;
															assign node38676 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node38679 = (inp[5]) ? node38695 : node38680;
												assign node38680 = (inp[12]) ? node38684 : node38681;
													assign node38681 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node38684 = (inp[1]) ? node38690 : node38685;
														assign node38685 = (inp[13]) ? node38687 : 4'b0110;
															assign node38687 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38690 = (inp[7]) ? 4'b0010 : node38691;
															assign node38691 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node38695 = (inp[12]) ? node38709 : node38696;
													assign node38696 = (inp[1]) ? node38704 : node38697;
														assign node38697 = (inp[7]) ? node38701 : node38698;
															assign node38698 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node38701 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node38704 = (inp[13]) ? 4'b0110 : node38705;
															assign node38705 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node38709 = (inp[1]) ? node38715 : node38710;
														assign node38710 = (inp[10]) ? node38712 : 4'b0110;
															assign node38712 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node38715 = (inp[7]) ? node38717 : 4'b0010;
															assign node38717 = (inp[13]) ? 4'b0010 : 4'b0011;
									assign node38720 = (inp[5]) ? node38782 : node38721;
										assign node38721 = (inp[0]) ? node38753 : node38722;
											assign node38722 = (inp[2]) ? node38738 : node38723;
												assign node38723 = (inp[12]) ? node38727 : node38724;
													assign node38724 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node38727 = (inp[1]) ? node38733 : node38728;
														assign node38728 = (inp[13]) ? node38730 : 4'b0110;
															assign node38730 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38733 = (inp[7]) ? 4'b0010 : node38734;
															assign node38734 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node38738 = (inp[12]) ? node38742 : node38739;
													assign node38739 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node38742 = (inp[1]) ? node38748 : node38743;
														assign node38743 = (inp[7]) ? node38745 : 4'b0111;
															assign node38745 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node38748 = (inp[13]) ? 4'b0011 : node38749;
															assign node38749 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node38753 = (inp[2]) ? node38767 : node38754;
												assign node38754 = (inp[12]) ? node38758 : node38755;
													assign node38755 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node38758 = (inp[1]) ? node38762 : node38759;
														assign node38759 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node38762 = (inp[13]) ? 4'b0011 : node38763;
															assign node38763 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node38767 = (inp[12]) ? node38771 : node38768;
													assign node38768 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node38771 = (inp[1]) ? node38777 : node38772;
														assign node38772 = (inp[13]) ? node38774 : 4'b0110;
															assign node38774 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node38777 = (inp[7]) ? 4'b0010 : node38778;
															assign node38778 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node38782 = (inp[10]) ? node38846 : node38783;
											assign node38783 = (inp[0]) ? node38807 : node38784;
												assign node38784 = (inp[7]) ? node38798 : node38785;
													assign node38785 = (inp[12]) ? node38791 : node38786;
														assign node38786 = (inp[13]) ? node38788 : 4'b0111;
															assign node38788 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node38791 = (inp[1]) ? 4'b0010 : node38792;
															assign node38792 = (inp[2]) ? 4'b0110 : node38793;
																assign node38793 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node38798 = (inp[12]) ? node38802 : node38799;
														assign node38799 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node38802 = (inp[1]) ? node38804 : 4'b0111;
															assign node38804 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node38807 = (inp[7]) ? node38829 : node38808;
													assign node38808 = (inp[2]) ? node38818 : node38809;
														assign node38809 = (inp[13]) ? node38811 : 4'b0011;
															assign node38811 = (inp[12]) ? node38815 : node38812;
																assign node38812 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node38815 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node38818 = (inp[13]) ? node38826 : node38819;
															assign node38819 = (inp[1]) ? node38823 : node38820;
																assign node38820 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node38823 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node38826 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node38829 = (inp[13]) ? node38841 : node38830;
														assign node38830 = (inp[2]) ? node38838 : node38831;
															assign node38831 = (inp[1]) ? node38835 : node38832;
																assign node38832 = (inp[12]) ? 4'b0111 : 4'b0010;
																assign node38835 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node38838 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node38841 = (inp[2]) ? 4'b0110 : node38842;
															assign node38842 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node38846 = (inp[7]) ? node38894 : node38847;
												assign node38847 = (inp[2]) ? node38873 : node38848;
													assign node38848 = (inp[0]) ? node38862 : node38849;
														assign node38849 = (inp[13]) ? node38855 : node38850;
															assign node38850 = (inp[12]) ? node38852 : 4'b0010;
																assign node38852 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node38855 = (inp[1]) ? node38859 : node38856;
																assign node38856 = (inp[12]) ? 4'b0111 : 4'b0011;
																assign node38859 = (inp[12]) ? 4'b0010 : 4'b0111;
														assign node38862 = (inp[13]) ? node38868 : node38863;
															assign node38863 = (inp[1]) ? node38865 : 4'b0111;
																assign node38865 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node38868 = (inp[12]) ? node38870 : 4'b0110;
																assign node38870 = (inp[1]) ? 4'b0011 : 4'b0110;
													assign node38873 = (inp[12]) ? node38887 : node38874;
														assign node38874 = (inp[1]) ? node38882 : node38875;
															assign node38875 = (inp[0]) ? node38879 : node38876;
																assign node38876 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node38879 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node38882 = (inp[0]) ? node38884 : 4'b0110;
																assign node38884 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node38887 = (inp[1]) ? node38891 : node38888;
															assign node38888 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node38891 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node38894 = (inp[2]) ? node38912 : node38895;
													assign node38895 = (inp[13]) ? node38905 : node38896;
														assign node38896 = (inp[0]) ? node38900 : node38897;
															assign node38897 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node38900 = (inp[12]) ? 4'b0010 : node38901;
																assign node38901 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node38905 = (inp[0]) ? 4'b0011 : node38906;
															assign node38906 = (inp[1]) ? node38908 : 4'b0010;
																assign node38908 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node38912 = (inp[1]) ? node38922 : node38913;
														assign node38913 = (inp[12]) ? 4'b0110 : node38914;
															assign node38914 = (inp[13]) ? node38918 : node38915;
																assign node38915 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node38918 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node38922 = (inp[12]) ? node38924 : 4'b0111;
															assign node38924 = (inp[13]) ? 4'b0010 : 4'b0011;
								assign node38927 = (inp[0]) ? node39093 : node38928;
									assign node38928 = (inp[2]) ? node39030 : node38929;
										assign node38929 = (inp[5]) ? node38977 : node38930;
											assign node38930 = (inp[7]) ? node38958 : node38931;
												assign node38931 = (inp[11]) ? node38941 : node38932;
													assign node38932 = (inp[1]) ? node38936 : node38933;
														assign node38933 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38936 = (inp[12]) ? node38938 : 4'b0110;
															assign node38938 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node38941 = (inp[13]) ? node38947 : node38942;
														assign node38942 = (inp[1]) ? 4'b0110 : node38943;
															assign node38943 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node38947 = (inp[10]) ? node38953 : node38948;
															assign node38948 = (inp[12]) ? 4'b0110 : node38949;
																assign node38949 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node38953 = (inp[1]) ? 4'b0010 : node38954;
																assign node38954 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node38958 = (inp[11]) ? node38966 : node38959;
													assign node38959 = (inp[1]) ? 4'b0010 : node38960;
														assign node38960 = (inp[12]) ? node38962 : 4'b0010;
															assign node38962 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node38966 = (inp[10]) ? node38972 : node38967;
														assign node38967 = (inp[12]) ? 4'b0010 : node38968;
															assign node38968 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node38972 = (inp[12]) ? 4'b0110 : node38973;
															assign node38973 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node38977 = (inp[12]) ? node39019 : node38978;
												assign node38978 = (inp[1]) ? node38998 : node38979;
													assign node38979 = (inp[11]) ? node38993 : node38980;
														assign node38980 = (inp[10]) ? node38986 : node38981;
															assign node38981 = (inp[13]) ? node38983 : 4'b0010;
																assign node38983 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node38986 = (inp[13]) ? node38990 : node38987;
																assign node38987 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node38990 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node38993 = (inp[7]) ? 4'b0011 : node38994;
															assign node38994 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node38998 = (inp[11]) ? node39008 : node38999;
														assign node38999 = (inp[10]) ? node39001 : 4'b0110;
															assign node39001 = (inp[7]) ? node39005 : node39002;
																assign node39002 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node39005 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node39008 = (inp[10]) ? node39014 : node39009;
															assign node39009 = (inp[13]) ? node39011 : 4'b0111;
																assign node39011 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39014 = (inp[7]) ? 4'b0111 : node39015;
																assign node39015 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node39019 = (inp[1]) ? node39025 : node39020;
													assign node39020 = (inp[7]) ? 4'b0110 : node39021;
														assign node39021 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node39025 = (inp[7]) ? node39027 : 4'b0010;
														assign node39027 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node39030 = (inp[5]) ? node39048 : node39031;
											assign node39031 = (inp[12]) ? node39035 : node39032;
												assign node39032 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node39035 = (inp[1]) ? node39043 : node39036;
													assign node39036 = (inp[11]) ? node39038 : 4'b0111;
														assign node39038 = (inp[7]) ? node39040 : 4'b0111;
															assign node39040 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node39043 = (inp[7]) ? 4'b0011 : node39044;
														assign node39044 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node39048 = (inp[12]) ? node39082 : node39049;
												assign node39049 = (inp[1]) ? node39067 : node39050;
													assign node39050 = (inp[10]) ? node39062 : node39051;
														assign node39051 = (inp[11]) ? node39057 : node39052;
															assign node39052 = (inp[13]) ? 4'b0010 : node39053;
																assign node39053 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node39057 = (inp[13]) ? node39059 : 4'b0010;
																assign node39059 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node39062 = (inp[7]) ? 4'b0011 : node39063;
															assign node39063 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node39067 = (inp[11]) ? node39073 : node39068;
														assign node39068 = (inp[13]) ? 4'b0111 : node39069;
															assign node39069 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39073 = (inp[10]) ? node39077 : node39074;
															assign node39074 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node39077 = (inp[13]) ? 4'b0110 : node39078;
																assign node39078 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39082 = (inp[1]) ? node39088 : node39083;
													assign node39083 = (inp[13]) ? node39085 : 4'b0111;
														assign node39085 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node39088 = (inp[13]) ? 4'b0011 : node39089;
														assign node39089 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node39093 = (inp[2]) ? node39143 : node39094;
										assign node39094 = (inp[5]) ? node39110 : node39095;
											assign node39095 = (inp[12]) ? node39099 : node39096;
												assign node39096 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node39099 = (inp[1]) ? node39105 : node39100;
													assign node39100 = (inp[13]) ? node39102 : 4'b0111;
														assign node39102 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node39105 = (inp[7]) ? 4'b0011 : node39106;
														assign node39106 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node39110 = (inp[12]) ? node39132 : node39111;
												assign node39111 = (inp[1]) ? node39119 : node39112;
													assign node39112 = (inp[7]) ? node39116 : node39113;
														assign node39113 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node39116 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node39119 = (inp[10]) ? node39127 : node39120;
														assign node39120 = (inp[7]) ? node39124 : node39121;
															assign node39121 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node39124 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node39127 = (inp[13]) ? node39129 : 4'b0110;
															assign node39129 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node39132 = (inp[1]) ? node39138 : node39133;
													assign node39133 = (inp[7]) ? 4'b0111 : node39134;
														assign node39134 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node39138 = (inp[13]) ? 4'b0011 : node39139;
														assign node39139 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node39143 = (inp[5]) ? node39159 : node39144;
											assign node39144 = (inp[12]) ? node39148 : node39145;
												assign node39145 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node39148 = (inp[1]) ? node39154 : node39149;
													assign node39149 = (inp[13]) ? node39151 : 4'b0110;
														assign node39151 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node39154 = (inp[7]) ? 4'b0010 : node39155;
														assign node39155 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node39159 = (inp[12]) ? node39191 : node39160;
												assign node39160 = (inp[1]) ? node39178 : node39161;
													assign node39161 = (inp[10]) ? node39171 : node39162;
														assign node39162 = (inp[11]) ? node39164 : 4'b0010;
															assign node39164 = (inp[7]) ? node39168 : node39165;
																assign node39165 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node39168 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node39171 = (inp[13]) ? node39175 : node39172;
															assign node39172 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node39175 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node39178 = (inp[10]) ? node39184 : node39179;
														assign node39179 = (inp[13]) ? node39181 : 4'b0111;
															assign node39181 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39184 = (inp[7]) ? node39188 : node39185;
															assign node39185 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node39188 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node39191 = (inp[1]) ? node39197 : node39192;
													assign node39192 = (inp[13]) ? node39194 : 4'b0110;
														assign node39194 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node39197 = (inp[13]) ? 4'b0010 : node39198;
														assign node39198 = (inp[7]) ? 4'b0011 : 4'b0010;
						assign node39202 = (inp[2]) ? node39662 : node39203;
							assign node39203 = (inp[0]) ? node39407 : node39204;
								assign node39204 = (inp[14]) ? node39354 : node39205;
									assign node39205 = (inp[12]) ? node39287 : node39206;
										assign node39206 = (inp[1]) ? node39260 : node39207;
											assign node39207 = (inp[11]) ? node39227 : node39208;
												assign node39208 = (inp[13]) ? node39216 : node39209;
													assign node39209 = (inp[7]) ? node39213 : node39210;
														assign node39210 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node39213 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node39216 = (inp[9]) ? node39222 : node39217;
														assign node39217 = (inp[7]) ? node39219 : 4'b0111;
															assign node39219 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node39222 = (inp[7]) ? node39224 : 4'b0011;
															assign node39224 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node39227 = (inp[13]) ? node39237 : node39228;
													assign node39228 = (inp[9]) ? 4'b0010 : node39229;
														assign node39229 = (inp[10]) ? 4'b0111 : node39230;
															assign node39230 = (inp[7]) ? 4'b0010 : node39231;
																assign node39231 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node39237 = (inp[10]) ? node39245 : node39238;
														assign node39238 = (inp[7]) ? node39242 : node39239;
															assign node39239 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node39242 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node39245 = (inp[9]) ? node39253 : node39246;
															assign node39246 = (inp[5]) ? node39250 : node39247;
																assign node39247 = (inp[7]) ? 4'b0110 : 4'b0010;
																assign node39250 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node39253 = (inp[5]) ? node39257 : node39254;
																assign node39254 = (inp[7]) ? 4'b0110 : 4'b0010;
																assign node39257 = (inp[7]) ? 4'b0010 : 4'b0110;
											assign node39260 = (inp[11]) ? node39274 : node39261;
												assign node39261 = (inp[7]) ? node39267 : node39262;
													assign node39262 = (inp[5]) ? node39264 : 4'b0110;
														assign node39264 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node39267 = (inp[5]) ? node39271 : node39268;
														assign node39268 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node39271 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node39274 = (inp[5]) ? node39280 : node39275;
													assign node39275 = (inp[7]) ? node39277 : 4'b0111;
														assign node39277 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node39280 = (inp[7]) ? node39284 : node39281;
														assign node39281 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node39284 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node39287 = (inp[5]) ? node39339 : node39288;
											assign node39288 = (inp[1]) ? node39324 : node39289;
												assign node39289 = (inp[10]) ? node39313 : node39290;
													assign node39290 = (inp[7]) ? node39306 : node39291;
														assign node39291 = (inp[9]) ? node39299 : node39292;
															assign node39292 = (inp[11]) ? node39296 : node39293;
																assign node39293 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node39296 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node39299 = (inp[13]) ? node39303 : node39300;
																assign node39300 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node39303 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node39306 = (inp[13]) ? node39310 : node39307;
															assign node39307 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node39310 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node39313 = (inp[11]) ? node39315 : 4'b0010;
														assign node39315 = (inp[9]) ? 4'b0011 : node39316;
															assign node39316 = (inp[7]) ? node39320 : node39317;
																assign node39317 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node39320 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node39324 = (inp[10]) ? node39332 : node39325;
													assign node39325 = (inp[7]) ? node39329 : node39326;
														assign node39326 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node39329 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node39332 = (inp[7]) ? node39336 : node39333;
														assign node39333 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node39336 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node39339 = (inp[1]) ? node39347 : node39340;
												assign node39340 = (inp[11]) ? node39344 : node39341;
													assign node39341 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node39344 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node39347 = (inp[11]) ? node39351 : node39348;
													assign node39348 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node39351 = (inp[13]) ? 4'b0010 : 4'b0011;
									assign node39354 = (inp[5]) ? node39392 : node39355;
										assign node39355 = (inp[13]) ? node39377 : node39356;
											assign node39356 = (inp[7]) ? node39370 : node39357;
												assign node39357 = (inp[10]) ? node39365 : node39358;
													assign node39358 = (inp[12]) ? node39362 : node39359;
														assign node39359 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node39362 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node39365 = (inp[1]) ? 4'b0110 : node39366;
														assign node39366 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node39370 = (inp[12]) ? node39374 : node39371;
													assign node39371 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node39374 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node39377 = (inp[7]) ? node39385 : node39378;
												assign node39378 = (inp[1]) ? node39382 : node39379;
													assign node39379 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node39382 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node39385 = (inp[12]) ? node39389 : node39386;
													assign node39386 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node39389 = (inp[1]) ? 4'b0010 : 4'b0110;
										assign node39392 = (inp[12]) ? node39404 : node39393;
											assign node39393 = (inp[1]) ? node39399 : node39394;
												assign node39394 = (inp[13]) ? node39396 : 4'b0010;
													assign node39396 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node39399 = (inp[13]) ? 4'b0110 : node39400;
													assign node39400 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node39404 = (inp[1]) ? 4'b0010 : 4'b0110;
								assign node39407 = (inp[14]) ? node39605 : node39408;
									assign node39408 = (inp[7]) ? node39462 : node39409;
										assign node39409 = (inp[11]) ? node39435 : node39410;
											assign node39410 = (inp[13]) ? node39422 : node39411;
												assign node39411 = (inp[1]) ? node39415 : node39412;
													assign node39412 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node39415 = (inp[5]) ? node39419 : node39416;
														assign node39416 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node39419 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node39422 = (inp[12]) ? node39428 : node39423;
													assign node39423 = (inp[1]) ? node39425 : 4'b0110;
														assign node39425 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node39428 = (inp[1]) ? node39432 : node39429;
														assign node39429 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node39432 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node39435 = (inp[13]) ? node39447 : node39436;
												assign node39436 = (inp[1]) ? node39440 : node39437;
													assign node39437 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node39440 = (inp[5]) ? node39444 : node39441;
														assign node39441 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node39444 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node39447 = (inp[12]) ? node39455 : node39448;
													assign node39448 = (inp[1]) ? node39452 : node39449;
														assign node39449 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node39452 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node39455 = (inp[1]) ? node39459 : node39456;
														assign node39456 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node39459 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node39462 = (inp[10]) ? node39516 : node39463;
											assign node39463 = (inp[12]) ? node39491 : node39464;
												assign node39464 = (inp[11]) ? node39482 : node39465;
													assign node39465 = (inp[13]) ? node39477 : node39466;
														assign node39466 = (inp[9]) ? node39472 : node39467;
															assign node39467 = (inp[1]) ? 4'b0111 : node39468;
																assign node39468 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node39472 = (inp[5]) ? node39474 : 4'b0010;
																assign node39474 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node39477 = (inp[1]) ? 4'b0110 : node39478;
															assign node39478 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node39482 = (inp[13]) ? node39488 : node39483;
														assign node39483 = (inp[5]) ? 4'b0110 : node39484;
															assign node39484 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node39488 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node39491 = (inp[11]) ? node39503 : node39492;
													assign node39492 = (inp[1]) ? node39498 : node39493;
														assign node39493 = (inp[5]) ? 4'b0110 : node39494;
															assign node39494 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node39498 = (inp[5]) ? node39500 : 4'b0111;
															assign node39500 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node39503 = (inp[1]) ? node39511 : node39504;
														assign node39504 = (inp[5]) ? node39508 : node39505;
															assign node39505 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node39508 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node39511 = (inp[5]) ? node39513 : 4'b0110;
															assign node39513 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node39516 = (inp[9]) ? node39566 : node39517;
												assign node39517 = (inp[13]) ? node39541 : node39518;
													assign node39518 = (inp[12]) ? node39534 : node39519;
														assign node39519 = (inp[1]) ? node39527 : node39520;
															assign node39520 = (inp[5]) ? node39524 : node39521;
																assign node39521 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node39524 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node39527 = (inp[5]) ? node39531 : node39528;
																assign node39528 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node39531 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node39534 = (inp[11]) ? node39536 : 4'b0111;
															assign node39536 = (inp[5]) ? 4'b0110 : node39537;
																assign node39537 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node39541 = (inp[5]) ? node39555 : node39542;
														assign node39542 = (inp[11]) ? node39548 : node39543;
															assign node39543 = (inp[1]) ? node39545 : 4'b0110;
																assign node39545 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node39548 = (inp[12]) ? node39552 : node39549;
																assign node39549 = (inp[1]) ? 4'b0010 : 4'b0111;
																assign node39552 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node39555 = (inp[11]) ? node39561 : node39556;
															assign node39556 = (inp[12]) ? 4'b0010 : node39557;
																assign node39557 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node39561 = (inp[12]) ? 4'b0011 : node39562;
																assign node39562 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node39566 = (inp[5]) ? node39588 : node39567;
													assign node39567 = (inp[12]) ? node39577 : node39568;
														assign node39568 = (inp[1]) ? 4'b0011 : node39569;
															assign node39569 = (inp[11]) ? node39573 : node39570;
																assign node39570 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node39573 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node39577 = (inp[1]) ? node39585 : node39578;
															assign node39578 = (inp[13]) ? node39582 : node39579;
																assign node39579 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node39582 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node39585 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node39588 = (inp[13]) ? node39602 : node39589;
														assign node39589 = (inp[11]) ? node39597 : node39590;
															assign node39590 = (inp[12]) ? node39594 : node39591;
																assign node39591 = (inp[1]) ? 4'b0111 : 4'b0010;
																assign node39594 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node39597 = (inp[12]) ? 4'b0110 : node39598;
																assign node39598 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node39602 = (inp[11]) ? 4'b0111 : 4'b0110;
									assign node39605 = (inp[5]) ? node39647 : node39606;
										assign node39606 = (inp[12]) ? node39618 : node39607;
											assign node39607 = (inp[1]) ? node39613 : node39608;
												assign node39608 = (inp[7]) ? 4'b0011 : node39609;
													assign node39609 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node39613 = (inp[7]) ? node39615 : 4'b0111;
													assign node39615 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node39618 = (inp[1]) ? node39626 : node39619;
												assign node39619 = (inp[7]) ? node39623 : node39620;
													assign node39620 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node39623 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node39626 = (inp[10]) ? node39640 : node39627;
													assign node39627 = (inp[9]) ? node39635 : node39628;
														assign node39628 = (inp[13]) ? node39632 : node39629;
															assign node39629 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node39632 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node39635 = (inp[7]) ? node39637 : 4'b0011;
															assign node39637 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node39640 = (inp[13]) ? node39644 : node39641;
														assign node39641 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node39644 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node39647 = (inp[12]) ? node39659 : node39648;
											assign node39648 = (inp[1]) ? node39654 : node39649;
												assign node39649 = (inp[13]) ? node39651 : 4'b0011;
													assign node39651 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node39654 = (inp[13]) ? 4'b0111 : node39655;
													assign node39655 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node39659 = (inp[1]) ? 4'b0011 : 4'b0111;
							assign node39662 = (inp[0]) ? node39792 : node39663;
								assign node39663 = (inp[14]) ? node39749 : node39664;
									assign node39664 = (inp[11]) ? node39702 : node39665;
										assign node39665 = (inp[5]) ? node39687 : node39666;
											assign node39666 = (inp[1]) ? node39672 : node39667;
												assign node39667 = (inp[7]) ? node39669 : 4'b0010;
													assign node39669 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node39672 = (inp[12]) ? node39678 : node39673;
													assign node39673 = (inp[7]) ? 4'b0011 : node39674;
														assign node39674 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node39678 = (inp[9]) ? node39680 : 4'b0110;
														assign node39680 = (inp[7]) ? node39684 : node39681;
															assign node39681 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node39684 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node39687 = (inp[1]) ? node39695 : node39688;
												assign node39688 = (inp[12]) ? 4'b0110 : node39689;
													assign node39689 = (inp[7]) ? node39691 : 4'b0110;
														assign node39691 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node39695 = (inp[7]) ? node39699 : node39696;
													assign node39696 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node39699 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node39702 = (inp[5]) ? node39736 : node39703;
											assign node39703 = (inp[1]) ? node39711 : node39704;
												assign node39704 = (inp[12]) ? node39708 : node39705;
													assign node39705 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node39708 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node39711 = (inp[12]) ? node39717 : node39712;
													assign node39712 = (inp[7]) ? 4'b0010 : node39713;
														assign node39713 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node39717 = (inp[10]) ? node39729 : node39718;
														assign node39718 = (inp[9]) ? node39724 : node39719;
															assign node39719 = (inp[13]) ? node39721 : 4'b0111;
																assign node39721 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39724 = (inp[13]) ? 4'b0111 : node39725;
																assign node39725 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39729 = (inp[13]) ? node39733 : node39730;
															assign node39730 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39733 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node39736 = (inp[12]) ? node39746 : node39737;
												assign node39737 = (inp[7]) ? node39741 : node39738;
													assign node39738 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node39741 = (inp[1]) ? 4'b0111 : node39742;
														assign node39742 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node39746 = (inp[1]) ? 4'b0011 : 4'b0111;
									assign node39749 = (inp[5]) ? node39777 : node39750;
										assign node39750 = (inp[12]) ? node39762 : node39751;
											assign node39751 = (inp[1]) ? node39757 : node39752;
												assign node39752 = (inp[13]) ? node39754 : 4'b0011;
													assign node39754 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node39757 = (inp[7]) ? node39759 : 4'b0111;
													assign node39759 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node39762 = (inp[1]) ? node39770 : node39763;
												assign node39763 = (inp[13]) ? node39767 : node39764;
													assign node39764 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node39767 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node39770 = (inp[7]) ? node39774 : node39771;
													assign node39771 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node39774 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node39777 = (inp[12]) ? node39789 : node39778;
											assign node39778 = (inp[1]) ? node39784 : node39779;
												assign node39779 = (inp[7]) ? node39781 : 4'b0011;
													assign node39781 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node39784 = (inp[13]) ? 4'b0111 : node39785;
													assign node39785 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node39789 = (inp[1]) ? 4'b0011 : 4'b0111;
								assign node39792 = (inp[14]) ? node39894 : node39793;
									assign node39793 = (inp[11]) ? node39837 : node39794;
										assign node39794 = (inp[1]) ? node39808 : node39795;
											assign node39795 = (inp[5]) ? node39801 : node39796;
												assign node39796 = (inp[7]) ? node39798 : 4'b0011;
													assign node39798 = (inp[12]) ? 4'b0010 : 4'b0111;
												assign node39801 = (inp[12]) ? 4'b0111 : node39802;
													assign node39802 = (inp[7]) ? node39804 : 4'b0111;
														assign node39804 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node39808 = (inp[5]) ? node39830 : node39809;
												assign node39809 = (inp[12]) ? node39815 : node39810;
													assign node39810 = (inp[7]) ? 4'b0010 : node39811;
														assign node39811 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node39815 = (inp[9]) ? node39823 : node39816;
														assign node39816 = (inp[13]) ? node39820 : node39817;
															assign node39817 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39820 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node39823 = (inp[13]) ? node39827 : node39824;
															assign node39824 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39827 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node39830 = (inp[7]) ? node39834 : node39831;
													assign node39831 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node39834 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node39837 = (inp[1]) ? node39853 : node39838;
											assign node39838 = (inp[5]) ? node39846 : node39839;
												assign node39839 = (inp[12]) ? node39843 : node39840;
													assign node39840 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node39843 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node39846 = (inp[7]) ? node39848 : 4'b0110;
													assign node39848 = (inp[12]) ? 4'b0110 : node39849;
														assign node39849 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node39853 = (inp[12]) ? node39877 : node39854;
												assign node39854 = (inp[13]) ? node39862 : node39855;
													assign node39855 = (inp[5]) ? node39859 : node39856;
														assign node39856 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node39859 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node39862 = (inp[9]) ? node39870 : node39863;
														assign node39863 = (inp[7]) ? node39867 : node39864;
															assign node39864 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node39867 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node39870 = (inp[7]) ? node39874 : node39871;
															assign node39871 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node39874 = (inp[5]) ? 4'b0110 : 4'b0011;
												assign node39877 = (inp[5]) ? 4'b0010 : node39878;
													assign node39878 = (inp[9]) ? node39880 : 4'b0110;
														assign node39880 = (inp[10]) ? node39888 : node39881;
															assign node39881 = (inp[13]) ? node39885 : node39882;
																assign node39882 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node39885 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39888 = (inp[7]) ? 4'b0110 : node39889;
																assign node39889 = (inp[13]) ? 4'b0111 : 4'b0110;
									assign node39894 = (inp[5]) ? node39942 : node39895;
										assign node39895 = (inp[12]) ? node39907 : node39896;
											assign node39896 = (inp[1]) ? node39902 : node39897;
												assign node39897 = (inp[7]) ? 4'b0010 : node39898;
													assign node39898 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node39902 = (inp[13]) ? 4'b0110 : node39903;
													assign node39903 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node39907 = (inp[1]) ? node39915 : node39908;
												assign node39908 = (inp[13]) ? node39912 : node39909;
													assign node39909 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node39912 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39915 = (inp[10]) ? node39935 : node39916;
													assign node39916 = (inp[11]) ? node39930 : node39917;
														assign node39917 = (inp[9]) ? node39925 : node39918;
															assign node39918 = (inp[7]) ? node39922 : node39919;
																assign node39919 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node39922 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node39925 = (inp[7]) ? node39927 : 4'b0010;
																assign node39927 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node39930 = (inp[9]) ? node39932 : 4'b0010;
															assign node39932 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node39935 = (inp[13]) ? node39939 : node39936;
														assign node39936 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node39939 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node39942 = (inp[12]) ? node39954 : node39943;
											assign node39943 = (inp[1]) ? node39949 : node39944;
												assign node39944 = (inp[7]) ? node39946 : 4'b0010;
													assign node39946 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node39949 = (inp[13]) ? 4'b0110 : node39950;
													assign node39950 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node39954 = (inp[1]) ? 4'b0010 : 4'b0110;
					assign node39957 = (inp[14]) ? node41033 : node39958;
						assign node39958 = (inp[15]) ? node40534 : node39959;
							assign node39959 = (inp[12]) ? node40231 : node39960;
								assign node39960 = (inp[1]) ? node40130 : node39961;
									assign node39961 = (inp[5]) ? node40067 : node39962;
										assign node39962 = (inp[7]) ? node40014 : node39963;
											assign node39963 = (inp[13]) ? node39999 : node39964;
												assign node39964 = (inp[9]) ? node39982 : node39965;
													assign node39965 = (inp[0]) ? node39975 : node39966;
														assign node39966 = (inp[10]) ? node39968 : 4'b0010;
															assign node39968 = (inp[2]) ? node39972 : node39969;
																assign node39969 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node39972 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node39975 = (inp[2]) ? node39979 : node39976;
															assign node39976 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node39979 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node39982 = (inp[11]) ? node39994 : node39983;
														assign node39983 = (inp[10]) ? node39989 : node39984;
															assign node39984 = (inp[0]) ? node39986 : 4'b0010;
																assign node39986 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node39989 = (inp[0]) ? 4'b0010 : node39990;
																assign node39990 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node39994 = (inp[2]) ? 4'b0011 : node39995;
															assign node39995 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node39999 = (inp[2]) ? node40007 : node40000;
													assign node40000 = (inp[11]) ? node40004 : node40001;
														assign node40001 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node40004 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node40007 = (inp[10]) ? 4'b0010 : node40008;
														assign node40008 = (inp[11]) ? 4'b0010 : node40009;
															assign node40009 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node40014 = (inp[10]) ? node40034 : node40015;
												assign node40015 = (inp[0]) ? node40027 : node40016;
													assign node40016 = (inp[11]) ? node40022 : node40017;
														assign node40017 = (inp[2]) ? node40019 : 4'b0010;
															assign node40019 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node40022 = (inp[13]) ? 4'b0011 : node40023;
															assign node40023 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node40027 = (inp[11]) ? node40029 : 4'b0011;
														assign node40029 = (inp[13]) ? 4'b0010 : node40030;
															assign node40030 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node40034 = (inp[13]) ? node40054 : node40035;
													assign node40035 = (inp[9]) ? node40047 : node40036;
														assign node40036 = (inp[11]) ? node40042 : node40037;
															assign node40037 = (inp[0]) ? node40039 : 4'b0010;
																assign node40039 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node40042 = (inp[0]) ? node40044 : 4'b0011;
																assign node40044 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node40047 = (inp[2]) ? 4'b0010 : node40048;
															assign node40048 = (inp[0]) ? node40050 : 4'b0010;
																assign node40050 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node40054 = (inp[9]) ? node40060 : node40055;
														assign node40055 = (inp[11]) ? 4'b0010 : node40056;
															assign node40056 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node40060 = (inp[11]) ? node40064 : node40061;
															assign node40061 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node40064 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node40067 = (inp[13]) ? node40089 : node40068;
											assign node40068 = (inp[11]) ? node40076 : node40069;
												assign node40069 = (inp[0]) ? node40073 : node40070;
													assign node40070 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node40073 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node40076 = (inp[10]) ? node40084 : node40077;
													assign node40077 = (inp[0]) ? node40081 : node40078;
														assign node40078 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node40081 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node40084 = (inp[7]) ? 4'b0110 : node40085;
														assign node40085 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node40089 = (inp[11]) ? node40113 : node40090;
												assign node40090 = (inp[2]) ? node40098 : node40091;
													assign node40091 = (inp[0]) ? node40095 : node40092;
														assign node40092 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node40095 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node40098 = (inp[9]) ? node40106 : node40099;
														assign node40099 = (inp[0]) ? node40103 : node40100;
															assign node40100 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node40103 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node40106 = (inp[7]) ? node40110 : node40107;
															assign node40107 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node40110 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node40113 = (inp[0]) ? node40121 : node40114;
													assign node40114 = (inp[7]) ? node40118 : node40115;
														assign node40115 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node40118 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node40121 = (inp[10]) ? node40127 : node40122;
														assign node40122 = (inp[7]) ? node40124 : 4'b0111;
															assign node40124 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node40127 = (inp[7]) ? 4'b0111 : 4'b0110;
									assign node40130 = (inp[5]) ? node40154 : node40131;
										assign node40131 = (inp[11]) ? node40143 : node40132;
											assign node40132 = (inp[0]) ? node40138 : node40133;
												assign node40133 = (inp[2]) ? node40135 : 4'b0110;
													assign node40135 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node40138 = (inp[13]) ? 4'b0111 : node40139;
													assign node40139 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node40143 = (inp[0]) ? node40149 : node40144;
												assign node40144 = (inp[13]) ? 4'b0111 : node40145;
													assign node40145 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node40149 = (inp[13]) ? 4'b0110 : node40150;
													assign node40150 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node40154 = (inp[2]) ? node40178 : node40155;
											assign node40155 = (inp[7]) ? node40163 : node40156;
												assign node40156 = (inp[0]) ? node40160 : node40157;
													assign node40157 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node40160 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node40163 = (inp[13]) ? node40171 : node40164;
													assign node40164 = (inp[0]) ? node40168 : node40165;
														assign node40165 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node40168 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node40171 = (inp[11]) ? node40175 : node40172;
														assign node40172 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node40175 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node40178 = (inp[7]) ? node40204 : node40179;
												assign node40179 = (inp[9]) ? node40191 : node40180;
													assign node40180 = (inp[11]) ? node40182 : 4'b0010;
														assign node40182 = (inp[10]) ? node40186 : node40183;
															assign node40183 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node40186 = (inp[0]) ? node40188 : 4'b0010;
																assign node40188 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node40191 = (inp[11]) ? node40199 : node40192;
														assign node40192 = (inp[13]) ? node40196 : node40193;
															assign node40193 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node40196 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node40199 = (inp[13]) ? 4'b0010 : node40200;
															assign node40200 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node40204 = (inp[10]) ? node40220 : node40205;
													assign node40205 = (inp[0]) ? node40211 : node40206;
														assign node40206 = (inp[13]) ? node40208 : 4'b0010;
															assign node40208 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node40211 = (inp[9]) ? node40213 : 4'b0011;
															assign node40213 = (inp[11]) ? node40217 : node40214;
																assign node40214 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node40217 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node40220 = (inp[9]) ? node40222 : 4'b0011;
														assign node40222 = (inp[11]) ? node40224 : 4'b0011;
															assign node40224 = (inp[13]) ? node40228 : node40225;
																assign node40225 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node40228 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node40231 = (inp[2]) ? node40379 : node40232;
									assign node40232 = (inp[7]) ? node40292 : node40233;
										assign node40233 = (inp[11]) ? node40253 : node40234;
											assign node40234 = (inp[1]) ? node40242 : node40235;
												assign node40235 = (inp[5]) ? node40239 : node40236;
													assign node40236 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node40239 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node40242 = (inp[5]) ? node40250 : node40243;
													assign node40243 = (inp[13]) ? node40247 : node40244;
														assign node40244 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node40247 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node40250 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node40253 = (inp[0]) ? node40271 : node40254;
												assign node40254 = (inp[13]) ? node40264 : node40255;
													assign node40255 = (inp[9]) ? node40257 : 4'b0010;
														assign node40257 = (inp[1]) ? node40261 : node40258;
															assign node40258 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node40261 = (inp[5]) ? 4'b0111 : 4'b0010;
													assign node40264 = (inp[5]) ? node40268 : node40265;
														assign node40265 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node40268 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node40271 = (inp[13]) ? node40285 : node40272;
													assign node40272 = (inp[9]) ? node40280 : node40273;
														assign node40273 = (inp[1]) ? node40277 : node40274;
															assign node40274 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node40277 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node40280 = (inp[1]) ? node40282 : 4'b0110;
															assign node40282 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node40285 = (inp[5]) ? node40289 : node40286;
														assign node40286 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node40289 = (inp[1]) ? 4'b0110 : 4'b0011;
										assign node40292 = (inp[1]) ? node40324 : node40293;
											assign node40293 = (inp[5]) ? node40309 : node40294;
												assign node40294 = (inp[13]) ? node40302 : node40295;
													assign node40295 = (inp[0]) ? node40299 : node40296;
														assign node40296 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node40299 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node40302 = (inp[0]) ? node40306 : node40303;
														assign node40303 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node40306 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node40309 = (inp[11]) ? node40317 : node40310;
													assign node40310 = (inp[0]) ? node40314 : node40311;
														assign node40311 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node40314 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node40317 = (inp[0]) ? node40321 : node40318;
														assign node40318 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node40321 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node40324 = (inp[5]) ? node40356 : node40325;
												assign node40325 = (inp[9]) ? node40339 : node40326;
													assign node40326 = (inp[10]) ? node40332 : node40327;
														assign node40327 = (inp[0]) ? node40329 : 4'b0110;
															assign node40329 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node40332 = (inp[0]) ? node40336 : node40333;
															assign node40333 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node40336 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node40339 = (inp[13]) ? node40347 : node40340;
														assign node40340 = (inp[0]) ? node40344 : node40341;
															assign node40341 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node40344 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node40347 = (inp[10]) ? 4'b0110 : node40348;
															assign node40348 = (inp[0]) ? node40352 : node40349;
																assign node40349 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node40352 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node40356 = (inp[10]) ? node40364 : node40357;
													assign node40357 = (inp[0]) ? node40361 : node40358;
														assign node40358 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node40361 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node40364 = (inp[9]) ? node40372 : node40365;
														assign node40365 = (inp[13]) ? node40367 : 4'b0011;
															assign node40367 = (inp[11]) ? node40369 : 4'b0011;
																assign node40369 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node40372 = (inp[0]) ? node40376 : node40373;
															assign node40373 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node40376 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node40379 = (inp[0]) ? node40477 : node40380;
										assign node40380 = (inp[13]) ? node40432 : node40381;
											assign node40381 = (inp[5]) ? node40395 : node40382;
												assign node40382 = (inp[11]) ? node40390 : node40383;
													assign node40383 = (inp[1]) ? node40387 : node40384;
														assign node40384 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node40387 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node40390 = (inp[7]) ? 4'b0011 : node40391;
														assign node40391 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node40395 = (inp[10]) ? node40409 : node40396;
													assign node40396 = (inp[1]) ? node40404 : node40397;
														assign node40397 = (inp[11]) ? node40401 : node40398;
															assign node40398 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node40401 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node40404 = (inp[7]) ? 4'b0011 : node40405;
															assign node40405 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node40409 = (inp[9]) ? node40419 : node40410;
														assign node40410 = (inp[11]) ? node40414 : node40411;
															assign node40411 = (inp[7]) ? 4'b0011 : 4'b0111;
															assign node40414 = (inp[1]) ? 4'b0010 : node40415;
																assign node40415 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node40419 = (inp[1]) ? node40427 : node40420;
															assign node40420 = (inp[7]) ? node40424 : node40421;
																assign node40421 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node40424 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node40427 = (inp[7]) ? node40429 : 4'b0110;
																assign node40429 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node40432 = (inp[11]) ? node40462 : node40433;
												assign node40433 = (inp[9]) ? node40445 : node40434;
													assign node40434 = (inp[7]) ? node40442 : node40435;
														assign node40435 = (inp[5]) ? node40439 : node40436;
															assign node40436 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node40439 = (inp[1]) ? 4'b0110 : 4'b0011;
														assign node40442 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node40445 = (inp[7]) ? node40453 : node40446;
														assign node40446 = (inp[10]) ? node40448 : 4'b0011;
															assign node40448 = (inp[1]) ? node40450 : 4'b0110;
																assign node40450 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node40453 = (inp[10]) ? node40455 : 4'b0110;
															assign node40455 = (inp[5]) ? node40459 : node40456;
																assign node40456 = (inp[1]) ? 4'b0110 : 4'b0011;
																assign node40459 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node40462 = (inp[7]) ? node40470 : node40463;
													assign node40463 = (inp[1]) ? node40467 : node40464;
														assign node40464 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node40467 = (inp[5]) ? 4'b0111 : 4'b0010;
													assign node40470 = (inp[1]) ? node40474 : node40471;
														assign node40471 = (inp[5]) ? 4'b0111 : 4'b0010;
														assign node40474 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node40477 = (inp[5]) ? node40505 : node40478;
											assign node40478 = (inp[11]) ? node40492 : node40479;
												assign node40479 = (inp[1]) ? node40487 : node40480;
													assign node40480 = (inp[7]) ? node40484 : node40481;
														assign node40481 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node40484 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node40487 = (inp[7]) ? node40489 : 4'b0010;
														assign node40489 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node40492 = (inp[7]) ? node40498 : node40493;
													assign node40493 = (inp[1]) ? 4'b0011 : node40494;
														assign node40494 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node40498 = (inp[1]) ? node40502 : node40499;
														assign node40499 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node40502 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node40505 = (inp[11]) ? node40519 : node40506;
												assign node40506 = (inp[7]) ? node40514 : node40507;
													assign node40507 = (inp[1]) ? node40511 : node40508;
														assign node40508 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node40511 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node40514 = (inp[1]) ? node40516 : 4'b0111;
														assign node40516 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node40519 = (inp[13]) ? node40527 : node40520;
													assign node40520 = (inp[1]) ? node40524 : node40521;
														assign node40521 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node40524 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node40527 = (inp[1]) ? node40531 : node40528;
														assign node40528 = (inp[7]) ? 4'b0110 : 4'b0011;
														assign node40531 = (inp[7]) ? 4'b0010 : 4'b0110;
							assign node40534 = (inp[5]) ? node40804 : node40535;
								assign node40535 = (inp[1]) ? node40675 : node40536;
									assign node40536 = (inp[12]) ? node40618 : node40537;
										assign node40537 = (inp[7]) ? node40593 : node40538;
											assign node40538 = (inp[10]) ? node40570 : node40539;
												assign node40539 = (inp[9]) ? node40557 : node40540;
													assign node40540 = (inp[0]) ? node40550 : node40541;
														assign node40541 = (inp[2]) ? node40547 : node40542;
															assign node40542 = (inp[11]) ? node40544 : 4'b0100;
																assign node40544 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node40547 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node40550 = (inp[13]) ? 4'b0100 : node40551;
															assign node40551 = (inp[11]) ? 4'b0100 : node40552;
																assign node40552 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node40557 = (inp[0]) ? node40565 : node40558;
														assign node40558 = (inp[11]) ? 4'b0100 : node40559;
															assign node40559 = (inp[2]) ? 4'b0101 : node40560;
																assign node40560 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node40565 = (inp[11]) ? 4'b0101 : node40566;
															assign node40566 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node40570 = (inp[2]) ? node40580 : node40571;
													assign node40571 = (inp[11]) ? node40573 : 4'b0100;
														assign node40573 = (inp[13]) ? node40577 : node40574;
															assign node40574 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node40577 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node40580 = (inp[9]) ? node40588 : node40581;
														assign node40581 = (inp[0]) ? node40585 : node40582;
															assign node40582 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node40585 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node40588 = (inp[13]) ? 4'b0100 : node40589;
															assign node40589 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node40593 = (inp[2]) ? node40601 : node40594;
												assign node40594 = (inp[11]) ? node40598 : node40595;
													assign node40595 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40598 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node40601 = (inp[13]) ? node40613 : node40602;
													assign node40602 = (inp[10]) ? node40608 : node40603;
														assign node40603 = (inp[11]) ? 4'b0001 : node40604;
															assign node40604 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node40608 = (inp[11]) ? 4'b0000 : node40609;
															assign node40609 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40613 = (inp[0]) ? 4'b0000 : node40614;
														assign node40614 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node40618 = (inp[7]) ? node40652 : node40619;
											assign node40619 = (inp[2]) ? node40627 : node40620;
												assign node40620 = (inp[11]) ? node40624 : node40621;
													assign node40621 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40624 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node40627 = (inp[0]) ? node40645 : node40628;
													assign node40628 = (inp[9]) ? node40638 : node40629;
														assign node40629 = (inp[10]) ? node40631 : 4'b0001;
															assign node40631 = (inp[11]) ? node40635 : node40632;
																assign node40632 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node40635 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node40638 = (inp[11]) ? node40642 : node40639;
															assign node40639 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node40642 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node40645 = (inp[11]) ? node40649 : node40646;
														assign node40646 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node40649 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node40652 = (inp[11]) ? node40664 : node40653;
												assign node40653 = (inp[0]) ? node40659 : node40654;
													assign node40654 = (inp[13]) ? node40656 : 4'b0001;
														assign node40656 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node40659 = (inp[13]) ? node40661 : 4'b0000;
														assign node40661 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node40664 = (inp[0]) ? node40670 : node40665;
													assign node40665 = (inp[13]) ? node40667 : 4'b0000;
														assign node40667 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node40670 = (inp[13]) ? node40672 : 4'b0001;
														assign node40672 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node40675 = (inp[7]) ? node40747 : node40676;
										assign node40676 = (inp[12]) ? node40724 : node40677;
											assign node40677 = (inp[10]) ? node40697 : node40678;
												assign node40678 = (inp[2]) ? node40690 : node40679;
													assign node40679 = (inp[9]) ? node40681 : 4'b0000;
														assign node40681 = (inp[11]) ? 4'b0000 : node40682;
															assign node40682 = (inp[0]) ? node40686 : node40683;
																assign node40683 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node40686 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node40690 = (inp[11]) ? node40694 : node40691;
														assign node40691 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node40694 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node40697 = (inp[13]) ? node40709 : node40698;
													assign node40698 = (inp[11]) ? node40704 : node40699;
														assign node40699 = (inp[2]) ? node40701 : 4'b0001;
															assign node40701 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node40704 = (inp[0]) ? 4'b0000 : node40705;
															assign node40705 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node40709 = (inp[9]) ? node40717 : node40710;
														assign node40710 = (inp[11]) ? node40714 : node40711;
															assign node40711 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node40714 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node40717 = (inp[0]) ? node40721 : node40718;
															assign node40718 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node40721 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node40724 = (inp[0]) ? node40736 : node40725;
												assign node40725 = (inp[11]) ? node40731 : node40726;
													assign node40726 = (inp[13]) ? 4'b0101 : node40727;
														assign node40727 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40731 = (inp[2]) ? 4'b0100 : node40732;
														assign node40732 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node40736 = (inp[11]) ? node40742 : node40737;
													assign node40737 = (inp[13]) ? 4'b0100 : node40738;
														assign node40738 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node40742 = (inp[13]) ? 4'b0101 : node40743;
														assign node40743 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node40747 = (inp[13]) ? node40789 : node40748;
											assign node40748 = (inp[0]) ? node40774 : node40749;
												assign node40749 = (inp[9]) ? node40767 : node40750;
													assign node40750 = (inp[10]) ? node40760 : node40751;
														assign node40751 = (inp[12]) ? 4'b0101 : node40752;
															assign node40752 = (inp[2]) ? node40756 : node40753;
																assign node40753 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node40756 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node40760 = (inp[11]) ? node40764 : node40761;
															assign node40761 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node40764 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40767 = (inp[11]) ? node40771 : node40768;
														assign node40768 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40771 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node40774 = (inp[10]) ? node40782 : node40775;
													assign node40775 = (inp[2]) ? node40779 : node40776;
														assign node40776 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node40779 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node40782 = (inp[11]) ? node40786 : node40783;
														assign node40783 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node40786 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node40789 = (inp[9]) ? node40797 : node40790;
												assign node40790 = (inp[11]) ? node40794 : node40791;
													assign node40791 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node40794 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node40797 = (inp[0]) ? node40801 : node40798;
													assign node40798 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node40801 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node40804 = (inp[1]) ? node40952 : node40805;
									assign node40805 = (inp[7]) ? node40859 : node40806;
										assign node40806 = (inp[12]) ? node40830 : node40807;
											assign node40807 = (inp[0]) ? node40819 : node40808;
												assign node40808 = (inp[11]) ? node40814 : node40809;
													assign node40809 = (inp[2]) ? 4'b0000 : node40810;
														assign node40810 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node40814 = (inp[13]) ? 4'b0001 : node40815;
														assign node40815 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node40819 = (inp[11]) ? node40825 : node40820;
													assign node40820 = (inp[2]) ? 4'b0001 : node40821;
														assign node40821 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node40825 = (inp[2]) ? 4'b0000 : node40826;
														assign node40826 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node40830 = (inp[13]) ? node40846 : node40831;
												assign node40831 = (inp[0]) ? node40839 : node40832;
													assign node40832 = (inp[2]) ? node40836 : node40833;
														assign node40833 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node40836 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node40839 = (inp[11]) ? node40843 : node40840;
														assign node40840 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node40843 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node40846 = (inp[2]) ? node40852 : node40847;
													assign node40847 = (inp[0]) ? node40849 : 4'b0101;
														assign node40849 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node40852 = (inp[0]) ? node40856 : node40853;
														assign node40853 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node40856 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node40859 = (inp[11]) ? node40899 : node40860;
											assign node40860 = (inp[2]) ? node40892 : node40861;
												assign node40861 = (inp[13]) ? node40875 : node40862;
													assign node40862 = (inp[10]) ? node40870 : node40863;
														assign node40863 = (inp[12]) ? node40867 : node40864;
															assign node40864 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node40867 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node40870 = (inp[12]) ? node40872 : 4'b0100;
															assign node40872 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40875 = (inp[10]) ? node40887 : node40876;
														assign node40876 = (inp[9]) ? node40882 : node40877;
															assign node40877 = (inp[12]) ? 4'b0100 : node40878;
																assign node40878 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node40882 = (inp[0]) ? 4'b0101 : node40883;
																assign node40883 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node40887 = (inp[9]) ? node40889 : 4'b0101;
															assign node40889 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node40892 = (inp[0]) ? node40896 : node40893;
													assign node40893 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node40896 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node40899 = (inp[10]) ? node40921 : node40900;
												assign node40900 = (inp[13]) ? node40914 : node40901;
													assign node40901 = (inp[0]) ? node40903 : 4'b0100;
														assign node40903 = (inp[9]) ? node40909 : node40904;
															assign node40904 = (inp[12]) ? node40906 : 4'b0100;
																assign node40906 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node40909 = (inp[12]) ? 4'b0100 : node40910;
																assign node40910 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40914 = (inp[12]) ? node40918 : node40915;
														assign node40915 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node40918 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node40921 = (inp[13]) ? node40945 : node40922;
													assign node40922 = (inp[9]) ? node40932 : node40923;
														assign node40923 = (inp[12]) ? node40925 : 4'b0101;
															assign node40925 = (inp[0]) ? node40929 : node40926;
																assign node40926 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node40929 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40932 = (inp[12]) ? node40938 : node40933;
															assign node40933 = (inp[0]) ? 4'b0100 : node40934;
																assign node40934 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node40938 = (inp[2]) ? node40942 : node40939;
																assign node40939 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node40942 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40945 = (inp[0]) ? node40949 : node40946;
														assign node40946 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node40949 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node40952 = (inp[12]) ? node41000 : node40953;
										assign node40953 = (inp[7]) ? node40977 : node40954;
											assign node40954 = (inp[0]) ? node40966 : node40955;
												assign node40955 = (inp[11]) ? node40961 : node40956;
													assign node40956 = (inp[2]) ? node40958 : 4'b0101;
														assign node40958 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node40961 = (inp[13]) ? node40963 : 4'b0100;
														assign node40963 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node40966 = (inp[11]) ? node40972 : node40967;
													assign node40967 = (inp[2]) ? node40969 : 4'b0100;
														assign node40969 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node40972 = (inp[2]) ? node40974 : 4'b0101;
														assign node40974 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node40977 = (inp[11]) ? node40989 : node40978;
												assign node40978 = (inp[0]) ? node40984 : node40979;
													assign node40979 = (inp[13]) ? 4'b0000 : node40980;
														assign node40980 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node40984 = (inp[13]) ? 4'b0001 : node40985;
														assign node40985 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node40989 = (inp[0]) ? node40995 : node40990;
													assign node40990 = (inp[2]) ? 4'b0001 : node40991;
														assign node40991 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node40995 = (inp[13]) ? 4'b0000 : node40996;
														assign node40996 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node41000 = (inp[13]) ? node41026 : node41001;
											assign node41001 = (inp[2]) ? node41009 : node41002;
												assign node41002 = (inp[0]) ? node41006 : node41003;
													assign node41003 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node41006 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node41009 = (inp[7]) ? node41019 : node41010;
													assign node41010 = (inp[9]) ? 4'b0001 : node41011;
														assign node41011 = (inp[11]) ? node41015 : node41012;
															assign node41012 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node41015 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node41019 = (inp[11]) ? node41023 : node41020;
														assign node41020 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41023 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node41026 = (inp[0]) ? node41030 : node41027;
												assign node41027 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node41030 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node41033 = (inp[1]) ? node41383 : node41034;
							assign node41034 = (inp[15]) ? node41152 : node41035;
								assign node41035 = (inp[7]) ? node41059 : node41036;
									assign node41036 = (inp[5]) ? node41048 : node41037;
										assign node41037 = (inp[0]) ? node41043 : node41038;
											assign node41038 = (inp[13]) ? node41040 : 4'b0000;
												assign node41040 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node41043 = (inp[13]) ? node41045 : 4'b0001;
												assign node41045 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node41048 = (inp[0]) ? node41054 : node41049;
											assign node41049 = (inp[12]) ? node41051 : 4'b0001;
												assign node41051 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node41054 = (inp[12]) ? node41056 : 4'b0000;
												assign node41056 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node41059 = (inp[9]) ? node41103 : node41060;
										assign node41060 = (inp[13]) ? node41076 : node41061;
											assign node41061 = (inp[11]) ? node41069 : node41062;
												assign node41062 = (inp[12]) ? node41066 : node41063;
													assign node41063 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node41066 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node41069 = (inp[12]) ? node41073 : node41070;
													assign node41070 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node41073 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node41076 = (inp[10]) ? node41092 : node41077;
												assign node41077 = (inp[5]) ? node41085 : node41078;
													assign node41078 = (inp[0]) ? node41082 : node41079;
														assign node41079 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node41082 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node41085 = (inp[12]) ? node41089 : node41086;
														assign node41086 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node41089 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node41092 = (inp[5]) ? 4'b0101 : node41093;
													assign node41093 = (inp[11]) ? 4'b0101 : node41094;
														assign node41094 = (inp[0]) ? node41098 : node41095;
															assign node41095 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node41098 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node41103 = (inp[2]) ? node41137 : node41104;
											assign node41104 = (inp[11]) ? node41112 : node41105;
												assign node41105 = (inp[0]) ? node41109 : node41106;
													assign node41106 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node41109 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node41112 = (inp[13]) ? node41120 : node41113;
													assign node41113 = (inp[12]) ? node41117 : node41114;
														assign node41114 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node41117 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node41120 = (inp[10]) ? node41128 : node41121;
														assign node41121 = (inp[12]) ? node41125 : node41122;
															assign node41122 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node41125 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node41128 = (inp[5]) ? node41130 : 4'b0100;
															assign node41130 = (inp[12]) ? node41134 : node41131;
																assign node41131 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node41134 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node41137 = (inp[5]) ? node41145 : node41138;
												assign node41138 = (inp[12]) ? node41142 : node41139;
													assign node41139 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node41142 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node41145 = (inp[12]) ? node41149 : node41146;
													assign node41146 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node41149 = (inp[0]) ? 4'b0100 : 4'b0101;
								assign node41152 = (inp[2]) ? node41308 : node41153;
									assign node41153 = (inp[9]) ? node41265 : node41154;
										assign node41154 = (inp[7]) ? node41200 : node41155;
											assign node41155 = (inp[10]) ? node41179 : node41156;
												assign node41156 = (inp[5]) ? node41168 : node41157;
													assign node41157 = (inp[0]) ? node41163 : node41158;
														assign node41158 = (inp[13]) ? node41160 : 4'b0100;
															assign node41160 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node41163 = (inp[13]) ? node41165 : 4'b0101;
															assign node41165 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node41168 = (inp[0]) ? node41174 : node41169;
														assign node41169 = (inp[13]) ? node41171 : 4'b0101;
															assign node41171 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node41174 = (inp[12]) ? 4'b0100 : node41175;
															assign node41175 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node41179 = (inp[13]) ? node41185 : node41180;
													assign node41180 = (inp[0]) ? node41182 : 4'b0100;
														assign node41182 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node41185 = (inp[0]) ? node41193 : node41186;
														assign node41186 = (inp[5]) ? node41190 : node41187;
															assign node41187 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node41190 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node41193 = (inp[11]) ? node41195 : 4'b0100;
															assign node41195 = (inp[5]) ? 4'b0100 : node41196;
																assign node41196 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node41200 = (inp[11]) ? node41236 : node41201;
												assign node41201 = (inp[10]) ? node41223 : node41202;
													assign node41202 = (inp[13]) ? node41212 : node41203;
														assign node41203 = (inp[5]) ? node41207 : node41204;
															assign node41204 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node41207 = (inp[12]) ? 4'b0101 : node41208;
																assign node41208 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node41212 = (inp[5]) ? node41218 : node41213;
															assign node41213 = (inp[12]) ? 4'b0101 : node41214;
																assign node41214 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node41218 = (inp[0]) ? 4'b0100 : node41219;
																assign node41219 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node41223 = (inp[5]) ? node41229 : node41224;
														assign node41224 = (inp[0]) ? node41226 : 4'b0100;
															assign node41226 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node41229 = (inp[0]) ? node41233 : node41230;
															assign node41230 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node41233 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node41236 = (inp[10]) ? node41248 : node41237;
													assign node41237 = (inp[5]) ? node41239 : 4'b0100;
														assign node41239 = (inp[13]) ? node41245 : node41240;
															assign node41240 = (inp[12]) ? node41242 : 4'b0100;
																assign node41242 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node41245 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node41248 = (inp[13]) ? node41258 : node41249;
														assign node41249 = (inp[5]) ? node41255 : node41250;
															assign node41250 = (inp[0]) ? node41252 : 4'b0101;
																assign node41252 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node41255 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node41258 = (inp[12]) ? node41262 : node41259;
															assign node41259 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node41262 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node41265 = (inp[5]) ? node41295 : node41266;
											assign node41266 = (inp[0]) ? node41276 : node41267;
												assign node41267 = (inp[12]) ? node41273 : node41268;
													assign node41268 = (inp[7]) ? 4'b0100 : node41269;
														assign node41269 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node41273 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node41276 = (inp[13]) ? node41282 : node41277;
													assign node41277 = (inp[7]) ? node41279 : 4'b0101;
														assign node41279 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node41282 = (inp[11]) ? node41288 : node41283;
														assign node41283 = (inp[12]) ? 4'b0101 : node41284;
															assign node41284 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node41288 = (inp[7]) ? node41292 : node41289;
															assign node41289 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node41292 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node41295 = (inp[0]) ? node41303 : node41296;
												assign node41296 = (inp[12]) ? 4'b0101 : node41297;
													assign node41297 = (inp[13]) ? 4'b0100 : node41298;
														assign node41298 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node41303 = (inp[12]) ? 4'b0100 : node41304;
													assign node41304 = (inp[13]) ? 4'b0101 : 4'b0100;
									assign node41308 = (inp[7]) ? node41332 : node41309;
										assign node41309 = (inp[5]) ? node41321 : node41310;
											assign node41310 = (inp[0]) ? node41316 : node41311;
												assign node41311 = (inp[12]) ? 4'b0100 : node41312;
													assign node41312 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node41316 = (inp[12]) ? 4'b0101 : node41317;
													assign node41317 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node41321 = (inp[0]) ? node41327 : node41322;
												assign node41322 = (inp[12]) ? 4'b0101 : node41323;
													assign node41323 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node41327 = (inp[12]) ? 4'b0100 : node41328;
													assign node41328 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node41332 = (inp[10]) ? node41340 : node41333;
											assign node41333 = (inp[0]) ? node41337 : node41334;
												assign node41334 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node41337 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node41340 = (inp[11]) ? node41362 : node41341;
												assign node41341 = (inp[5]) ? node41355 : node41342;
													assign node41342 = (inp[9]) ? node41348 : node41343;
														assign node41343 = (inp[0]) ? node41345 : 4'b0101;
															assign node41345 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node41348 = (inp[0]) ? node41352 : node41349;
															assign node41349 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node41352 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node41355 = (inp[0]) ? node41359 : node41356;
														assign node41356 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node41359 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node41362 = (inp[5]) ? node41374 : node41363;
													assign node41363 = (inp[13]) ? node41369 : node41364;
														assign node41364 = (inp[0]) ? 4'b0100 : node41365;
															assign node41365 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node41369 = (inp[0]) ? 4'b0101 : node41370;
															assign node41370 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node41374 = (inp[13]) ? node41376 : 4'b0101;
														assign node41376 = (inp[9]) ? node41378 : 4'b0100;
															assign node41378 = (inp[0]) ? node41380 : 4'b0101;
																assign node41380 = (inp[12]) ? 4'b0100 : 4'b0101;
							assign node41383 = (inp[7]) ? node41581 : node41384;
								assign node41384 = (inp[15]) ? node41408 : node41385;
									assign node41385 = (inp[0]) ? node41397 : node41386;
										assign node41386 = (inp[5]) ? node41392 : node41387;
											assign node41387 = (inp[13]) ? 4'b0100 : node41388;
												assign node41388 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node41392 = (inp[13]) ? 4'b0101 : node41393;
												assign node41393 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node41397 = (inp[5]) ? node41403 : node41398;
											assign node41398 = (inp[13]) ? 4'b0101 : node41399;
												assign node41399 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node41403 = (inp[12]) ? node41405 : 4'b0100;
												assign node41405 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node41408 = (inp[2]) ? node41502 : node41409;
										assign node41409 = (inp[10]) ? node41465 : node41410;
											assign node41410 = (inp[9]) ? node41438 : node41411;
												assign node41411 = (inp[11]) ? node41433 : node41412;
													assign node41412 = (inp[12]) ? node41422 : node41413;
														assign node41413 = (inp[13]) ? 4'b0000 : node41414;
															assign node41414 = (inp[0]) ? node41418 : node41415;
																assign node41415 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node41418 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node41422 = (inp[13]) ? node41428 : node41423;
															assign node41423 = (inp[0]) ? node41425 : 4'b0001;
																assign node41425 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node41428 = (inp[5]) ? 4'b0001 : node41429;
																assign node41429 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node41433 = (inp[0]) ? 4'b0001 : node41434;
														assign node41434 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node41438 = (inp[12]) ? node41452 : node41439;
													assign node41439 = (inp[13]) ? node41445 : node41440;
														assign node41440 = (inp[5]) ? node41442 : 4'b0001;
															assign node41442 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41445 = (inp[5]) ? node41449 : node41446;
															assign node41446 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node41449 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node41452 = (inp[11]) ? node41458 : node41453;
														assign node41453 = (inp[5]) ? node41455 : 4'b0001;
															assign node41455 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node41458 = (inp[13]) ? 4'b0000 : node41459;
															assign node41459 = (inp[0]) ? 4'b0000 : node41460;
																assign node41460 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node41465 = (inp[9]) ? node41489 : node41466;
												assign node41466 = (inp[12]) ? node41482 : node41467;
													assign node41467 = (inp[0]) ? node41475 : node41468;
														assign node41468 = (inp[13]) ? node41472 : node41469;
															assign node41469 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node41472 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node41475 = (inp[13]) ? node41479 : node41476;
															assign node41476 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node41479 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node41482 = (inp[5]) ? node41486 : node41483;
														assign node41483 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41486 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node41489 = (inp[13]) ? node41495 : node41490;
													assign node41490 = (inp[0]) ? 4'b0001 : node41491;
														assign node41491 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node41495 = (inp[0]) ? node41499 : node41496;
														assign node41496 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node41499 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node41502 = (inp[13]) ? node41542 : node41503;
											assign node41503 = (inp[11]) ? node41521 : node41504;
												assign node41504 = (inp[5]) ? node41510 : node41505;
													assign node41505 = (inp[0]) ? node41507 : 4'b0000;
														assign node41507 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node41510 = (inp[9]) ? node41516 : node41511;
														assign node41511 = (inp[12]) ? node41513 : 4'b0000;
															assign node41513 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node41516 = (inp[12]) ? node41518 : 4'b0001;
															assign node41518 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node41521 = (inp[12]) ? node41535 : node41522;
													assign node41522 = (inp[9]) ? node41530 : node41523;
														assign node41523 = (inp[0]) ? node41527 : node41524;
															assign node41524 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node41527 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node41530 = (inp[0]) ? node41532 : 4'b0000;
															assign node41532 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node41535 = (inp[0]) ? node41539 : node41536;
														assign node41536 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node41539 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node41542 = (inp[11]) ? node41558 : node41543;
												assign node41543 = (inp[9]) ? node41551 : node41544;
													assign node41544 = (inp[5]) ? node41548 : node41545;
														assign node41545 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41548 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node41551 = (inp[5]) ? node41555 : node41552;
														assign node41552 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41555 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node41558 = (inp[9]) ? node41566 : node41559;
													assign node41559 = (inp[5]) ? node41563 : node41560;
														assign node41560 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node41563 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node41566 = (inp[12]) ? node41574 : node41567;
														assign node41567 = (inp[5]) ? node41571 : node41568;
															assign node41568 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node41571 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node41574 = (inp[0]) ? node41578 : node41575;
															assign node41575 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41578 = (inp[5]) ? 4'b0000 : 4'b0001;
								assign node41581 = (inp[0]) ? node41587 : node41582;
									assign node41582 = (inp[15]) ? 4'b0001 : node41583;
										assign node41583 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node41587 = (inp[15]) ? 4'b0000 : node41588;
										assign node41588 = (inp[13]) ? 4'b0000 : 4'b0001;
				assign node41592 = (inp[15]) ? node43496 : node41593;
					assign node41593 = (inp[14]) ? node42849 : node41594;
						assign node41594 = (inp[5]) ? node42374 : node41595;
							assign node41595 = (inp[7]) ? node41991 : node41596;
								assign node41596 = (inp[9]) ? node41780 : node41597;
									assign node41597 = (inp[1]) ? node41671 : node41598;
										assign node41598 = (inp[0]) ? node41646 : node41599;
											assign node41599 = (inp[10]) ? node41617 : node41600;
												assign node41600 = (inp[11]) ? node41610 : node41601;
													assign node41601 = (inp[13]) ? node41603 : 4'b0010;
														assign node41603 = (inp[4]) ? node41605 : 4'b0011;
															assign node41605 = (inp[12]) ? 4'b0011 : node41606;
																assign node41606 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node41610 = (inp[13]) ? node41612 : 4'b0011;
														assign node41612 = (inp[4]) ? node41614 : 4'b0010;
															assign node41614 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node41617 = (inp[12]) ? node41631 : node41618;
													assign node41618 = (inp[11]) ? node41626 : node41619;
														assign node41619 = (inp[13]) ? 4'b0011 : node41620;
															assign node41620 = (inp[4]) ? node41622 : 4'b0010;
																assign node41622 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node41626 = (inp[13]) ? 4'b0010 : node41627;
															assign node41627 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node41631 = (inp[4]) ? node41639 : node41632;
														assign node41632 = (inp[13]) ? node41636 : node41633;
															assign node41633 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node41636 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41639 = (inp[13]) ? node41643 : node41640;
															assign node41640 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node41643 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node41646 = (inp[2]) ? node41654 : node41647;
												assign node41647 = (inp[13]) ? node41651 : node41648;
													assign node41648 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node41651 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node41654 = (inp[11]) ? node41666 : node41655;
													assign node41655 = (inp[13]) ? node41661 : node41656;
														assign node41656 = (inp[4]) ? node41658 : 4'b0010;
															assign node41658 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node41661 = (inp[4]) ? node41663 : 4'b0011;
															assign node41663 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node41666 = (inp[13]) ? node41668 : 4'b0011;
														assign node41668 = (inp[12]) ? 4'b0010 : 4'b0011;
										assign node41671 = (inp[4]) ? node41743 : node41672;
											assign node41672 = (inp[11]) ? node41704 : node41673;
												assign node41673 = (inp[10]) ? node41689 : node41674;
													assign node41674 = (inp[2]) ? node41680 : node41675;
														assign node41675 = (inp[13]) ? node41677 : 4'b0010;
															assign node41677 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node41680 = (inp[0]) ? 4'b0011 : node41681;
															assign node41681 = (inp[12]) ? node41685 : node41682;
																assign node41682 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41685 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node41689 = (inp[2]) ? node41697 : node41690;
														assign node41690 = (inp[12]) ? node41694 : node41691;
															assign node41691 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node41694 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node41697 = (inp[12]) ? node41701 : node41698;
															assign node41698 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node41701 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node41704 = (inp[13]) ? node41720 : node41705;
													assign node41705 = (inp[10]) ? node41713 : node41706;
														assign node41706 = (inp[12]) ? node41710 : node41707;
															assign node41707 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node41710 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node41713 = (inp[2]) ? node41717 : node41714;
															assign node41714 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node41717 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node41720 = (inp[0]) ? node41734 : node41721;
														assign node41721 = (inp[10]) ? node41727 : node41722;
															assign node41722 = (inp[2]) ? node41724 : 4'b0011;
																assign node41724 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node41727 = (inp[12]) ? node41731 : node41728;
																assign node41728 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node41731 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node41734 = (inp[10]) ? 4'b0010 : node41735;
															assign node41735 = (inp[12]) ? node41739 : node41736;
																assign node41736 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node41739 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node41743 = (inp[10]) ? node41761 : node41744;
												assign node41744 = (inp[13]) ? node41752 : node41745;
													assign node41745 = (inp[11]) ? node41747 : 4'b0010;
														assign node41747 = (inp[2]) ? node41749 : 4'b0011;
															assign node41749 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node41752 = (inp[11]) ? node41758 : node41753;
														assign node41753 = (inp[12]) ? node41755 : 4'b0011;
															assign node41755 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node41758 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node41761 = (inp[13]) ? node41771 : node41762;
													assign node41762 = (inp[11]) ? node41766 : node41763;
														assign node41763 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node41766 = (inp[12]) ? node41768 : 4'b0011;
															assign node41768 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node41771 = (inp[11]) ? node41775 : node41772;
														assign node41772 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node41775 = (inp[2]) ? node41777 : 4'b0010;
															assign node41777 = (inp[12]) ? 4'b0011 : 4'b0010;
									assign node41780 = (inp[10]) ? node41912 : node41781;
										assign node41781 = (inp[0]) ? node41853 : node41782;
											assign node41782 = (inp[4]) ? node41828 : node41783;
												assign node41783 = (inp[1]) ? node41809 : node41784;
													assign node41784 = (inp[2]) ? node41800 : node41785;
														assign node41785 = (inp[12]) ? node41793 : node41786;
															assign node41786 = (inp[13]) ? node41790 : node41787;
																assign node41787 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41790 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node41793 = (inp[13]) ? node41797 : node41794;
																assign node41794 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41797 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41800 = (inp[12]) ? node41802 : 4'b0011;
															assign node41802 = (inp[13]) ? node41806 : node41803;
																assign node41803 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41806 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node41809 = (inp[12]) ? node41819 : node41810;
														assign node41810 = (inp[2]) ? 4'b0010 : node41811;
															assign node41811 = (inp[13]) ? node41815 : node41812;
																assign node41812 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41815 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node41819 = (inp[13]) ? 4'b0011 : node41820;
															assign node41820 = (inp[2]) ? node41824 : node41821;
																assign node41821 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node41824 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node41828 = (inp[1]) ? node41840 : node41829;
													assign node41829 = (inp[11]) ? node41831 : 4'b0010;
														assign node41831 = (inp[12]) ? 4'b0011 : node41832;
															assign node41832 = (inp[2]) ? node41836 : node41833;
																assign node41833 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node41836 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node41840 = (inp[11]) ? node41842 : 4'b0011;
														assign node41842 = (inp[13]) ? node41848 : node41843;
															assign node41843 = (inp[12]) ? node41845 : 4'b0011;
																assign node41845 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node41848 = (inp[2]) ? node41850 : 4'b0010;
																assign node41850 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node41853 = (inp[13]) ? node41881 : node41854;
												assign node41854 = (inp[11]) ? node41872 : node41855;
													assign node41855 = (inp[2]) ? node41863 : node41856;
														assign node41856 = (inp[4]) ? 4'b0010 : node41857;
															assign node41857 = (inp[1]) ? node41859 : 4'b0010;
																assign node41859 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node41863 = (inp[4]) ? node41865 : 4'b0010;
															assign node41865 = (inp[1]) ? node41869 : node41866;
																assign node41866 = (inp[12]) ? 4'b0010 : 4'b0011;
																assign node41869 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node41872 = (inp[1]) ? node41874 : 4'b0011;
														assign node41874 = (inp[12]) ? node41876 : 4'b0011;
															assign node41876 = (inp[2]) ? 4'b0010 : node41877;
																assign node41877 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node41881 = (inp[11]) ? node41895 : node41882;
													assign node41882 = (inp[2]) ? node41884 : 4'b0011;
														assign node41884 = (inp[4]) ? node41890 : node41885;
															assign node41885 = (inp[12]) ? 4'b0011 : node41886;
																assign node41886 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node41890 = (inp[12]) ? 4'b0010 : node41891;
																assign node41891 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node41895 = (inp[2]) ? node41901 : node41896;
														assign node41896 = (inp[12]) ? node41898 : 4'b0010;
															assign node41898 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node41901 = (inp[12]) ? node41907 : node41902;
															assign node41902 = (inp[1]) ? node41904 : 4'b0011;
																assign node41904 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node41907 = (inp[4]) ? node41909 : 4'b0010;
																assign node41909 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node41912 = (inp[1]) ? node41944 : node41913;
											assign node41913 = (inp[11]) ? node41929 : node41914;
												assign node41914 = (inp[13]) ? node41922 : node41915;
													assign node41915 = (inp[2]) ? node41917 : 4'b0010;
														assign node41917 = (inp[12]) ? 4'b0010 : node41918;
															assign node41918 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node41922 = (inp[2]) ? node41924 : 4'b0011;
														assign node41924 = (inp[12]) ? 4'b0011 : node41925;
															assign node41925 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node41929 = (inp[13]) ? node41937 : node41930;
													assign node41930 = (inp[4]) ? node41932 : 4'b0011;
														assign node41932 = (inp[12]) ? 4'b0011 : node41933;
															assign node41933 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node41937 = (inp[12]) ? 4'b0010 : node41938;
														assign node41938 = (inp[4]) ? node41940 : 4'b0010;
															assign node41940 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node41944 = (inp[4]) ? node41972 : node41945;
												assign node41945 = (inp[13]) ? node41965 : node41946;
													assign node41946 = (inp[0]) ? node41958 : node41947;
														assign node41947 = (inp[12]) ? node41953 : node41948;
															assign node41948 = (inp[11]) ? 4'b0010 : node41949;
																assign node41949 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node41953 = (inp[11]) ? 4'b0011 : node41954;
																assign node41954 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node41958 = (inp[12]) ? node41960 : 4'b0010;
															assign node41960 = (inp[11]) ? 4'b0010 : node41961;
																assign node41961 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node41965 = (inp[2]) ? 4'b0010 : node41966;
														assign node41966 = (inp[12]) ? 4'b0010 : node41967;
															assign node41967 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node41972 = (inp[11]) ? node41984 : node41973;
													assign node41973 = (inp[13]) ? node41979 : node41974;
														assign node41974 = (inp[12]) ? node41976 : 4'b0010;
															assign node41976 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node41979 = (inp[2]) ? node41981 : 4'b0011;
															assign node41981 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node41984 = (inp[13]) ? node41986 : 4'b0011;
														assign node41986 = (inp[12]) ? node41988 : 4'b0010;
															assign node41988 = (inp[2]) ? 4'b0011 : 4'b0010;
								assign node41991 = (inp[9]) ? node42229 : node41992;
									assign node41992 = (inp[10]) ? node42098 : node41993;
										assign node41993 = (inp[4]) ? node42055 : node41994;
											assign node41994 = (inp[0]) ? node42018 : node41995;
												assign node41995 = (inp[2]) ? node42003 : node41996;
													assign node41996 = (inp[13]) ? node42000 : node41997;
														assign node41997 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42000 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42003 = (inp[13]) ? node42007 : node42004;
														assign node42004 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42007 = (inp[1]) ? node42013 : node42008;
															assign node42008 = (inp[12]) ? 4'b0111 : node42009;
																assign node42009 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42013 = (inp[11]) ? node42015 : 4'b0110;
																assign node42015 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node42018 = (inp[2]) ? node42038 : node42019;
													assign node42019 = (inp[1]) ? node42027 : node42020;
														assign node42020 = (inp[13]) ? node42024 : node42021;
															assign node42021 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42024 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42027 = (inp[12]) ? node42033 : node42028;
															assign node42028 = (inp[13]) ? 4'b0110 : node42029;
																assign node42029 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42033 = (inp[13]) ? node42035 : 4'b0110;
																assign node42035 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42038 = (inp[11]) ? node42050 : node42039;
														assign node42039 = (inp[13]) ? node42045 : node42040;
															assign node42040 = (inp[12]) ? 4'b0110 : node42041;
																assign node42041 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42045 = (inp[1]) ? node42047 : 4'b0111;
																assign node42047 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node42050 = (inp[12]) ? 4'b0111 : node42051;
															assign node42051 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node42055 = (inp[12]) ? node42083 : node42056;
												assign node42056 = (inp[0]) ? node42074 : node42057;
													assign node42057 = (inp[1]) ? node42069 : node42058;
														assign node42058 = (inp[2]) ? node42064 : node42059;
															assign node42059 = (inp[11]) ? node42061 : 4'b0111;
																assign node42061 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node42064 = (inp[13]) ? node42066 : 4'b0110;
																assign node42066 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42069 = (inp[13]) ? 4'b0110 : node42070;
															assign node42070 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node42074 = (inp[1]) ? 4'b0111 : node42075;
														assign node42075 = (inp[2]) ? 4'b0111 : node42076;
															assign node42076 = (inp[13]) ? node42078 : 4'b0110;
																assign node42078 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42083 = (inp[13]) ? node42089 : node42084;
													assign node42084 = (inp[11]) ? node42086 : 4'b0110;
														assign node42086 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node42089 = (inp[11]) ? node42093 : node42090;
														assign node42090 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42093 = (inp[1]) ? 4'b0110 : node42094;
															assign node42094 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node42098 = (inp[0]) ? node42162 : node42099;
											assign node42099 = (inp[12]) ? node42135 : node42100;
												assign node42100 = (inp[1]) ? node42116 : node42101;
													assign node42101 = (inp[13]) ? node42111 : node42102;
														assign node42102 = (inp[2]) ? node42106 : node42103;
															assign node42103 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42106 = (inp[11]) ? 4'b0110 : node42107;
																assign node42107 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node42111 = (inp[11]) ? 4'b0110 : node42112;
															assign node42112 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node42116 = (inp[11]) ? node42124 : node42117;
														assign node42117 = (inp[13]) ? 4'b0111 : node42118;
															assign node42118 = (inp[2]) ? node42120 : 4'b0110;
																assign node42120 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node42124 = (inp[13]) ? node42130 : node42125;
															assign node42125 = (inp[2]) ? node42127 : 4'b0111;
																assign node42127 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node42130 = (inp[4]) ? 4'b0110 : node42131;
																assign node42131 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node42135 = (inp[13]) ? node42145 : node42136;
													assign node42136 = (inp[11]) ? 4'b0111 : node42137;
														assign node42137 = (inp[1]) ? 4'b0110 : node42138;
															assign node42138 = (inp[2]) ? node42140 : 4'b0111;
																assign node42140 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node42145 = (inp[11]) ? node42155 : node42146;
														assign node42146 = (inp[1]) ? 4'b0111 : node42147;
															assign node42147 = (inp[4]) ? node42151 : node42148;
																assign node42148 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node42151 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node42155 = (inp[1]) ? 4'b0110 : node42156;
															assign node42156 = (inp[2]) ? node42158 : 4'b0111;
																assign node42158 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node42162 = (inp[4]) ? node42198 : node42163;
												assign node42163 = (inp[12]) ? node42183 : node42164;
													assign node42164 = (inp[13]) ? node42174 : node42165;
														assign node42165 = (inp[1]) ? node42167 : 4'b0110;
															assign node42167 = (inp[11]) ? node42171 : node42168;
																assign node42168 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node42171 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node42174 = (inp[11]) ? node42180 : node42175;
															assign node42175 = (inp[2]) ? node42177 : 4'b0111;
																assign node42177 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node42180 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node42183 = (inp[1]) ? node42191 : node42184;
														assign node42184 = (inp[11]) ? node42186 : 4'b0110;
															assign node42186 = (inp[2]) ? 4'b0110 : node42187;
																assign node42187 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node42191 = (inp[11]) ? node42195 : node42192;
															assign node42192 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node42195 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node42198 = (inp[12]) ? node42216 : node42199;
													assign node42199 = (inp[1]) ? node42209 : node42200;
														assign node42200 = (inp[2]) ? 4'b0110 : node42201;
															assign node42201 = (inp[13]) ? node42205 : node42202;
																assign node42202 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node42205 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42209 = (inp[13]) ? node42213 : node42210;
															assign node42210 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42213 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42216 = (inp[1]) ? node42224 : node42217;
														assign node42217 = (inp[2]) ? 4'b0111 : node42218;
															assign node42218 = (inp[11]) ? node42220 : 4'b0111;
																assign node42220 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node42224 = (inp[11]) ? node42226 : 4'b0110;
															assign node42226 = (inp[13]) ? 4'b0110 : 4'b0111;
									assign node42229 = (inp[4]) ? node42329 : node42230;
										assign node42230 = (inp[0]) ? node42272 : node42231;
											assign node42231 = (inp[12]) ? node42251 : node42232;
												assign node42232 = (inp[11]) ? node42242 : node42233;
													assign node42233 = (inp[13]) ? node42237 : node42234;
														assign node42234 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42237 = (inp[1]) ? node42239 : 4'b0111;
															assign node42239 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node42242 = (inp[10]) ? 4'b0111 : node42243;
														assign node42243 = (inp[2]) ? node42245 : 4'b0111;
															assign node42245 = (inp[13]) ? 4'b0111 : node42246;
																assign node42246 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node42251 = (inp[11]) ? node42263 : node42252;
													assign node42252 = (inp[13]) ? node42258 : node42253;
														assign node42253 = (inp[10]) ? 4'b0110 : node42254;
															assign node42254 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node42258 = (inp[2]) ? node42260 : 4'b0111;
															assign node42260 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node42263 = (inp[13]) ? node42267 : node42264;
														assign node42264 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42267 = (inp[2]) ? node42269 : 4'b0110;
															assign node42269 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node42272 = (inp[10]) ? node42302 : node42273;
												assign node42273 = (inp[12]) ? node42287 : node42274;
													assign node42274 = (inp[1]) ? node42276 : 4'b0111;
														assign node42276 = (inp[11]) ? node42282 : node42277;
															assign node42277 = (inp[2]) ? node42279 : 4'b0111;
																assign node42279 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node42282 = (inp[13]) ? node42284 : 4'b0110;
																assign node42284 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node42287 = (inp[1]) ? node42295 : node42288;
														assign node42288 = (inp[13]) ? node42290 : 4'b0110;
															assign node42290 = (inp[2]) ? 4'b0110 : node42291;
																assign node42291 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42295 = (inp[13]) ? node42299 : node42296;
															assign node42296 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42299 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42302 = (inp[12]) ? node42314 : node42303;
													assign node42303 = (inp[1]) ? 4'b0110 : node42304;
														assign node42304 = (inp[2]) ? node42310 : node42305;
															assign node42305 = (inp[13]) ? 4'b0110 : node42306;
																assign node42306 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42310 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42314 = (inp[13]) ? node42322 : node42315;
														assign node42315 = (inp[1]) ? node42319 : node42316;
															assign node42316 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42319 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42322 = (inp[11]) ? node42326 : node42323;
															assign node42323 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42326 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node42329 = (inp[11]) ? node42349 : node42330;
											assign node42330 = (inp[13]) ? node42340 : node42331;
												assign node42331 = (inp[1]) ? 4'b0110 : node42332;
													assign node42332 = (inp[2]) ? node42336 : node42333;
														assign node42333 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node42336 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node42340 = (inp[1]) ? 4'b0111 : node42341;
													assign node42341 = (inp[2]) ? node42345 : node42342;
														assign node42342 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node42345 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node42349 = (inp[13]) ? node42365 : node42350;
												assign node42350 = (inp[1]) ? 4'b0111 : node42351;
													assign node42351 = (inp[0]) ? node42359 : node42352;
														assign node42352 = (inp[12]) ? node42356 : node42353;
															assign node42353 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node42356 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node42359 = (inp[12]) ? node42361 : 4'b0111;
															assign node42361 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node42365 = (inp[1]) ? 4'b0110 : node42366;
													assign node42366 = (inp[12]) ? node42370 : node42367;
														assign node42367 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node42370 = (inp[2]) ? 4'b0110 : 4'b0111;
							assign node42374 = (inp[7]) ? node42708 : node42375;
								assign node42375 = (inp[2]) ? node42583 : node42376;
									assign node42376 = (inp[0]) ? node42480 : node42377;
										assign node42377 = (inp[1]) ? node42423 : node42378;
											assign node42378 = (inp[4]) ? node42386 : node42379;
												assign node42379 = (inp[11]) ? node42383 : node42380;
													assign node42380 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node42383 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node42386 = (inp[11]) ? node42398 : node42387;
													assign node42387 = (inp[10]) ? node42389 : 4'b0110;
														assign node42389 = (inp[9]) ? node42395 : node42390;
															assign node42390 = (inp[13]) ? 4'b0110 : node42391;
																assign node42391 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node42395 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node42398 = (inp[9]) ? node42408 : node42399;
														assign node42399 = (inp[10]) ? 4'b0110 : node42400;
															assign node42400 = (inp[12]) ? node42404 : node42401;
																assign node42401 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node42404 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node42408 = (inp[10]) ? node42416 : node42409;
															assign node42409 = (inp[13]) ? node42413 : node42410;
																assign node42410 = (inp[12]) ? 4'b0110 : 4'b0111;
																assign node42413 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node42416 = (inp[12]) ? node42420 : node42417;
																assign node42417 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node42420 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node42423 = (inp[10]) ? node42455 : node42424;
												assign node42424 = (inp[12]) ? node42430 : node42425;
													assign node42425 = (inp[9]) ? 4'b0111 : node42426;
														assign node42426 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node42430 = (inp[9]) ? node42440 : node42431;
														assign node42431 = (inp[13]) ? node42433 : 4'b0111;
															assign node42433 = (inp[11]) ? node42437 : node42434;
																assign node42434 = (inp[4]) ? 4'b0111 : 4'b0110;
																assign node42437 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node42440 = (inp[13]) ? node42448 : node42441;
															assign node42441 = (inp[11]) ? node42445 : node42442;
																assign node42442 = (inp[4]) ? 4'b0110 : 4'b0111;
																assign node42445 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node42448 = (inp[4]) ? node42452 : node42449;
																assign node42449 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node42452 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42455 = (inp[4]) ? node42469 : node42456;
													assign node42456 = (inp[12]) ? node42464 : node42457;
														assign node42457 = (inp[11]) ? node42461 : node42458;
															assign node42458 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node42461 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node42464 = (inp[13]) ? 4'b0110 : node42465;
															assign node42465 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42469 = (inp[12]) ? node42475 : node42470;
														assign node42470 = (inp[13]) ? 4'b0110 : node42471;
															assign node42471 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42475 = (inp[11]) ? 4'b0111 : node42476;
															assign node42476 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node42480 = (inp[10]) ? node42536 : node42481;
											assign node42481 = (inp[12]) ? node42503 : node42482;
												assign node42482 = (inp[4]) ? node42490 : node42483;
													assign node42483 = (inp[13]) ? node42487 : node42484;
														assign node42484 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42487 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42490 = (inp[11]) ? node42496 : node42491;
														assign node42491 = (inp[1]) ? node42493 : 4'b0111;
															assign node42493 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node42496 = (inp[9]) ? node42498 : 4'b0111;
															assign node42498 = (inp[1]) ? node42500 : 4'b0110;
																assign node42500 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node42503 = (inp[13]) ? node42519 : node42504;
													assign node42504 = (inp[11]) ? node42512 : node42505;
														assign node42505 = (inp[1]) ? node42509 : node42506;
															assign node42506 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node42509 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node42512 = (inp[4]) ? node42516 : node42513;
															assign node42513 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node42516 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node42519 = (inp[1]) ? node42527 : node42520;
														assign node42520 = (inp[4]) ? node42524 : node42521;
															assign node42521 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42524 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42527 = (inp[9]) ? node42531 : node42528;
															assign node42528 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node42531 = (inp[4]) ? 4'b0110 : node42532;
																assign node42532 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node42536 = (inp[13]) ? node42558 : node42537;
												assign node42537 = (inp[1]) ? node42549 : node42538;
													assign node42538 = (inp[11]) ? node42544 : node42539;
														assign node42539 = (inp[4]) ? node42541 : 4'b0110;
															assign node42541 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node42544 = (inp[4]) ? node42546 : 4'b0111;
															assign node42546 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node42549 = (inp[11]) ? node42551 : 4'b0111;
														assign node42551 = (inp[12]) ? node42555 : node42552;
															assign node42552 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node42555 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node42558 = (inp[11]) ? node42572 : node42559;
													assign node42559 = (inp[4]) ? node42561 : 4'b0111;
														assign node42561 = (inp[9]) ? node42567 : node42562;
															assign node42562 = (inp[1]) ? 4'b0111 : node42563;
																assign node42563 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node42567 = (inp[12]) ? 4'b0111 : node42568;
																assign node42568 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node42572 = (inp[12]) ? node42578 : node42573;
														assign node42573 = (inp[4]) ? node42575 : 4'b0110;
															assign node42575 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42578 = (inp[9]) ? 4'b0111 : node42579;
															assign node42579 = (inp[4]) ? 4'b0110 : 4'b0111;
									assign node42583 = (inp[9]) ? node42617 : node42584;
										assign node42584 = (inp[11]) ? node42598 : node42585;
											assign node42585 = (inp[13]) ? node42593 : node42586;
												assign node42586 = (inp[4]) ? 4'b0110 : node42587;
													assign node42587 = (inp[12]) ? 4'b0110 : node42588;
														assign node42588 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node42593 = (inp[4]) ? 4'b0111 : node42594;
													assign node42594 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node42598 = (inp[13]) ? node42608 : node42599;
												assign node42599 = (inp[1]) ? node42601 : 4'b0111;
													assign node42601 = (inp[10]) ? 4'b0111 : node42602;
														assign node42602 = (inp[4]) ? 4'b0111 : node42603;
															assign node42603 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node42608 = (inp[4]) ? 4'b0110 : node42609;
													assign node42609 = (inp[0]) ? node42611 : 4'b0110;
														assign node42611 = (inp[12]) ? 4'b0110 : node42612;
															assign node42612 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node42617 = (inp[4]) ? node42659 : node42618;
											assign node42618 = (inp[1]) ? node42626 : node42619;
												assign node42619 = (inp[13]) ? node42623 : node42620;
													assign node42620 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node42623 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42626 = (inp[10]) ? node42638 : node42627;
													assign node42627 = (inp[0]) ? node42629 : 4'b0110;
														assign node42629 = (inp[12]) ? node42631 : 4'b0111;
															assign node42631 = (inp[13]) ? node42635 : node42632;
																assign node42632 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node42635 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42638 = (inp[0]) ? node42652 : node42639;
														assign node42639 = (inp[12]) ? node42647 : node42640;
															assign node42640 = (inp[13]) ? node42644 : node42641;
																assign node42641 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node42644 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42647 = (inp[13]) ? node42649 : 4'b0110;
																assign node42649 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42652 = (inp[13]) ? 4'b0110 : node42653;
															assign node42653 = (inp[11]) ? node42655 : 4'b0110;
																assign node42655 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node42659 = (inp[10]) ? node42687 : node42660;
												assign node42660 = (inp[1]) ? node42680 : node42661;
													assign node42661 = (inp[12]) ? node42675 : node42662;
														assign node42662 = (inp[0]) ? node42668 : node42663;
															assign node42663 = (inp[11]) ? node42665 : 4'b0110;
																assign node42665 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node42668 = (inp[11]) ? node42672 : node42669;
																assign node42669 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node42672 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node42675 = (inp[13]) ? node42677 : 4'b0110;
															assign node42677 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42680 = (inp[13]) ? node42684 : node42681;
														assign node42681 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42684 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node42687 = (inp[0]) ? node42701 : node42688;
													assign node42688 = (inp[12]) ? node42696 : node42689;
														assign node42689 = (inp[13]) ? node42693 : node42690;
															assign node42690 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node42693 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node42696 = (inp[13]) ? node42698 : 4'b0111;
															assign node42698 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node42701 = (inp[13]) ? node42705 : node42702;
														assign node42702 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42705 = (inp[11]) ? 4'b0110 : 4'b0111;
								assign node42708 = (inp[13]) ? node42776 : node42709;
									assign node42709 = (inp[11]) ? node42753 : node42710;
										assign node42710 = (inp[2]) ? node42746 : node42711;
											assign node42711 = (inp[12]) ? node42717 : node42712;
												assign node42712 = (inp[1]) ? 4'b0010 : node42713;
													assign node42713 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node42717 = (inp[0]) ? node42733 : node42718;
													assign node42718 = (inp[10]) ? 4'b0011 : node42719;
														assign node42719 = (inp[9]) ? node42725 : node42720;
															assign node42720 = (inp[4]) ? 4'b0011 : node42721;
																assign node42721 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node42725 = (inp[1]) ? node42729 : node42726;
																assign node42726 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node42729 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node42733 = (inp[10]) ? node42741 : node42734;
														assign node42734 = (inp[1]) ? node42738 : node42735;
															assign node42735 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node42738 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node42741 = (inp[4]) ? node42743 : 4'b0010;
															assign node42743 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node42746 = (inp[4]) ? node42748 : 4'b0010;
												assign node42748 = (inp[12]) ? 4'b0010 : node42749;
													assign node42749 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node42753 = (inp[1]) ? node42767 : node42754;
											assign node42754 = (inp[4]) ? node42760 : node42755;
												assign node42755 = (inp[12]) ? 4'b0011 : node42756;
													assign node42756 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node42760 = (inp[2]) ? node42764 : node42761;
													assign node42761 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node42764 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node42767 = (inp[4]) ? 4'b0011 : node42768;
												assign node42768 = (inp[9]) ? 4'b0011 : node42769;
													assign node42769 = (inp[12]) ? node42771 : 4'b0011;
														assign node42771 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node42776 = (inp[11]) ? node42806 : node42777;
										assign node42777 = (inp[1]) ? node42799 : node42778;
											assign node42778 = (inp[12]) ? node42794 : node42779;
												assign node42779 = (inp[9]) ? node42787 : node42780;
													assign node42780 = (inp[2]) ? node42784 : node42781;
														assign node42781 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node42784 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node42787 = (inp[4]) ? node42791 : node42788;
														assign node42788 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node42791 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node42794 = (inp[4]) ? node42796 : 4'b0011;
													assign node42796 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node42799 = (inp[12]) ? node42801 : 4'b0011;
												assign node42801 = (inp[4]) ? 4'b0011 : node42802;
													assign node42802 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node42806 = (inp[1]) ? node42842 : node42807;
											assign node42807 = (inp[4]) ? node42813 : node42808;
												assign node42808 = (inp[2]) ? 4'b0010 : node42809;
													assign node42809 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node42813 = (inp[9]) ? node42835 : node42814;
													assign node42814 = (inp[0]) ? node42822 : node42815;
														assign node42815 = (inp[2]) ? node42819 : node42816;
															assign node42816 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node42819 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node42822 = (inp[10]) ? node42830 : node42823;
															assign node42823 = (inp[12]) ? node42827 : node42824;
																assign node42824 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node42827 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node42830 = (inp[2]) ? 4'b0011 : node42831;
																assign node42831 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node42835 = (inp[2]) ? node42839 : node42836;
														assign node42836 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node42839 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node42842 = (inp[2]) ? 4'b0010 : node42843;
												assign node42843 = (inp[12]) ? node42845 : 4'b0010;
													assign node42845 = (inp[4]) ? 4'b0010 : 4'b0011;
						assign node42849 = (inp[7]) ? node43209 : node42850;
							assign node42850 = (inp[4]) ? node43040 : node42851;
								assign node42851 = (inp[12]) ? node43017 : node42852;
									assign node42852 = (inp[1]) ? node42938 : node42853;
										assign node42853 = (inp[9]) ? node42901 : node42854;
											assign node42854 = (inp[10]) ? node42888 : node42855;
												assign node42855 = (inp[11]) ? node42869 : node42856;
													assign node42856 = (inp[5]) ? node42862 : node42857;
														assign node42857 = (inp[0]) ? node42859 : 4'b0001;
															assign node42859 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node42862 = (inp[13]) ? node42866 : node42863;
															assign node42863 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node42866 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node42869 = (inp[5]) ? node42881 : node42870;
														assign node42870 = (inp[0]) ? node42876 : node42871;
															assign node42871 = (inp[13]) ? 4'b0000 : node42872;
																assign node42872 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node42876 = (inp[13]) ? node42878 : 4'b0000;
																assign node42878 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node42881 = (inp[2]) ? node42885 : node42882;
															assign node42882 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node42885 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node42888 = (inp[5]) ? node42896 : node42889;
													assign node42889 = (inp[13]) ? node42893 : node42890;
														assign node42890 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node42893 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node42896 = (inp[13]) ? node42898 : 4'b0000;
														assign node42898 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node42901 = (inp[11]) ? node42931 : node42902;
												assign node42902 = (inp[10]) ? node42916 : node42903;
													assign node42903 = (inp[5]) ? node42911 : node42904;
														assign node42904 = (inp[0]) ? 4'b0000 : node42905;
															assign node42905 = (inp[13]) ? 4'b0001 : node42906;
																assign node42906 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node42911 = (inp[0]) ? node42913 : 4'b0000;
															assign node42913 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node42916 = (inp[0]) ? node42924 : node42917;
														assign node42917 = (inp[13]) ? node42921 : node42918;
															assign node42918 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node42921 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node42924 = (inp[13]) ? node42928 : node42925;
															assign node42925 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node42928 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node42931 = (inp[13]) ? node42935 : node42932;
													assign node42932 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node42935 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node42938 = (inp[5]) ? node42966 : node42939;
											assign node42939 = (inp[9]) ? node42959 : node42940;
												assign node42940 = (inp[11]) ? node42952 : node42941;
													assign node42941 = (inp[10]) ? node42947 : node42942;
														assign node42942 = (inp[13]) ? 4'b0000 : node42943;
															assign node42943 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node42947 = (inp[2]) ? 4'b0001 : node42948;
															assign node42948 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node42952 = (inp[13]) ? node42956 : node42953;
														assign node42953 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node42956 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node42959 = (inp[13]) ? node42963 : node42960;
													assign node42960 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node42963 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node42966 = (inp[9]) ? node42974 : node42967;
												assign node42967 = (inp[13]) ? node42971 : node42968;
													assign node42968 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node42971 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node42974 = (inp[10]) ? node43002 : node42975;
													assign node42975 = (inp[11]) ? node42989 : node42976;
														assign node42976 = (inp[0]) ? node42984 : node42977;
															assign node42977 = (inp[13]) ? node42981 : node42978;
																assign node42978 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node42981 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node42984 = (inp[13]) ? 4'b0000 : node42985;
																assign node42985 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node42989 = (inp[0]) ? node42997 : node42990;
															assign node42990 = (inp[2]) ? node42994 : node42991;
																assign node42991 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node42994 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node42997 = (inp[13]) ? node42999 : 4'b0001;
																assign node42999 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node43002 = (inp[11]) ? node43010 : node43003;
														assign node43003 = (inp[0]) ? 4'b0001 : node43004;
															assign node43004 = (inp[13]) ? 4'b0001 : node43005;
																assign node43005 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node43010 = (inp[13]) ? node43014 : node43011;
															assign node43011 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node43014 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node43017 = (inp[2]) ? node43029 : node43018;
										assign node43018 = (inp[13]) ? node43024 : node43019;
											assign node43019 = (inp[5]) ? 4'b0100 : node43020;
												assign node43020 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node43024 = (inp[5]) ? 4'b0101 : node43025;
												assign node43025 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node43029 = (inp[13]) ? node43035 : node43030;
											assign node43030 = (inp[1]) ? node43032 : 4'b0101;
												assign node43032 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node43035 = (inp[5]) ? 4'b0100 : node43036;
												assign node43036 = (inp[1]) ? 4'b0101 : 4'b0100;
								assign node43040 = (inp[2]) ? node43106 : node43041;
									assign node43041 = (inp[10]) ? node43049 : node43042;
										assign node43042 = (inp[5]) ? node43046 : node43043;
											assign node43043 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node43046 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node43049 = (inp[11]) ? node43081 : node43050;
											assign node43050 = (inp[0]) ? node43066 : node43051;
												assign node43051 = (inp[1]) ? node43059 : node43052;
													assign node43052 = (inp[13]) ? node43056 : node43053;
														assign node43053 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43056 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node43059 = (inp[5]) ? node43063 : node43060;
														assign node43060 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43063 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node43066 = (inp[12]) ? node43074 : node43067;
													assign node43067 = (inp[13]) ? node43071 : node43068;
														assign node43068 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43071 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node43074 = (inp[5]) ? node43078 : node43075;
														assign node43075 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43078 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node43081 = (inp[9]) ? node43089 : node43082;
												assign node43082 = (inp[5]) ? node43086 : node43083;
													assign node43083 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node43086 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node43089 = (inp[1]) ? node43097 : node43090;
													assign node43090 = (inp[5]) ? node43094 : node43091;
														assign node43091 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43094 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node43097 = (inp[12]) ? node43099 : 4'b0100;
														assign node43099 = (inp[5]) ? node43103 : node43100;
															assign node43100 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node43103 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node43106 = (inp[10]) ? node43114 : node43107;
										assign node43107 = (inp[13]) ? node43111 : node43108;
											assign node43108 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node43111 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node43114 = (inp[9]) ? node43170 : node43115;
											assign node43115 = (inp[0]) ? node43143 : node43116;
												assign node43116 = (inp[12]) ? node43122 : node43117;
													assign node43117 = (inp[13]) ? 4'b0101 : node43118;
														assign node43118 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node43122 = (inp[11]) ? node43134 : node43123;
														assign node43123 = (inp[1]) ? node43129 : node43124;
															assign node43124 = (inp[5]) ? node43126 : 4'b0101;
																assign node43126 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node43129 = (inp[13]) ? 4'b0101 : node43130;
																assign node43130 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43134 = (inp[1]) ? 4'b0100 : node43135;
															assign node43135 = (inp[13]) ? node43139 : node43136;
																assign node43136 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node43139 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node43143 = (inp[12]) ? node43159 : node43144;
													assign node43144 = (inp[1]) ? node43152 : node43145;
														assign node43145 = (inp[13]) ? node43149 : node43146;
															assign node43146 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node43149 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node43152 = (inp[5]) ? node43156 : node43153;
															assign node43153 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node43156 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node43159 = (inp[1]) ? node43165 : node43160;
														assign node43160 = (inp[5]) ? 4'b0101 : node43161;
															assign node43161 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43165 = (inp[13]) ? node43167 : 4'b0101;
															assign node43167 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node43170 = (inp[0]) ? node43194 : node43171;
												assign node43171 = (inp[1]) ? node43179 : node43172;
													assign node43172 = (inp[13]) ? node43176 : node43173;
														assign node43173 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43176 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node43179 = (inp[11]) ? node43187 : node43180;
														assign node43180 = (inp[5]) ? node43184 : node43181;
															assign node43181 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node43184 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node43187 = (inp[5]) ? node43191 : node43188;
															assign node43188 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node43191 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node43194 = (inp[12]) ? node43202 : node43195;
													assign node43195 = (inp[5]) ? node43199 : node43196;
														assign node43196 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43199 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node43202 = (inp[13]) ? node43206 : node43203;
														assign node43203 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43206 = (inp[5]) ? 4'b0100 : 4'b0101;
							assign node43209 = (inp[12]) ? node43469 : node43210;
								assign node43210 = (inp[4]) ? node43392 : node43211;
									assign node43211 = (inp[9]) ? node43331 : node43212;
										assign node43212 = (inp[1]) ? node43266 : node43213;
											assign node43213 = (inp[0]) ? node43243 : node43214;
												assign node43214 = (inp[10]) ? node43230 : node43215;
													assign node43215 = (inp[2]) ? node43223 : node43216;
														assign node43216 = (inp[13]) ? node43220 : node43217;
															assign node43217 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node43220 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node43223 = (inp[5]) ? node43227 : node43224;
															assign node43224 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node43227 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node43230 = (inp[2]) ? node43236 : node43231;
														assign node43231 = (inp[13]) ? 4'b0101 : node43232;
															assign node43232 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43236 = (inp[13]) ? node43240 : node43237;
															assign node43237 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node43240 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node43243 = (inp[10]) ? node43257 : node43244;
													assign node43244 = (inp[11]) ? node43254 : node43245;
														assign node43245 = (inp[5]) ? node43247 : 4'b0101;
															assign node43247 = (inp[2]) ? node43251 : node43248;
																assign node43248 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node43251 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43254 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node43257 = (inp[2]) ? 4'b0100 : node43258;
														assign node43258 = (inp[5]) ? node43262 : node43259;
															assign node43259 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node43262 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node43266 = (inp[0]) ? node43296 : node43267;
												assign node43267 = (inp[10]) ? node43281 : node43268;
													assign node43268 = (inp[5]) ? node43276 : node43269;
														assign node43269 = (inp[13]) ? node43273 : node43270;
															assign node43270 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node43273 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43276 = (inp[2]) ? 4'b0101 : node43277;
															assign node43277 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node43281 = (inp[11]) ? node43289 : node43282;
														assign node43282 = (inp[13]) ? node43286 : node43283;
															assign node43283 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node43286 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43289 = (inp[13]) ? node43293 : node43290;
															assign node43290 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node43293 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node43296 = (inp[10]) ? node43316 : node43297;
													assign node43297 = (inp[5]) ? node43303 : node43298;
														assign node43298 = (inp[13]) ? node43300 : 4'b0101;
															assign node43300 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43303 = (inp[11]) ? node43311 : node43304;
															assign node43304 = (inp[2]) ? node43308 : node43305;
																assign node43305 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node43308 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node43311 = (inp[13]) ? 4'b0100 : node43312;
																assign node43312 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node43316 = (inp[11]) ? node43324 : node43317;
														assign node43317 = (inp[5]) ? node43319 : 4'b0101;
															assign node43319 = (inp[13]) ? node43321 : 4'b0101;
																assign node43321 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43324 = (inp[5]) ? 4'b0101 : node43325;
															assign node43325 = (inp[13]) ? 4'b0101 : node43326;
																assign node43326 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node43331 = (inp[1]) ? node43385 : node43332;
											assign node43332 = (inp[2]) ? node43358 : node43333;
												assign node43333 = (inp[11]) ? node43347 : node43334;
													assign node43334 = (inp[10]) ? node43340 : node43335;
														assign node43335 = (inp[5]) ? 4'b0101 : node43336;
															assign node43336 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node43340 = (inp[13]) ? node43344 : node43341;
															assign node43341 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node43344 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node43347 = (inp[0]) ? 4'b0101 : node43348;
														assign node43348 = (inp[10]) ? node43354 : node43349;
															assign node43349 = (inp[13]) ? 4'b0101 : node43350;
																assign node43350 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node43354 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node43358 = (inp[0]) ? node43366 : node43359;
													assign node43359 = (inp[13]) ? node43363 : node43360;
														assign node43360 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node43363 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node43366 = (inp[10]) ? node43372 : node43367;
														assign node43367 = (inp[13]) ? node43369 : 4'b0101;
															assign node43369 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node43372 = (inp[11]) ? node43380 : node43373;
															assign node43373 = (inp[13]) ? node43377 : node43374;
																assign node43374 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node43377 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node43380 = (inp[13]) ? 4'b0100 : node43381;
																assign node43381 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node43385 = (inp[13]) ? node43389 : node43386;
												assign node43386 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node43389 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node43392 = (inp[10]) ? node43408 : node43393;
										assign node43393 = (inp[0]) ? node43401 : node43394;
											assign node43394 = (inp[13]) ? node43398 : node43395;
												assign node43395 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node43398 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node43401 = (inp[1]) ? node43405 : node43402;
												assign node43402 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node43405 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node43408 = (inp[0]) ? node43454 : node43409;
											assign node43409 = (inp[5]) ? node43439 : node43410;
												assign node43410 = (inp[11]) ? node43432 : node43411;
													assign node43411 = (inp[9]) ? node43425 : node43412;
														assign node43412 = (inp[2]) ? node43420 : node43413;
															assign node43413 = (inp[13]) ? node43417 : node43414;
																assign node43414 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node43417 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node43420 = (inp[13]) ? 4'b0001 : node43421;
																assign node43421 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node43425 = (inp[13]) ? node43429 : node43426;
															assign node43426 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node43429 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node43432 = (inp[1]) ? node43436 : node43433;
														assign node43433 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node43436 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node43439 = (inp[11]) ? node43447 : node43440;
													assign node43440 = (inp[1]) ? node43444 : node43441;
														assign node43441 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node43444 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node43447 = (inp[1]) ? node43451 : node43448;
														assign node43448 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node43451 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node43454 = (inp[5]) ? node43462 : node43455;
												assign node43455 = (inp[13]) ? node43459 : node43456;
													assign node43456 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node43459 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node43462 = (inp[1]) ? node43466 : node43463;
													assign node43463 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node43466 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node43469 = (inp[13]) ? node43483 : node43470;
									assign node43470 = (inp[4]) ? 4'b0001 : node43471;
										assign node43471 = (inp[2]) ? node43477 : node43472;
											assign node43472 = (inp[5]) ? 4'b0000 : node43473;
												assign node43473 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node43477 = (inp[5]) ? 4'b0001 : node43478;
												assign node43478 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node43483 = (inp[4]) ? 4'b0000 : node43484;
										assign node43484 = (inp[2]) ? node43490 : node43485;
											assign node43485 = (inp[1]) ? 4'b0001 : node43486;
												assign node43486 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node43490 = (inp[5]) ? 4'b0000 : node43491;
												assign node43491 = (inp[1]) ? 4'b0000 : 4'b0001;
					assign node43496 = (inp[5]) ? node43836 : node43497;
						assign node43497 = (inp[14]) ? node43749 : node43498;
							assign node43498 = (inp[4]) ? node43664 : node43499;
								assign node43499 = (inp[12]) ? node43591 : node43500;
									assign node43500 = (inp[0]) ? node43568 : node43501;
										assign node43501 = (inp[9]) ? node43529 : node43502;
											assign node43502 = (inp[7]) ? node43510 : node43503;
												assign node43503 = (inp[11]) ? node43507 : node43504;
													assign node43504 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node43507 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node43510 = (inp[1]) ? node43518 : node43511;
													assign node43511 = (inp[11]) ? node43515 : node43512;
														assign node43512 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node43515 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node43518 = (inp[10]) ? node43524 : node43519;
														assign node43519 = (inp[2]) ? 4'b0000 : node43520;
															assign node43520 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node43524 = (inp[2]) ? node43526 : 4'b0000;
															assign node43526 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node43529 = (inp[7]) ? node43537 : node43530;
												assign node43530 = (inp[11]) ? node43534 : node43531;
													assign node43531 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node43534 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node43537 = (inp[11]) ? node43555 : node43538;
													assign node43538 = (inp[10]) ? node43548 : node43539;
														assign node43539 = (inp[13]) ? node43541 : 4'b0000;
															assign node43541 = (inp[1]) ? node43545 : node43542;
																assign node43542 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node43545 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node43548 = (inp[1]) ? node43552 : node43549;
															assign node43549 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node43552 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node43555 = (inp[13]) ? 4'b0001 : node43556;
														assign node43556 = (inp[10]) ? node43562 : node43557;
															assign node43557 = (inp[1]) ? 4'b0001 : node43558;
																assign node43558 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node43562 = (inp[2]) ? 4'b0001 : node43563;
																assign node43563 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node43568 = (inp[1]) ? node43580 : node43569;
											assign node43569 = (inp[11]) ? node43575 : node43570;
												assign node43570 = (inp[7]) ? node43572 : 4'b0000;
													assign node43572 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node43575 = (inp[7]) ? node43577 : 4'b0001;
													assign node43577 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node43580 = (inp[11]) ? node43586 : node43581;
												assign node43581 = (inp[2]) ? node43583 : 4'b0001;
													assign node43583 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node43586 = (inp[2]) ? node43588 : 4'b0000;
													assign node43588 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node43591 = (inp[0]) ? node43657 : node43592;
										assign node43592 = (inp[13]) ? node43650 : node43593;
											assign node43593 = (inp[1]) ? node43623 : node43594;
												assign node43594 = (inp[10]) ? node43616 : node43595;
													assign node43595 = (inp[2]) ? node43609 : node43596;
														assign node43596 = (inp[9]) ? node43604 : node43597;
															assign node43597 = (inp[7]) ? node43601 : node43598;
																assign node43598 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node43601 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node43604 = (inp[7]) ? 4'b0100 : node43605;
																assign node43605 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node43609 = (inp[9]) ? node43611 : 4'b0100;
															assign node43611 = (inp[7]) ? node43613 : 4'b0100;
																assign node43613 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node43616 = (inp[11]) ? node43620 : node43617;
														assign node43617 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node43620 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node43623 = (inp[2]) ? node43643 : node43624;
													assign node43624 = (inp[9]) ? node43632 : node43625;
														assign node43625 = (inp[7]) ? node43629 : node43626;
															assign node43626 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node43629 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node43632 = (inp[10]) ? node43638 : node43633;
															assign node43633 = (inp[7]) ? 4'b0100 : node43634;
																assign node43634 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node43638 = (inp[11]) ? 4'b0100 : node43639;
																assign node43639 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node43643 = (inp[11]) ? node43647 : node43644;
														assign node43644 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node43647 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node43650 = (inp[11]) ? node43654 : node43651;
												assign node43651 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node43654 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node43657 = (inp[11]) ? node43661 : node43658;
											assign node43658 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node43661 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node43664 = (inp[7]) ? node43738 : node43665;
									assign node43665 = (inp[11]) ? node43675 : node43666;
										assign node43666 = (inp[12]) ? 4'b0100 : node43667;
											assign node43667 = (inp[2]) ? node43671 : node43668;
												assign node43668 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node43671 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node43675 = (inp[12]) ? 4'b0101 : node43676;
											assign node43676 = (inp[9]) ? node43700 : node43677;
												assign node43677 = (inp[0]) ? node43693 : node43678;
													assign node43678 = (inp[10]) ? node43686 : node43679;
														assign node43679 = (inp[1]) ? node43683 : node43680;
															assign node43680 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node43683 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node43686 = (inp[1]) ? node43690 : node43687;
															assign node43687 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node43690 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node43693 = (inp[2]) ? node43697 : node43694;
														assign node43694 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node43697 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node43700 = (inp[10]) ? node43720 : node43701;
													assign node43701 = (inp[0]) ? node43713 : node43702;
														assign node43702 = (inp[13]) ? node43708 : node43703;
															assign node43703 = (inp[1]) ? node43705 : 4'b0100;
																assign node43705 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node43708 = (inp[1]) ? node43710 : 4'b0101;
																assign node43710 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node43713 = (inp[13]) ? 4'b0100 : node43714;
															assign node43714 = (inp[2]) ? node43716 : 4'b0100;
																assign node43716 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node43720 = (inp[0]) ? node43728 : node43721;
														assign node43721 = (inp[2]) ? node43725 : node43722;
															assign node43722 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node43725 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node43728 = (inp[13]) ? node43732 : node43729;
															assign node43729 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node43732 = (inp[2]) ? 4'b0101 : node43733;
																assign node43733 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node43738 = (inp[11]) ? node43744 : node43739;
										assign node43739 = (inp[12]) ? 4'b0101 : node43740;
											assign node43740 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node43744 = (inp[12]) ? 4'b0100 : node43745;
											assign node43745 = (inp[1]) ? 4'b0100 : 4'b0101;
							assign node43749 = (inp[12]) ? node43825 : node43750;
								assign node43750 = (inp[4]) ? node43758 : node43751;
									assign node43751 = (inp[1]) ? node43755 : node43752;
										assign node43752 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node43755 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node43758 = (inp[0]) ? node43766 : node43759;
										assign node43759 = (inp[1]) ? node43763 : node43760;
											assign node43760 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node43763 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node43766 = (inp[2]) ? node43774 : node43767;
											assign node43767 = (inp[7]) ? node43771 : node43768;
												assign node43768 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node43771 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node43774 = (inp[10]) ? node43796 : node43775;
												assign node43775 = (inp[13]) ? node43783 : node43776;
													assign node43776 = (inp[7]) ? node43780 : node43777;
														assign node43777 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node43780 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node43783 = (inp[9]) ? node43789 : node43784;
														assign node43784 = (inp[7]) ? node43786 : 4'b0001;
															assign node43786 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node43789 = (inp[11]) ? node43791 : 4'b0000;
															assign node43791 = (inp[7]) ? node43793 : 4'b0001;
																assign node43793 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node43796 = (inp[9]) ? node43808 : node43797;
													assign node43797 = (inp[11]) ? node43803 : node43798;
														assign node43798 = (inp[7]) ? node43800 : 4'b0001;
															assign node43800 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node43803 = (inp[7]) ? 4'b0001 : node43804;
															assign node43804 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node43808 = (inp[11]) ? node43814 : node43809;
														assign node43809 = (inp[7]) ? 4'b0001 : node43810;
															assign node43810 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node43814 = (inp[13]) ? node43820 : node43815;
															assign node43815 = (inp[7]) ? 4'b0000 : node43816;
																assign node43816 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node43820 = (inp[7]) ? node43822 : 4'b0001;
																assign node43822 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node43825 = (inp[7]) ? node43831 : node43826;
									assign node43826 = (inp[2]) ? 4'b0001 : node43827;
										assign node43827 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node43831 = (inp[4]) ? 4'b0000 : node43832;
										assign node43832 = (inp[2]) ? 4'b0000 : 4'b0001;
						assign node43836 = (inp[4]) ? node44062 : node43837;
							assign node43837 = (inp[12]) ? node44051 : node43838;
								assign node43838 = (inp[0]) ? node43998 : node43839;
									assign node43839 = (inp[10]) ? node43883 : node43840;
										assign node43840 = (inp[2]) ? node43872 : node43841;
											assign node43841 = (inp[1]) ? node43851 : node43842;
												assign node43842 = (inp[14]) ? 4'b0100 : node43843;
													assign node43843 = (inp[11]) ? node43847 : node43844;
														assign node43844 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node43847 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node43851 = (inp[14]) ? 4'b0101 : node43852;
													assign node43852 = (inp[9]) ? node43862 : node43853;
														assign node43853 = (inp[13]) ? node43855 : 4'b0100;
															assign node43855 = (inp[11]) ? node43859 : node43856;
																assign node43856 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node43859 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node43862 = (inp[13]) ? node43864 : 4'b0101;
															assign node43864 = (inp[7]) ? node43868 : node43865;
																assign node43865 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node43868 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node43872 = (inp[1]) ? node43878 : node43873;
												assign node43873 = (inp[11]) ? 4'b0101 : node43874;
													assign node43874 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node43878 = (inp[14]) ? 4'b0100 : node43879;
													assign node43879 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node43883 = (inp[13]) ? node43935 : node43884;
											assign node43884 = (inp[14]) ? node43920 : node43885;
												assign node43885 = (inp[9]) ? node43905 : node43886;
													assign node43886 = (inp[7]) ? node43896 : node43887;
														assign node43887 = (inp[2]) ? node43889 : 4'b0101;
															assign node43889 = (inp[1]) ? node43893 : node43890;
																assign node43890 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node43893 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node43896 = (inp[2]) ? node43898 : 4'b0100;
															assign node43898 = (inp[11]) ? node43902 : node43899;
																assign node43899 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node43902 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node43905 = (inp[7]) ? node43911 : node43906;
														assign node43906 = (inp[1]) ? node43908 : 4'b0100;
															assign node43908 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node43911 = (inp[2]) ? node43913 : 4'b0100;
															assign node43913 = (inp[11]) ? node43917 : node43914;
																assign node43914 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node43917 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node43920 = (inp[9]) ? node43928 : node43921;
													assign node43921 = (inp[2]) ? node43925 : node43922;
														assign node43922 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node43925 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node43928 = (inp[2]) ? node43932 : node43929;
														assign node43929 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node43932 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node43935 = (inp[9]) ? node43969 : node43936;
												assign node43936 = (inp[14]) ? node43952 : node43937;
													assign node43937 = (inp[1]) ? node43943 : node43938;
														assign node43938 = (inp[11]) ? 4'b0101 : node43939;
															assign node43939 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43943 = (inp[11]) ? node43949 : node43944;
															assign node43944 = (inp[2]) ? 4'b0101 : node43945;
																assign node43945 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node43949 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node43952 = (inp[11]) ? node43962 : node43953;
														assign node43953 = (inp[7]) ? node43955 : 4'b0101;
															assign node43955 = (inp[1]) ? node43959 : node43956;
																assign node43956 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node43959 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node43962 = (inp[7]) ? 4'b0101 : node43963;
															assign node43963 = (inp[1]) ? node43965 : 4'b0100;
																assign node43965 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node43969 = (inp[11]) ? node43987 : node43970;
													assign node43970 = (inp[1]) ? node43978 : node43971;
														assign node43971 = (inp[7]) ? node43973 : 4'b0100;
															assign node43973 = (inp[2]) ? 4'b0101 : node43974;
																assign node43974 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node43978 = (inp[7]) ? node43984 : node43979;
															assign node43979 = (inp[2]) ? node43981 : 4'b0101;
																assign node43981 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node43984 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node43987 = (inp[1]) ? node43993 : node43988;
														assign node43988 = (inp[2]) ? 4'b0101 : node43989;
															assign node43989 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node43993 = (inp[2]) ? 4'b0100 : node43994;
															assign node43994 = (inp[14]) ? 4'b0101 : 4'b0100;
									assign node43998 = (inp[7]) ? node44022 : node43999;
										assign node43999 = (inp[11]) ? node44011 : node44000;
											assign node44000 = (inp[1]) ? node44006 : node44001;
												assign node44001 = (inp[14]) ? node44003 : 4'b0100;
													assign node44003 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node44006 = (inp[14]) ? node44008 : 4'b0101;
													assign node44008 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node44011 = (inp[1]) ? node44017 : node44012;
												assign node44012 = (inp[14]) ? node44014 : 4'b0101;
													assign node44014 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node44017 = (inp[2]) ? 4'b0100 : node44018;
													assign node44018 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node44022 = (inp[11]) ? node44036 : node44023;
											assign node44023 = (inp[1]) ? node44029 : node44024;
												assign node44024 = (inp[2]) ? node44026 : 4'b0100;
													assign node44026 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node44029 = (inp[2]) ? node44033 : node44030;
													assign node44030 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node44033 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node44036 = (inp[10]) ? node44044 : node44037;
												assign node44037 = (inp[2]) ? node44041 : node44038;
													assign node44038 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node44041 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node44044 = (inp[1]) ? node44048 : node44045;
													assign node44045 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44048 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node44051 = (inp[2]) ? node44057 : node44052;
									assign node44052 = (inp[14]) ? 4'b0001 : node44053;
										assign node44053 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node44057 = (inp[14]) ? 4'b0000 : node44058;
										assign node44058 = (inp[11]) ? 4'b0000 : 4'b0001;
							assign node44062 = (inp[11]) ? node44082 : node44063;
								assign node44063 = (inp[14]) ? node44077 : node44064;
									assign node44064 = (inp[12]) ? 4'b0001 : node44065;
										assign node44065 = (inp[1]) ? node44071 : node44066;
											assign node44066 = (inp[7]) ? 4'b0000 : node44067;
												assign node44067 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node44071 = (inp[2]) ? 4'b0001 : node44072;
												assign node44072 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node44077 = (inp[1]) ? 4'b0000 : node44078;
										assign node44078 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node44082 = (inp[12]) ? 4'b0000 : node44083;
									assign node44083 = (inp[1]) ? node44091 : node44084;
										assign node44084 = (inp[2]) ? 4'b0001 : node44085;
											assign node44085 = (inp[7]) ? 4'b0001 : node44086;
												assign node44086 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node44091 = (inp[2]) ? 4'b0000 : node44092;
											assign node44092 = (inp[14]) ? 4'b0000 : node44093;
												assign node44093 = (inp[7]) ? 4'b0000 : 4'b0001;

endmodule