module dtc_split125_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node15;
	wire [4-1:0] node17;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node23;
	wire [4-1:0] node27;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node43;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node69;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node81;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node89;
	wire [4-1:0] node92;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node101;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node116;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node122;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node160;
	wire [4-1:0] node163;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node182;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node215;
	wire [4-1:0] node218;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node231;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node239;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node251;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node267;
	wire [4-1:0] node270;
	wire [4-1:0] node271;
	wire [4-1:0] node274;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node280;
	wire [4-1:0] node284;
	wire [4-1:0] node285;
	wire [4-1:0] node287;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node317;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node331;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node356;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node396;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node417;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node423;
	wire [4-1:0] node427;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node458;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node461;
	wire [4-1:0] node462;
	wire [4-1:0] node467;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node484;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node503;
	wire [4-1:0] node505;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node512;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node532;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node543;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node560;
	wire [4-1:0] node563;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node576;
	wire [4-1:0] node578;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node594;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node604;
	wire [4-1:0] node607;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node619;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node630;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node637;
	wire [4-1:0] node640;
	wire [4-1:0] node642;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node667;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node676;
	wire [4-1:0] node679;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node692;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node705;
	wire [4-1:0] node708;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node713;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node738;
	wire [4-1:0] node740;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node750;
	wire [4-1:0] node752;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node817;
	wire [4-1:0] node819;
	wire [4-1:0] node822;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node855;
	wire [4-1:0] node857;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node907;
	wire [4-1:0] node909;
	wire [4-1:0] node911;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node921;
	wire [4-1:0] node924;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node947;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node964;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node972;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node996;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1004;
	wire [4-1:0] node1007;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1019;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1034;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1040;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1076;
	wire [4-1:0] node1079;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1093;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1100;
	wire [4-1:0] node1103;
	wire [4-1:0] node1106;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1133;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1148;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1163;
	wire [4-1:0] node1164;
	wire [4-1:0] node1166;
	wire [4-1:0] node1170;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1174;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1189;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1196;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1214;
	wire [4-1:0] node1217;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1229;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1244;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1254;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1268;
	wire [4-1:0] node1269;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1316;
	wire [4-1:0] node1319;
	wire [4-1:0] node1321;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1337;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1359;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1374;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1384;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1412;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1433;
	wire [4-1:0] node1437;
	wire [4-1:0] node1438;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1447;
	wire [4-1:0] node1450;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1470;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1487;
	wire [4-1:0] node1489;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1508;
	wire [4-1:0] node1510;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1527;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1544;
	wire [4-1:0] node1546;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1564;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1584;
	wire [4-1:0] node1587;
	wire [4-1:0] node1590;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1602;
	wire [4-1:0] node1604;
	wire [4-1:0] node1607;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1624;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1629;
	wire [4-1:0] node1630;
	wire [4-1:0] node1634;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1661;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1673;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1678;
	wire [4-1:0] node1683;
	wire [4-1:0] node1684;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1691;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1712;
	wire [4-1:0] node1715;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1722;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1733;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1740;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1773;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1801;
	wire [4-1:0] node1804;
	wire [4-1:0] node1806;
	wire [4-1:0] node1809;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1816;
	wire [4-1:0] node1818;
	wire [4-1:0] node1821;
	wire [4-1:0] node1822;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1834;
	wire [4-1:0] node1835;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1839;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1847;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1860;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1870;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1888;
	wire [4-1:0] node1890;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1897;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1901;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1911;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1918;
	wire [4-1:0] node1920;
	wire [4-1:0] node1923;
	wire [4-1:0] node1924;
	wire [4-1:0] node1927;
	wire [4-1:0] node1930;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1939;
	wire [4-1:0] node1941;
	wire [4-1:0] node1944;
	wire [4-1:0] node1946;
	wire [4-1:0] node1948;
	wire [4-1:0] node1950;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1958;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1966;
	wire [4-1:0] node1968;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1983;
	wire [4-1:0] node1984;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1991;
	wire [4-1:0] node1996;
	wire [4-1:0] node1998;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2011;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2016;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2030;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2036;
	wire [4-1:0] node2037;
	wire [4-1:0] node2039;
	wire [4-1:0] node2041;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2059;
	wire [4-1:0] node2061;
	wire [4-1:0] node2062;
	wire [4-1:0] node2066;
	wire [4-1:0] node2067;
	wire [4-1:0] node2068;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2075;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2085;
	wire [4-1:0] node2087;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2101;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2112;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2119;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2127;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2130;
	wire [4-1:0] node2132;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2147;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2154;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2160;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2172;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2181;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2187;
	wire [4-1:0] node2190;
	wire [4-1:0] node2191;
	wire [4-1:0] node2194;
	wire [4-1:0] node2197;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2204;
	wire [4-1:0] node2206;
	wire [4-1:0] node2208;
	wire [4-1:0] node2209;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2221;
	wire [4-1:0] node2222;
	wire [4-1:0] node2224;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2240;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2245;
	wire [4-1:0] node2246;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2265;
	wire [4-1:0] node2267;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2274;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2279;
	wire [4-1:0] node2281;
	wire [4-1:0] node2285;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2294;
	wire [4-1:0] node2295;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2311;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2317;
	wire [4-1:0] node2322;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2328;
	wire [4-1:0] node2331;
	wire [4-1:0] node2332;
	wire [4-1:0] node2334;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2340;
	wire [4-1:0] node2343;
	wire [4-1:0] node2344;
	wire [4-1:0] node2347;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2360;
	wire [4-1:0] node2363;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2370;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2378;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2384;
	wire [4-1:0] node2386;
	wire [4-1:0] node2389;
	wire [4-1:0] node2390;
	wire [4-1:0] node2393;
	wire [4-1:0] node2396;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2402;
	wire [4-1:0] node2404;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2411;
	wire [4-1:0] node2414;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2424;
	wire [4-1:0] node2427;
	wire [4-1:0] node2430;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2434;
	wire [4-1:0] node2437;
	wire [4-1:0] node2438;
	wire [4-1:0] node2439;
	wire [4-1:0] node2443;
	wire [4-1:0] node2446;
	wire [4-1:0] node2447;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2452;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2460;
	wire [4-1:0] node2461;
	wire [4-1:0] node2462;
	wire [4-1:0] node2464;
	wire [4-1:0] node2466;
	wire [4-1:0] node2469;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2476;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2482;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2489;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2494;
	wire [4-1:0] node2497;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2502;
	wire [4-1:0] node2503;
	wire [4-1:0] node2504;
	wire [4-1:0] node2506;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2515;
	wire [4-1:0] node2516;
	wire [4-1:0] node2518;
	wire [4-1:0] node2521;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2534;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2545;
	wire [4-1:0] node2547;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2562;
	wire [4-1:0] node2564;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2572;
	wire [4-1:0] node2573;
	wire [4-1:0] node2577;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2584;
	wire [4-1:0] node2587;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2596;
	wire [4-1:0] node2598;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2613;
	wire [4-1:0] node2615;
	wire [4-1:0] node2616;
	wire [4-1:0] node2619;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2627;
	wire [4-1:0] node2628;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2634;
	wire [4-1:0] node2638;
	wire [4-1:0] node2639;
	wire [4-1:0] node2641;
	wire [4-1:0] node2643;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2650;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2660;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2666;
	wire [4-1:0] node2669;
	wire [4-1:0] node2671;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2686;
	wire [4-1:0] node2687;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2699;
	wire [4-1:0] node2701;
	wire [4-1:0] node2704;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2727;
	wire [4-1:0] node2729;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2743;
	wire [4-1:0] node2744;
	wire [4-1:0] node2748;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2752;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2763;
	wire [4-1:0] node2765;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2773;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2786;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2791;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2820;
	wire [4-1:0] node2823;
	wire [4-1:0] node2825;
	wire [4-1:0] node2828;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2839;
	wire [4-1:0] node2841;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2847;
	wire [4-1:0] node2848;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2861;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2867;
	wire [4-1:0] node2869;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2875;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2881;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2887;
	wire [4-1:0] node2891;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2899;
	wire [4-1:0] node2902;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2909;
	wire [4-1:0] node2911;
	wire [4-1:0] node2913;
	wire [4-1:0] node2916;
	wire [4-1:0] node2917;
	wire [4-1:0] node2918;
	wire [4-1:0] node2920;
	wire [4-1:0] node2922;
	wire [4-1:0] node2924;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2935;
	wire [4-1:0] node2939;
	wire [4-1:0] node2940;
	wire [4-1:0] node2941;
	wire [4-1:0] node2945;
	wire [4-1:0] node2947;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2960;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2970;
	wire [4-1:0] node2974;
	wire [4-1:0] node2975;
	wire [4-1:0] node2976;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2982;
	wire [4-1:0] node2986;
	wire [4-1:0] node2987;
	wire [4-1:0] node2988;
	wire [4-1:0] node2993;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2996;
	wire [4-1:0] node2997;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3011;
	wire [4-1:0] node3012;
	wire [4-1:0] node3014;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3023;
	wire [4-1:0] node3027;
	wire [4-1:0] node3030;
	wire [4-1:0] node3031;
	wire [4-1:0] node3032;
	wire [4-1:0] node3034;
	wire [4-1:0] node3037;
	wire [4-1:0] node3038;
	wire [4-1:0] node3039;
	wire [4-1:0] node3044;
	wire [4-1:0] node3045;
	wire [4-1:0] node3046;
	wire [4-1:0] node3047;
	wire [4-1:0] node3049;
	wire [4-1:0] node3053;
	wire [4-1:0] node3054;
	wire [4-1:0] node3057;
	wire [4-1:0] node3060;
	wire [4-1:0] node3062;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3072;
	wire [4-1:0] node3075;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3084;
	wire [4-1:0] node3085;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3091;
	wire [4-1:0] node3094;
	wire [4-1:0] node3096;
	wire [4-1:0] node3098;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3104;
	wire [4-1:0] node3106;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3114;
	wire [4-1:0] node3116;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3130;
	wire [4-1:0] node3134;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3152;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3171;
	wire [4-1:0] node3172;
	wire [4-1:0] node3174;
	wire [4-1:0] node3176;
	wire [4-1:0] node3178;
	wire [4-1:0] node3181;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3185;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3197;
	wire [4-1:0] node3198;
	wire [4-1:0] node3202;
	wire [4-1:0] node3203;
	wire [4-1:0] node3205;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3216;
	wire [4-1:0] node3219;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3223;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3231;
	wire [4-1:0] node3233;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3239;
	wire [4-1:0] node3240;
	wire [4-1:0] node3242;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3256;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3259;
	wire [4-1:0] node3263;
	wire [4-1:0] node3265;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3275;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3282;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3295;
	wire [4-1:0] node3298;
	wire [4-1:0] node3299;
	wire [4-1:0] node3300;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3307;
	wire [4-1:0] node3311;
	wire [4-1:0] node3314;
	wire [4-1:0] node3315;
	wire [4-1:0] node3316;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3327;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3331;
	wire [4-1:0] node3333;
	wire [4-1:0] node3337;
	wire [4-1:0] node3339;
	wire [4-1:0] node3341;
	wire [4-1:0] node3344;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3350;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3357;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3367;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3381;
	wire [4-1:0] node3384;
	wire [4-1:0] node3387;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3395;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3400;
	wire [4-1:0] node3403;
	wire [4-1:0] node3406;
	wire [4-1:0] node3407;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3420;
	wire [4-1:0] node3424;
	wire [4-1:0] node3425;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3434;
	wire [4-1:0] node3436;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3443;
	wire [4-1:0] node3446;
	wire [4-1:0] node3448;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3458;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3464;
	wire [4-1:0] node3467;
	wire [4-1:0] node3470;
	wire [4-1:0] node3471;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3487;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3492;
	wire [4-1:0] node3493;
	wire [4-1:0] node3497;
	wire [4-1:0] node3498;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3506;
	wire [4-1:0] node3507;
	wire [4-1:0] node3509;
	wire [4-1:0] node3510;
	wire [4-1:0] node3512;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3526;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3532;
	wire [4-1:0] node3535;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3553;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3560;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3571;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3589;
	wire [4-1:0] node3590;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3596;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3613;
	wire [4-1:0] node3614;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3630;
	wire [4-1:0] node3633;
	wire [4-1:0] node3634;
	wire [4-1:0] node3638;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3642;
	wire [4-1:0] node3645;
	wire [4-1:0] node3647;
	wire [4-1:0] node3649;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3661;
	wire [4-1:0] node3665;
	wire [4-1:0] node3666;
	wire [4-1:0] node3667;
	wire [4-1:0] node3668;
	wire [4-1:0] node3670;
	wire [4-1:0] node3673;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3684;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3697;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3702;
	wire [4-1:0] node3707;
	wire [4-1:0] node3709;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3715;
	wire [4-1:0] node3716;
	wire [4-1:0] node3717;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3726;
	wire [4-1:0] node3729;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3734;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3741;
	wire [4-1:0] node3744;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3756;
	wire [4-1:0] node3757;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3761;
	wire [4-1:0] node3764;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3771;
	wire [4-1:0] node3772;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3780;
	wire [4-1:0] node3783;
	wire [4-1:0] node3785;
	wire [4-1:0] node3788;
	wire [4-1:0] node3790;
	wire [4-1:0] node3792;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3798;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3804;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3818;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3825;
	wire [4-1:0] node3829;
	wire [4-1:0] node3831;
	wire [4-1:0] node3833;
	wire [4-1:0] node3834;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3840;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3845;
	wire [4-1:0] node3848;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3855;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3867;
	wire [4-1:0] node3870;
	wire [4-1:0] node3871;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3881;
	wire [4-1:0] node3884;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3891;
	wire [4-1:0] node3892;
	wire [4-1:0] node3893;
	wire [4-1:0] node3894;
	wire [4-1:0] node3896;
	wire [4-1:0] node3899;
	wire [4-1:0] node3900;
	wire [4-1:0] node3902;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3910;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3918;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3925;
	wire [4-1:0] node3928;
	wire [4-1:0] node3930;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3939;
	wire [4-1:0] node3942;
	wire [4-1:0] node3945;
	wire [4-1:0] node3948;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3957;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3964;
	wire [4-1:0] node3966;
	wire [4-1:0] node3969;
	wire [4-1:0] node3970;
	wire [4-1:0] node3972;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3988;
	wire [4-1:0] node3991;
	wire [4-1:0] node3992;
	wire [4-1:0] node3994;
	wire [4-1:0] node3998;
	wire [4-1:0] node4000;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4007;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4012;
	wire [4-1:0] node4015;
	wire [4-1:0] node4017;
	wire [4-1:0] node4020;
	wire [4-1:0] node4021;
	wire [4-1:0] node4022;
	wire [4-1:0] node4023;
	wire [4-1:0] node4024;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4035;
	wire [4-1:0] node4038;
	wire [4-1:0] node4039;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4048;
	wire [4-1:0] node4051;
	wire [4-1:0] node4054;
	wire [4-1:0] node4056;
	wire [4-1:0] node4058;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4063;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4074;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4082;
	wire [4-1:0] node4083;
	wire [4-1:0] node4085;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4090;
	wire [4-1:0] node4092;
	wire [4-1:0] node4095;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4107;
	wire [4-1:0] node4110;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4121;
	wire [4-1:0] node4122;
	wire [4-1:0] node4123;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4137;
	wire [4-1:0] node4138;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4144;
	wire [4-1:0] node4145;
	wire [4-1:0] node4146;
	wire [4-1:0] node4147;
	wire [4-1:0] node4149;
	wire [4-1:0] node4152;
	wire [4-1:0] node4155;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4159;
	wire [4-1:0] node4163;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4168;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4175;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4181;
	wire [4-1:0] node4184;
	wire [4-1:0] node4185;
	wire [4-1:0] node4188;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4193;
	wire [4-1:0] node4194;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4201;
	wire [4-1:0] node4204;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4212;
	wire [4-1:0] node4215;
	wire [4-1:0] node4216;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4228;
	wire [4-1:0] node4229;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4236;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4244;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4258;
	wire [4-1:0] node4259;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4267;
	wire [4-1:0] node4268;
	wire [4-1:0] node4271;
	wire [4-1:0] node4274;
	wire [4-1:0] node4275;
	wire [4-1:0] node4276;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4282;
	wire [4-1:0] node4286;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4292;
	wire [4-1:0] node4295;
	wire [4-1:0] node4297;
	wire [4-1:0] node4300;
	wire [4-1:0] node4301;
	wire [4-1:0] node4304;
	wire [4-1:0] node4305;
	wire [4-1:0] node4306;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4316;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4324;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4330;
	wire [4-1:0] node4334;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4344;
	wire [4-1:0] node4346;
	wire [4-1:0] node4347;
	wire [4-1:0] node4351;
	wire [4-1:0] node4352;
	wire [4-1:0] node4353;
	wire [4-1:0] node4355;
	wire [4-1:0] node4357;
	wire [4-1:0] node4358;
	wire [4-1:0] node4361;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4368;
	wire [4-1:0] node4370;
	wire [4-1:0] node4373;
	wire [4-1:0] node4377;
	wire [4-1:0] node4380;
	wire [4-1:0] node4381;
	wire [4-1:0] node4382;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4386;
	wire [4-1:0] node4389;
	wire [4-1:0] node4391;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4398;
	wire [4-1:0] node4401;
	wire [4-1:0] node4402;
	wire [4-1:0] node4404;
	wire [4-1:0] node4406;
	wire [4-1:0] node4410;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4416;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4423;
	wire [4-1:0] node4427;
	wire [4-1:0] node4428;
	wire [4-1:0] node4430;
	wire [4-1:0] node4434;
	wire [4-1:0] node4435;
	wire [4-1:0] node4437;
	wire [4-1:0] node4440;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4444;
	wire [4-1:0] node4449;
	wire [4-1:0] node4450;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4455;
	wire [4-1:0] node4456;
	wire [4-1:0] node4457;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4466;
	wire [4-1:0] node4467;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4473;
	wire [4-1:0] node4475;
	wire [4-1:0] node4477;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4498;
	wire [4-1:0] node4499;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4508;
	wire [4-1:0] node4511;
	wire [4-1:0] node4512;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4518;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4530;
	wire [4-1:0] node4531;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4540;
	wire [4-1:0] node4542;
	wire [4-1:0] node4545;
	wire [4-1:0] node4548;
	wire [4-1:0] node4549;
	wire [4-1:0] node4550;
	wire [4-1:0] node4552;
	wire [4-1:0] node4554;
	wire [4-1:0] node4557;
	wire [4-1:0] node4559;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4570;
	wire [4-1:0] node4572;
	wire [4-1:0] node4575;
	wire [4-1:0] node4576;
	wire [4-1:0] node4577;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4585;
	wire [4-1:0] node4586;
	wire [4-1:0] node4589;
	wire [4-1:0] node4592;
	wire [4-1:0] node4593;
	wire [4-1:0] node4594;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4603;
	wire [4-1:0] node4604;
	wire [4-1:0] node4608;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4611;
	wire [4-1:0] node4617;
	wire [4-1:0] node4618;
	wire [4-1:0] node4619;
	wire [4-1:0] node4622;
	wire [4-1:0] node4625;
	wire [4-1:0] node4628;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4638;
	wire [4-1:0] node4639;
	wire [4-1:0] node4640;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4649;
	wire [4-1:0] node4650;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4656;
	wire [4-1:0] node4658;
	wire [4-1:0] node4660;
	wire [4-1:0] node4664;
	wire [4-1:0] node4666;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4671;
	wire [4-1:0] node4672;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4677;
	wire [4-1:0] node4679;
	wire [4-1:0] node4682;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4689;
	wire [4-1:0] node4690;
	wire [4-1:0] node4692;
	wire [4-1:0] node4695;
	wire [4-1:0] node4697;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4714;
	wire [4-1:0] node4716;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4725;
	wire [4-1:0] node4726;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4731;
	wire [4-1:0] node4733;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4745;
	wire [4-1:0] node4748;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4754;
	wire [4-1:0] node4757;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4766;
	wire [4-1:0] node4769;
	wire [4-1:0] node4771;
	wire [4-1:0] node4774;
	wire [4-1:0] node4775;
	wire [4-1:0] node4776;
	wire [4-1:0] node4777;
	wire [4-1:0] node4778;
	wire [4-1:0] node4783;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4790;
	wire [4-1:0] node4792;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4797;
	wire [4-1:0] node4799;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4805;
	wire [4-1:0] node4809;
	wire [4-1:0] node4810;
	wire [4-1:0] node4814;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4821;
	wire [4-1:0] node4822;
	wire [4-1:0] node4826;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4830;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4838;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4849;
	wire [4-1:0] node4855;
	wire [4-1:0] node4856;
	wire [4-1:0] node4857;
	wire [4-1:0] node4860;
	wire [4-1:0] node4862;
	wire [4-1:0] node4865;
	wire [4-1:0] node4867;
	wire [4-1:0] node4870;
	wire [4-1:0] node4871;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4878;
	wire [4-1:0] node4883;
	wire [4-1:0] node4886;
	wire [4-1:0] node4888;
	wire [4-1:0] node4889;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4896;
	wire [4-1:0] node4898;
	wire [4-1:0] node4901;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4905;
	wire [4-1:0] node4906;
	wire [4-1:0] node4907;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4922;
	wire [4-1:0] node4927;
	wire [4-1:0] node4929;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4934;
	wire [4-1:0] node4936;
	wire [4-1:0] node4939;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4945;
	wire [4-1:0] node4946;
	wire [4-1:0] node4948;
	wire [4-1:0] node4950;
	wire [4-1:0] node4952;
	wire [4-1:0] node4955;
	wire [4-1:0] node4956;
	wire [4-1:0] node4958;
	wire [4-1:0] node4961;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4967;
	wire [4-1:0] node4969;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4975;
	wire [4-1:0] node4980;
	wire [4-1:0] node4983;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4988;
	wire [4-1:0] node4991;
	wire [4-1:0] node4993;
	wire [4-1:0] node4994;
	wire [4-1:0] node4995;
	wire [4-1:0] node4998;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5005;
	wire [4-1:0] node5007;
	wire [4-1:0] node5011;
	wire [4-1:0] node5013;
	wire [4-1:0] node5014;
	wire [4-1:0] node5017;
	wire [4-1:0] node5020;
	wire [4-1:0] node5021;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5029;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5036;
	wire [4-1:0] node5037;
	wire [4-1:0] node5038;
	wire [4-1:0] node5041;
	wire [4-1:0] node5046;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5053;
	wire [4-1:0] node5054;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5062;
	wire [4-1:0] node5065;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5072;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5078;
	wire [4-1:0] node5080;
	wire [4-1:0] node5083;
	wire [4-1:0] node5085;
	wire [4-1:0] node5088;
	wire [4-1:0] node5089;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5096;
	wire [4-1:0] node5097;
	wire [4-1:0] node5099;
	wire [4-1:0] node5102;
	wire [4-1:0] node5105;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5109;
	wire [4-1:0] node5110;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5125;
	wire [4-1:0] node5128;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5134;
	wire [4-1:0] node5136;
	wire [4-1:0] node5139;
	wire [4-1:0] node5140;
	wire [4-1:0] node5142;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5166;
	wire [4-1:0] node5167;
	wire [4-1:0] node5169;
	wire [4-1:0] node5170;
	wire [4-1:0] node5174;
	wire [4-1:0] node5177;
	wire [4-1:0] node5178;
	wire [4-1:0] node5179;
	wire [4-1:0] node5181;
	wire [4-1:0] node5184;
	wire [4-1:0] node5186;
	wire [4-1:0] node5189;
	wire [4-1:0] node5190;
	wire [4-1:0] node5191;
	wire [4-1:0] node5192;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5203;
	wire [4-1:0] node5207;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5214;
	wire [4-1:0] node5215;
	wire [4-1:0] node5216;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5224;
	wire [4-1:0] node5225;
	wire [4-1:0] node5226;
	wire [4-1:0] node5230;
	wire [4-1:0] node5231;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5237;
	wire [4-1:0] node5238;
	wire [4-1:0] node5239;
	wire [4-1:0] node5241;
	wire [4-1:0] node5242;
	wire [4-1:0] node5244;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5250;
	wire [4-1:0] node5253;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5261;
	wire [4-1:0] node5262;
	wire [4-1:0] node5263;
	wire [4-1:0] node5264;
	wire [4-1:0] node5268;
	wire [4-1:0] node5269;
	wire [4-1:0] node5272;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5278;
	wire [4-1:0] node5283;
	wire [4-1:0] node5285;
	wire [4-1:0] node5286;
	wire [4-1:0] node5287;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5294;
	wire [4-1:0] node5297;
	wire [4-1:0] node5300;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5303;
	wire [4-1:0] node5307;
	wire [4-1:0] node5308;
	wire [4-1:0] node5311;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5318;
	wire [4-1:0] node5321;
	wire [4-1:0] node5322;
	wire [4-1:0] node5323;
	wire [4-1:0] node5324;
	wire [4-1:0] node5327;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5335;
	wire [4-1:0] node5338;
	wire [4-1:0] node5339;
	wire [4-1:0] node5341;
	wire [4-1:0] node5343;
	wire [4-1:0] node5346;
	wire [4-1:0] node5348;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5355;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5366;
	wire [4-1:0] node5367;
	wire [4-1:0] node5368;
	wire [4-1:0] node5369;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5379;
	wire [4-1:0] node5382;
	wire [4-1:0] node5385;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5390;
	wire [4-1:0] node5391;
	wire [4-1:0] node5395;
	wire [4-1:0] node5397;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5407;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5410;
	wire [4-1:0] node5414;
	wire [4-1:0] node5416;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5425;
	wire [4-1:0] node5426;
	wire [4-1:0] node5430;
	wire [4-1:0] node5432;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5437;
	wire [4-1:0] node5438;
	wire [4-1:0] node5442;
	wire [4-1:0] node5445;
	wire [4-1:0] node5446;
	wire [4-1:0] node5450;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5455;
	wire [4-1:0] node5457;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5469;
	wire [4-1:0] node5472;
	wire [4-1:0] node5473;
	wire [4-1:0] node5476;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5484;
	wire [4-1:0] node5487;
	wire [4-1:0] node5490;
	wire [4-1:0] node5492;
	wire [4-1:0] node5495;
	wire [4-1:0] node5496;
	wire [4-1:0] node5499;
	wire [4-1:0] node5500;
	wire [4-1:0] node5502;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5508;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5516;
	wire [4-1:0] node5517;
	wire [4-1:0] node5518;
	wire [4-1:0] node5522;
	wire [4-1:0] node5524;
	wire [4-1:0] node5527;
	wire [4-1:0] node5528;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5545;
	wire [4-1:0] node5546;
	wire [4-1:0] node5549;
	wire [4-1:0] node5550;
	wire [4-1:0] node5554;
	wire [4-1:0] node5556;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5564;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5574;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5577;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5598;
	wire [4-1:0] node5599;
	wire [4-1:0] node5600;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5608;
	wire [4-1:0] node5609;
	wire [4-1:0] node5611;
	wire [4-1:0] node5612;
	wire [4-1:0] node5617;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5621;
	wire [4-1:0] node5623;
	wire [4-1:0] node5624;
	wire [4-1:0] node5627;
	wire [4-1:0] node5630;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5637;
	wire [4-1:0] node5638;
	wire [4-1:0] node5639;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5647;
	wire [4-1:0] node5648;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5658;
	wire [4-1:0] node5662;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5668;
	wire [4-1:0] node5670;
	wire [4-1:0] node5673;
	wire [4-1:0] node5675;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5682;
	wire [4-1:0] node5683;
	wire [4-1:0] node5689;
	wire [4-1:0] node5691;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5700;
	wire [4-1:0] node5703;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5709;
	wire [4-1:0] node5713;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5719;
	wire [4-1:0] node5720;
	wire [4-1:0] node5725;
	wire [4-1:0] node5726;
	wire [4-1:0] node5728;
	wire [4-1:0] node5731;
	wire [4-1:0] node5732;
	wire [4-1:0] node5735;
	wire [4-1:0] node5738;
	wire [4-1:0] node5739;
	wire [4-1:0] node5740;
	wire [4-1:0] node5742;
	wire [4-1:0] node5743;
	wire [4-1:0] node5748;
	wire [4-1:0] node5749;
	wire [4-1:0] node5750;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5760;
	wire [4-1:0] node5763;
	wire [4-1:0] node5765;
	wire [4-1:0] node5768;
	wire [4-1:0] node5769;
	wire [4-1:0] node5770;
	wire [4-1:0] node5773;
	wire [4-1:0] node5776;
	wire [4-1:0] node5778;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5788;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5794;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5802;
	wire [4-1:0] node5803;
	wire [4-1:0] node5806;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5816;
	wire [4-1:0] node5819;
	wire [4-1:0] node5821;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5830;
	wire [4-1:0] node5834;
	wire [4-1:0] node5836;
	wire [4-1:0] node5838;
	wire [4-1:0] node5841;
	wire [4-1:0] node5842;
	wire [4-1:0] node5843;
	wire [4-1:0] node5845;
	wire [4-1:0] node5849;
	wire [4-1:0] node5851;
	wire [4-1:0] node5853;
	wire [4-1:0] node5856;
	wire [4-1:0] node5857;
	wire [4-1:0] node5858;
	wire [4-1:0] node5859;
	wire [4-1:0] node5860;
	wire [4-1:0] node5864;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5871;
	wire [4-1:0] node5872;
	wire [4-1:0] node5874;
	wire [4-1:0] node5877;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5888;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5894;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5903;
	wire [4-1:0] node5906;
	wire [4-1:0] node5907;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5913;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5918;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5926;
	wire [4-1:0] node5928;
	wire [4-1:0] node5931;
	wire [4-1:0] node5932;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5936;
	wire [4-1:0] node5940;
	wire [4-1:0] node5941;
	wire [4-1:0] node5945;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5951;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5957;
	wire [4-1:0] node5958;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5961;
	wire [4-1:0] node5967;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5972;
	wire [4-1:0] node5976;
	wire [4-1:0] node5977;
	wire [4-1:0] node5979;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5989;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5997;
	wire [4-1:0] node5998;
	wire [4-1:0] node5999;
	wire [4-1:0] node6000;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6007;
	wire [4-1:0] node6009;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6020;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6027;
	wire [4-1:0] node6028;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6031;
	wire [4-1:0] node6037;
	wire [4-1:0] node6038;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6045;
	wire [4-1:0] node6047;
	wire [4-1:0] node6048;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6059;
	wire [4-1:0] node6060;
	wire [4-1:0] node6063;
	wire [4-1:0] node6066;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6075;
	wire [4-1:0] node6079;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6086;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6091;
	wire [4-1:0] node6092;
	wire [4-1:0] node6095;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6101;
	wire [4-1:0] node6103;
	wire [4-1:0] node6106;
	wire [4-1:0] node6109;
	wire [4-1:0] node6110;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6114;
	wire [4-1:0] node6119;
	wire [4-1:0] node6122;
	wire [4-1:0] node6123;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6130;
	wire [4-1:0] node6132;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6141;
	wire [4-1:0] node6144;
	wire [4-1:0] node6145;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6152;
	wire [4-1:0] node6155;
	wire [4-1:0] node6158;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6165;
	wire [4-1:0] node6167;
	wire [4-1:0] node6168;
	wire [4-1:0] node6172;
	wire [4-1:0] node6173;
	wire [4-1:0] node6176;
	wire [4-1:0] node6178;
	wire [4-1:0] node6181;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6187;
	wire [4-1:0] node6188;
	wire [4-1:0] node6190;
	wire [4-1:0] node6193;
	wire [4-1:0] node6194;
	wire [4-1:0] node6195;
	wire [4-1:0] node6198;
	wire [4-1:0] node6202;
	wire [4-1:0] node6203;
	wire [4-1:0] node6204;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6211;
	wire [4-1:0] node6213;
	wire [4-1:0] node6216;
	wire [4-1:0] node6217;
	wire [4-1:0] node6218;
	wire [4-1:0] node6219;
	wire [4-1:0] node6222;
	wire [4-1:0] node6225;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6230;
	wire [4-1:0] node6231;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6241;
	wire [4-1:0] node6242;
	wire [4-1:0] node6245;
	wire [4-1:0] node6247;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6254;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6265;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6272;
	wire [4-1:0] node6273;
	wire [4-1:0] node6274;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6278;
	wire [4-1:0] node6281;
	wire [4-1:0] node6283;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6291;
	wire [4-1:0] node6293;
	wire [4-1:0] node6296;
	wire [4-1:0] node6297;
	wire [4-1:0] node6299;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6307;
	wire [4-1:0] node6311;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6314;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6319;
	wire [4-1:0] node6322;
	wire [4-1:0] node6324;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6330;
	wire [4-1:0] node6333;
	wire [4-1:0] node6336;
	wire [4-1:0] node6337;
	wire [4-1:0] node6338;
	wire [4-1:0] node6339;
	wire [4-1:0] node6343;
	wire [4-1:0] node6345;
	wire [4-1:0] node6347;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6365;
	wire [4-1:0] node6368;
	wire [4-1:0] node6371;
	wire [4-1:0] node6374;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6379;
	wire [4-1:0] node6382;
	wire [4-1:0] node6385;
	wire [4-1:0] node6387;
	wire [4-1:0] node6390;
	wire [4-1:0] node6391;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6395;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6402;
	wire [4-1:0] node6404;
	wire [4-1:0] node6407;
	wire [4-1:0] node6408;
	wire [4-1:0] node6409;
	wire [4-1:0] node6412;
	wire [4-1:0] node6413;
	wire [4-1:0] node6417;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6422;
	wire [4-1:0] node6423;
	wire [4-1:0] node6428;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6431;
	wire [4-1:0] node6432;
	wire [4-1:0] node6434;
	wire [4-1:0] node6437;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6451;
	wire [4-1:0] node6453;
	wire [4-1:0] node6456;
	wire [4-1:0] node6457;
	wire [4-1:0] node6458;
	wire [4-1:0] node6462;
	wire [4-1:0] node6463;
	wire [4-1:0] node6464;
	wire [4-1:0] node6467;
	wire [4-1:0] node6471;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6476;
	wire [4-1:0] node6477;
	wire [4-1:0] node6478;
	wire [4-1:0] node6483;
	wire [4-1:0] node6485;
	wire [4-1:0] node6486;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6493;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6498;
	wire [4-1:0] node6501;
	wire [4-1:0] node6503;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6510;
	wire [4-1:0] node6511;
	wire [4-1:0] node6513;
	wire [4-1:0] node6516;
	wire [4-1:0] node6518;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6527;
	wire [4-1:0] node6530;
	wire [4-1:0] node6531;
	wire [4-1:0] node6536;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6542;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6548;
	wire [4-1:0] node6553;
	wire [4-1:0] node6554;
	wire [4-1:0] node6555;
	wire [4-1:0] node6559;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6564;
	wire [4-1:0] node6565;
	wire [4-1:0] node6566;
	wire [4-1:0] node6568;
	wire [4-1:0] node6571;
	wire [4-1:0] node6573;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6582;
	wire [4-1:0] node6583;
	wire [4-1:0] node6585;
	wire [4-1:0] node6589;
	wire [4-1:0] node6592;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6599;
	wire [4-1:0] node6600;
	wire [4-1:0] node6601;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6606;
	wire [4-1:0] node6610;
	wire [4-1:0] node6612;
	wire [4-1:0] node6615;
	wire [4-1:0] node6616;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6622;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6630;
	wire [4-1:0] node6632;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6644;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6652;
	wire [4-1:0] node6656;
	wire [4-1:0] node6659;
	wire [4-1:0] node6661;
	wire [4-1:0] node6662;
	wire [4-1:0] node6666;
	wire [4-1:0] node6667;
	wire [4-1:0] node6668;
	wire [4-1:0] node6669;
	wire [4-1:0] node6673;
	wire [4-1:0] node6674;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6684;
	wire [4-1:0] node6686;
	wire [4-1:0] node6689;
	wire [4-1:0] node6691;
	wire [4-1:0] node6693;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6699;
	wire [4-1:0] node6702;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6711;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6718;
	wire [4-1:0] node6721;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6726;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6733;
	wire [4-1:0] node6735;
	wire [4-1:0] node6738;
	wire [4-1:0] node6739;
	wire [4-1:0] node6740;
	wire [4-1:0] node6742;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6749;
	wire [4-1:0] node6750;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6762;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6767;
	wire [4-1:0] node6770;
	wire [4-1:0] node6772;
	wire [4-1:0] node6773;
	wire [4-1:0] node6777;
	wire [4-1:0] node6778;
	wire [4-1:0] node6780;
	wire [4-1:0] node6783;
	wire [4-1:0] node6784;
	wire [4-1:0] node6786;
	wire [4-1:0] node6790;
	wire [4-1:0] node6791;
	wire [4-1:0] node6792;
	wire [4-1:0] node6793;
	wire [4-1:0] node6795;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6801;
	wire [4-1:0] node6803;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6810;
	wire [4-1:0] node6812;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6818;
	wire [4-1:0] node6821;
	wire [4-1:0] node6823;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6838;
	wire [4-1:0] node6841;
	wire [4-1:0] node6842;
	wire [4-1:0] node6844;
	wire [4-1:0] node6847;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6854;
	wire [4-1:0] node6857;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6865;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6872;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6877;
	wire [4-1:0] node6881;
	wire [4-1:0] node6883;
	wire [4-1:0] node6886;
	wire [4-1:0] node6887;
	wire [4-1:0] node6891;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6895;
	wire [4-1:0] node6899;
	wire [4-1:0] node6902;
	wire [4-1:0] node6903;
	wire [4-1:0] node6905;
	wire [4-1:0] node6909;
	wire [4-1:0] node6910;
	wire [4-1:0] node6913;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6928;
	wire [4-1:0] node6930;
	wire [4-1:0] node6933;
	wire [4-1:0] node6934;
	wire [4-1:0] node6935;
	wire [4-1:0] node6938;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6945;
	wire [4-1:0] node6947;
	wire [4-1:0] node6951;
	wire [4-1:0] node6952;
	wire [4-1:0] node6953;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6958;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6967;
	wire [4-1:0] node6969;
	wire [4-1:0] node6971;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6977;
	wire [4-1:0] node6980;
	wire [4-1:0] node6982;
	wire [4-1:0] node6985;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6989;
	wire [4-1:0] node6992;
	wire [4-1:0] node6994;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node6999;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7007;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7013;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7024;
	wire [4-1:0] node7025;
	wire [4-1:0] node7027;
	wire [4-1:0] node7028;
	wire [4-1:0] node7031;
	wire [4-1:0] node7034;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7041;
	wire [4-1:0] node7042;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7055;
	wire [4-1:0] node7058;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7066;
	wire [4-1:0] node7068;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7074;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7080;
	wire [4-1:0] node7084;
	wire [4-1:0] node7085;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7097;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7100;
	wire [4-1:0] node7101;
	wire [4-1:0] node7102;
	wire [4-1:0] node7106;
	wire [4-1:0] node7108;
	wire [4-1:0] node7109;
	wire [4-1:0] node7113;
	wire [4-1:0] node7114;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7120;
	wire [4-1:0] node7123;
	wire [4-1:0] node7126;
	wire [4-1:0] node7128;
	wire [4-1:0] node7129;
	wire [4-1:0] node7131;
	wire [4-1:0] node7134;
	wire [4-1:0] node7137;
	wire [4-1:0] node7138;
	wire [4-1:0] node7139;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7153;
	wire [4-1:0] node7154;
	wire [4-1:0] node7156;
	wire [4-1:0] node7158;
	wire [4-1:0] node7159;
	wire [4-1:0] node7164;
	wire [4-1:0] node7165;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7174;
	wire [4-1:0] node7176;
	wire [4-1:0] node7179;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7187;
	wire [4-1:0] node7190;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7196;
	wire [4-1:0] node7199;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7206;
	wire [4-1:0] node7207;
	wire [4-1:0] node7211;
	wire [4-1:0] node7212;
	wire [4-1:0] node7213;
	wire [4-1:0] node7214;
	wire [4-1:0] node7216;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7221;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7232;
	wire [4-1:0] node7235;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7243;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7254;
	wire [4-1:0] node7257;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7275;
	wire [4-1:0] node7278;
	wire [4-1:0] node7281;
	wire [4-1:0] node7282;
	wire [4-1:0] node7284;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7293;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7300;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7308;
	wire [4-1:0] node7311;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7314;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7317;
	wire [4-1:0] node7319;
	wire [4-1:0] node7321;
	wire [4-1:0] node7322;
	wire [4-1:0] node7326;
	wire [4-1:0] node7328;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7339;
	wire [4-1:0] node7341;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7348;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7355;
	wire [4-1:0] node7357;
	wire [4-1:0] node7359;
	wire [4-1:0] node7362;
	wire [4-1:0] node7365;
	wire [4-1:0] node7366;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7371;
	wire [4-1:0] node7376;
	wire [4-1:0] node7377;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7383;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7390;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7395;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7408;
	wire [4-1:0] node7409;
	wire [4-1:0] node7412;
	wire [4-1:0] node7413;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7419;
	wire [4-1:0] node7422;
	wire [4-1:0] node7425;
	wire [4-1:0] node7426;
	wire [4-1:0] node7429;
	wire [4-1:0] node7431;
	wire [4-1:0] node7434;
	wire [4-1:0] node7435;
	wire [4-1:0] node7436;
	wire [4-1:0] node7437;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7442;
	wire [4-1:0] node7445;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7461;
	wire [4-1:0] node7465;
	wire [4-1:0] node7467;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7474;
	wire [4-1:0] node7476;
	wire [4-1:0] node7478;
	wire [4-1:0] node7482;
	wire [4-1:0] node7483;
	wire [4-1:0] node7484;
	wire [4-1:0] node7487;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7494;
	wire [4-1:0] node7497;
	wire [4-1:0] node7498;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7501;
	wire [4-1:0] node7502;
	wire [4-1:0] node7505;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7512;
	wire [4-1:0] node7514;
	wire [4-1:0] node7515;
	wire [4-1:0] node7518;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7528;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7534;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7544;
	wire [4-1:0] node7550;
	wire [4-1:0] node7551;
	wire [4-1:0] node7554;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7559;
	wire [4-1:0] node7560;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7566;
	wire [4-1:0] node7567;
	wire [4-1:0] node7568;
	wire [4-1:0] node7573;
	wire [4-1:0] node7574;
	wire [4-1:0] node7576;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7586;
	wire [4-1:0] node7587;
	wire [4-1:0] node7589;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7595;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7603;
	wire [4-1:0] node7607;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7618;
	wire [4-1:0] node7619;
	wire [4-1:0] node7620;
	wire [4-1:0] node7621;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7626;
	wire [4-1:0] node7627;
	wire [4-1:0] node7628;
	wire [4-1:0] node7631;
	wire [4-1:0] node7634;
	wire [4-1:0] node7636;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7644;
	wire [4-1:0] node7647;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7653;
	wire [4-1:0] node7656;
	wire [4-1:0] node7657;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7664;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7669;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7673;
	wire [4-1:0] node7678;
	wire [4-1:0] node7680;
	wire [4-1:0] node7681;
	wire [4-1:0] node7683;
	wire [4-1:0] node7687;
	wire [4-1:0] node7688;
	wire [4-1:0] node7690;
	wire [4-1:0] node7692;
	wire [4-1:0] node7695;
	wire [4-1:0] node7697;
	wire [4-1:0] node7699;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7708;
	wire [4-1:0] node7710;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7715;
	wire [4-1:0] node7718;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7724;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7733;
	wire [4-1:0] node7735;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7743;
	wire [4-1:0] node7744;
	wire [4-1:0] node7746;
	wire [4-1:0] node7747;
	wire [4-1:0] node7750;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7758;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7768;
	wire [4-1:0] node7770;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7777;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7784;
	wire [4-1:0] node7785;
	wire [4-1:0] node7788;
	wire [4-1:0] node7791;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7800;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7811;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7815;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7818;
	wire [4-1:0] node7822;
	wire [4-1:0] node7825;
	wire [4-1:0] node7826;
	wire [4-1:0] node7829;
	wire [4-1:0] node7830;
	wire [4-1:0] node7834;
	wire [4-1:0] node7836;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7841;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7849;
	wire [4-1:0] node7851;
	wire [4-1:0] node7854;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7861;
	wire [4-1:0] node7862;
	wire [4-1:0] node7865;
	wire [4-1:0] node7868;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7873;
	wire [4-1:0] node7876;
	wire [4-1:0] node7877;
	wire [4-1:0] node7879;
	wire [4-1:0] node7883;
	wire [4-1:0] node7884;
	wire [4-1:0] node7887;
	wire [4-1:0] node7888;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7904;
	wire [4-1:0] node7905;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7914;
	wire [4-1:0] node7917;
	wire [4-1:0] node7918;
	wire [4-1:0] node7919;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7925;
	wire [4-1:0] node7928;
	wire [4-1:0] node7929;
	wire [4-1:0] node7930;
	wire [4-1:0] node7933;
	wire [4-1:0] node7935;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7955;
	wire [4-1:0] node7956;
	wire [4-1:0] node7958;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7966;
	wire [4-1:0] node7969;
	wire [4-1:0] node7970;
	wire [4-1:0] node7971;
	wire [4-1:0] node7972;
	wire [4-1:0] node7976;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7986;
	wire [4-1:0] node7989;
	wire [4-1:0] node7991;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node7997;
	wire [4-1:0] node7998;
	wire [4-1:0] node7999;
	wire [4-1:0] node8000;
	wire [4-1:0] node8002;
	wire [4-1:0] node8006;
	wire [4-1:0] node8008;
	wire [4-1:0] node8010;
	wire [4-1:0] node8012;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8017;
	wire [4-1:0] node8020;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8025;
	wire [4-1:0] node8027;
	wire [4-1:0] node8031;
	wire [4-1:0] node8032;
	wire [4-1:0] node8033;
	wire [4-1:0] node8037;
	wire [4-1:0] node8040;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8045;
	wire [4-1:0] node8046;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8058;
	wire [4-1:0] node8060;
	wire [4-1:0] node8063;
	wire [4-1:0] node8066;
	wire [4-1:0] node8067;
	wire [4-1:0] node8068;
	wire [4-1:0] node8072;
	wire [4-1:0] node8074;
	wire [4-1:0] node8076;
	wire [4-1:0] node8077;
	wire [4-1:0] node8080;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8086;
	wire [4-1:0] node8087;
	wire [4-1:0] node8088;
	wire [4-1:0] node8092;
	wire [4-1:0] node8093;
	wire [4-1:0] node8096;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8103;
	wire [4-1:0] node8104;
	wire [4-1:0] node8105;
	wire [4-1:0] node8108;
	wire [4-1:0] node8111;
	wire [4-1:0] node8114;
	wire [4-1:0] node8115;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8128;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8135;
	wire [4-1:0] node8137;
	wire [4-1:0] node8140;
	wire [4-1:0] node8142;
	wire [4-1:0] node8145;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8148;
	wire [4-1:0] node8151;
	wire [4-1:0] node8153;
	wire [4-1:0] node8155;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8161;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8171;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8175;
	wire [4-1:0] node8178;
	wire [4-1:0] node8180;
	wire [4-1:0] node8182;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8190;
	wire [4-1:0] node8191;
	wire [4-1:0] node8192;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8195;
	wire [4-1:0] node8197;
	wire [4-1:0] node8199;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8209;
	wire [4-1:0] node8210;
	wire [4-1:0] node8211;
	wire [4-1:0] node8215;
	wire [4-1:0] node8218;
	wire [4-1:0] node8219;
	wire [4-1:0] node8221;
	wire [4-1:0] node8224;
	wire [4-1:0] node8225;
	wire [4-1:0] node8227;
	wire [4-1:0] node8231;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8243;
	wire [4-1:0] node8244;
	wire [4-1:0] node8246;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8256;
	wire [4-1:0] node8259;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8267;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8275;
	wire [4-1:0] node8276;
	wire [4-1:0] node8281;
	wire [4-1:0] node8282;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8288;
	wire [4-1:0] node8291;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8297;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8309;
	wire [4-1:0] node8312;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8319;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8326;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8334;
	wire [4-1:0] node8335;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8351;
	wire [4-1:0] node8356;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8361;
	wire [4-1:0] node8364;
	wire [4-1:0] node8367;
	wire [4-1:0] node8368;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8372;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8381;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8392;
	wire [4-1:0] node8395;
	wire [4-1:0] node8396;
	wire [4-1:0] node8398;
	wire [4-1:0] node8402;
	wire [4-1:0] node8403;
	wire [4-1:0] node8404;
	wire [4-1:0] node8406;
	wire [4-1:0] node8408;
	wire [4-1:0] node8411;
	wire [4-1:0] node8412;
	wire [4-1:0] node8413;
	wire [4-1:0] node8415;
	wire [4-1:0] node8418;
	wire [4-1:0] node8419;
	wire [4-1:0] node8423;
	wire [4-1:0] node8426;
	wire [4-1:0] node8427;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8432;
	wire [4-1:0] node8433;
	wire [4-1:0] node8438;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8451;
	wire [4-1:0] node8452;
	wire [4-1:0] node8456;
	wire [4-1:0] node8459;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8467;
	wire [4-1:0] node8469;
	wire [4-1:0] node8472;
	wire [4-1:0] node8473;
	wire [4-1:0] node8474;
	wire [4-1:0] node8477;
	wire [4-1:0] node8479;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8484;
	wire [4-1:0] node8486;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8494;
	wire [4-1:0] node8497;
	wire [4-1:0] node8498;
	wire [4-1:0] node8499;
	wire [4-1:0] node8500;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8512;
	wire [4-1:0] node8513;
	wire [4-1:0] node8516;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8528;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8536;
	wire [4-1:0] node8539;
	wire [4-1:0] node8540;
	wire [4-1:0] node8542;
	wire [4-1:0] node8545;
	wire [4-1:0] node8547;
	wire [4-1:0] node8550;
	wire [4-1:0] node8551;
	wire [4-1:0] node8552;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8559;
	wire [4-1:0] node8562;
	wire [4-1:0] node8565;
	wire [4-1:0] node8566;
	wire [4-1:0] node8569;
	wire [4-1:0] node8571;
	wire [4-1:0] node8573;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8578;
	wire [4-1:0] node8581;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8588;
	wire [4-1:0] node8589;
	wire [4-1:0] node8592;
	wire [4-1:0] node8594;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8601;
	wire [4-1:0] node8604;
	wire [4-1:0] node8605;
	wire [4-1:0] node8606;
	wire [4-1:0] node8609;
	wire [4-1:0] node8611;
	wire [4-1:0] node8614;
	wire [4-1:0] node8615;
	wire [4-1:0] node8619;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8629;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8637;
	wire [4-1:0] node8639;
	wire [4-1:0] node8642;
	wire [4-1:0] node8643;
	wire [4-1:0] node8644;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8649;
	wire [4-1:0] node8651;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8668;
	wire [4-1:0] node8669;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8677;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8682;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8689;
	wire [4-1:0] node8693;
	wire [4-1:0] node8694;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8702;
	wire [4-1:0] node8703;
	wire [4-1:0] node8706;
	wire [4-1:0] node8708;
	wire [4-1:0] node8711;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8715;
	wire [4-1:0] node8716;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8723;
	wire [4-1:0] node8725;
	wire [4-1:0] node8726;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8734;
	wire [4-1:0] node8737;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8746;
	wire [4-1:0] node8748;
	wire [4-1:0] node8751;
	wire [4-1:0] node8753;
	wire [4-1:0] node8757;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8761;
	wire [4-1:0] node8764;
	wire [4-1:0] node8765;
	wire [4-1:0] node8767;
	wire [4-1:0] node8768;
	wire [4-1:0] node8772;
	wire [4-1:0] node8774;
	wire [4-1:0] node8777;
	wire [4-1:0] node8778;
	wire [4-1:0] node8780;
	wire [4-1:0] node8783;
	wire [4-1:0] node8784;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8795;
	wire [4-1:0] node8796;
	wire [4-1:0] node8798;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8809;
	wire [4-1:0] node8810;
	wire [4-1:0] node8813;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8819;
	wire [4-1:0] node8821;
	wire [4-1:0] node8825;
	wire [4-1:0] node8827;
	wire [4-1:0] node8828;
	wire [4-1:0] node8830;
	wire [4-1:0] node8834;
	wire [4-1:0] node8835;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8842;
	wire [4-1:0] node8844;
	wire [4-1:0] node8845;
	wire [4-1:0] node8848;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8856;
	wire [4-1:0] node8858;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8865;
	wire [4-1:0] node8867;
	wire [4-1:0] node8871;
	wire [4-1:0] node8872;
	wire [4-1:0] node8873;
	wire [4-1:0] node8876;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8886;
	wire [4-1:0] node8890;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8908;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8918;
	wire [4-1:0] node8920;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8930;
	wire [4-1:0] node8932;
	wire [4-1:0] node8935;
	wire [4-1:0] node8936;
	wire [4-1:0] node8938;
	wire [4-1:0] node8939;
	wire [4-1:0] node8942;
	wire [4-1:0] node8943;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8950;
	wire [4-1:0] node8951;
	wire [4-1:0] node8955;
	wire [4-1:0] node8956;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8964;
	wire [4-1:0] node8968;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8976;
	wire [4-1:0] node8978;
	wire [4-1:0] node8979;
	wire [4-1:0] node8983;
	wire [4-1:0] node8986;
	wire [4-1:0] node8987;
	wire [4-1:0] node8988;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9007;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9013;
	wire [4-1:0] node9017;
	wire [4-1:0] node9019;
	wire [4-1:0] node9021;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9027;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9035;
	wire [4-1:0] node9038;
	wire [4-1:0] node9041;
	wire [4-1:0] node9043;
	wire [4-1:0] node9047;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9050;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9062;
	wire [4-1:0] node9063;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9072;
	wire [4-1:0] node9076;
	wire [4-1:0] node9078;
	wire [4-1:0] node9081;
	wire [4-1:0] node9082;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9090;
	wire [4-1:0] node9092;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9100;
	wire [4-1:0] node9101;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9104;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9111;
	wire [4-1:0] node9113;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9119;
	wire [4-1:0] node9122;
	wire [4-1:0] node9123;
	wire [4-1:0] node9125;
	wire [4-1:0] node9129;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9135;
	wire [4-1:0] node9141;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9147;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9153;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9160;
	wire [4-1:0] node9163;
	wire [4-1:0] node9165;
	wire [4-1:0] node9168;
	wire [4-1:0] node9169;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9173;
	wire [4-1:0] node9174;
	wire [4-1:0] node9176;
	wire [4-1:0] node9179;
	wire [4-1:0] node9180;
	wire [4-1:0] node9184;
	wire [4-1:0] node9185;
	wire [4-1:0] node9187;
	wire [4-1:0] node9190;
	wire [4-1:0] node9191;
	wire [4-1:0] node9193;
	wire [4-1:0] node9197;
	wire [4-1:0] node9198;
	wire [4-1:0] node9200;
	wire [4-1:0] node9202;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9210;
	wire [4-1:0] node9214;
	wire [4-1:0] node9215;
	wire [4-1:0] node9216;
	wire [4-1:0] node9219;
	wire [4-1:0] node9221;
	wire [4-1:0] node9222;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9228;
	wire [4-1:0] node9229;
	wire [4-1:0] node9235;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9242;
	wire [4-1:0] node9243;
	wire [4-1:0] node9249;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9255;
	wire [4-1:0] node9256;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9266;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9271;
	wire [4-1:0] node9272;
	wire [4-1:0] node9276;
	wire [4-1:0] node9278;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9285;
	wire [4-1:0] node9289;
	wire [4-1:0] node9290;
	wire [4-1:0] node9292;
	wire [4-1:0] node9294;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9302;
	wire [4-1:0] node9305;
	wire [4-1:0] node9306;
	wire [4-1:0] node9309;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9315;
	wire [4-1:0] node9317;
	wire [4-1:0] node9320;
	wire [4-1:0] node9321;
	wire [4-1:0] node9323;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9333;
	wire [4-1:0] node9337;
	wire [4-1:0] node9340;
	wire [4-1:0] node9341;
	wire [4-1:0] node9342;
	wire [4-1:0] node9343;
	wire [4-1:0] node9345;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9352;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9360;
	wire [4-1:0] node9362;
	wire [4-1:0] node9365;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9369;
	wire [4-1:0] node9372;
	wire [4-1:0] node9374;
	wire [4-1:0] node9375;
	wire [4-1:0] node9377;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9388;
	wire [4-1:0] node9390;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9400;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9405;
	wire [4-1:0] node9407;
	wire [4-1:0] node9412;
	wire [4-1:0] node9413;
	wire [4-1:0] node9415;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9427;
	wire [4-1:0] node9428;
	wire [4-1:0] node9429;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9435;
	wire [4-1:0] node9439;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9454;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9457;
	wire [4-1:0] node9460;
	wire [4-1:0] node9462;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9470;
	wire [4-1:0] node9472;
	wire [4-1:0] node9475;
	wire [4-1:0] node9476;
	wire [4-1:0] node9480;
	wire [4-1:0] node9481;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9490;
	wire [4-1:0] node9493;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9501;
	wire [4-1:0] node9502;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9509;
	wire [4-1:0] node9510;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9518;
	wire [4-1:0] node9519;
	wire [4-1:0] node9521;
	wire [4-1:0] node9526;
	wire [4-1:0] node9527;
	wire [4-1:0] node9528;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9537;
	wire [4-1:0] node9538;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9543;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9555;
	wire [4-1:0] node9556;
	wire [4-1:0] node9558;
	wire [4-1:0] node9560;
	wire [4-1:0] node9563;
	wire [4-1:0] node9565;
	wire [4-1:0] node9566;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9578;
	wire [4-1:0] node9581;
	wire [4-1:0] node9582;
	wire [4-1:0] node9583;
	wire [4-1:0] node9588;
	wire [4-1:0] node9589;
	wire [4-1:0] node9591;
	wire [4-1:0] node9593;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9616;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9622;
	wire [4-1:0] node9624;
	wire [4-1:0] node9626;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9633;
	wire [4-1:0] node9634;
	wire [4-1:0] node9637;
	wire [4-1:0] node9640;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9647;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9665;
	wire [4-1:0] node9666;
	wire [4-1:0] node9670;
	wire [4-1:0] node9671;

	assign outp = (inp[3]) ? node5366 : node1;
		assign node1 = (inp[6]) ? node2993 : node2;
			assign node2 = (inp[8]) ? node1492 : node3;
				assign node3 = (inp[14]) ? node757 : node4;
					assign node4 = (inp[9]) ? node388 : node5;
						assign node5 = (inp[0]) ? node185 : node6;
							assign node6 = (inp[13]) ? node104 : node7;
								assign node7 = (inp[2]) ? node51 : node8;
									assign node8 = (inp[4]) ? node20 : node9;
										assign node9 = (inp[10]) ? node15 : node10;
											assign node10 = (inp[5]) ? 4'b0000 : node11;
												assign node11 = (inp[7]) ? 4'b0001 : 4'b0010;
											assign node15 = (inp[5]) ? node17 : 4'b0001;
												assign node17 = (inp[11]) ? 4'b0001 : 4'b0100;
										assign node20 = (inp[7]) ? node38 : node21;
											assign node21 = (inp[11]) ? node27 : node22;
												assign node22 = (inp[5]) ? 4'b0001 : node23;
													assign node23 = (inp[1]) ? 4'b0001 : 4'b0011;
												assign node27 = (inp[10]) ? node35 : node28;
													assign node28 = (inp[5]) ? node32 : node29;
														assign node29 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node32 = (inp[12]) ? 4'b0111 : 4'b0101;
													assign node35 = (inp[12]) ? 4'b0111 : 4'b0000;
											assign node38 = (inp[1]) ? node40 : 4'b0111;
												assign node40 = (inp[10]) ? node46 : node41;
													assign node41 = (inp[12]) ? node43 : 4'b0100;
														assign node43 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node46 = (inp[12]) ? 4'b0011 : node47;
														assign node47 = (inp[11]) ? 4'b0011 : 4'b0000;
									assign node51 = (inp[4]) ? node85 : node52;
										assign node52 = (inp[15]) ? node72 : node53;
											assign node53 = (inp[5]) ? node65 : node54;
												assign node54 = (inp[10]) ? node60 : node55;
													assign node55 = (inp[12]) ? 4'b0111 : node56;
														assign node56 = (inp[7]) ? 4'b0110 : 4'b0100;
													assign node60 = (inp[1]) ? node62 : 4'b0111;
														assign node62 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node65 = (inp[11]) ? node69 : node66;
													assign node66 = (inp[12]) ? 4'b0001 : 4'b0011;
													assign node69 = (inp[10]) ? 4'b0101 : 4'b0111;
											assign node72 = (inp[10]) ? 4'b0010 : node73;
												assign node73 = (inp[12]) ? node77 : node74;
													assign node74 = (inp[7]) ? 4'b0110 : 4'b0100;
													assign node77 = (inp[7]) ? node81 : node78;
														assign node78 = (inp[11]) ? 4'b0010 : 4'b0110;
														assign node81 = (inp[5]) ? 4'b0100 : 4'b0001;
										assign node85 = (inp[5]) ? node95 : node86;
											assign node86 = (inp[11]) ? node92 : node87;
												assign node87 = (inp[1]) ? node89 : 4'b0011;
													assign node89 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node92 = (inp[7]) ? 4'b0001 : 4'b0010;
											assign node95 = (inp[1]) ? node101 : node96;
												assign node96 = (inp[10]) ? 4'b0100 : node97;
													assign node97 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node101 = (inp[10]) ? 4'b0001 : 4'b0000;
								assign node104 = (inp[2]) ? node134 : node105;
									assign node105 = (inp[5]) ? node119 : node106;
										assign node106 = (inp[1]) ? node112 : node107;
											assign node107 = (inp[4]) ? 4'b0010 : node108;
												assign node108 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node112 = (inp[11]) ? node116 : node113;
												assign node113 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node116 = (inp[4]) ? 4'b0010 : 4'b0100;
										assign node119 = (inp[12]) ? node125 : node120;
											assign node120 = (inp[1]) ? node122 : 4'b0010;
												assign node122 = (inp[11]) ? 4'b0010 : 4'b0000;
											assign node125 = (inp[11]) ? 4'b0101 : node126;
												assign node126 = (inp[1]) ? 4'b0000 : node127;
													assign node127 = (inp[10]) ? 4'b0100 : node128;
														assign node128 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node134 = (inp[1]) ? node166 : node135;
										assign node135 = (inp[12]) ? node151 : node136;
											assign node136 = (inp[10]) ? node146 : node137;
												assign node137 = (inp[5]) ? node141 : node138;
													assign node138 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node141 = (inp[15]) ? 4'b0000 : node142;
														assign node142 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node146 = (inp[11]) ? 4'b0010 : node147;
													assign node147 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node151 = (inp[4]) ? node157 : node152;
												assign node152 = (inp[11]) ? node154 : 4'b0010;
													assign node154 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node157 = (inp[7]) ? node163 : node158;
													assign node158 = (inp[10]) ? node160 : 4'b0111;
														assign node160 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node163 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node166 = (inp[5]) ? node178 : node167;
											assign node167 = (inp[11]) ? node171 : node168;
												assign node168 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node171 = (inp[12]) ? node175 : node172;
													assign node172 = (inp[15]) ? 4'b0110 : 4'b0011;
													assign node175 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node178 = (inp[11]) ? node182 : node179;
												assign node179 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node182 = (inp[4]) ? 4'b0010 : 4'b0110;
							assign node185 = (inp[1]) ? node295 : node186;
								assign node186 = (inp[4]) ? node234 : node187;
									assign node187 = (inp[2]) ? node221 : node188;
										assign node188 = (inp[13]) ? node206 : node189;
											assign node189 = (inp[7]) ? node197 : node190;
												assign node190 = (inp[12]) ? node194 : node191;
													assign node191 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node194 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node197 = (inp[12]) ? node201 : node198;
													assign node198 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node201 = (inp[5]) ? 4'b0100 : node202;
														assign node202 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node206 = (inp[11]) ? node212 : node207;
												assign node207 = (inp[12]) ? 4'b0101 : node208;
													assign node208 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node212 = (inp[15]) ? node218 : node213;
													assign node213 = (inp[10]) ? node215 : 4'b0111;
														assign node215 = (inp[12]) ? 4'b0100 : 4'b0100;
													assign node218 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node221 = (inp[10]) ? node227 : node222;
											assign node222 = (inp[11]) ? 4'b0010 : node223;
												assign node223 = (inp[13]) ? 4'b0010 : 4'b0100;
											assign node227 = (inp[7]) ? node231 : node228;
												assign node228 = (inp[13]) ? 4'b0010 : 4'b0101;
												assign node231 = (inp[12]) ? 4'b0100 : 4'b0110;
									assign node234 = (inp[12]) ? node262 : node235;
										assign node235 = (inp[5]) ? node251 : node236;
											assign node236 = (inp[11]) ? node242 : node237;
												assign node237 = (inp[13]) ? node239 : 4'b0000;
													assign node239 = (inp[10]) ? 4'b0110 : 4'b0100;
												assign node242 = (inp[10]) ? node246 : node243;
													assign node243 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node246 = (inp[2]) ? node248 : 4'b0110;
														assign node248 = (inp[15]) ? 4'b0101 : 4'b0001;
											assign node251 = (inp[2]) ? node253 : 4'b0000;
												assign node253 = (inp[13]) ? 4'b0010 : node254;
													assign node254 = (inp[11]) ? node258 : node255;
														assign node255 = (inp[7]) ? 4'b0101 : 4'b0010;
														assign node258 = (inp[10]) ? 4'b0110 : 4'b0100;
										assign node262 = (inp[2]) ? node284 : node263;
											assign node263 = (inp[10]) ? node277 : node264;
												assign node264 = (inp[7]) ? node270 : node265;
													assign node265 = (inp[5]) ? node267 : 4'b0011;
														assign node267 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node270 = (inp[15]) ? node274 : node271;
														assign node271 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node274 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node277 = (inp[5]) ? 4'b0110 : node278;
													assign node278 = (inp[13]) ? node280 : 4'b0000;
														assign node280 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node284 = (inp[5]) ? node290 : node285;
												assign node285 = (inp[15]) ? node287 : 4'b0100;
													assign node287 = (inp[13]) ? 4'b0110 : 4'b0100;
												assign node290 = (inp[7]) ? 4'b0011 : node291;
													assign node291 = (inp[10]) ? 4'b0010 : 4'b0011;
								assign node295 = (inp[5]) ? node347 : node296;
									assign node296 = (inp[15]) ? node326 : node297;
										assign node297 = (inp[4]) ? node307 : node298;
											assign node298 = (inp[2]) ? 4'b0011 : node299;
												assign node299 = (inp[13]) ? 4'b0110 : node300;
													assign node300 = (inp[12]) ? 4'b0101 : node301;
														assign node301 = (inp[10]) ? 4'b0010 : 4'b0001;
											assign node307 = (inp[7]) ? node315 : node308;
												assign node308 = (inp[12]) ? 4'b0111 : node309;
													assign node309 = (inp[13]) ? node311 : 4'b0100;
														assign node311 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node315 = (inp[12]) ? node321 : node316;
													assign node316 = (inp[13]) ? 4'b0110 : node317;
														assign node317 = (inp[11]) ? 4'b0010 : 4'b0110;
													assign node321 = (inp[2]) ? node323 : 4'b0101;
														assign node323 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node326 = (inp[2]) ? node334 : node327;
											assign node327 = (inp[13]) ? node331 : node328;
												assign node328 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node331 = (inp[7]) ? 4'b0100 : 4'b0110;
											assign node334 = (inp[11]) ? node340 : node335;
												assign node335 = (inp[4]) ? 4'b0010 : node336;
													assign node336 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node340 = (inp[4]) ? 4'b0101 : node341;
													assign node341 = (inp[13]) ? 4'b0111 : node342;
														assign node342 = (inp[7]) ? 4'b0010 : 4'b0110;
									assign node347 = (inp[10]) ? node369 : node348;
										assign node348 = (inp[15]) ? node356 : node349;
											assign node349 = (inp[2]) ? node353 : node350;
												assign node350 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node353 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node356 = (inp[7]) ? node364 : node357;
												assign node357 = (inp[13]) ? 4'b0101 : node358;
													assign node358 = (inp[2]) ? node360 : 4'b0110;
														assign node360 = (inp[4]) ? 4'b0000 : 4'b0000;
												assign node364 = (inp[13]) ? 4'b0010 : node365;
													assign node365 = (inp[11]) ? 4'b0100 : 4'b0110;
										assign node369 = (inp[4]) ? node377 : node370;
											assign node370 = (inp[15]) ? node374 : node371;
												assign node371 = (inp[12]) ? 4'b0011 : 4'b0100;
												assign node374 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node377 = (inp[12]) ? node381 : node378;
												assign node378 = (inp[13]) ? 4'b0010 : 4'b0000;
												assign node381 = (inp[11]) ? 4'b0111 : node382;
													assign node382 = (inp[7]) ? 4'b0010 : node383;
														assign node383 = (inp[2]) ? 4'b0110 : 4'b0011;
						assign node388 = (inp[15]) ? node586 : node389;
							assign node389 = (inp[4]) ? node477 : node390;
								assign node390 = (inp[5]) ? node434 : node391;
									assign node391 = (inp[2]) ? node413 : node392;
										assign node392 = (inp[13]) ? node404 : node393;
											assign node393 = (inp[1]) ? node399 : node394;
												assign node394 = (inp[7]) ? node396 : 4'b0010;
													assign node396 = (inp[12]) ? 4'b0001 : 4'b0011;
												assign node399 = (inp[7]) ? 4'b0011 : node400;
													assign node400 = (inp[10]) ? 4'b0011 : 4'b0001;
											assign node404 = (inp[12]) ? node408 : node405;
												assign node405 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node408 = (inp[0]) ? 4'b0111 : node409;
													assign node409 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node413 = (inp[13]) ? node427 : node414;
											assign node414 = (inp[12]) ? node420 : node415;
												assign node415 = (inp[7]) ? node417 : 4'b0100;
													assign node417 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node420 = (inp[11]) ? 4'b0111 : node421;
													assign node421 = (inp[10]) ? node423 : 4'b0110;
														assign node423 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node427 = (inp[7]) ? node429 : 4'b0000;
												assign node429 = (inp[12]) ? node431 : 4'b0011;
													assign node431 = (inp[10]) ? 4'b0101 : 4'b0001;
									assign node434 = (inp[7]) ? node458 : node435;
										assign node435 = (inp[12]) ? node445 : node436;
											assign node436 = (inp[13]) ? node442 : node437;
												assign node437 = (inp[10]) ? 4'b0100 : node438;
													assign node438 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node442 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node445 = (inp[1]) ? node449 : node446;
												assign node446 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node449 = (inp[0]) ? node453 : node450;
													assign node450 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node453 = (inp[2]) ? 4'b0110 : node454;
														assign node454 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node458 = (inp[12]) ? node470 : node459;
											assign node459 = (inp[1]) ? node467 : node460;
												assign node460 = (inp[13]) ? 4'b0111 : node461;
													assign node461 = (inp[2]) ? 4'b0111 : node462;
														assign node462 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node467 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node470 = (inp[10]) ? node472 : 4'b0101;
												assign node472 = (inp[13]) ? 4'b0001 : node473;
													assign node473 = (inp[2]) ? 4'b0000 : 4'b0100;
								assign node477 = (inp[0]) ? node535 : node478;
									assign node478 = (inp[11]) ? node508 : node479;
										assign node479 = (inp[2]) ? node491 : node480;
											assign node480 = (inp[7]) ? node484 : node481;
												assign node481 = (inp[13]) ? 4'b0010 : 4'b0000;
												assign node484 = (inp[12]) ? node486 : 4'b0010;
													assign node486 = (inp[13]) ? 4'b0101 : node487;
														assign node487 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node491 = (inp[5]) ? node499 : node492;
												assign node492 = (inp[1]) ? node494 : 4'b0101;
													assign node494 = (inp[12]) ? node496 : 4'b0111;
														assign node496 = (inp[7]) ? 4'b0101 : 4'b0111;
												assign node499 = (inp[1]) ? node503 : node500;
													assign node500 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node503 = (inp[7]) ? node505 : 4'b0111;
														assign node505 = (inp[13]) ? 4'b0111 : 4'b0011;
										assign node508 = (inp[5]) ? node522 : node509;
											assign node509 = (inp[10]) ? node517 : node510;
												assign node510 = (inp[2]) ? 4'b0001 : node511;
													assign node511 = (inp[1]) ? 4'b0111 : node512;
														assign node512 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node517 = (inp[1]) ? 4'b0101 : node518;
													assign node518 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node522 = (inp[2]) ? node526 : node523;
												assign node523 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node526 = (inp[13]) ? node532 : node527;
													assign node527 = (inp[10]) ? 4'b0100 : node528;
														assign node528 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node532 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node535 = (inp[2]) ? node555 : node536;
										assign node536 = (inp[10]) ? node538 : 4'b0111;
											assign node538 = (inp[5]) ? node546 : node539;
												assign node539 = (inp[7]) ? node543 : node540;
													assign node540 = (inp[11]) ? 4'b0111 : 4'b0011;
													assign node543 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node546 = (inp[7]) ? node552 : node547;
													assign node547 = (inp[12]) ? node549 : 4'b0001;
														assign node549 = (inp[11]) ? 4'b0011 : 4'b0111;
													assign node552 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node555 = (inp[10]) ? node573 : node556;
											assign node556 = (inp[7]) ? node568 : node557;
												assign node557 = (inp[12]) ? node563 : node558;
													assign node558 = (inp[11]) ? node560 : 4'b0001;
														assign node560 = (inp[1]) ? 4'b0000 : 4'b0101;
													assign node563 = (inp[13]) ? node565 : 4'b0011;
														assign node565 = (inp[5]) ? 4'b0011 : 4'b0110;
												assign node568 = (inp[12]) ? 4'b0001 : node569;
													assign node569 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node573 = (inp[13]) ? node581 : node574;
												assign node574 = (inp[1]) ? node576 : 4'b0111;
													assign node576 = (inp[5]) ? node578 : 4'b0101;
														assign node578 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node581 = (inp[5]) ? node583 : 4'b0000;
													assign node583 = (inp[1]) ? 4'b0001 : 4'b0000;
							assign node586 = (inp[7]) ? node670 : node587;
								assign node587 = (inp[4]) ? node627 : node588;
									assign node588 = (inp[12]) ? node616 : node589;
										assign node589 = (inp[11]) ? node607 : node590;
											assign node590 = (inp[2]) ? node598 : node591;
												assign node591 = (inp[5]) ? 4'b0101 : node592;
													assign node592 = (inp[10]) ? node594 : 4'b0100;
														assign node594 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node598 = (inp[13]) ? node604 : node599;
													assign node599 = (inp[10]) ? 4'b0101 : node600;
														assign node600 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node604 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node607 = (inp[2]) ? node609 : 4'b0001;
												assign node609 = (inp[0]) ? 4'b0100 : node610;
													assign node610 = (inp[13]) ? 4'b0001 : node611;
														assign node611 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node616 = (inp[13]) ? node622 : node617;
											assign node617 = (inp[10]) ? node619 : 4'b0110;
												assign node619 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node622 = (inp[11]) ? node624 : 4'b0011;
												assign node624 = (inp[0]) ? 4'b0011 : 4'b0110;
									assign node627 = (inp[12]) ? node649 : node628;
										assign node628 = (inp[13]) ? node634 : node629;
											assign node629 = (inp[2]) ? 4'b0010 : node630;
												assign node630 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node634 = (inp[2]) ? node640 : node635;
												assign node635 = (inp[10]) ? node637 : 4'b0110;
													assign node637 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node640 = (inp[1]) ? node642 : 4'b0111;
													assign node642 = (inp[11]) ? node646 : node643;
														assign node643 = (inp[5]) ? 4'b0110 : 4'b0110;
														assign node646 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node649 = (inp[5]) ? node655 : node650;
											assign node650 = (inp[13]) ? 4'b0001 : node651;
												assign node651 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node655 = (inp[13]) ? node661 : node656;
												assign node656 = (inp[1]) ? 4'b0100 : node657;
													assign node657 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node661 = (inp[2]) ? node667 : node662;
													assign node662 = (inp[1]) ? 4'b0001 : node663;
														assign node663 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node667 = (inp[1]) ? 4'b0100 : 4'b0000;
								assign node670 = (inp[0]) ? node724 : node671;
									assign node671 = (inp[4]) ? node699 : node672;
										assign node672 = (inp[12]) ? node686 : node673;
											assign node673 = (inp[10]) ? node679 : node674;
												assign node674 = (inp[13]) ? node676 : 4'b0010;
													assign node676 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node679 = (inp[1]) ? node681 : 4'b0111;
													assign node681 = (inp[13]) ? 4'b0010 : node682;
														assign node682 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node686 = (inp[10]) ? node692 : node687;
												assign node687 = (inp[2]) ? 4'b0000 : node688;
													assign node688 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node692 = (inp[11]) ? node694 : 4'b0001;
													assign node694 = (inp[13]) ? 4'b0001 : node695;
														assign node695 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node699 = (inp[12]) ? node711 : node700;
											assign node700 = (inp[13]) ? node702 : 4'b0000;
												assign node702 = (inp[5]) ? node708 : node703;
													assign node703 = (inp[2]) ? node705 : 4'b0100;
														assign node705 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node708 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node711 = (inp[11]) ? node717 : node712;
												assign node712 = (inp[1]) ? 4'b0010 : node713;
													assign node713 = (inp[5]) ? 4'b0111 : 4'b0010;
												assign node717 = (inp[2]) ? 4'b0011 : node718;
													assign node718 = (inp[10]) ? 4'b0111 : node719;
														assign node719 = (inp[5]) ? 4'b0111 : 4'b0011;
									assign node724 = (inp[1]) ? node750 : node725;
										assign node725 = (inp[11]) ? node735 : node726;
											assign node726 = (inp[12]) ? node732 : node727;
												assign node727 = (inp[4]) ? node729 : 4'b0110;
													assign node729 = (inp[10]) ? 4'b0101 : 4'b0000;
												assign node732 = (inp[4]) ? 4'b0111 : 4'b0001;
											assign node735 = (inp[5]) ? node743 : node736;
												assign node736 = (inp[2]) ? node738 : 4'b0001;
													assign node738 = (inp[12]) ? node740 : 4'b0010;
														assign node740 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node743 = (inp[10]) ? 4'b0011 : node744;
													assign node744 = (inp[12]) ? 4'b0110 : node745;
														assign node745 = (inp[4]) ? 4'b0101 : 4'b0011;
										assign node750 = (inp[13]) ? node752 : 4'b0011;
											assign node752 = (inp[4]) ? node754 : 4'b0111;
												assign node754 = (inp[11]) ? 4'b0110 : 4'b0111;
					assign node757 = (inp[7]) ? node1121 : node758;
						assign node758 = (inp[12]) ? node914 : node759;
							assign node759 = (inp[4]) ? node833 : node760;
								assign node760 = (inp[15]) ? node802 : node761;
									assign node761 = (inp[1]) ? node777 : node762;
										assign node762 = (inp[13]) ? node770 : node763;
											assign node763 = (inp[9]) ? node767 : node764;
												assign node764 = (inp[11]) ? 4'b1000 : 4'b1100;
												assign node767 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node770 = (inp[10]) ? node772 : 4'b1101;
												assign node772 = (inp[11]) ? node774 : 4'b1101;
													assign node774 = (inp[0]) ? 4'b1101 : 4'b1001;
										assign node777 = (inp[9]) ? node793 : node778;
											assign node778 = (inp[5]) ? node784 : node779;
												assign node779 = (inp[13]) ? node781 : 4'b1100;
													assign node781 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node784 = (inp[11]) ? node790 : node785;
													assign node785 = (inp[0]) ? 4'b1101 : node786;
														assign node786 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node790 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node793 = (inp[11]) ? node795 : 4'b1000;
												assign node795 = (inp[5]) ? node799 : node796;
													assign node796 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node799 = (inp[10]) ? 4'b1100 : 4'b1101;
									assign node802 = (inp[1]) ? node822 : node803;
										assign node803 = (inp[11]) ? node817 : node804;
											assign node804 = (inp[0]) ? node808 : node805;
												assign node805 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node808 = (inp[2]) ? node812 : node809;
													assign node809 = (inp[10]) ? 4'b1010 : 4'b1111;
													assign node812 = (inp[13]) ? 4'b1110 : node813;
														assign node813 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node817 = (inp[10]) ? node819 : 4'b1010;
												assign node819 = (inp[9]) ? 4'b1110 : 4'b1010;
										assign node822 = (inp[5]) ? node824 : 4'b1010;
											assign node824 = (inp[2]) ? node826 : 4'b1110;
												assign node826 = (inp[13]) ? node828 : 4'b1111;
													assign node828 = (inp[0]) ? 4'b1011 : node829;
														assign node829 = (inp[11]) ? 4'b1011 : 4'b1010;
								assign node833 = (inp[5]) ? node877 : node834;
									assign node834 = (inp[0]) ? node860 : node835;
										assign node835 = (inp[11]) ? node849 : node836;
											assign node836 = (inp[15]) ? node844 : node837;
												assign node837 = (inp[10]) ? node839 : 4'b1101;
													assign node839 = (inp[2]) ? 4'b1101 : node840;
														assign node840 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node844 = (inp[2]) ? node846 : 4'b1001;
													assign node846 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node849 = (inp[10]) ? node855 : node850;
												assign node850 = (inp[1]) ? 4'b1101 : node851;
													assign node851 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node855 = (inp[15]) ? node857 : 4'b1000;
													assign node857 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node860 = (inp[13]) ? node866 : node861;
											assign node861 = (inp[11]) ? node863 : 4'b1001;
												assign node863 = (inp[15]) ? 4'b1101 : 4'b1001;
											assign node866 = (inp[11]) ? 4'b1001 : node867;
												assign node867 = (inp[1]) ? 4'b1000 : node868;
													assign node868 = (inp[9]) ? node872 : node869;
														assign node869 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node872 = (inp[2]) ? 4'b1000 : 4'b1001;
									assign node877 = (inp[10]) ? node907 : node878;
										assign node878 = (inp[15]) ? node888 : node879;
											assign node879 = (inp[11]) ? 4'b1001 : node880;
												assign node880 = (inp[2]) ? node882 : 4'b1100;
													assign node882 = (inp[13]) ? 4'b1101 : node883;
														assign node883 = (inp[1]) ? 4'b1101 : 4'b1001;
											assign node888 = (inp[9]) ? node898 : node889;
												assign node889 = (inp[2]) ? node893 : node890;
													assign node890 = (inp[13]) ? 4'b1100 : 4'b1001;
													assign node893 = (inp[13]) ? node895 : 4'b1100;
														assign node895 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node898 = (inp[0]) ? 4'b1100 : node899;
													assign node899 = (inp[1]) ? node903 : node900;
														assign node900 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node903 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node907 = (inp[9]) ? node909 : 4'b1101;
											assign node909 = (inp[13]) ? node911 : 4'b1100;
												assign node911 = (inp[15]) ? 4'b1100 : 4'b1000;
							assign node914 = (inp[4]) ? node1012 : node915;
								assign node915 = (inp[15]) ? node951 : node916;
									assign node916 = (inp[2]) ? node942 : node917;
										assign node917 = (inp[13]) ? node931 : node918;
											assign node918 = (inp[5]) ? node924 : node919;
												assign node919 = (inp[1]) ? node921 : 4'b1010;
													assign node921 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node924 = (inp[10]) ? node926 : 4'b1011;
													assign node926 = (inp[9]) ? node928 : 4'b1011;
														assign node928 = (inp[0]) ? 4'b1010 : 4'b1010;
											assign node931 = (inp[11]) ? 4'b1110 : node932;
												assign node932 = (inp[1]) ? node938 : node933;
													assign node933 = (inp[0]) ? 4'b1111 : node934;
														assign node934 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node938 = (inp[0]) ? 4'b1110 : 4'b1011;
										assign node942 = (inp[13]) ? 4'b1011 : node943;
											assign node943 = (inp[1]) ? node947 : node944;
												assign node944 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node947 = (inp[0]) ? 4'b1011 : 4'b1010;
									assign node951 = (inp[10]) ? node981 : node952;
										assign node952 = (inp[13]) ? node972 : node953;
											assign node953 = (inp[2]) ? node961 : node954;
												assign node954 = (inp[5]) ? node956 : 4'b1100;
													assign node956 = (inp[11]) ? 4'b1101 : node957;
														assign node957 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node961 = (inp[9]) ? node967 : node962;
													assign node962 = (inp[11]) ? node964 : 4'b1001;
														assign node964 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node967 = (inp[0]) ? 4'b1000 : node968;
														assign node968 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node972 = (inp[2]) ? node974 : 4'b1001;
												assign node974 = (inp[0]) ? 4'b1101 : node975;
													assign node975 = (inp[5]) ? 4'b1000 : node976;
														assign node976 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node981 = (inp[0]) ? node1001 : node982;
											assign node982 = (inp[5]) ? node990 : node983;
												assign node983 = (inp[11]) ? node985 : 4'b1101;
													assign node985 = (inp[9]) ? 4'b1001 : node986;
														assign node986 = (inp[13]) ? 4'b1100 : 4'b1001;
												assign node990 = (inp[2]) ? node996 : node991;
													assign node991 = (inp[9]) ? node993 : 4'b1100;
														assign node993 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node996 = (inp[1]) ? node998 : 4'b1000;
														assign node998 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node1001 = (inp[9]) ? node1007 : node1002;
												assign node1002 = (inp[5]) ? node1004 : 4'b1000;
													assign node1004 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node1007 = (inp[13]) ? node1009 : 4'b1100;
													assign node1009 = (inp[1]) ? 4'b1100 : 4'b1001;
								assign node1012 = (inp[11]) ? node1082 : node1013;
									assign node1013 = (inp[1]) ? node1043 : node1014;
										assign node1014 = (inp[5]) ? node1026 : node1015;
											assign node1015 = (inp[2]) ? node1019 : node1016;
												assign node1016 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node1019 = (inp[10]) ? node1021 : 4'b1011;
													assign node1021 = (inp[9]) ? node1023 : 4'b1010;
														assign node1023 = (inp[0]) ? 4'b1010 : 4'b1110;
											assign node1026 = (inp[0]) ? node1034 : node1027;
												assign node1027 = (inp[9]) ? node1029 : 4'b1011;
													assign node1029 = (inp[13]) ? 4'b1010 : node1030;
														assign node1030 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node1034 = (inp[15]) ? node1036 : 4'b1011;
													assign node1036 = (inp[2]) ? node1040 : node1037;
														assign node1037 = (inp[9]) ? 4'b1010 : 4'b1010;
														assign node1040 = (inp[13]) ? 4'b1010 : 4'b1110;
										assign node1043 = (inp[2]) ? node1063 : node1044;
											assign node1044 = (inp[13]) ? node1052 : node1045;
												assign node1045 = (inp[15]) ? node1049 : node1046;
													assign node1046 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node1049 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node1052 = (inp[10]) ? node1058 : node1053;
													assign node1053 = (inp[9]) ? 4'b1010 : node1054;
														assign node1054 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node1058 = (inp[0]) ? node1060 : 4'b1111;
														assign node1060 = (inp[15]) ? 4'b1111 : 4'b1010;
											assign node1063 = (inp[15]) ? node1071 : node1064;
												assign node1064 = (inp[13]) ? node1068 : node1065;
													assign node1065 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node1068 = (inp[5]) ? 4'b1111 : 4'b1011;
												assign node1071 = (inp[10]) ? node1079 : node1072;
													assign node1072 = (inp[9]) ? node1076 : node1073;
														assign node1073 = (inp[0]) ? 4'b1111 : 4'b1010;
														assign node1076 = (inp[5]) ? 4'b1011 : 4'b1011;
													assign node1079 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node1082 = (inp[2]) ? node1096 : node1083;
										assign node1083 = (inp[10]) ? node1091 : node1084;
											assign node1084 = (inp[13]) ? node1088 : node1085;
												assign node1085 = (inp[5]) ? 4'b1010 : 4'b1111;
												assign node1088 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node1091 = (inp[13]) ? node1093 : 4'b1011;
												assign node1093 = (inp[1]) ? 4'b1111 : 4'b1011;
										assign node1096 = (inp[9]) ? node1110 : node1097;
											assign node1097 = (inp[1]) ? 4'b1110 : node1098;
												assign node1098 = (inp[5]) ? node1106 : node1099;
													assign node1099 = (inp[0]) ? node1103 : node1100;
														assign node1100 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node1103 = (inp[15]) ? 4'b1011 : 4'b1011;
													assign node1106 = (inp[15]) ? 4'b1110 : 4'b1111;
											assign node1110 = (inp[13]) ? 4'b1110 : node1111;
												assign node1111 = (inp[10]) ? node1115 : node1112;
													assign node1112 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node1115 = (inp[15]) ? 4'b1110 : node1116;
														assign node1116 = (inp[0]) ? 4'b1010 : 4'b1110;
						assign node1121 = (inp[12]) ? node1303 : node1122;
							assign node1122 = (inp[15]) ? node1224 : node1123;
								assign node1123 = (inp[10]) ? node1183 : node1124;
									assign node1124 = (inp[9]) ? node1160 : node1125;
										assign node1125 = (inp[11]) ? node1143 : node1126;
											assign node1126 = (inp[0]) ? node1136 : node1127;
												assign node1127 = (inp[1]) ? node1129 : 4'b1011;
													assign node1129 = (inp[2]) ? node1133 : node1130;
														assign node1130 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node1133 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node1136 = (inp[13]) ? 4'b1010 : node1137;
													assign node1137 = (inp[5]) ? 4'b1110 : node1138;
														assign node1138 = (inp[2]) ? 4'b1110 : 4'b1010;
											assign node1143 = (inp[2]) ? node1151 : node1144;
												assign node1144 = (inp[0]) ? node1148 : node1145;
													assign node1145 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node1148 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node1151 = (inp[13]) ? 4'b1011 : node1152;
													assign node1152 = (inp[1]) ? node1156 : node1153;
														assign node1153 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node1156 = (inp[4]) ? 4'b1111 : 4'b1110;
										assign node1160 = (inp[11]) ? node1170 : node1161;
											assign node1161 = (inp[5]) ? node1163 : 4'b1111;
												assign node1163 = (inp[4]) ? 4'b1011 : node1164;
													assign node1164 = (inp[2]) ? node1166 : 4'b1110;
														assign node1166 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node1170 = (inp[13]) ? node1172 : 4'b1111;
												assign node1172 = (inp[4]) ? node1180 : node1173;
													assign node1173 = (inp[5]) ? node1177 : node1174;
														assign node1174 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node1177 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node1180 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node1183 = (inp[9]) ? node1205 : node1184;
										assign node1184 = (inp[2]) ? node1192 : node1185;
											assign node1185 = (inp[0]) ? node1189 : node1186;
												assign node1186 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node1189 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node1192 = (inp[0]) ? node1200 : node1193;
												assign node1193 = (inp[4]) ? 4'b1110 : node1194;
													assign node1194 = (inp[1]) ? node1196 : 4'b1111;
														assign node1196 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node1200 = (inp[1]) ? 4'b1110 : node1201;
													assign node1201 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node1205 = (inp[13]) ? node1217 : node1206;
											assign node1206 = (inp[5]) ? node1208 : 4'b1110;
												assign node1208 = (inp[2]) ? node1214 : node1209;
													assign node1209 = (inp[4]) ? 4'b1010 : node1210;
														assign node1210 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node1214 = (inp[1]) ? 4'b1111 : 4'b1010;
											assign node1217 = (inp[5]) ? node1219 : 4'b1011;
												assign node1219 = (inp[11]) ? 4'b1010 : node1220;
													assign node1220 = (inp[1]) ? 4'b1110 : 4'b1010;
								assign node1224 = (inp[4]) ? node1268 : node1225;
									assign node1225 = (inp[10]) ? node1247 : node1226;
										assign node1226 = (inp[2]) ? node1236 : node1227;
											assign node1227 = (inp[1]) ? node1229 : 4'b1001;
												assign node1229 = (inp[0]) ? node1231 : 4'b1100;
													assign node1231 = (inp[11]) ? 4'b1101 : node1232;
														assign node1232 = (inp[5]) ? 4'b1001 : 4'b1101;
											assign node1236 = (inp[5]) ? node1240 : node1237;
												assign node1237 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node1240 = (inp[0]) ? node1244 : node1241;
													assign node1241 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node1244 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node1247 = (inp[0]) ? node1257 : node1248;
											assign node1248 = (inp[1]) ? node1254 : node1249;
												assign node1249 = (inp[5]) ? node1251 : 4'b1101;
													assign node1251 = (inp[2]) ? 4'b1101 : 4'b1000;
												assign node1254 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node1257 = (inp[1]) ? node1263 : node1258;
												assign node1258 = (inp[2]) ? node1260 : 4'b1000;
													assign node1260 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node1263 = (inp[5]) ? 4'b1101 : node1264;
													assign node1264 = (inp[2]) ? 4'b1000 : 4'b1101;
									assign node1268 = (inp[9]) ? node1286 : node1269;
										assign node1269 = (inp[0]) ? node1275 : node1270;
											assign node1270 = (inp[11]) ? 4'b1110 : node1271;
												assign node1271 = (inp[5]) ? 4'b1010 : 4'b1110;
											assign node1275 = (inp[10]) ? node1281 : node1276;
												assign node1276 = (inp[13]) ? node1278 : 4'b1010;
													assign node1278 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node1281 = (inp[11]) ? 4'b1111 : node1282;
													assign node1282 = (inp[1]) ? 4'b1110 : 4'b1010;
										assign node1286 = (inp[11]) ? node1300 : node1287;
											assign node1287 = (inp[2]) ? node1297 : node1288;
												assign node1288 = (inp[1]) ? node1292 : node1289;
													assign node1289 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node1292 = (inp[0]) ? 4'b1011 : node1293;
														assign node1293 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node1297 = (inp[13]) ? 4'b1011 : 4'b1111;
											assign node1300 = (inp[2]) ? 4'b1010 : 4'b1110;
							assign node1303 = (inp[15]) ? node1401 : node1304;
								assign node1304 = (inp[13]) ? node1362 : node1305;
									assign node1305 = (inp[0]) ? node1333 : node1306;
										assign node1306 = (inp[11]) ? node1324 : node1307;
											assign node1307 = (inp[1]) ? node1311 : node1308;
												assign node1308 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node1311 = (inp[10]) ? node1319 : node1312;
													assign node1312 = (inp[2]) ? node1316 : node1313;
														assign node1313 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node1316 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node1319 = (inp[4]) ? node1321 : 4'b1101;
														assign node1321 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node1324 = (inp[9]) ? node1328 : node1325;
												assign node1325 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node1328 = (inp[2]) ? 4'b1000 : node1329;
													assign node1329 = (inp[1]) ? 4'b1100 : 4'b1101;
										assign node1333 = (inp[5]) ? node1345 : node1334;
											assign node1334 = (inp[10]) ? node1342 : node1335;
												assign node1335 = (inp[9]) ? node1337 : 4'b1101;
													assign node1337 = (inp[4]) ? node1339 : 4'b1100;
														assign node1339 = (inp[11]) ? 4'b1001 : 4'b1100;
												assign node1342 = (inp[9]) ? 4'b1101 : 4'b1001;
											assign node1345 = (inp[11]) ? node1349 : node1346;
												assign node1346 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node1349 = (inp[4]) ? node1355 : node1350;
													assign node1350 = (inp[1]) ? 4'b1000 : node1351;
														assign node1351 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node1355 = (inp[2]) ? node1359 : node1356;
														assign node1356 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node1359 = (inp[1]) ? 4'b1101 : 4'b1000;
									assign node1362 = (inp[10]) ? node1388 : node1363;
										assign node1363 = (inp[0]) ? node1377 : node1364;
											assign node1364 = (inp[4]) ? node1374 : node1365;
												assign node1365 = (inp[2]) ? node1367 : 4'b1100;
													assign node1367 = (inp[9]) ? node1371 : node1368;
														assign node1368 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node1371 = (inp[11]) ? 4'b1100 : 4'b1100;
												assign node1374 = (inp[1]) ? 4'b1000 : 4'b1101;
											assign node1377 = (inp[11]) ? 4'b1100 : node1378;
												assign node1378 = (inp[5]) ? node1380 : 4'b1000;
													assign node1380 = (inp[9]) ? node1384 : node1381;
														assign node1381 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node1384 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node1388 = (inp[4]) ? node1396 : node1389;
											assign node1389 = (inp[1]) ? node1391 : 4'b1000;
												assign node1391 = (inp[2]) ? 4'b1101 : node1392;
													assign node1392 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node1396 = (inp[2]) ? 4'b1000 : node1397;
												assign node1397 = (inp[1]) ? 4'b1100 : 4'b1101;
								assign node1401 = (inp[4]) ? node1453 : node1402;
									assign node1402 = (inp[9]) ? node1428 : node1403;
										assign node1403 = (inp[0]) ? node1417 : node1404;
											assign node1404 = (inp[13]) ? node1408 : node1405;
												assign node1405 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node1408 = (inp[2]) ? node1412 : node1409;
													assign node1409 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node1412 = (inp[1]) ? node1414 : 4'b1111;
														assign node1414 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node1417 = (inp[1]) ? node1421 : node1418;
												assign node1418 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node1421 = (inp[2]) ? node1425 : node1422;
													assign node1422 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node1425 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node1428 = (inp[2]) ? node1442 : node1429;
											assign node1429 = (inp[1]) ? node1437 : node1430;
												assign node1430 = (inp[11]) ? 4'b1111 : node1431;
													assign node1431 = (inp[10]) ? node1433 : 4'b1010;
														assign node1433 = (inp[0]) ? 4'b1011 : 4'b1110;
												assign node1437 = (inp[10]) ? 4'b1010 : node1438;
													assign node1438 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node1442 = (inp[10]) ? node1444 : 4'b1010;
												assign node1444 = (inp[13]) ? node1450 : node1445;
													assign node1445 = (inp[11]) ? node1447 : 4'b1111;
														assign node1447 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node1450 = (inp[0]) ? 4'b1110 : 4'b1010;
									assign node1453 = (inp[2]) ? node1473 : node1454;
										assign node1454 = (inp[13]) ? node1460 : node1455;
											assign node1455 = (inp[1]) ? 4'b1000 : node1456;
												assign node1456 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node1460 = (inp[0]) ? node1466 : node1461;
												assign node1461 = (inp[10]) ? 4'b1101 : node1462;
													assign node1462 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node1466 = (inp[1]) ? node1470 : node1467;
													assign node1467 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node1470 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node1473 = (inp[13]) ? node1487 : node1474;
											assign node1474 = (inp[10]) ? 4'b1100 : node1475;
												assign node1475 = (inp[0]) ? node1481 : node1476;
													assign node1476 = (inp[5]) ? 4'b1101 : node1477;
														assign node1477 = (inp[11]) ? 4'b1100 : 4'b1100;
													assign node1481 = (inp[1]) ? 4'b1101 : node1482;
														assign node1482 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node1487 = (inp[0]) ? node1489 : 4'b1000;
												assign node1489 = (inp[10]) ? 4'b1100 : 4'b1001;
				assign node1492 = (inp[9]) ? node2256 : node1493;
					assign node1493 = (inp[14]) ? node1893 : node1494;
						assign node1494 = (inp[2]) ? node1694 : node1495;
							assign node1495 = (inp[1]) ? node1593 : node1496;
								assign node1496 = (inp[0]) ? node1538 : node1497;
									assign node1497 = (inp[10]) ? node1513 : node1498;
										assign node1498 = (inp[11]) ? node1508 : node1499;
											assign node1499 = (inp[15]) ? node1501 : 4'b1010;
												assign node1501 = (inp[4]) ? 4'b1001 : node1502;
													assign node1502 = (inp[12]) ? node1504 : 4'b1000;
														assign node1504 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node1508 = (inp[7]) ? node1510 : 4'b1000;
												assign node1510 = (inp[5]) ? 4'b1010 : 4'b1001;
										assign node1513 = (inp[15]) ? node1527 : node1514;
											assign node1514 = (inp[5]) ? node1520 : node1515;
												assign node1515 = (inp[12]) ? 4'b1101 : node1516;
													assign node1516 = (inp[11]) ? 4'b1011 : 4'b1001;
												assign node1520 = (inp[7]) ? 4'b1111 : node1521;
													assign node1521 = (inp[11]) ? 4'b1000 : node1522;
														assign node1522 = (inp[12]) ? 4'b1000 : 4'b1010;
											assign node1527 = (inp[5]) ? node1529 : 4'b1011;
												assign node1529 = (inp[7]) ? node1533 : node1530;
													assign node1530 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node1533 = (inp[12]) ? node1535 : 4'b1000;
														assign node1535 = (inp[4]) ? 4'b1000 : 4'b1011;
									assign node1538 = (inp[7]) ? node1564 : node1539;
										assign node1539 = (inp[5]) ? node1549 : node1540;
											assign node1540 = (inp[12]) ? node1544 : node1541;
												assign node1541 = (inp[4]) ? 4'b1011 : 4'b1000;
												assign node1544 = (inp[15]) ? node1546 : 4'b1011;
													assign node1546 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node1549 = (inp[12]) ? node1557 : node1550;
												assign node1550 = (inp[4]) ? node1552 : 4'b1001;
													assign node1552 = (inp[15]) ? 4'b1111 : node1553;
														assign node1553 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node1557 = (inp[11]) ? node1559 : 4'b1000;
													assign node1559 = (inp[15]) ? 4'b1001 : node1560;
														assign node1560 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node1564 = (inp[11]) ? node1578 : node1565;
											assign node1565 = (inp[12]) ? node1569 : node1566;
												assign node1566 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node1569 = (inp[5]) ? node1573 : node1570;
													assign node1570 = (inp[4]) ? 4'b1101 : 4'b1110;
													assign node1573 = (inp[15]) ? 4'b1000 : node1574;
														assign node1574 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node1578 = (inp[12]) ? node1590 : node1579;
												assign node1579 = (inp[4]) ? node1587 : node1580;
													assign node1580 = (inp[13]) ? node1584 : node1581;
														assign node1581 = (inp[15]) ? 4'b1000 : 4'b1101;
														assign node1584 = (inp[15]) ? 4'b1101 : 4'b1000;
													assign node1587 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node1590 = (inp[13]) ? 4'b1011 : 4'b1111;
								assign node1593 = (inp[13]) ? node1637 : node1594;
									assign node1594 = (inp[12]) ? node1614 : node1595;
										assign node1595 = (inp[4]) ? node1607 : node1596;
											assign node1596 = (inp[7]) ? node1602 : node1597;
												assign node1597 = (inp[0]) ? 4'b1101 : node1598;
													assign node1598 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node1602 = (inp[15]) ? node1604 : 4'b1001;
													assign node1604 = (inp[0]) ? 4'b1001 : 4'b1101;
											assign node1607 = (inp[5]) ? node1609 : 4'b1111;
												assign node1609 = (inp[7]) ? 4'b1010 : node1610;
													assign node1610 = (inp[15]) ? 4'b1011 : 4'b1111;
										assign node1614 = (inp[4]) ? node1624 : node1615;
											assign node1615 = (inp[5]) ? node1619 : node1616;
												assign node1616 = (inp[7]) ? 4'b1011 : 4'b1111;
												assign node1619 = (inp[0]) ? 4'b1110 : node1620;
													assign node1620 = (inp[7]) ? 4'b1010 : 4'b1110;
											assign node1624 = (inp[5]) ? node1634 : node1625;
												assign node1625 = (inp[10]) ? node1629 : node1626;
													assign node1626 = (inp[11]) ? 4'b1001 : 4'b1100;
													assign node1629 = (inp[7]) ? 4'b1100 : node1630;
														assign node1630 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node1634 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node1637 = (inp[5]) ? node1665 : node1638;
										assign node1638 = (inp[11]) ? node1654 : node1639;
											assign node1639 = (inp[0]) ? node1647 : node1640;
												assign node1640 = (inp[10]) ? 4'b1111 : node1641;
													assign node1641 = (inp[12]) ? 4'b1111 : node1642;
														assign node1642 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node1647 = (inp[12]) ? node1651 : node1648;
													assign node1648 = (inp[7]) ? 4'b1110 : 4'b1100;
													assign node1651 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node1654 = (inp[15]) ? node1658 : node1655;
												assign node1655 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node1658 = (inp[0]) ? 4'b1110 : node1659;
													assign node1659 = (inp[4]) ? node1661 : 4'b1001;
														assign node1661 = (inp[7]) ? 4'b1111 : 4'b1101;
										assign node1665 = (inp[11]) ? node1683 : node1666;
											assign node1666 = (inp[12]) ? node1676 : node1667;
												assign node1667 = (inp[4]) ? node1669 : 4'b1001;
													assign node1669 = (inp[7]) ? node1673 : node1670;
														assign node1670 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node1673 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node1676 = (inp[4]) ? 4'b1101 : node1677;
													assign node1677 = (inp[7]) ? 4'b1111 : node1678;
														assign node1678 = (inp[15]) ? 4'b1110 : 4'b1111;
											assign node1683 = (inp[0]) ? node1691 : node1684;
												assign node1684 = (inp[7]) ? 4'b1010 : node1685;
													assign node1685 = (inp[4]) ? 4'b1010 : node1686;
														assign node1686 = (inp[12]) ? 4'b1110 : 4'b1100;
												assign node1691 = (inp[7]) ? 4'b1100 : 4'b1110;
							assign node1694 = (inp[1]) ? node1790 : node1695;
								assign node1695 = (inp[0]) ? node1733 : node1696;
									assign node1696 = (inp[7]) ? node1708 : node1697;
										assign node1697 = (inp[12]) ? 4'b1110 : node1698;
											assign node1698 = (inp[4]) ? node1702 : node1699;
												assign node1699 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node1702 = (inp[10]) ? 4'b1110 : node1703;
													assign node1703 = (inp[13]) ? 4'b1110 : 4'b1111;
										assign node1708 = (inp[4]) ? node1722 : node1709;
											assign node1709 = (inp[12]) ? node1715 : node1710;
												assign node1710 = (inp[15]) ? node1712 : 4'b1101;
													assign node1712 = (inp[13]) ? 4'b1101 : 4'b1000;
												assign node1715 = (inp[10]) ? node1717 : 4'b1110;
													assign node1717 = (inp[11]) ? 4'b1011 : node1718;
														assign node1718 = (inp[5]) ? 4'b1110 : 4'b1011;
											assign node1722 = (inp[12]) ? node1726 : node1723;
												assign node1723 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node1726 = (inp[15]) ? 4'b1100 : node1727;
													assign node1727 = (inp[10]) ? 4'b1101 : node1728;
														assign node1728 = (inp[5]) ? 4'b1100 : 4'b1100;
									assign node1733 = (inp[5]) ? node1769 : node1734;
										assign node1734 = (inp[15]) ? node1752 : node1735;
											assign node1735 = (inp[10]) ? node1743 : node1736;
												assign node1736 = (inp[13]) ? node1740 : node1737;
													assign node1737 = (inp[4]) ? 4'b1000 : 4'b1111;
													assign node1740 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node1743 = (inp[11]) ? node1747 : node1744;
													assign node1744 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node1747 = (inp[4]) ? 4'b1111 : node1748;
														assign node1748 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node1752 = (inp[7]) ? node1756 : node1753;
												assign node1753 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node1756 = (inp[4]) ? node1764 : node1757;
													assign node1757 = (inp[12]) ? node1761 : node1758;
														assign node1758 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node1761 = (inp[10]) ? 4'b1010 : 4'b1010;
													assign node1764 = (inp[11]) ? 4'b1000 : node1765;
														assign node1765 = (inp[10]) ? 4'b1111 : 4'b1110;
										assign node1769 = (inp[11]) ? node1779 : node1770;
											assign node1770 = (inp[7]) ? node1776 : node1771;
												assign node1771 = (inp[12]) ? node1773 : 4'b1110;
													assign node1773 = (inp[4]) ? 4'b1101 : 4'b1111;
												assign node1776 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node1779 = (inp[4]) ? node1787 : node1780;
												assign node1780 = (inp[15]) ? node1782 : 4'b1011;
													assign node1782 = (inp[12]) ? node1784 : 4'b1101;
														assign node1784 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node1787 = (inp[7]) ? 4'b1111 : 4'b1101;
								assign node1790 = (inp[10]) ? node1834 : node1791;
									assign node1791 = (inp[13]) ? node1809 : node1792;
										assign node1792 = (inp[5]) ? node1804 : node1793;
											assign node1793 = (inp[7]) ? node1799 : node1794;
												assign node1794 = (inp[11]) ? node1796 : 4'b1001;
													assign node1796 = (inp[15]) ? 4'b1001 : 4'b1100;
												assign node1799 = (inp[15]) ? node1801 : 4'b1010;
													assign node1801 = (inp[12]) ? 4'b1111 : 4'b1101;
											assign node1804 = (inp[11]) ? node1806 : 4'b1000;
												assign node1806 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node1809 = (inp[0]) ? node1821 : node1810;
											assign node1810 = (inp[7]) ? node1816 : node1811;
												assign node1811 = (inp[11]) ? 4'b1010 : node1812;
													assign node1812 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node1816 = (inp[12]) ? node1818 : 4'b1100;
													assign node1818 = (inp[4]) ? 4'b1000 : 4'b1010;
											assign node1821 = (inp[15]) ? node1825 : node1822;
												assign node1822 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node1825 = (inp[11]) ? node1829 : node1826;
													assign node1826 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node1829 = (inp[5]) ? 4'b1011 : node1830;
														assign node1830 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node1834 = (inp[11]) ? node1860 : node1835;
										assign node1835 = (inp[13]) ? node1851 : node1836;
											assign node1836 = (inp[15]) ? node1844 : node1837;
												assign node1837 = (inp[0]) ? node1839 : 4'b1010;
													assign node1839 = (inp[7]) ? node1841 : 4'b1011;
														assign node1841 = (inp[4]) ? 4'b1111 : 4'b1101;
												assign node1844 = (inp[0]) ? 4'b1010 : node1845;
													assign node1845 = (inp[5]) ? node1847 : 4'b1101;
														assign node1847 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node1851 = (inp[7]) ? node1855 : node1852;
												assign node1852 = (inp[12]) ? 4'b1001 : 4'b1111;
												assign node1855 = (inp[0]) ? 4'b1100 : node1856;
													assign node1856 = (inp[4]) ? 4'b1100 : 4'b1101;
										assign node1860 = (inp[15]) ? node1878 : node1861;
											assign node1861 = (inp[4]) ? node1865 : node1862;
												assign node1862 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node1865 = (inp[12]) ? node1873 : node1866;
													assign node1866 = (inp[5]) ? node1870 : node1867;
														assign node1867 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node1870 = (inp[0]) ? 4'b1010 : 4'b1110;
													assign node1873 = (inp[13]) ? 4'b1101 : node1874;
														assign node1874 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node1878 = (inp[13]) ? node1886 : node1879;
												assign node1879 = (inp[12]) ? node1883 : node1880;
													assign node1880 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node1883 = (inp[0]) ? 4'b1010 : 4'b1110;
												assign node1886 = (inp[0]) ? node1888 : 4'b1000;
													assign node1888 = (inp[7]) ? node1890 : 4'b1010;
														assign node1890 = (inp[12]) ? 4'b1110 : 4'b1010;
						assign node1893 = (inp[1]) ? node2079 : node1894;
							assign node1894 = (inp[2]) ? node1974 : node1895;
								assign node1895 = (inp[7]) ? node1937 : node1896;
									assign node1896 = (inp[4]) ? node1914 : node1897;
										assign node1897 = (inp[12]) ? node1905 : node1898;
											assign node1898 = (inp[13]) ? 4'b1001 : node1899;
												assign node1899 = (inp[15]) ? node1901 : 4'b1100;
													assign node1901 = (inp[5]) ? 4'b1001 : 4'b1000;
											assign node1905 = (inp[15]) ? node1911 : node1906;
												assign node1906 = (inp[13]) ? 4'b1011 : node1907;
													assign node1907 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node1911 = (inp[5]) ? 4'b1011 : 4'b1111;
										assign node1914 = (inp[12]) ? node1930 : node1915;
											assign node1915 = (inp[0]) ? node1923 : node1916;
												assign node1916 = (inp[15]) ? node1918 : 4'b1111;
													assign node1918 = (inp[5]) ? node1920 : 4'b1111;
														assign node1920 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node1923 = (inp[13]) ? node1927 : node1924;
													assign node1924 = (inp[11]) ? 4'b1010 : 4'b1110;
													assign node1927 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node1930 = (inp[11]) ? 4'b1101 : node1931;
												assign node1931 = (inp[15]) ? 4'b1100 : node1932;
													assign node1932 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node1937 = (inp[13]) ? node1953 : node1938;
										assign node1938 = (inp[11]) ? node1944 : node1939;
											assign node1939 = (inp[5]) ? node1941 : 4'b1011;
												assign node1941 = (inp[15]) ? 4'b1010 : 4'b1011;
											assign node1944 = (inp[5]) ? node1946 : 4'b1010;
												assign node1946 = (inp[12]) ? node1948 : 4'b1101;
													assign node1948 = (inp[10]) ? node1950 : 4'b1001;
														assign node1950 = (inp[15]) ? 4'b1010 : 4'b1011;
										assign node1953 = (inp[4]) ? node1963 : node1954;
											assign node1954 = (inp[12]) ? 4'b1110 : node1955;
												assign node1955 = (inp[11]) ? 4'b1000 : node1956;
													assign node1956 = (inp[10]) ? node1958 : 4'b1100;
														assign node1958 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node1963 = (inp[12]) ? node1971 : node1964;
												assign node1964 = (inp[11]) ? node1966 : 4'b1011;
													assign node1966 = (inp[5]) ? node1968 : 4'b1010;
														assign node1968 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node1971 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node1974 = (inp[7]) ? node2034 : node1975;
									assign node1975 = (inp[4]) ? node2001 : node1976;
										assign node1976 = (inp[12]) ? node1988 : node1977;
											assign node1977 = (inp[11]) ? node1983 : node1978;
												assign node1978 = (inp[5]) ? 4'b1101 : node1979;
													assign node1979 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node1983 = (inp[10]) ? 4'b1101 : node1984;
													assign node1984 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node1988 = (inp[13]) ? node1996 : node1989;
												assign node1989 = (inp[11]) ? 4'b1111 : node1990;
													assign node1990 = (inp[15]) ? 4'b1010 : node1991;
														assign node1991 = (inp[0]) ? 4'b1110 : 4'b1110;
												assign node1996 = (inp[10]) ? node1998 : 4'b1110;
													assign node1998 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node2001 = (inp[12]) ? node2021 : node2002;
											assign node2002 = (inp[0]) ? node2014 : node2003;
												assign node2003 = (inp[13]) ? node2009 : node2004;
													assign node2004 = (inp[5]) ? node2006 : 4'b1010;
														assign node2006 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node2009 = (inp[15]) ? node2011 : 4'b1110;
														assign node2011 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node2014 = (inp[13]) ? 4'b1011 : node2015;
													assign node2015 = (inp[15]) ? 4'b1110 : node2016;
														assign node2016 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node2021 = (inp[11]) ? 4'b1100 : node2022;
												assign node2022 = (inp[13]) ? node2026 : node2023;
													assign node2023 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node2026 = (inp[15]) ? node2030 : node2027;
														assign node2027 = (inp[0]) ? 4'b1100 : 4'b1000;
														assign node2030 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node2034 = (inp[15]) ? node2056 : node2035;
										assign node2035 = (inp[13]) ? node2045 : node2036;
											assign node2036 = (inp[10]) ? 4'b1111 : node2037;
												assign node2037 = (inp[5]) ? node2039 : 4'b1101;
													assign node2039 = (inp[4]) ? node2041 : 4'b1100;
														assign node2041 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node2045 = (inp[4]) ? node2053 : node2046;
												assign node2046 = (inp[10]) ? node2048 : 4'b1100;
													assign node2048 = (inp[5]) ? 4'b1101 : node2049;
														assign node2049 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node2053 = (inp[11]) ? 4'b1111 : 4'b1101;
										assign node2056 = (inp[5]) ? node2066 : node2057;
											assign node2057 = (inp[12]) ? node2059 : 4'b1110;
												assign node2059 = (inp[4]) ? node2061 : 4'b1110;
													assign node2061 = (inp[0]) ? 4'b1100 : node2062;
														assign node2062 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node2066 = (inp[12]) ? node2072 : node2067;
												assign node2067 = (inp[0]) ? 4'b1110 : node2068;
													assign node2068 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node2072 = (inp[4]) ? 4'b1101 : node2073;
													assign node2073 = (inp[0]) ? node2075 : 4'b1111;
														assign node2075 = (inp[11]) ? 4'b1111 : 4'b1110;
							assign node2079 = (inp[2]) ? node2157 : node2080;
								assign node2080 = (inp[7]) ? node2126 : node2081;
									assign node2081 = (inp[4]) ? node2105 : node2082;
										assign node2082 = (inp[12]) ? node2090 : node2083;
											assign node2083 = (inp[0]) ? node2085 : 4'b1100;
												assign node2085 = (inp[10]) ? node2087 : 4'b1101;
													assign node2087 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node2090 = (inp[10]) ? node2098 : node2091;
												assign node2091 = (inp[5]) ? node2093 : 4'b1011;
													assign node2093 = (inp[0]) ? 4'b1111 : node2094;
														assign node2094 = (inp[13]) ? 4'b1110 : 4'b1110;
												assign node2098 = (inp[11]) ? 4'b1110 : node2099;
													assign node2099 = (inp[5]) ? node2101 : 4'b1110;
														assign node2101 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node2105 = (inp[12]) ? node2115 : node2106;
											assign node2106 = (inp[11]) ? node2108 : 4'b1010;
												assign node2108 = (inp[10]) ? node2112 : node2109;
													assign node2109 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node2112 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node2115 = (inp[15]) ? node2123 : node2116;
												assign node2116 = (inp[5]) ? 4'b1001 : node2117;
													assign node2117 = (inp[0]) ? node2119 : 4'b1100;
														assign node2119 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node2123 = (inp[5]) ? 4'b1100 : 4'b1000;
									assign node2126 = (inp[12]) ? node2144 : node2127;
										assign node2127 = (inp[4]) ? node2139 : node2128;
											assign node2128 = (inp[15]) ? node2136 : node2129;
												assign node2129 = (inp[5]) ? 4'b1100 : node2130;
													assign node2130 = (inp[13]) ? node2132 : 4'b1101;
														assign node2132 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node2136 = (inp[5]) ? 4'b1001 : 4'b1100;
											assign node2139 = (inp[10]) ? 4'b1110 : node2140;
												assign node2140 = (inp[15]) ? 4'b1111 : 4'b1110;
										assign node2144 = (inp[4]) ? node2152 : node2145;
											assign node2145 = (inp[13]) ? node2147 : 4'b1111;
												assign node2147 = (inp[15]) ? node2149 : 4'b1111;
													assign node2149 = (inp[5]) ? 4'b1110 : 4'b1111;
											assign node2152 = (inp[13]) ? node2154 : 4'b1101;
												assign node2154 = (inp[15]) ? 4'b1100 : 4'b1101;
								assign node2157 = (inp[7]) ? node2213 : node2158;
									assign node2158 = (inp[10]) ? node2184 : node2159;
										assign node2159 = (inp[12]) ? node2175 : node2160;
											assign node2160 = (inp[4]) ? node2168 : node2161;
												assign node2161 = (inp[11]) ? node2165 : node2162;
													assign node2162 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node2165 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node2168 = (inp[13]) ? node2172 : node2169;
													assign node2169 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node2172 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node2175 = (inp[4]) ? node2181 : node2176;
												assign node2176 = (inp[5]) ? 4'b1011 : node2177;
													assign node2177 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node2181 = (inp[5]) ? 4'b1001 : 4'b1101;
										assign node2184 = (inp[11]) ? node2204 : node2185;
											assign node2185 = (inp[4]) ? node2197 : node2186;
												assign node2186 = (inp[12]) ? node2190 : node2187;
													assign node2187 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node2190 = (inp[0]) ? node2194 : node2191;
														assign node2191 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node2194 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node2197 = (inp[12]) ? node2199 : 4'b1011;
													assign node2199 = (inp[0]) ? 4'b1000 : node2200;
														assign node2200 = (inp[15]) ? 4'b1101 : 4'b1000;
											assign node2204 = (inp[0]) ? node2206 : 4'b1100;
												assign node2206 = (inp[4]) ? node2208 : 4'b1010;
													assign node2208 = (inp[5]) ? 4'b1110 : node2209;
														assign node2209 = (inp[15]) ? 4'b1110 : 4'b1011;
									assign node2213 = (inp[11]) ? node2233 : node2214;
										assign node2214 = (inp[12]) ? node2228 : node2215;
											assign node2215 = (inp[4]) ? node2221 : node2216;
												assign node2216 = (inp[5]) ? 4'b1001 : node2217;
													assign node2217 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node2221 = (inp[10]) ? 4'b1011 : node2222;
													assign node2222 = (inp[15]) ? node2224 : 4'b1010;
														assign node2224 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node2228 = (inp[4]) ? node2230 : 4'b1010;
												assign node2230 = (inp[5]) ? 4'b1000 : 4'b1001;
										assign node2233 = (inp[12]) ? node2243 : node2234;
											assign node2234 = (inp[4]) ? node2238 : node2235;
												assign node2235 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node2238 = (inp[5]) ? node2240 : 4'b1010;
													assign node2240 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node2243 = (inp[4]) ? node2253 : node2244;
												assign node2244 = (inp[0]) ? node2250 : node2245;
													assign node2245 = (inp[15]) ? 4'b1011 : node2246;
														assign node2246 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node2250 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node2253 = (inp[0]) ? 4'b1001 : 4'b1000;
					assign node2256 = (inp[5]) ? node2622 : node2257;
						assign node2257 = (inp[12]) ? node2457 : node2258;
							assign node2258 = (inp[4]) ? node2354 : node2259;
								assign node2259 = (inp[1]) ? node2307 : node2260;
									assign node2260 = (inp[2]) ? node2290 : node2261;
										assign node2261 = (inp[14]) ? node2277 : node2262;
											assign node2262 = (inp[15]) ? node2270 : node2263;
												assign node2263 = (inp[11]) ? node2265 : 4'b1000;
													assign node2265 = (inp[7]) ? node2267 : 4'b1000;
														assign node2267 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node2270 = (inp[7]) ? node2274 : node2271;
													assign node2271 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node2274 = (inp[13]) ? 4'b1100 : 4'b1101;
											assign node2277 = (inp[11]) ? node2285 : node2278;
												assign node2278 = (inp[13]) ? 4'b1001 : node2279;
													assign node2279 = (inp[0]) ? node2281 : 4'b1000;
														assign node2281 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node2285 = (inp[13]) ? node2287 : 4'b1000;
													assign node2287 = (inp[15]) ? 4'b1000 : 4'b1001;
										assign node2290 = (inp[14]) ? 4'b1100 : node2291;
											assign node2291 = (inp[15]) ? node2299 : node2292;
												assign node2292 = (inp[11]) ? node2294 : 4'b1101;
													assign node2294 = (inp[0]) ? 4'b1101 : node2295;
														assign node2295 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node2299 = (inp[7]) ? 4'b1000 : node2300;
													assign node2300 = (inp[0]) ? 4'b1100 : node2301;
														assign node2301 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node2307 = (inp[2]) ? node2331 : node2308;
										assign node2308 = (inp[0]) ? node2322 : node2309;
											assign node2309 = (inp[10]) ? node2315 : node2310;
												assign node2310 = (inp[14]) ? 4'b1100 : node2311;
													assign node2311 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node2315 = (inp[14]) ? 4'b1101 : node2316;
													assign node2316 = (inp[7]) ? 4'b1000 : node2317;
														assign node2317 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node2322 = (inp[13]) ? node2324 : 4'b1101;
												assign node2324 = (inp[10]) ? node2328 : node2325;
													assign node2325 = (inp[14]) ? 4'b1101 : 4'b1000;
													assign node2328 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node2331 = (inp[13]) ? node2343 : node2332;
											assign node2332 = (inp[0]) ? node2334 : 4'b1001;
												assign node2334 = (inp[7]) ? node2336 : 4'b1001;
													assign node2336 = (inp[14]) ? node2340 : node2337;
														assign node2337 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node2340 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node2343 = (inp[14]) ? node2347 : node2344;
												assign node2344 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node2347 = (inp[15]) ? node2349 : 4'b1000;
													assign node2349 = (inp[11]) ? 4'b1001 : node2350;
														assign node2350 = (inp[0]) ? 4'b1000 : 4'b1000;
								assign node2354 = (inp[11]) ? node2408 : node2355;
									assign node2355 = (inp[13]) ? node2381 : node2356;
										assign node2356 = (inp[15]) ? node2370 : node2357;
											assign node2357 = (inp[7]) ? node2363 : node2358;
												assign node2358 = (inp[2]) ? node2360 : 4'b1010;
													assign node2360 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node2363 = (inp[2]) ? node2365 : 4'b1011;
													assign node2365 = (inp[10]) ? 4'b1010 : node2366;
														assign node2366 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node2370 = (inp[0]) ? node2378 : node2371;
												assign node2371 = (inp[10]) ? 4'b1011 : node2372;
													assign node2372 = (inp[7]) ? 4'b1010 : node2373;
														assign node2373 = (inp[1]) ? 4'b1110 : 4'b1010;
												assign node2378 = (inp[2]) ? 4'b1110 : 4'b1010;
										assign node2381 = (inp[10]) ? node2399 : node2382;
											assign node2382 = (inp[15]) ? node2396 : node2383;
												assign node2383 = (inp[1]) ? node2389 : node2384;
													assign node2384 = (inp[2]) ? node2386 : 4'b1011;
														assign node2386 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node2389 = (inp[0]) ? node2393 : node2390;
														assign node2390 = (inp[7]) ? 4'b1010 : 4'b1110;
														assign node2393 = (inp[7]) ? 4'b1111 : 4'b1011;
												assign node2396 = (inp[14]) ? 4'b1111 : 4'b1011;
											assign node2399 = (inp[15]) ? 4'b1010 : node2400;
												assign node2400 = (inp[0]) ? node2402 : 4'b1111;
													assign node2402 = (inp[7]) ? node2404 : 4'b1010;
														assign node2404 = (inp[2]) ? 4'b1110 : 4'b1010;
									assign node2408 = (inp[13]) ? node2430 : node2409;
										assign node2409 = (inp[7]) ? node2417 : node2410;
											assign node2410 = (inp[0]) ? node2414 : node2411;
												assign node2411 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node2414 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node2417 = (inp[10]) ? node2427 : node2418;
												assign node2418 = (inp[0]) ? node2424 : node2419;
													assign node2419 = (inp[14]) ? 4'b1111 : node2420;
														assign node2420 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node2424 = (inp[15]) ? 4'b1110 : 4'b1010;
												assign node2427 = (inp[15]) ? 4'b1010 : 4'b1110;
										assign node2430 = (inp[10]) ? node2446 : node2431;
											assign node2431 = (inp[15]) ? node2437 : node2432;
												assign node2432 = (inp[0]) ? node2434 : 4'b1110;
													assign node2434 = (inp[7]) ? 4'b1111 : 4'b1011;
												assign node2437 = (inp[1]) ? node2443 : node2438;
													assign node2438 = (inp[2]) ? 4'b1011 : node2439;
														assign node2439 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node2443 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node2446 = (inp[1]) ? node2450 : node2447;
												assign node2447 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node2450 = (inp[2]) ? 4'b1010 : node2451;
													assign node2451 = (inp[7]) ? 4'b1110 : node2452;
														assign node2452 = (inp[15]) ? 4'b1010 : 4'b1110;
							assign node2457 = (inp[4]) ? node2553 : node2458;
								assign node2458 = (inp[1]) ? node2500 : node2459;
									assign node2459 = (inp[2]) ? node2479 : node2460;
										assign node2460 = (inp[0]) ? node2474 : node2461;
											assign node2461 = (inp[10]) ? node2469 : node2462;
												assign node2462 = (inp[11]) ? node2464 : 4'b1010;
													assign node2464 = (inp[15]) ? node2466 : 4'b1011;
														assign node2466 = (inp[7]) ? 4'b1010 : 4'b1111;
												assign node2469 = (inp[7]) ? node2471 : 4'b1011;
													assign node2471 = (inp[13]) ? 4'b1011 : 4'b1111;
											assign node2474 = (inp[11]) ? node2476 : 4'b1011;
												assign node2476 = (inp[7]) ? 4'b1011 : 4'b1010;
										assign node2479 = (inp[14]) ? node2489 : node2480;
											assign node2480 = (inp[11]) ? node2482 : 4'b1110;
												assign node2482 = (inp[0]) ? node2484 : 4'b1111;
													assign node2484 = (inp[10]) ? 4'b1111 : node2485;
														assign node2485 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node2489 = (inp[7]) ? node2491 : 4'b1010;
												assign node2491 = (inp[15]) ? node2497 : node2492;
													assign node2492 = (inp[10]) ? node2494 : 4'b1010;
														assign node2494 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node2497 = (inp[13]) ? 4'b1111 : 4'b1110;
									assign node2500 = (inp[2]) ? node2530 : node2501;
										assign node2501 = (inp[10]) ? node2515 : node2502;
											assign node2502 = (inp[11]) ? node2510 : node2503;
												assign node2503 = (inp[15]) ? 4'b1111 : node2504;
													assign node2504 = (inp[13]) ? node2506 : 4'b1110;
														assign node2506 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node2510 = (inp[15]) ? 4'b1110 : node2511;
													assign node2511 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node2515 = (inp[15]) ? node2521 : node2516;
												assign node2516 = (inp[14]) ? node2518 : 4'b1111;
													assign node2518 = (inp[11]) ? 4'b1010 : 4'b1111;
												assign node2521 = (inp[13]) ? node2523 : 4'b1110;
													assign node2523 = (inp[11]) ? node2527 : node2524;
														assign node2524 = (inp[0]) ? 4'b1010 : 4'b1111;
														assign node2527 = (inp[7]) ? 4'b1011 : 4'b1011;
										assign node2530 = (inp[7]) ? node2542 : node2531;
											assign node2531 = (inp[14]) ? node2539 : node2532;
												assign node2532 = (inp[11]) ? node2534 : 4'b1010;
													assign node2534 = (inp[13]) ? node2536 : 4'b1011;
														assign node2536 = (inp[10]) ? 4'b1010 : 4'b1010;
												assign node2539 = (inp[0]) ? 4'b1011 : 4'b1111;
											assign node2542 = (inp[0]) ? node2550 : node2543;
												assign node2543 = (inp[10]) ? node2545 : 4'b1010;
													assign node2545 = (inp[15]) ? node2547 : 4'b1111;
														assign node2547 = (inp[14]) ? 4'b1011 : 4'b1111;
												assign node2550 = (inp[10]) ? 4'b1110 : 4'b1111;
								assign node2553 = (inp[11]) ? node2587 : node2554;
									assign node2554 = (inp[13]) ? node2568 : node2555;
										assign node2555 = (inp[7]) ? node2559 : node2556;
											assign node2556 = (inp[15]) ? 4'b1001 : 4'b1101;
											assign node2559 = (inp[14]) ? 4'b1101 : node2560;
												assign node2560 = (inp[10]) ? node2562 : 4'b1101;
													assign node2562 = (inp[1]) ? node2564 : 4'b1100;
														assign node2564 = (inp[2]) ? 4'b1100 : 4'b1000;
										assign node2568 = (inp[1]) ? node2580 : node2569;
											assign node2569 = (inp[2]) ? node2577 : node2570;
												assign node2570 = (inp[0]) ? node2572 : 4'b1000;
													assign node2572 = (inp[10]) ? 4'b1001 : node2573;
														assign node2573 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node2577 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node2580 = (inp[14]) ? node2584 : node2581;
												assign node2581 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node2584 = (inp[2]) ? 4'b1000 : 4'b1100;
									assign node2587 = (inp[2]) ? node2601 : node2588;
										assign node2588 = (inp[0]) ? node2596 : node2589;
											assign node2589 = (inp[10]) ? node2591 : 4'b1000;
												assign node2591 = (inp[14]) ? 4'b1100 : node2592;
													assign node2592 = (inp[15]) ? 4'b1001 : 4'b1101;
											assign node2596 = (inp[14]) ? node2598 : 4'b1100;
												assign node2598 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node2601 = (inp[13]) ? node2607 : node2602;
											assign node2602 = (inp[10]) ? 4'b1100 : node2603;
												assign node2603 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node2607 = (inp[1]) ? node2613 : node2608;
												assign node2608 = (inp[7]) ? 4'b1101 : node2609;
													assign node2609 = (inp[0]) ? 4'b1000 : 4'b1100;
												assign node2613 = (inp[10]) ? node2615 : 4'b1001;
													assign node2615 = (inp[7]) ? node2619 : node2616;
														assign node2616 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node2619 = (inp[0]) ? 4'b1000 : 4'b1001;
						assign node2622 = (inp[4]) ? node2812 : node2623;
							assign node2623 = (inp[12]) ? node2717 : node2624;
								assign node2624 = (inp[0]) ? node2674 : node2625;
									assign node2625 = (inp[13]) ? node2647 : node2626;
										assign node2626 = (inp[7]) ? node2638 : node2627;
											assign node2627 = (inp[10]) ? node2631 : node2628;
												assign node2628 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node2631 = (inp[15]) ? 4'b1001 : node2632;
													assign node2632 = (inp[14]) ? node2634 : 4'b1001;
														assign node2634 = (inp[1]) ? 4'b1001 : 4'b1100;
											assign node2638 = (inp[10]) ? 4'b1000 : node2639;
												assign node2639 = (inp[1]) ? node2641 : 4'b1001;
													assign node2641 = (inp[15]) ? node2643 : 4'b1000;
														assign node2643 = (inp[14]) ? 4'b1000 : 4'b1000;
										assign node2647 = (inp[11]) ? node2653 : node2648;
											assign node2648 = (inp[1]) ? node2650 : 4'b1100;
												assign node2650 = (inp[10]) ? 4'b1100 : 4'b1000;
											assign node2653 = (inp[15]) ? node2663 : node2654;
												assign node2654 = (inp[1]) ? node2660 : node2655;
													assign node2655 = (inp[14]) ? 4'b1001 : node2656;
														assign node2656 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node2660 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node2663 = (inp[14]) ? node2669 : node2664;
													assign node2664 = (inp[10]) ? node2666 : 4'b1100;
														assign node2666 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node2669 = (inp[1]) ? node2671 : 4'b1100;
														assign node2671 = (inp[2]) ? 4'b1101 : 4'b1001;
									assign node2674 = (inp[10]) ? node2704 : node2675;
										assign node2675 = (inp[14]) ? node2695 : node2676;
											assign node2676 = (inp[1]) ? node2686 : node2677;
												assign node2677 = (inp[11]) ? node2681 : node2678;
													assign node2678 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node2681 = (inp[7]) ? 4'b1001 : node2682;
														assign node2682 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node2686 = (inp[7]) ? node2690 : node2687;
													assign node2687 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node2690 = (inp[15]) ? 4'b1001 : node2691;
														assign node2691 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node2695 = (inp[2]) ? node2699 : node2696;
												assign node2696 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node2699 = (inp[7]) ? node2701 : 4'b1000;
													assign node2701 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node2704 = (inp[7]) ? node2712 : node2705;
											assign node2705 = (inp[14]) ? node2709 : node2706;
												assign node2706 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node2709 = (inp[11]) ? 4'b1001 : 4'b1101;
											assign node2712 = (inp[14]) ? node2714 : 4'b1000;
												assign node2714 = (inp[13]) ? 4'b1100 : 4'b1000;
								assign node2717 = (inp[13]) ? node2773 : node2718;
									assign node2718 = (inp[14]) ? node2748 : node2719;
										assign node2719 = (inp[2]) ? node2733 : node2720;
											assign node2720 = (inp[0]) ? 4'b1010 : node2721;
												assign node2721 = (inp[15]) ? node2727 : node2722;
													assign node2722 = (inp[10]) ? 4'b1110 : node2723;
														assign node2723 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node2727 = (inp[10]) ? node2729 : 4'b1010;
														assign node2729 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node2733 = (inp[1]) ? node2743 : node2734;
												assign node2734 = (inp[0]) ? node2740 : node2735;
													assign node2735 = (inp[7]) ? node2737 : 4'b1110;
														assign node2737 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node2740 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node2743 = (inp[10]) ? 4'b1010 : node2744;
													assign node2744 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node2748 = (inp[1]) ? node2760 : node2749;
											assign node2749 = (inp[2]) ? node2755 : node2750;
												assign node2750 = (inp[0]) ? node2752 : 4'b1011;
													assign node2752 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node2755 = (inp[7]) ? 4'b1111 : node2756;
													assign node2756 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node2760 = (inp[2]) ? node2768 : node2761;
												assign node2761 = (inp[10]) ? node2763 : 4'b1110;
													assign node2763 = (inp[7]) ? node2765 : 4'b1111;
														assign node2765 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node2768 = (inp[0]) ? 4'b1010 : node2769;
													assign node2769 = (inp[7]) ? 4'b1011 : 4'b1010;
									assign node2773 = (inp[15]) ? node2795 : node2774;
										assign node2774 = (inp[7]) ? node2786 : node2775;
											assign node2775 = (inp[2]) ? node2779 : node2776;
												assign node2776 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node2779 = (inp[1]) ? node2781 : 4'b1111;
													assign node2781 = (inp[0]) ? 4'b1010 : node2782;
														assign node2782 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node2786 = (inp[14]) ? node2788 : 4'b1010;
												assign node2788 = (inp[2]) ? 4'b1011 : node2789;
													assign node2789 = (inp[0]) ? node2791 : 4'b1010;
														assign node2791 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node2795 = (inp[2]) ? node2807 : node2796;
											assign node2796 = (inp[1]) ? node2802 : node2797;
												assign node2797 = (inp[10]) ? 4'b1010 : node2798;
													assign node2798 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node2802 = (inp[10]) ? 4'b1111 : node2803;
													assign node2803 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node2807 = (inp[1]) ? 4'b1011 : node2808;
												assign node2808 = (inp[0]) ? 4'b1111 : 4'b1110;
							assign node2812 = (inp[12]) ? node2916 : node2813;
								assign node2813 = (inp[0]) ? node2879 : node2814;
									assign node2814 = (inp[15]) ? node2844 : node2815;
										assign node2815 = (inp[13]) ? node2835 : node2816;
											assign node2816 = (inp[10]) ? node2828 : node2817;
												assign node2817 = (inp[7]) ? node2823 : node2818;
													assign node2818 = (inp[11]) ? node2820 : 4'b1010;
														assign node2820 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node2823 = (inp[2]) ? node2825 : 4'b1010;
														assign node2825 = (inp[11]) ? 4'b1011 : 4'b1111;
												assign node2828 = (inp[2]) ? node2830 : 4'b1111;
													assign node2830 = (inp[11]) ? 4'b1011 : node2831;
														assign node2831 = (inp[7]) ? 4'b1011 : 4'b1111;
											assign node2835 = (inp[14]) ? node2839 : node2836;
												assign node2836 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node2839 = (inp[7]) ? node2841 : 4'b1011;
													assign node2841 = (inp[2]) ? 4'b1011 : 4'b1111;
										assign node2844 = (inp[14]) ? node2864 : node2845;
											assign node2845 = (inp[2]) ? node2855 : node2846;
												assign node2846 = (inp[7]) ? node2852 : node2847;
													assign node2847 = (inp[10]) ? 4'b1010 : node2848;
														assign node2848 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node2852 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node2855 = (inp[13]) ? node2857 : 4'b1111;
													assign node2857 = (inp[11]) ? node2861 : node2858;
														assign node2858 = (inp[7]) ? 4'b1010 : 4'b1111;
														assign node2861 = (inp[10]) ? 4'b1110 : 4'b1010;
											assign node2864 = (inp[11]) ? node2872 : node2865;
												assign node2865 = (inp[10]) ? node2867 : 4'b1011;
													assign node2867 = (inp[7]) ? node2869 : 4'b1111;
														assign node2869 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node2872 = (inp[2]) ? 4'b1111 : node2873;
													assign node2873 = (inp[1]) ? node2875 : 4'b1010;
														assign node2875 = (inp[7]) ? 4'b1110 : 4'b1111;
									assign node2879 = (inp[14]) ? node2895 : node2880;
										assign node2880 = (inp[15]) ? node2884 : node2881;
											assign node2881 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node2884 = (inp[11]) ? 4'b1010 : node2885;
												assign node2885 = (inp[7]) ? node2891 : node2886;
													assign node2886 = (inp[13]) ? 4'b1110 : node2887;
														assign node2887 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node2891 = (inp[13]) ? 4'b1111 : 4'b1110;
										assign node2895 = (inp[15]) ? node2905 : node2896;
											assign node2896 = (inp[10]) ? node2902 : node2897;
												assign node2897 = (inp[7]) ? node2899 : 4'b1110;
													assign node2899 = (inp[1]) ? 4'b1110 : 4'b1011;
												assign node2902 = (inp[2]) ? 4'b1110 : 4'b1010;
											assign node2905 = (inp[1]) ? node2909 : node2906;
												assign node2906 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node2909 = (inp[2]) ? node2911 : 4'b1111;
													assign node2911 = (inp[11]) ? node2913 : 4'b1010;
														assign node2913 = (inp[13]) ? 4'b1011 : 4'b1010;
								assign node2916 = (inp[14]) ? node2950 : node2917;
									assign node2917 = (inp[15]) ? node2927 : node2918;
										assign node2918 = (inp[11]) ? node2920 : 4'b1101;
											assign node2920 = (inp[0]) ? node2922 : 4'b1000;
												assign node2922 = (inp[7]) ? node2924 : 4'b1100;
													assign node2924 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node2927 = (inp[2]) ? node2939 : node2928;
											assign node2928 = (inp[1]) ? node2932 : node2929;
												assign node2929 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node2932 = (inp[13]) ? 4'b1101 : node2933;
													assign node2933 = (inp[11]) ? node2935 : 4'b1100;
														assign node2935 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node2939 = (inp[1]) ? node2945 : node2940;
												assign node2940 = (inp[10]) ? 4'b1101 : node2941;
													assign node2941 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node2945 = (inp[11]) ? node2947 : 4'b1001;
													assign node2947 = (inp[10]) ? 4'b1000 : 4'b1001;
									assign node2950 = (inp[11]) ? node2974 : node2951;
										assign node2951 = (inp[1]) ? node2967 : node2952;
											assign node2952 = (inp[2]) ? node2960 : node2953;
												assign node2953 = (inp[7]) ? 4'b1001 : node2954;
													assign node2954 = (inp[13]) ? 4'b1000 : node2955;
														assign node2955 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node2960 = (inp[15]) ? node2964 : node2961;
													assign node2961 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node2964 = (inp[13]) ? 4'b1101 : 4'b1100;
											assign node2967 = (inp[15]) ? 4'b1000 : node2968;
												assign node2968 = (inp[13]) ? node2970 : 4'b1000;
													assign node2970 = (inp[0]) ? 4'b1100 : 4'b1000;
										assign node2974 = (inp[0]) ? node2986 : node2975;
											assign node2975 = (inp[10]) ? 4'b1101 : node2976;
												assign node2976 = (inp[13]) ? node2978 : 4'b1100;
													assign node2978 = (inp[1]) ? node2982 : node2979;
														assign node2979 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node2982 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node2986 = (inp[10]) ? 4'b1000 : node2987;
												assign node2987 = (inp[15]) ? 4'b1101 : node2988;
													assign node2988 = (inp[7]) ? 4'b1001 : 4'b1101;
			assign node2993 = (inp[14]) ? node4313 : node2994;
				assign node2994 = (inp[8]) ? node3610 : node2995;
					assign node2995 = (inp[7]) ? node3279 : node2996;
						assign node2996 = (inp[15]) ? node3134 : node2997;
							assign node2997 = (inp[4]) ? node3067 : node2998;
								assign node2998 = (inp[1]) ? node3030 : node2999;
									assign node2999 = (inp[5]) ? node3009 : node3000;
										assign node3000 = (inp[13]) ? 4'b1101 : node3001;
											assign node3001 = (inp[12]) ? node3003 : 4'b1000;
												assign node3003 = (inp[10]) ? 4'b1001 : node3004;
													assign node3004 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node3009 = (inp[13]) ? node3019 : node3010;
											assign node3010 = (inp[10]) ? 4'b1100 : node3011;
												assign node3011 = (inp[9]) ? 4'b1101 : node3012;
													assign node3012 = (inp[11]) ? node3014 : 4'b1100;
														assign node3014 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node3019 = (inp[10]) ? node3027 : node3020;
												assign node3020 = (inp[11]) ? 4'b1001 : node3021;
													assign node3021 = (inp[0]) ? node3023 : 4'b1000;
														assign node3023 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node3027 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node3030 = (inp[2]) ? node3044 : node3031;
										assign node3031 = (inp[0]) ? node3037 : node3032;
											assign node3032 = (inp[13]) ? node3034 : 4'b1000;
												assign node3034 = (inp[12]) ? 4'b1001 : 4'b1100;
											assign node3037 = (inp[11]) ? 4'b1001 : node3038;
												assign node3038 = (inp[12]) ? 4'b1101 : node3039;
													assign node3039 = (inp[5]) ? 4'b1101 : 4'b1001;
										assign node3044 = (inp[5]) ? node3060 : node3045;
											assign node3045 = (inp[9]) ? node3053 : node3046;
												assign node3046 = (inp[11]) ? 4'b1100 : node3047;
													assign node3047 = (inp[0]) ? node3049 : 4'b1000;
														assign node3049 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node3053 = (inp[10]) ? node3057 : node3054;
													assign node3054 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node3057 = (inp[0]) ? 4'b1000 : 4'b1100;
											assign node3060 = (inp[11]) ? node3062 : 4'b1000;
												assign node3062 = (inp[10]) ? node3064 : 4'b1001;
													assign node3064 = (inp[13]) ? 4'b1100 : 4'b1001;
								assign node3067 = (inp[13]) ? node3101 : node3068;
									assign node3068 = (inp[5]) ? node3084 : node3069;
										assign node3069 = (inp[2]) ? node3075 : node3070;
											assign node3070 = (inp[0]) ? node3072 : 4'b1001;
												assign node3072 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node3075 = (inp[0]) ? node3077 : 4'b1000;
												assign node3077 = (inp[1]) ? 4'b1001 : node3078;
													assign node3078 = (inp[12]) ? 4'b1100 : node3079;
														assign node3079 = (inp[9]) ? 4'b1000 : 4'b1000;
										assign node3084 = (inp[1]) ? node3094 : node3085;
											assign node3085 = (inp[12]) ? node3089 : node3086;
												assign node3086 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node3089 = (inp[10]) ? node3091 : 4'b1000;
													assign node3091 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node3094 = (inp[0]) ? node3096 : 4'b1101;
												assign node3096 = (inp[12]) ? node3098 : 4'b1100;
													assign node3098 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node3101 = (inp[5]) ? node3121 : node3102;
										assign node3102 = (inp[1]) ? node3112 : node3103;
											assign node3103 = (inp[12]) ? node3109 : node3104;
												assign node3104 = (inp[9]) ? node3106 : 4'b1101;
													assign node3106 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node3109 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node3112 = (inp[11]) ? 4'b1100 : node3113;
												assign node3113 = (inp[0]) ? 4'b1100 : node3114;
													assign node3114 = (inp[2]) ? node3116 : 4'b1100;
														assign node3116 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node3121 = (inp[1]) ? node3127 : node3122;
											assign node3122 = (inp[12]) ? node3124 : 4'b1000;
												assign node3124 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node3127 = (inp[11]) ? 4'b1001 : node3128;
												assign node3128 = (inp[0]) ? node3130 : 4'b1000;
													assign node3130 = (inp[2]) ? 4'b1001 : 4'b1000;
							assign node3134 = (inp[13]) ? node3194 : node3135;
								assign node3135 = (inp[5]) ? node3171 : node3136;
									assign node3136 = (inp[1]) ? node3158 : node3137;
										assign node3137 = (inp[0]) ? node3149 : node3138;
											assign node3138 = (inp[4]) ? node3142 : node3139;
												assign node3139 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node3142 = (inp[11]) ? 4'b1011 : node3143;
													assign node3143 = (inp[2]) ? 4'b1011 : node3144;
														assign node3144 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node3149 = (inp[2]) ? 4'b1010 : node3150;
												assign node3150 = (inp[11]) ? 4'b1010 : node3151;
													assign node3151 = (inp[9]) ? 4'b1011 : node3152;
														assign node3152 = (inp[4]) ? 4'b1011 : 4'b1010;
										assign node3158 = (inp[10]) ? node3168 : node3159;
											assign node3159 = (inp[2]) ? node3161 : 4'b1010;
												assign node3161 = (inp[0]) ? node3165 : node3162;
													assign node3162 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node3165 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node3168 = (inp[2]) ? 4'b1011 : 4'b1111;
									assign node3171 = (inp[1]) ? node3181 : node3172;
										assign node3172 = (inp[0]) ? node3174 : 4'b1111;
											assign node3174 = (inp[11]) ? node3176 : 4'b1111;
												assign node3176 = (inp[4]) ? node3178 : 4'b1110;
													assign node3178 = (inp[2]) ? 4'b1111 : 4'b1110;
										assign node3181 = (inp[12]) ? node3189 : node3182;
											assign node3182 = (inp[4]) ? 4'b1010 : node3183;
												assign node3183 = (inp[11]) ? node3185 : 4'b1110;
													assign node3185 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node3189 = (inp[4]) ? 4'b1111 : node3190;
												assign node3190 = (inp[11]) ? 4'b1011 : 4'b1010;
								assign node3194 = (inp[5]) ? node3236 : node3195;
									assign node3195 = (inp[1]) ? node3213 : node3196;
										assign node3196 = (inp[10]) ? node3202 : node3197;
											assign node3197 = (inp[11]) ? 4'b1110 : node3198;
												assign node3198 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node3202 = (inp[0]) ? node3208 : node3203;
												assign node3203 = (inp[9]) ? node3205 : 4'b1110;
													assign node3205 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node3208 = (inp[12]) ? 4'b1111 : node3209;
													assign node3209 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node3213 = (inp[10]) ? node3219 : node3214;
											assign node3214 = (inp[4]) ? node3216 : 4'b1010;
												assign node3216 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node3219 = (inp[2]) ? node3227 : node3220;
												assign node3220 = (inp[12]) ? 4'b1111 : node3221;
													assign node3221 = (inp[11]) ? node3223 : 4'b1011;
														assign node3223 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node3227 = (inp[0]) ? node3231 : node3228;
													assign node3228 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node3231 = (inp[9]) ? node3233 : 4'b1110;
														assign node3233 = (inp[12]) ? 4'b1111 : 4'b1110;
									assign node3236 = (inp[1]) ? node3256 : node3237;
										assign node3237 = (inp[11]) ? node3239 : 4'b1010;
											assign node3239 = (inp[12]) ? node3245 : node3240;
												assign node3240 = (inp[4]) ? node3242 : 4'b1011;
													assign node3242 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node3245 = (inp[0]) ? node3251 : node3246;
													assign node3246 = (inp[9]) ? 4'b1010 : node3247;
														assign node3247 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node3251 = (inp[9]) ? 4'b1011 : node3252;
														assign node3252 = (inp[4]) ? 4'b1010 : 4'b1011;
										assign node3256 = (inp[11]) ? node3268 : node3257;
											assign node3257 = (inp[4]) ? node3263 : node3258;
												assign node3258 = (inp[9]) ? 4'b1011 : node3259;
													assign node3259 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node3263 = (inp[2]) ? node3265 : 4'b1111;
													assign node3265 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node3268 = (inp[10]) ? 4'b1110 : node3269;
												assign node3269 = (inp[12]) ? node3275 : node3270;
													assign node3270 = (inp[4]) ? 4'b1111 : node3271;
														assign node3271 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node3275 = (inp[4]) ? 4'b1010 : 4'b1110;
						assign node3279 = (inp[15]) ? node3451 : node3280;
							assign node3280 = (inp[9]) ? node3360 : node3281;
								assign node3281 = (inp[1]) ? node3327 : node3282;
									assign node3282 = (inp[10]) ? node3314 : node3283;
										assign node3283 = (inp[0]) ? node3305 : node3284;
											assign node3284 = (inp[11]) ? node3298 : node3285;
												assign node3285 = (inp[4]) ? node3291 : node3286;
													assign node3286 = (inp[12]) ? 4'b1111 : node3287;
														assign node3287 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node3291 = (inp[13]) ? node3295 : node3292;
														assign node3292 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node3295 = (inp[12]) ? 4'b1010 : 4'b1011;
												assign node3298 = (inp[5]) ? 4'b1110 : node3299;
													assign node3299 = (inp[2]) ? 4'b1111 : node3300;
														assign node3300 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node3305 = (inp[5]) ? node3311 : node3306;
												assign node3306 = (inp[12]) ? 4'b1111 : node3307;
													assign node3307 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node3311 = (inp[13]) ? 4'b1011 : 4'b1110;
										assign node3314 = (inp[2]) ? node3320 : node3315;
											assign node3315 = (inp[11]) ? 4'b1111 : node3316;
												assign node3316 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node3320 = (inp[11]) ? 4'b1011 : node3321;
												assign node3321 = (inp[13]) ? 4'b1111 : node3322;
													assign node3322 = (inp[5]) ? 4'b1111 : 4'b1011;
									assign node3327 = (inp[11]) ? node3353 : node3328;
										assign node3328 = (inp[13]) ? node3344 : node3329;
											assign node3329 = (inp[10]) ? node3337 : node3330;
												assign node3330 = (inp[5]) ? 4'b1111 : node3331;
													assign node3331 = (inp[4]) ? node3333 : 4'b1111;
														assign node3333 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node3337 = (inp[5]) ? node3339 : 4'b1110;
													assign node3339 = (inp[4]) ? node3341 : 4'b1011;
														assign node3341 = (inp[12]) ? 4'b1111 : 4'b1110;
											assign node3344 = (inp[0]) ? node3350 : node3345;
												assign node3345 = (inp[10]) ? 4'b1010 : node3346;
													assign node3346 = (inp[5]) ? 4'b1011 : 4'b1010;
												assign node3350 = (inp[12]) ? 4'b1010 : 4'b1110;
										assign node3353 = (inp[2]) ? node3357 : node3354;
											assign node3354 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node3357 = (inp[0]) ? 4'b1011 : 4'b1010;
								assign node3360 = (inp[5]) ? node3406 : node3361;
									assign node3361 = (inp[13]) ? node3387 : node3362;
										assign node3362 = (inp[12]) ? node3374 : node3363;
											assign node3363 = (inp[2]) ? node3367 : node3364;
												assign node3364 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node3367 = (inp[11]) ? node3369 : 4'b1010;
													assign node3369 = (inp[4]) ? 4'b1011 : node3370;
														assign node3370 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node3374 = (inp[11]) ? node3378 : node3375;
												assign node3375 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node3378 = (inp[0]) ? node3384 : node3379;
													assign node3379 = (inp[1]) ? node3381 : 4'b1110;
														assign node3381 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node3384 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node3387 = (inp[1]) ? node3395 : node3388;
											assign node3388 = (inp[2]) ? 4'b1111 : node3389;
												assign node3389 = (inp[12]) ? 4'b1011 : node3390;
													assign node3390 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node3395 = (inp[4]) ? node3397 : 4'b1010;
												assign node3397 = (inp[11]) ? node3403 : node3398;
													assign node3398 = (inp[10]) ? node3400 : 4'b1111;
														assign node3400 = (inp[12]) ? 4'b1111 : 4'b1110;
													assign node3403 = (inp[2]) ? 4'b1111 : 4'b1110;
									assign node3406 = (inp[13]) ? node3424 : node3407;
										assign node3407 = (inp[4]) ? 4'b1110 : node3408;
											assign node3408 = (inp[12]) ? node3416 : node3409;
												assign node3409 = (inp[10]) ? node3411 : 4'b1111;
													assign node3411 = (inp[1]) ? 4'b1110 : node3412;
														assign node3412 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node3416 = (inp[1]) ? node3420 : node3417;
													assign node3417 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node3420 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node3424 = (inp[12]) ? node3432 : node3425;
											assign node3425 = (inp[10]) ? node3427 : 4'b1010;
												assign node3427 = (inp[4]) ? 4'b1010 : node3428;
													assign node3428 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node3432 = (inp[4]) ? node3440 : node3433;
												assign node3433 = (inp[10]) ? 4'b1110 : node3434;
													assign node3434 = (inp[0]) ? node3436 : 4'b1111;
														assign node3436 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node3440 = (inp[1]) ? node3446 : node3441;
													assign node3441 = (inp[2]) ? node3443 : 4'b1111;
														assign node3443 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node3446 = (inp[10]) ? node3448 : 4'b1011;
														assign node3448 = (inp[11]) ? 4'b1010 : 4'b1010;
							assign node3451 = (inp[10]) ? node3523 : node3452;
								assign node3452 = (inp[2]) ? node3490 : node3453;
									assign node3453 = (inp[4]) ? node3475 : node3454;
										assign node3454 = (inp[0]) ? node3470 : node3455;
											assign node3455 = (inp[12]) ? node3461 : node3456;
												assign node3456 = (inp[11]) ? node3458 : 4'b1101;
													assign node3458 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node3461 = (inp[1]) ? node3467 : node3462;
													assign node3462 = (inp[5]) ? node3464 : 4'b1001;
														assign node3464 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node3467 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node3470 = (inp[11]) ? 4'b1001 : node3471;
												assign node3471 = (inp[12]) ? 4'b1000 : 4'b1001;
										assign node3475 = (inp[12]) ? node3481 : node3476;
											assign node3476 = (inp[11]) ? 4'b1000 : node3477;
												assign node3477 = (inp[1]) ? 4'b1000 : 4'b1100;
											assign node3481 = (inp[9]) ? node3487 : node3482;
												assign node3482 = (inp[5]) ? 4'b1001 : node3483;
													assign node3483 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node3487 = (inp[5]) ? 4'b1100 : 4'b1101;
									assign node3490 = (inp[5]) ? node3506 : node3491;
										assign node3491 = (inp[13]) ? node3497 : node3492;
											assign node3492 = (inp[11]) ? 4'b1001 : node3493;
												assign node3493 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node3497 = (inp[11]) ? node3501 : node3498;
												assign node3498 = (inp[4]) ? 4'b1100 : 4'b1101;
												assign node3501 = (inp[9]) ? 4'b1101 : node3502;
													assign node3502 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node3506 = (inp[13]) ? node3518 : node3507;
											assign node3507 = (inp[11]) ? node3509 : 4'b1101;
												assign node3509 = (inp[9]) ? node3515 : node3510;
													assign node3510 = (inp[0]) ? node3512 : 4'b1101;
														assign node3512 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node3515 = (inp[0]) ? 4'b1000 : 4'b1100;
											assign node3518 = (inp[0]) ? 4'b1001 : node3519;
												assign node3519 = (inp[9]) ? 4'b1000 : 4'b1001;
								assign node3523 = (inp[12]) ? node3575 : node3524;
									assign node3524 = (inp[5]) ? node3550 : node3525;
										assign node3525 = (inp[13]) ? node3535 : node3526;
											assign node3526 = (inp[4]) ? node3532 : node3527;
												assign node3527 = (inp[1]) ? 4'b1000 : node3528;
													assign node3528 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node3532 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node3535 = (inp[1]) ? node3537 : 4'b1100;
												assign node3537 = (inp[4]) ? node3543 : node3538;
													assign node3538 = (inp[9]) ? node3540 : 4'b1100;
														assign node3540 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node3543 = (inp[2]) ? node3547 : node3544;
														assign node3544 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node3547 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node3550 = (inp[13]) ? node3564 : node3551;
											assign node3551 = (inp[4]) ? node3557 : node3552;
												assign node3552 = (inp[1]) ? 4'b1101 : node3553;
													assign node3553 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node3557 = (inp[11]) ? 4'b1101 : node3558;
													assign node3558 = (inp[9]) ? node3560 : 4'b1100;
														assign node3560 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node3564 = (inp[1]) ? 4'b1000 : node3565;
												assign node3565 = (inp[4]) ? node3571 : node3566;
													assign node3566 = (inp[9]) ? 4'b1101 : node3567;
														assign node3567 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node3571 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node3575 = (inp[2]) ? node3589 : node3576;
										assign node3576 = (inp[11]) ? node3584 : node3577;
											assign node3577 = (inp[0]) ? 4'b1001 : node3578;
												assign node3578 = (inp[9]) ? 4'b1101 : node3579;
													assign node3579 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node3584 = (inp[1]) ? 4'b1100 : node3585;
												assign node3585 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node3589 = (inp[5]) ? node3599 : node3590;
											assign node3590 = (inp[0]) ? node3596 : node3591;
												assign node3591 = (inp[9]) ? 4'b1101 : node3592;
													assign node3592 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node3596 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node3599 = (inp[13]) ? node3605 : node3600;
												assign node3600 = (inp[4]) ? 4'b1001 : node3601;
													assign node3601 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node3605 = (inp[9]) ? 4'b1100 : node3606;
													assign node3606 = (inp[0]) ? 4'b1001 : 4'b1000;
					assign node3610 = (inp[13]) ? node3980 : node3611;
						assign node3611 = (inp[11]) ? node3797 : node3612;
							assign node3612 = (inp[10]) ? node3712 : node3613;
								assign node3613 = (inp[9]) ? node3665 : node3614;
									assign node3614 = (inp[4]) ? node3638 : node3615;
										assign node3615 = (inp[15]) ? node3623 : node3616;
											assign node3616 = (inp[1]) ? node3618 : 4'b0100;
												assign node3618 = (inp[7]) ? 4'b0000 : node3619;
													assign node3619 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node3623 = (inp[2]) ? node3627 : node3624;
												assign node3624 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node3627 = (inp[5]) ? node3633 : node3628;
													assign node3628 = (inp[7]) ? node3630 : 4'b0110;
														assign node3630 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node3633 = (inp[0]) ? 4'b0011 : node3634;
														assign node3634 = (inp[7]) ? 4'b0110 : 4'b0010;
										assign node3638 = (inp[15]) ? node3652 : node3639;
											assign node3639 = (inp[5]) ? node3645 : node3640;
												assign node3640 = (inp[0]) ? node3642 : 4'b0010;
													assign node3642 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node3645 = (inp[1]) ? node3647 : 4'b0111;
													assign node3647 = (inp[7]) ? node3649 : 4'b0011;
														assign node3649 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node3652 = (inp[12]) ? node3656 : node3653;
												assign node3653 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node3656 = (inp[0]) ? 4'b0000 : node3657;
													assign node3657 = (inp[1]) ? node3661 : node3658;
														assign node3658 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node3661 = (inp[2]) ? 4'b0000 : 4'b0100;
									assign node3665 = (inp[1]) ? node3687 : node3666;
										assign node3666 = (inp[2]) ? node3682 : node3667;
											assign node3667 = (inp[5]) ? node3673 : node3668;
												assign node3668 = (inp[12]) ? node3670 : 4'b0000;
													assign node3670 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node3673 = (inp[0]) ? node3675 : 4'b0110;
													assign node3675 = (inp[12]) ? node3679 : node3676;
														assign node3676 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node3679 = (inp[15]) ? 4'b0100 : 4'b0001;
											assign node3682 = (inp[5]) ? node3684 : 4'b0011;
												assign node3684 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node3687 = (inp[7]) ? node3707 : node3688;
											assign node3688 = (inp[12]) ? node3700 : node3689;
												assign node3689 = (inp[5]) ? node3693 : node3690;
													assign node3690 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node3693 = (inp[15]) ? node3697 : node3694;
														assign node3694 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node3697 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node3700 = (inp[15]) ? 4'b0001 : node3701;
													assign node3701 = (inp[0]) ? 4'b0100 : node3702;
														assign node3702 = (inp[5]) ? 4'b0111 : 4'b0101;
											assign node3707 = (inp[15]) ? node3709 : 4'b0100;
												assign node3709 = (inp[0]) ? 4'b0010 : 4'b0011;
								assign node3712 = (inp[15]) ? node3756 : node3713;
									assign node3713 = (inp[4]) ? node3729 : node3714;
										assign node3714 = (inp[12]) ? node3722 : node3715;
											assign node3715 = (inp[9]) ? 4'b0101 : node3716;
												assign node3716 = (inp[1]) ? 4'b0001 : node3717;
													assign node3717 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node3722 = (inp[5]) ? node3726 : node3723;
												assign node3723 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node3726 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node3729 = (inp[0]) ? node3747 : node3730;
											assign node3730 = (inp[2]) ? node3738 : node3731;
												assign node3731 = (inp[1]) ? 4'b0110 : node3732;
													assign node3732 = (inp[7]) ? node3734 : 4'b0110;
														assign node3734 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node3738 = (inp[12]) ? node3744 : node3739;
													assign node3739 = (inp[5]) ? node3741 : 4'b0111;
														assign node3741 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node3744 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node3747 = (inp[1]) ? 4'b0110 : node3748;
												assign node3748 = (inp[9]) ? node3750 : 4'b0010;
													assign node3750 = (inp[12]) ? 4'b0111 : node3751;
														assign node3751 = (inp[5]) ? 4'b0110 : 4'b0010;
									assign node3756 = (inp[4]) ? node3788 : node3757;
										assign node3757 = (inp[0]) ? node3771 : node3758;
											assign node3758 = (inp[7]) ? node3764 : node3759;
												assign node3759 = (inp[9]) ? node3761 : 4'b0110;
													assign node3761 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node3764 = (inp[12]) ? 4'b0010 : node3765;
													assign node3765 = (inp[1]) ? 4'b0011 : node3766;
														assign node3766 = (inp[5]) ? 4'b0011 : 4'b0110;
											assign node3771 = (inp[9]) ? node3777 : node3772;
												assign node3772 = (inp[2]) ? node3774 : 4'b0111;
													assign node3774 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node3777 = (inp[1]) ? node3783 : node3778;
													assign node3778 = (inp[7]) ? node3780 : 4'b0011;
														assign node3780 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node3783 = (inp[7]) ? node3785 : 4'b0110;
														assign node3785 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node3788 = (inp[5]) ? node3790 : 4'b0001;
											assign node3790 = (inp[1]) ? node3792 : 4'b0100;
												assign node3792 = (inp[9]) ? node3794 : 4'b0000;
													assign node3794 = (inp[7]) ? 4'b0001 : 4'b0000;
							assign node3797 = (inp[0]) ? node3891 : node3798;
								assign node3798 = (inp[12]) ? node3838 : node3799;
									assign node3799 = (inp[2]) ? node3821 : node3800;
										assign node3800 = (inp[1]) ? node3816 : node3801;
											assign node3801 = (inp[5]) ? node3809 : node3802;
												assign node3802 = (inp[9]) ? 4'b0001 : node3803;
													assign node3803 = (inp[4]) ? 4'b0011 : node3804;
														assign node3804 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node3809 = (inp[7]) ? node3813 : node3810;
													assign node3810 = (inp[10]) ? 4'b0111 : 4'b0101;
													assign node3813 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node3816 = (inp[10]) ? node3818 : 4'b0100;
												assign node3818 = (inp[7]) ? 4'b0000 : 4'b0010;
										assign node3821 = (inp[1]) ? node3829 : node3822;
											assign node3822 = (inp[7]) ? 4'b0001 : node3823;
												assign node3823 = (inp[10]) ? node3825 : 4'b0001;
													assign node3825 = (inp[5]) ? 4'b0001 : 4'b0100;
											assign node3829 = (inp[9]) ? node3831 : 4'b0101;
												assign node3831 = (inp[4]) ? node3833 : 4'b0000;
													assign node3833 = (inp[15]) ? 4'b0001 : node3834;
														assign node3834 = (inp[10]) ? 4'b0011 : 4'b0110;
									assign node3838 = (inp[7]) ? node3870 : node3839;
										assign node3839 = (inp[1]) ? node3851 : node3840;
											assign node3840 = (inp[5]) ? node3842 : 4'b0001;
												assign node3842 = (inp[9]) ? node3848 : node3843;
													assign node3843 = (inp[15]) ? node3845 : 4'b0101;
														assign node3845 = (inp[2]) ? 4'b0101 : 4'b0111;
													assign node3848 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node3851 = (inp[5]) ? node3863 : node3852;
												assign node3852 = (inp[10]) ? node3858 : node3853;
													assign node3853 = (inp[4]) ? node3855 : 4'b0100;
														assign node3855 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node3858 = (inp[4]) ? 4'b0100 : node3859;
														assign node3859 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node3863 = (inp[4]) ? node3867 : node3864;
													assign node3864 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node3867 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node3870 = (inp[1]) ? node3878 : node3871;
											assign node3871 = (inp[2]) ? node3873 : 4'b0001;
												assign node3873 = (inp[5]) ? 4'b0111 : node3874;
													assign node3874 = (inp[15]) ? 4'b0010 : 4'b0011;
											assign node3878 = (inp[5]) ? node3884 : node3879;
												assign node3879 = (inp[2]) ? node3881 : 4'b0111;
													assign node3881 = (inp[15]) ? 4'b0101 : 4'b0001;
												assign node3884 = (inp[15]) ? node3888 : node3885;
													assign node3885 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node3888 = (inp[2]) ? 4'b0001 : 4'b0000;
								assign node3891 = (inp[1]) ? node3933 : node3892;
									assign node3892 = (inp[4]) ? node3914 : node3893;
										assign node3893 = (inp[15]) ? node3899 : node3894;
											assign node3894 = (inp[10]) ? node3896 : 4'b0100;
												assign node3896 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node3899 = (inp[9]) ? node3905 : node3900;
												assign node3900 = (inp[5]) ? node3902 : 4'b0010;
													assign node3902 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node3905 = (inp[12]) ? 4'b0110 : node3906;
													assign node3906 = (inp[10]) ? node3910 : node3907;
														assign node3907 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node3910 = (inp[7]) ? 4'b0110 : 4'b0010;
										assign node3914 = (inp[15]) ? node3928 : node3915;
											assign node3915 = (inp[5]) ? node3921 : node3916;
												assign node3916 = (inp[2]) ? node3918 : 4'b0010;
													assign node3918 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node3921 = (inp[12]) ? node3925 : node3922;
													assign node3922 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node3925 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node3928 = (inp[10]) ? node3930 : 4'b0100;
												assign node3930 = (inp[12]) ? 4'b0100 : 4'b0000;
									assign node3933 = (inp[9]) ? node3961 : node3934;
										assign node3934 = (inp[4]) ? node3948 : node3935;
											assign node3935 = (inp[15]) ? node3945 : node3936;
												assign node3936 = (inp[2]) ? node3942 : node3937;
													assign node3937 = (inp[5]) ? node3939 : 4'b0000;
														assign node3939 = (inp[7]) ? 4'b0001 : 4'b0001;
													assign node3942 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node3945 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node3948 = (inp[15]) ? node3954 : node3949;
												assign node3949 = (inp[10]) ? 4'b0010 : node3950;
													assign node3950 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node3954 = (inp[2]) ? 4'b0100 : node3955;
													assign node3955 = (inp[5]) ? node3957 : 4'b0101;
														assign node3957 = (inp[12]) ? 4'b0001 : 4'b0001;
										assign node3961 = (inp[15]) ? node3969 : node3962;
											assign node3962 = (inp[4]) ? node3964 : 4'b0101;
												assign node3964 = (inp[2]) ? node3966 : 4'b0110;
													assign node3966 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node3969 = (inp[4]) ? node3975 : node3970;
												assign node3970 = (inp[10]) ? node3972 : 4'b0110;
													assign node3972 = (inp[12]) ? 4'b0110 : 4'b0011;
												assign node3975 = (inp[5]) ? 4'b0000 : node3976;
													assign node3976 = (inp[12]) ? 4'b0101 : 4'b0100;
						assign node3980 = (inp[0]) ? node4142 : node3981;
							assign node3981 = (inp[12]) ? node4061 : node3982;
								assign node3982 = (inp[11]) ? node4020 : node3983;
									assign node3983 = (inp[4]) ? node4007 : node3984;
										assign node3984 = (inp[15]) ? node3998 : node3985;
											assign node3985 = (inp[2]) ? node3991 : node3986;
												assign node3986 = (inp[5]) ? node3988 : 4'b0000;
													assign node3988 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node3991 = (inp[7]) ? 4'b0101 : node3992;
													assign node3992 = (inp[1]) ? node3994 : 4'b0001;
														assign node3994 = (inp[5]) ? 4'b0001 : 4'b0101;
											assign node3998 = (inp[5]) ? node4000 : 4'b0110;
												assign node4000 = (inp[1]) ? 4'b0110 : node4001;
													assign node4001 = (inp[7]) ? 4'b0011 : node4002;
														assign node4002 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node4007 = (inp[15]) ? node4015 : node4008;
											assign node4008 = (inp[5]) ? node4012 : node4009;
												assign node4009 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node4012 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node4015 = (inp[9]) ? node4017 : 4'b0000;
												assign node4017 = (inp[5]) ? 4'b0000 : 4'b0101;
									assign node4020 = (inp[7]) ? node4044 : node4021;
										assign node4021 = (inp[2]) ? node4033 : node4022;
											assign node4022 = (inp[15]) ? node4028 : node4023;
												assign node4023 = (inp[4]) ? 4'b0111 : node4024;
													assign node4024 = (inp[1]) ? 4'b0101 : 4'b0001;
												assign node4028 = (inp[4]) ? 4'b0001 : node4029;
													assign node4029 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node4033 = (inp[10]) ? 4'b0111 : node4034;
												assign node4034 = (inp[4]) ? node4038 : node4035;
													assign node4035 = (inp[15]) ? 4'b0111 : 4'b0100;
													assign node4038 = (inp[15]) ? 4'b0100 : node4039;
														assign node4039 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node4044 = (inp[4]) ? node4054 : node4045;
											assign node4045 = (inp[15]) ? node4051 : node4046;
												assign node4046 = (inp[5]) ? node4048 : 4'b0100;
													assign node4048 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node4051 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node4054 = (inp[1]) ? node4056 : 4'b0100;
												assign node4056 = (inp[9]) ? node4058 : 4'b0001;
													assign node4058 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node4061 = (inp[2]) ? node4103 : node4062;
									assign node4062 = (inp[15]) ? node4082 : node4063;
										assign node4063 = (inp[4]) ? node4069 : node4064;
											assign node4064 = (inp[10]) ? 4'b0100 : node4065;
												assign node4065 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node4069 = (inp[5]) ? node4077 : node4070;
												assign node4070 = (inp[7]) ? node4074 : node4071;
													assign node4071 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node4074 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node4077 = (inp[9]) ? 4'b0011 : node4078;
													assign node4078 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node4082 = (inp[4]) ? node4088 : node4083;
											assign node4083 = (inp[1]) ? node4085 : 4'b0011;
												assign node4085 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node4088 = (inp[5]) ? node4098 : node4089;
												assign node4089 = (inp[1]) ? node4095 : node4090;
													assign node4090 = (inp[7]) ? node4092 : 4'b0000;
														assign node4092 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node4095 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node4098 = (inp[1]) ? 4'b0001 : node4099;
													assign node4099 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node4103 = (inp[15]) ? node4119 : node4104;
										assign node4104 = (inp[4]) ? node4110 : node4105;
											assign node4105 = (inp[11]) ? node4107 : 4'b0001;
												assign node4107 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node4110 = (inp[11]) ? node4116 : node4111;
												assign node4111 = (inp[9]) ? 4'b0110 : node4112;
													assign node4112 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node4116 = (inp[9]) ? 4'b0010 : 4'b0111;
										assign node4119 = (inp[4]) ? node4135 : node4120;
											assign node4120 = (inp[1]) ? node4128 : node4121;
												assign node4121 = (inp[5]) ? 4'b0111 : node4122;
													assign node4122 = (inp[11]) ? 4'b0010 : node4123;
														assign node4123 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node4128 = (inp[9]) ? node4132 : node4129;
													assign node4129 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node4132 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node4135 = (inp[10]) ? node4137 : 4'b0000;
												assign node4137 = (inp[9]) ? 4'b0101 : node4138;
													assign node4138 = (inp[11]) ? 4'b0001 : 4'b0101;
							assign node4142 = (inp[2]) ? node4228 : node4143;
								assign node4143 = (inp[7]) ? node4191 : node4144;
									assign node4144 = (inp[5]) ? node4166 : node4145;
										assign node4145 = (inp[1]) ? node4155 : node4146;
											assign node4146 = (inp[11]) ? node4152 : node4147;
												assign node4147 = (inp[4]) ? node4149 : 4'b0001;
													assign node4149 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node4152 = (inp[15]) ? 4'b0101 : 4'b0000;
											assign node4155 = (inp[10]) ? node4163 : node4156;
												assign node4156 = (inp[9]) ? 4'b0101 : node4157;
													assign node4157 = (inp[11]) ? node4159 : 4'b0011;
														assign node4159 = (inp[12]) ? 4'b0101 : 4'b0110;
												assign node4163 = (inp[15]) ? 4'b0100 : 4'b0010;
										assign node4166 = (inp[1]) ? node4178 : node4167;
											assign node4167 = (inp[10]) ? node4175 : node4168;
												assign node4168 = (inp[4]) ? node4172 : node4169;
													assign node4169 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node4172 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node4175 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node4178 = (inp[11]) ? node4184 : node4179;
												assign node4179 = (inp[15]) ? node4181 : 4'b0010;
													assign node4181 = (inp[4]) ? 4'b0100 : 4'b0010;
												assign node4184 = (inp[15]) ? node4188 : node4185;
													assign node4185 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node4188 = (inp[12]) ? 4'b0011 : 4'b0010;
									assign node4191 = (inp[5]) ? node4209 : node4192;
										assign node4192 = (inp[9]) ? node4198 : node4193;
											assign node4193 = (inp[15]) ? 4'b0100 : node4194;
												assign node4194 = (inp[4]) ? 4'b0010 : 4'b0000;
											assign node4198 = (inp[15]) ? node4204 : node4199;
												assign node4199 = (inp[4]) ? node4201 : 4'b0001;
													assign node4201 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node4204 = (inp[4]) ? node4206 : 4'b0010;
													assign node4206 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node4209 = (inp[12]) ? node4215 : node4210;
											assign node4210 = (inp[1]) ? node4212 : 4'b0101;
												assign node4212 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node4215 = (inp[1]) ? node4219 : node4216;
												assign node4216 = (inp[9]) ? 4'b0100 : 4'b0110;
												assign node4219 = (inp[4]) ? node4223 : node4220;
													assign node4220 = (inp[15]) ? 4'b0010 : 4'b0100;
													assign node4223 = (inp[9]) ? 4'b0010 : node4224;
														assign node4224 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node4228 = (inp[10]) ? node4274 : node4229;
									assign node4229 = (inp[15]) ? node4247 : node4230;
										assign node4230 = (inp[4]) ? node4244 : node4231;
											assign node4231 = (inp[12]) ? node4235 : node4232;
												assign node4232 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node4235 = (inp[7]) ? node4239 : node4236;
													assign node4236 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node4239 = (inp[11]) ? 4'b0001 : node4240;
														assign node4240 = (inp[1]) ? 4'b0000 : 4'b0000;
											assign node4244 = (inp[12]) ? 4'b0111 : 4'b0010;
										assign node4247 = (inp[4]) ? node4263 : node4248;
											assign node4248 = (inp[7]) ? node4254 : node4249;
												assign node4249 = (inp[9]) ? node4251 : 4'b0011;
													assign node4251 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node4254 = (inp[9]) ? node4258 : node4255;
													assign node4255 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node4258 = (inp[11]) ? 4'b0011 : node4259;
														assign node4259 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node4263 = (inp[5]) ? node4267 : node4264;
												assign node4264 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node4267 = (inp[1]) ? node4271 : node4268;
													assign node4268 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node4271 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node4274 = (inp[12]) ? node4300 : node4275;
										assign node4275 = (inp[11]) ? node4289 : node4276;
											assign node4276 = (inp[4]) ? node4280 : node4277;
												assign node4277 = (inp[15]) ? 4'b0111 : 4'b0100;
												assign node4280 = (inp[15]) ? node4286 : node4281;
													assign node4281 = (inp[9]) ? 4'b0110 : node4282;
														assign node4282 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node4286 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node4289 = (inp[1]) ? node4295 : node4290;
												assign node4290 = (inp[7]) ? node4292 : 4'b0101;
													assign node4292 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node4295 = (inp[4]) ? node4297 : 4'b0101;
													assign node4297 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node4300 = (inp[5]) ? node4304 : node4301;
											assign node4301 = (inp[7]) ? 4'b0101 : 4'b0111;
											assign node4304 = (inp[11]) ? node4310 : node4305;
												assign node4305 = (inp[15]) ? 4'b0001 : node4306;
													assign node4306 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node4310 = (inp[1]) ? 4'b0000 : 4'b0100;
				assign node4313 = (inp[4]) ? node4901 : node4314;
					assign node4314 = (inp[7]) ? node4592 : node4315;
						assign node4315 = (inp[8]) ? node4449 : node4316;
							assign node4316 = (inp[13]) ? node4380 : node4317;
								assign node4317 = (inp[12]) ? node4351 : node4318;
									assign node4318 = (inp[1]) ? node4334 : node4319;
										assign node4319 = (inp[5]) ? node4327 : node4320;
											assign node4320 = (inp[2]) ? node4324 : node4321;
												assign node4321 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node4324 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node4327 = (inp[0]) ? 4'b0000 : node4328;
												assign node4328 = (inp[2]) ? node4330 : 4'b0001;
													assign node4330 = (inp[15]) ? 4'b0000 : 4'b0001;
										assign node4334 = (inp[15]) ? node4336 : 4'b0001;
											assign node4336 = (inp[11]) ? node4344 : node4337;
												assign node4337 = (inp[5]) ? 4'b0101 : node4338;
													assign node4338 = (inp[2]) ? 4'b0101 : node4339;
														assign node4339 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node4344 = (inp[10]) ? node4346 : 4'b0101;
													assign node4346 = (inp[2]) ? 4'b0100 : node4347;
														assign node4347 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node4351 = (inp[15]) ? node4365 : node4352;
										assign node4352 = (inp[0]) ? 4'b0100 : node4353;
											assign node4353 = (inp[11]) ? node4355 : 4'b0101;
												assign node4355 = (inp[9]) ? node4357 : 4'b0100;
													assign node4357 = (inp[5]) ? node4361 : node4358;
														assign node4358 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node4361 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node4365 = (inp[1]) ? node4377 : node4366;
											assign node4366 = (inp[5]) ? 4'b0101 : node4367;
												assign node4367 = (inp[0]) ? node4373 : node4368;
													assign node4368 = (inp[9]) ? node4370 : 4'b0101;
														assign node4370 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node4373 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node4377 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node4380 = (inp[12]) ? node4410 : node4381;
									assign node4381 = (inp[15]) ? node4395 : node4382;
										assign node4382 = (inp[11]) ? 4'b0101 : node4383;
											assign node4383 = (inp[0]) ? node4389 : node4384;
												assign node4384 = (inp[1]) ? node4386 : 4'b0101;
													assign node4386 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node4389 = (inp[1]) ? node4391 : 4'b0100;
													assign node4391 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node4395 = (inp[1]) ? node4401 : node4396;
											assign node4396 = (inp[9]) ? node4398 : 4'b0101;
												assign node4398 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node4401 = (inp[10]) ? 4'b0001 : node4402;
												assign node4402 = (inp[11]) ? node4404 : 4'b0000;
													assign node4404 = (inp[2]) ? node4406 : 4'b0001;
														assign node4406 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node4410 = (inp[15]) ? node4434 : node4411;
										assign node4411 = (inp[5]) ? node4427 : node4412;
											assign node4412 = (inp[11]) ? node4420 : node4413;
												assign node4413 = (inp[2]) ? 4'b0000 : node4414;
													assign node4414 = (inp[10]) ? node4416 : 4'b0000;
														assign node4416 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node4420 = (inp[9]) ? 4'b0001 : node4421;
													assign node4421 = (inp[2]) ? node4423 : 4'b0000;
														assign node4423 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node4427 = (inp[11]) ? 4'b0000 : node4428;
												assign node4428 = (inp[1]) ? node4430 : 4'b0000;
													assign node4430 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node4434 = (inp[1]) ? node4440 : node4435;
											assign node4435 = (inp[9]) ? node4437 : 4'b0001;
												assign node4437 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node4440 = (inp[10]) ? node4442 : 4'b0101;
												assign node4442 = (inp[5]) ? 4'b0100 : node4443;
													assign node4443 = (inp[0]) ? 4'b0101 : node4444;
														assign node4444 = (inp[2]) ? 4'b0101 : 4'b0100;
							assign node4449 = (inp[5]) ? node4535 : node4450;
								assign node4450 = (inp[13]) ? node4498 : node4451;
									assign node4451 = (inp[15]) ? node4471 : node4452;
										assign node4452 = (inp[9]) ? node4462 : node4453;
											assign node4453 = (inp[0]) ? node4455 : 4'b0010;
												assign node4455 = (inp[11]) ? 4'b0011 : node4456;
													assign node4456 = (inp[2]) ? 4'b0010 : node4457;
														assign node4457 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node4462 = (inp[11]) ? node4466 : node4463;
												assign node4463 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node4466 = (inp[10]) ? 4'b0010 : node4467;
													assign node4467 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node4471 = (inp[10]) ? node4481 : node4472;
											assign node4472 = (inp[0]) ? 4'b0010 : node4473;
												assign node4473 = (inp[2]) ? node4475 : 4'b0110;
													assign node4475 = (inp[12]) ? node4477 : 4'b0011;
														assign node4477 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node4481 = (inp[11]) ? node4491 : node4482;
												assign node4482 = (inp[2]) ? node4488 : node4483;
													assign node4483 = (inp[0]) ? node4485 : 4'b0010;
														assign node4485 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node4488 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node4491 = (inp[9]) ? 4'b0011 : node4492;
													assign node4492 = (inp[1]) ? 4'b0111 : node4493;
														assign node4493 = (inp[12]) ? 4'b0111 : 4'b0011;
									assign node4498 = (inp[0]) ? node4516 : node4499;
										assign node4499 = (inp[15]) ? node4505 : node4500;
											assign node4500 = (inp[12]) ? 4'b0110 : node4501;
												assign node4501 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node4505 = (inp[12]) ? node4511 : node4506;
												assign node4506 = (inp[1]) ? node4508 : 4'b0011;
													assign node4508 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node4511 = (inp[2]) ? 4'b0010 : node4512;
													assign node4512 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node4516 = (inp[2]) ? node4530 : node4517;
											assign node4517 = (inp[15]) ? node4525 : node4518;
												assign node4518 = (inp[1]) ? node4522 : node4519;
													assign node4519 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node4522 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node4525 = (inp[12]) ? 4'b0010 : node4526;
													assign node4526 = (inp[1]) ? 4'b0111 : 4'b0010;
											assign node4530 = (inp[9]) ? 4'b0110 : node4531;
												assign node4531 = (inp[15]) ? 4'b0011 : 4'b0110;
								assign node4535 = (inp[12]) ? node4575 : node4536;
									assign node4536 = (inp[1]) ? node4548 : node4537;
										assign node4537 = (inp[0]) ? node4545 : node4538;
											assign node4538 = (inp[2]) ? node4540 : 4'b0010;
												assign node4540 = (inp[13]) ? node4542 : 4'b0011;
													assign node4542 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node4545 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node4548 = (inp[11]) ? node4564 : node4549;
											assign node4549 = (inp[0]) ? node4557 : node4550;
												assign node4550 = (inp[13]) ? node4552 : 4'b0110;
													assign node4552 = (inp[15]) ? node4554 : 4'b0111;
														assign node4554 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node4557 = (inp[9]) ? node4559 : 4'b0111;
													assign node4559 = (inp[13]) ? node4561 : 4'b0111;
														assign node4561 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node4564 = (inp[9]) ? node4566 : 4'b0110;
												assign node4566 = (inp[13]) ? node4570 : node4567;
													assign node4567 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node4570 = (inp[0]) ? node4572 : 4'b0111;
														assign node4572 = (inp[15]) ? 4'b0110 : 4'b0110;
									assign node4575 = (inp[1]) ? node4585 : node4576;
										assign node4576 = (inp[15]) ? node4580 : node4577;
											assign node4577 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node4580 = (inp[9]) ? 4'b0110 : node4581;
												assign node4581 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node4585 = (inp[2]) ? node4589 : node4586;
											assign node4586 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node4589 = (inp[0]) ? 4'b0010 : 4'b0011;
						assign node4592 = (inp[0]) ? node4760 : node4593;
							assign node4593 = (inp[2]) ? node4669 : node4594;
								assign node4594 = (inp[11]) ? node4628 : node4595;
									assign node4595 = (inp[13]) ? node4617 : node4596;
										assign node4596 = (inp[12]) ? node4608 : node4597;
											assign node4597 = (inp[15]) ? node4603 : node4598;
												assign node4598 = (inp[5]) ? 4'b0010 : node4599;
													assign node4599 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node4603 = (inp[8]) ? 4'b0010 : node4604;
													assign node4604 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node4608 = (inp[10]) ? 4'b0110 : node4609;
												assign node4609 = (inp[5]) ? 4'b0011 : node4610;
													assign node4610 = (inp[15]) ? 4'b0111 : node4611;
														assign node4611 = (inp[8]) ? 4'b0110 : 4'b0110;
										assign node4617 = (inp[12]) ? node4625 : node4618;
											assign node4618 = (inp[1]) ? node4622 : node4619;
												assign node4619 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node4622 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node4625 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node4628 = (inp[12]) ? node4654 : node4629;
										assign node4629 = (inp[1]) ? node4637 : node4630;
											assign node4630 = (inp[5]) ? node4634 : node4631;
												assign node4631 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node4634 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node4637 = (inp[10]) ? node4645 : node4638;
												assign node4638 = (inp[15]) ? 4'b0111 : node4639;
													assign node4639 = (inp[8]) ? 4'b0110 : node4640;
														assign node4640 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node4645 = (inp[8]) ? node4649 : node4646;
													assign node4646 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node4649 = (inp[9]) ? 4'b0110 : node4650;
														assign node4650 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node4654 = (inp[1]) ? node4664 : node4655;
											assign node4655 = (inp[8]) ? 4'b0110 : node4656;
												assign node4656 = (inp[15]) ? node4658 : 4'b0010;
													assign node4658 = (inp[13]) ? node4660 : 4'b0010;
														assign node4660 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node4664 = (inp[13]) ? node4666 : 4'b0110;
												assign node4666 = (inp[8]) ? 4'b0010 : 4'b0011;
								assign node4669 = (inp[8]) ? node4725 : node4670;
									assign node4670 = (inp[11]) ? node4700 : node4671;
										assign node4671 = (inp[13]) ? node4687 : node4672;
											assign node4672 = (inp[12]) ? node4682 : node4673;
												assign node4673 = (inp[10]) ? node4677 : node4674;
													assign node4674 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node4677 = (inp[9]) ? node4679 : 4'b0011;
														assign node4679 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node4682 = (inp[9]) ? node4684 : 4'b0111;
													assign node4684 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node4687 = (inp[12]) ? node4689 : 4'b0111;
												assign node4689 = (inp[1]) ? node4695 : node4690;
													assign node4690 = (inp[5]) ? node4692 : 4'b0011;
														assign node4692 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node4695 = (inp[5]) ? node4697 : 4'b0010;
														assign node4697 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node4700 = (inp[9]) ? node4712 : node4701;
											assign node4701 = (inp[12]) ? node4703 : 4'b0010;
												assign node4703 = (inp[1]) ? node4709 : node4704;
													assign node4704 = (inp[13]) ? node4706 : 4'b0011;
														assign node4706 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node4709 = (inp[15]) ? 4'b0010 : 4'b0110;
											assign node4712 = (inp[10]) ? 4'b0010 : node4713;
												assign node4713 = (inp[12]) ? node4719 : node4714;
													assign node4714 = (inp[13]) ? node4716 : 4'b0011;
														assign node4716 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node4719 = (inp[13]) ? 4'b0010 : node4720;
														assign node4720 = (inp[15]) ? 4'b0110 : 4'b0111;
									assign node4725 = (inp[13]) ? node4751 : node4726;
										assign node4726 = (inp[10]) ? node4736 : node4727;
											assign node4727 = (inp[12]) ? node4731 : node4728;
												assign node4728 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node4731 = (inp[15]) ? node4733 : 4'b0010;
													assign node4733 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node4736 = (inp[1]) ? node4740 : node4737;
												assign node4737 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node4740 = (inp[12]) ? node4748 : node4741;
													assign node4741 = (inp[9]) ? node4745 : node4742;
														assign node4742 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node4745 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node4748 = (inp[15]) ? 4'b0010 : 4'b0011;
										assign node4751 = (inp[1]) ? node4757 : node4752;
											assign node4752 = (inp[12]) ? node4754 : 4'b0011;
												assign node4754 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node4757 = (inp[12]) ? 4'b0011 : 4'b0111;
							assign node4760 = (inp[2]) ? node4814 : node4761;
								assign node4761 = (inp[8]) ? node4795 : node4762;
									assign node4762 = (inp[1]) ? node4774 : node4763;
										assign node4763 = (inp[11]) ? node4769 : node4764;
											assign node4764 = (inp[15]) ? node4766 : 4'b0110;
												assign node4766 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node4769 = (inp[9]) ? node4771 : 4'b0110;
												assign node4771 = (inp[12]) ? 4'b0110 : 4'b0111;
										assign node4774 = (inp[11]) ? node4786 : node4775;
											assign node4775 = (inp[13]) ? node4783 : node4776;
												assign node4776 = (inp[10]) ? 4'b0111 : node4777;
													assign node4777 = (inp[9]) ? 4'b0110 : node4778;
														assign node4778 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node4783 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node4786 = (inp[13]) ? node4790 : node4787;
												assign node4787 = (inp[12]) ? 4'b0111 : 4'b0010;
												assign node4790 = (inp[12]) ? node4792 : 4'b0111;
													assign node4792 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node4795 = (inp[15]) ? node4809 : node4796;
										assign node4796 = (inp[12]) ? node4804 : node4797;
											assign node4797 = (inp[1]) ? node4799 : 4'b0011;
												assign node4799 = (inp[5]) ? node4801 : 4'b0111;
													assign node4801 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node4804 = (inp[1]) ? 4'b0011 : node4805;
												assign node4805 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node4809 = (inp[12]) ? 4'b0111 : node4810;
											assign node4810 = (inp[1]) ? 4'b0111 : 4'b0011;
								assign node4814 = (inp[8]) ? node4870 : node4815;
									assign node4815 = (inp[9]) ? node4845 : node4816;
										assign node4816 = (inp[5]) ? node4826 : node4817;
											assign node4817 = (inp[12]) ? node4821 : node4818;
												assign node4818 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node4821 = (inp[15]) ? 4'b0010 : node4822;
													assign node4822 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node4826 = (inp[11]) ? node4838 : node4827;
												assign node4827 = (inp[15]) ? node4833 : node4828;
													assign node4828 = (inp[1]) ? node4830 : 4'b0111;
														assign node4830 = (inp[12]) ? 4'b0011 : 4'b0011;
													assign node4833 = (inp[13]) ? 4'b0111 : node4834;
														assign node4834 = (inp[10]) ? 4'b0010 : 4'b0111;
												assign node4838 = (inp[15]) ? 4'b0111 : node4839;
													assign node4839 = (inp[13]) ? 4'b0010 : node4840;
														assign node4840 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node4845 = (inp[11]) ? node4855 : node4846;
											assign node4846 = (inp[15]) ? 4'b0110 : node4847;
												assign node4847 = (inp[1]) ? 4'b0010 : node4848;
													assign node4848 = (inp[12]) ? 4'b0110 : node4849;
														assign node4849 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node4855 = (inp[13]) ? node4865 : node4856;
												assign node4856 = (inp[5]) ? node4860 : node4857;
													assign node4857 = (inp[15]) ? 4'b0011 : 4'b0111;
													assign node4860 = (inp[12]) ? node4862 : 4'b0010;
														assign node4862 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node4865 = (inp[5]) ? node4867 : 4'b0110;
													assign node4867 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node4870 = (inp[10]) ? node4886 : node4871;
										assign node4871 = (inp[1]) ? node4883 : node4872;
											assign node4872 = (inp[12]) ? node4876 : node4873;
												assign node4873 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node4876 = (inp[5]) ? 4'b0110 : node4877;
													assign node4877 = (inp[11]) ? 4'b0111 : node4878;
														assign node4878 = (inp[15]) ? 4'b0110 : 4'b0110;
											assign node4883 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node4886 = (inp[5]) ? node4888 : 4'b0010;
											assign node4888 = (inp[1]) ? node4892 : node4889;
												assign node4889 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node4892 = (inp[12]) ? node4896 : node4893;
													assign node4893 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node4896 = (inp[9]) ? node4898 : 4'b0010;
														assign node4898 = (inp[15]) ? 4'b0010 : 4'b0011;
					assign node4901 = (inp[7]) ? node5235 : node4902;
						assign node4902 = (inp[8]) ? node5072 : node4903;
							assign node4903 = (inp[11]) ? node4983 : node4904;
								assign node4904 = (inp[1]) ? node4944 : node4905;
									assign node4905 = (inp[9]) ? node4927 : node4906;
										assign node4906 = (inp[12]) ? node4914 : node4907;
											assign node4907 = (inp[5]) ? node4909 : 4'b0110;
												assign node4909 = (inp[13]) ? 4'b0111 : node4910;
													assign node4910 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node4914 = (inp[13]) ? node4920 : node4915;
												assign node4915 = (inp[0]) ? 4'b0010 : node4916;
													assign node4916 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node4920 = (inp[15]) ? 4'b0010 : node4921;
													assign node4921 = (inp[5]) ? 4'b0110 : node4922;
														assign node4922 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node4927 = (inp[0]) ? node4929 : 4'b0010;
											assign node4929 = (inp[2]) ? node4939 : node4930;
												assign node4930 = (inp[10]) ? node4934 : node4931;
													assign node4931 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node4934 = (inp[5]) ? node4936 : 4'b0111;
														assign node4936 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node4939 = (inp[12]) ? node4941 : 4'b0011;
													assign node4941 = (inp[10]) ? 4'b0010 : 4'b0110;
									assign node4944 = (inp[15]) ? node4964 : node4945;
										assign node4945 = (inp[13]) ? node4955 : node4946;
											assign node4946 = (inp[12]) ? node4948 : 4'b0010;
												assign node4948 = (inp[0]) ? node4950 : 4'b0010;
													assign node4950 = (inp[5]) ? node4952 : 4'b0011;
														assign node4952 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node4955 = (inp[9]) ? node4961 : node4956;
												assign node4956 = (inp[5]) ? node4958 : 4'b0110;
													assign node4958 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node4961 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node4964 = (inp[13]) ? node4972 : node4965;
											assign node4965 = (inp[10]) ? node4967 : 4'b0111;
												assign node4967 = (inp[0]) ? node4969 : 4'b0110;
													assign node4969 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node4972 = (inp[5]) ? node4980 : node4973;
												assign node4973 = (inp[2]) ? 4'b0010 : node4974;
													assign node4974 = (inp[9]) ? 4'b0011 : node4975;
														assign node4975 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node4980 = (inp[9]) ? 4'b0010 : 4'b0011;
								assign node4983 = (inp[10]) ? node5033 : node4984;
									assign node4984 = (inp[12]) ? node5002 : node4985;
										assign node4985 = (inp[0]) ? node4991 : node4986;
											assign node4986 = (inp[5]) ? node4988 : 4'b0111;
												assign node4988 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node4991 = (inp[1]) ? node4993 : 4'b0010;
												assign node4993 = (inp[9]) ? 4'b0110 : node4994;
													assign node4994 = (inp[15]) ? node4998 : node4995;
														assign node4995 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node4998 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node5002 = (inp[15]) ? node5020 : node5003;
											assign node5003 = (inp[13]) ? node5011 : node5004;
												assign node5004 = (inp[2]) ? 4'b0011 : node5005;
													assign node5005 = (inp[5]) ? node5007 : 4'b0010;
														assign node5007 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node5011 = (inp[0]) ? node5013 : 4'b0111;
													assign node5013 = (inp[5]) ? node5017 : node5014;
														assign node5014 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node5017 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node5020 = (inp[13]) ? node5026 : node5021;
												assign node5021 = (inp[9]) ? node5023 : 4'b0111;
													assign node5023 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node5026 = (inp[9]) ? 4'b0010 : node5027;
													assign node5027 = (inp[5]) ? node5029 : 4'b0010;
														assign node5029 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node5033 = (inp[0]) ? node5049 : node5034;
										assign node5034 = (inp[1]) ? node5046 : node5035;
											assign node5035 = (inp[9]) ? 4'b0010 : node5036;
												assign node5036 = (inp[12]) ? 4'b0011 : node5037;
													assign node5037 = (inp[15]) ? node5041 : node5038;
														assign node5038 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node5041 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node5046 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node5049 = (inp[15]) ? node5059 : node5050;
											assign node5050 = (inp[13]) ? 4'b0111 : node5051;
												assign node5051 = (inp[12]) ? node5053 : 4'b0011;
													assign node5053 = (inp[9]) ? 4'b0011 : node5054;
														assign node5054 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node5059 = (inp[13]) ? node5065 : node5060;
												assign node5060 = (inp[5]) ? node5062 : 4'b0111;
													assign node5062 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node5065 = (inp[2]) ? node5067 : 4'b0010;
													assign node5067 = (inp[9]) ? node5069 : 4'b0011;
														assign node5069 = (inp[5]) ? 4'b0010 : 4'b0011;
							assign node5072 = (inp[2]) ? node5154 : node5073;
								assign node5073 = (inp[0]) ? node5105 : node5074;
									assign node5074 = (inp[5]) ? node5088 : node5075;
										assign node5075 = (inp[12]) ? node5083 : node5076;
											assign node5076 = (inp[15]) ? node5078 : 4'b0000;
												assign node5078 = (inp[11]) ? node5080 : 4'b0101;
													assign node5080 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node5083 = (inp[10]) ? node5085 : 4'b0100;
												assign node5085 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node5088 = (inp[12]) ? node5096 : node5089;
											assign node5089 = (inp[15]) ? node5093 : node5090;
												assign node5090 = (inp[1]) ? 4'b0101 : 4'b0001;
												assign node5093 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node5096 = (inp[15]) ? node5102 : node5097;
												assign node5097 = (inp[10]) ? node5099 : 4'b0001;
													assign node5099 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node5102 = (inp[1]) ? 4'b0001 : 4'b0101;
									assign node5105 = (inp[9]) ? node5139 : node5106;
										assign node5106 = (inp[10]) ? node5128 : node5107;
											assign node5107 = (inp[13]) ? node5119 : node5108;
												assign node5108 = (inp[1]) ? node5114 : node5109;
													assign node5109 = (inp[15]) ? 4'b0100 : node5110;
														assign node5110 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node5114 = (inp[5]) ? 4'b0101 : node5115;
														assign node5115 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node5119 = (inp[11]) ? node5125 : node5120;
													assign node5120 = (inp[5]) ? 4'b0001 : node5121;
														assign node5121 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node5125 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node5128 = (inp[12]) ? node5130 : 4'b0101;
												assign node5130 = (inp[13]) ? node5134 : node5131;
													assign node5131 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node5134 = (inp[11]) ? node5136 : 4'b0000;
														assign node5136 = (inp[5]) ? 4'b0000 : 4'b0101;
										assign node5139 = (inp[12]) ? node5145 : node5140;
											assign node5140 = (inp[15]) ? node5142 : 4'b0001;
												assign node5142 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node5145 = (inp[5]) ? node5149 : node5146;
												assign node5146 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node5149 = (inp[13]) ? 4'b0100 : node5150;
													assign node5150 = (inp[15]) ? 4'b0100 : 4'b0101;
								assign node5154 = (inp[10]) ? node5198 : node5155;
									assign node5155 = (inp[11]) ? node5177 : node5156;
										assign node5156 = (inp[12]) ? node5166 : node5157;
											assign node5157 = (inp[9]) ? 4'b0100 : node5158;
												assign node5158 = (inp[1]) ? 4'b0000 : node5159;
													assign node5159 = (inp[5]) ? 4'b0000 : node5160;
														assign node5160 = (inp[15]) ? 4'b0101 : 4'b0001;
											assign node5166 = (inp[1]) ? node5174 : node5167;
												assign node5167 = (inp[15]) ? node5169 : 4'b0001;
													assign node5169 = (inp[5]) ? 4'b0101 : node5170;
														assign node5170 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node5174 = (inp[15]) ? 4'b0001 : 4'b0101;
										assign node5177 = (inp[12]) ? node5189 : node5178;
											assign node5178 = (inp[13]) ? node5184 : node5179;
												assign node5179 = (inp[1]) ? node5181 : 4'b0101;
													assign node5181 = (inp[0]) ? 4'b0001 : 4'b0101;
												assign node5184 = (inp[0]) ? node5186 : 4'b0000;
													assign node5186 = (inp[15]) ? 4'b0100 : 4'b0001;
											assign node5189 = (inp[5]) ? 4'b0000 : node5190;
												assign node5190 = (inp[0]) ? 4'b0001 : node5191;
													assign node5191 = (inp[15]) ? 4'b0100 : node5192;
														assign node5192 = (inp[9]) ? 4'b0001 : 4'b0000;
									assign node5198 = (inp[1]) ? node5214 : node5199;
										assign node5199 = (inp[15]) ? node5201 : 4'b0001;
											assign node5201 = (inp[13]) ? node5207 : node5202;
												assign node5202 = (inp[0]) ? 4'b0101 : node5203;
													assign node5203 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node5207 = (inp[0]) ? 4'b0100 : node5208;
													assign node5208 = (inp[11]) ? 4'b0101 : node5209;
														assign node5209 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node5214 = (inp[15]) ? node5224 : node5215;
											assign node5215 = (inp[5]) ? node5219 : node5216;
												assign node5216 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node5219 = (inp[0]) ? 4'b0100 : node5220;
													assign node5220 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node5224 = (inp[9]) ? node5230 : node5225;
												assign node5225 = (inp[5]) ? 4'b0001 : node5226;
													assign node5226 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node5230 = (inp[5]) ? 4'b0000 : node5231;
													assign node5231 = (inp[11]) ? 4'b0001 : 4'b0000;
						assign node5235 = (inp[1]) ? node5321 : node5236;
							assign node5236 = (inp[8]) ? node5292 : node5237;
								assign node5237 = (inp[13]) ? node5261 : node5238;
									assign node5238 = (inp[11]) ? node5248 : node5239;
										assign node5239 = (inp[10]) ? node5241 : 4'b0000;
											assign node5241 = (inp[15]) ? 4'b0000 : node5242;
												assign node5242 = (inp[0]) ? node5244 : 4'b0001;
													assign node5244 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node5248 = (inp[0]) ? node5256 : node5249;
											assign node5249 = (inp[12]) ? node5253 : node5250;
												assign node5250 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node5253 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node5256 = (inp[10]) ? 4'b0001 : node5257;
												assign node5257 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node5261 = (inp[15]) ? node5275 : node5262;
										assign node5262 = (inp[5]) ? node5268 : node5263;
											assign node5263 = (inp[12]) ? 4'b0100 : node5264;
												assign node5264 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node5268 = (inp[12]) ? node5272 : node5269;
												assign node5269 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node5272 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node5275 = (inp[12]) ? node5283 : node5276;
											assign node5276 = (inp[5]) ? 4'b0100 : node5277;
												assign node5277 = (inp[2]) ? 4'b0101 : node5278;
													assign node5278 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node5283 = (inp[5]) ? node5285 : 4'b0100;
												assign node5285 = (inp[11]) ? 4'b0101 : node5286;
													assign node5286 = (inp[0]) ? 4'b0100 : node5287;
														assign node5287 = (inp[9]) ? 4'b0101 : 4'b0100;
								assign node5292 = (inp[2]) ? node5300 : node5293;
									assign node5293 = (inp[12]) ? node5297 : node5294;
										assign node5294 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node5297 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node5300 = (inp[13]) ? node5314 : node5301;
										assign node5301 = (inp[9]) ? node5307 : node5302;
											assign node5302 = (inp[0]) ? 4'b0100 : node5303;
												assign node5303 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node5307 = (inp[0]) ? node5311 : node5308;
												assign node5308 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node5311 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node5314 = (inp[0]) ? node5318 : node5315;
											assign node5315 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node5318 = (inp[12]) ? 4'b0100 : 4'b0101;
							assign node5321 = (inp[13]) ? node5355 : node5322;
								assign node5322 = (inp[8]) ? node5330 : node5323;
									assign node5323 = (inp[15]) ? node5327 : node5324;
										assign node5324 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node5327 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node5330 = (inp[12]) ? node5338 : node5331;
										assign node5331 = (inp[15]) ? node5335 : node5332;
											assign node5332 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node5335 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node5338 = (inp[9]) ? node5346 : node5339;
											assign node5339 = (inp[5]) ? node5341 : 4'b0000;
												assign node5341 = (inp[0]) ? node5343 : 4'b0000;
													assign node5343 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node5346 = (inp[10]) ? node5348 : 4'b0000;
												assign node5348 = (inp[11]) ? node5350 : 4'b0001;
													assign node5350 = (inp[0]) ? 4'b0000 : node5351;
														assign node5351 = (inp[15]) ? 4'b0001 : 4'b0000;
								assign node5355 = (inp[0]) ? node5361 : node5356;
									assign node5356 = (inp[9]) ? 4'b0001 : node5357;
										assign node5357 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node5361 = (inp[9]) ? 4'b0000 : node5362;
										assign node5362 = (inp[8]) ? 4'b0000 : 4'b0001;
		assign node5366 = (inp[14]) ? node7618 : node5367;
			assign node5367 = (inp[8]) ? node6705 : node5368;
				assign node5368 = (inp[5]) ? node6052 : node5369;
					assign node5369 = (inp[13]) ? node5713 : node5370;
						assign node5370 = (inp[6]) ? node5572 : node5371;
							assign node5371 = (inp[9]) ? node5479 : node5372;
								assign node5372 = (inp[11]) ? node5420 : node5373;
									assign node5373 = (inp[1]) ? node5401 : node5374;
										assign node5374 = (inp[4]) ? node5388 : node5375;
											assign node5375 = (inp[15]) ? node5385 : node5376;
												assign node5376 = (inp[2]) ? node5382 : node5377;
													assign node5377 = (inp[10]) ? node5379 : 4'b1010;
														assign node5379 = (inp[7]) ? 4'b1010 : 4'b1001;
													assign node5382 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node5385 = (inp[0]) ? 4'b1011 : 4'b1111;
											assign node5388 = (inp[7]) ? 4'b1111 : node5389;
												assign node5389 = (inp[15]) ? node5395 : node5390;
													assign node5390 = (inp[12]) ? 4'b1100 : node5391;
														assign node5391 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node5395 = (inp[10]) ? node5397 : 4'b1010;
														assign node5397 = (inp[2]) ? 4'b1000 : 4'b1101;
										assign node5401 = (inp[4]) ? node5407 : node5402;
											assign node5402 = (inp[10]) ? 4'b1101 : node5403;
												assign node5403 = (inp[15]) ? 4'b1100 : 4'b1000;
											assign node5407 = (inp[10]) ? 4'b1001 : node5408;
												assign node5408 = (inp[0]) ? node5414 : node5409;
													assign node5409 = (inp[7]) ? 4'b1101 : node5410;
														assign node5410 = (inp[2]) ? 4'b1011 : 4'b1110;
													assign node5414 = (inp[7]) ? node5416 : 4'b1101;
														assign node5416 = (inp[12]) ? 4'b1111 : 4'b1101;
									assign node5420 = (inp[10]) ? node5450 : node5421;
										assign node5421 = (inp[0]) ? node5435 : node5422;
											assign node5422 = (inp[12]) ? node5430 : node5423;
												assign node5423 = (inp[1]) ? node5425 : 4'b1010;
													assign node5425 = (inp[2]) ? 4'b1010 : node5426;
														assign node5426 = (inp[15]) ? 4'b1111 : 4'b1011;
												assign node5430 = (inp[4]) ? node5432 : 4'b1010;
													assign node5432 = (inp[1]) ? 4'b1100 : 4'b1110;
											assign node5435 = (inp[4]) ? node5445 : node5436;
												assign node5436 = (inp[2]) ? node5442 : node5437;
													assign node5437 = (inp[15]) ? 4'b1000 : node5438;
														assign node5438 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node5442 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node5445 = (inp[12]) ? 4'b1001 : node5446;
													assign node5446 = (inp[7]) ? 4'b1000 : 4'b1010;
										assign node5450 = (inp[1]) ? node5460 : node5451;
											assign node5451 = (inp[2]) ? node5455 : node5452;
												assign node5452 = (inp[12]) ? 4'b1010 : 4'b1001;
												assign node5455 = (inp[4]) ? node5457 : 4'b1111;
													assign node5457 = (inp[15]) ? 4'b1111 : 4'b1001;
											assign node5460 = (inp[2]) ? node5464 : node5461;
												assign node5461 = (inp[12]) ? 4'b1110 : 4'b1101;
												assign node5464 = (inp[7]) ? node5472 : node5465;
													assign node5465 = (inp[15]) ? node5469 : node5466;
														assign node5466 = (inp[4]) ? 4'b1000 : 4'b1000;
														assign node5469 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node5472 = (inp[4]) ? node5476 : node5473;
														assign node5473 = (inp[12]) ? 4'b1101 : 4'b1110;
														assign node5476 = (inp[12]) ? 4'b1010 : 4'b1111;
								assign node5479 = (inp[2]) ? node5527 : node5480;
									assign node5480 = (inp[1]) ? node5506 : node5481;
										assign node5481 = (inp[11]) ? node5495 : node5482;
											assign node5482 = (inp[7]) ? node5490 : node5483;
												assign node5483 = (inp[12]) ? node5487 : node5484;
													assign node5484 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node5487 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node5490 = (inp[15]) ? node5492 : 4'b1101;
													assign node5492 = (inp[12]) ? 4'b1001 : 4'b1010;
											assign node5495 = (inp[10]) ? node5499 : node5496;
												assign node5496 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node5499 = (inp[12]) ? 4'b1100 : node5500;
													assign node5500 = (inp[7]) ? node5502 : 4'b1000;
														assign node5502 = (inp[0]) ? 4'b1110 : 4'b1010;
										assign node5506 = (inp[7]) ? node5516 : node5507;
											assign node5507 = (inp[10]) ? 4'b1100 : node5508;
												assign node5508 = (inp[11]) ? node5510 : 4'b1111;
													assign node5510 = (inp[12]) ? 4'b1100 : node5511;
														assign node5511 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node5516 = (inp[15]) ? node5522 : node5517;
												assign node5517 = (inp[12]) ? 4'b1000 : node5518;
													assign node5518 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node5522 = (inp[12]) ? node5524 : 4'b1111;
													assign node5524 = (inp[4]) ? 4'b1100 : 4'b1101;
									assign node5527 = (inp[1]) ? node5543 : node5528;
										assign node5528 = (inp[7]) ? node5534 : node5529;
											assign node5529 = (inp[12]) ? 4'b1001 : node5530;
												assign node5530 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node5534 = (inp[10]) ? node5538 : node5535;
												assign node5535 = (inp[11]) ? 4'b1111 : 4'b1101;
												assign node5538 = (inp[11]) ? 4'b1011 : node5539;
													assign node5539 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node5543 = (inp[10]) ? node5561 : node5544;
											assign node5544 = (inp[0]) ? node5554 : node5545;
												assign node5545 = (inp[15]) ? node5549 : node5546;
													assign node5546 = (inp[11]) ? 4'b1000 : 4'b1010;
													assign node5549 = (inp[11]) ? 4'b1000 : node5550;
														assign node5550 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node5554 = (inp[7]) ? node5556 : 4'b1001;
													assign node5556 = (inp[4]) ? node5558 : 4'b1010;
														assign node5558 = (inp[11]) ? 4'b1010 : 4'b1100;
											assign node5561 = (inp[11]) ? node5569 : node5562;
												assign node5562 = (inp[4]) ? node5564 : 4'b1011;
													assign node5564 = (inp[12]) ? node5566 : 4'b1101;
														assign node5566 = (inp[7]) ? 4'b1011 : 4'b1000;
												assign node5569 = (inp[7]) ? 4'b1010 : 4'b1001;
							assign node5572 = (inp[12]) ? node5652 : node5573;
								assign node5573 = (inp[15]) ? node5617 : node5574;
									assign node5574 = (inp[7]) ? node5598 : node5575;
										assign node5575 = (inp[11]) ? node5585 : node5576;
											assign node5576 = (inp[4]) ? node5580 : node5577;
												assign node5577 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node5580 = (inp[9]) ? 4'b1001 : node5581;
													assign node5581 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node5585 = (inp[10]) ? node5591 : node5586;
												assign node5586 = (inp[0]) ? 4'b1000 : node5587;
													assign node5587 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node5591 = (inp[9]) ? 4'b1000 : node5592;
													assign node5592 = (inp[1]) ? 4'b1001 : node5593;
														assign node5593 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node5598 = (inp[4]) ? node5608 : node5599;
											assign node5599 = (inp[2]) ? node5603 : node5600;
												assign node5600 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5603 = (inp[9]) ? 4'b1011 : node5604;
													assign node5604 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node5608 = (inp[1]) ? 4'b1011 : node5609;
												assign node5609 = (inp[0]) ? node5611 : 4'b1111;
													assign node5611 = (inp[9]) ? 4'b1111 : node5612;
														assign node5612 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node5617 = (inp[7]) ? node5637 : node5618;
										assign node5618 = (inp[4]) ? node5630 : node5619;
											assign node5619 = (inp[1]) ? node5621 : 4'b1011;
												assign node5621 = (inp[0]) ? node5623 : 4'b1111;
													assign node5623 = (inp[2]) ? node5627 : node5624;
														assign node5624 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node5627 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node5630 = (inp[1]) ? node5632 : 4'b1110;
												assign node5632 = (inp[9]) ? 4'b1011 : node5633;
													assign node5633 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node5637 = (inp[4]) ? node5647 : node5638;
											assign node5638 = (inp[1]) ? 4'b1101 : node5639;
												assign node5639 = (inp[9]) ? node5641 : 4'b1001;
													assign node5641 = (inp[0]) ? 4'b1000 : node5642;
														assign node5642 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node5647 = (inp[1]) ? 4'b1000 : node5648;
												assign node5648 = (inp[2]) ? 4'b1101 : 4'b1100;
								assign node5652 = (inp[15]) ? node5678 : node5653;
									assign node5653 = (inp[7]) ? node5665 : node5654;
										assign node5654 = (inp[0]) ? node5662 : node5655;
											assign node5655 = (inp[11]) ? 4'b1000 : node5656;
												assign node5656 = (inp[9]) ? node5658 : 4'b1000;
													assign node5658 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node5662 = (inp[1]) ? 4'b1101 : 4'b1000;
										assign node5665 = (inp[1]) ? node5673 : node5666;
											assign node5666 = (inp[4]) ? node5668 : 4'b1111;
												assign node5668 = (inp[9]) ? node5670 : 4'b1011;
													assign node5670 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node5673 = (inp[11]) ? node5675 : 4'b1010;
												assign node5675 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node5678 = (inp[7]) ? node5698 : node5679;
										assign node5679 = (inp[4]) ? node5689 : node5680;
											assign node5680 = (inp[1]) ? 4'b1010 : node5681;
												assign node5681 = (inp[0]) ? 4'b1011 : node5682;
													assign node5682 = (inp[11]) ? 4'b1010 : node5683;
														assign node5683 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node5689 = (inp[2]) ? node5691 : 4'b1011;
												assign node5691 = (inp[11]) ? node5693 : 4'b1011;
													assign node5693 = (inp[9]) ? 4'b1010 : node5694;
														assign node5694 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node5698 = (inp[0]) ? node5706 : node5699;
											assign node5699 = (inp[9]) ? node5703 : node5700;
												assign node5700 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node5703 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node5706 = (inp[1]) ? 4'b1001 : node5707;
												assign node5707 = (inp[4]) ? node5709 : 4'b1001;
													assign node5709 = (inp[11]) ? 4'b1001 : 4'b1000;
						assign node5713 = (inp[6]) ? node5911 : node5714;
							assign node5714 = (inp[10]) ? node5810 : node5715;
								assign node5715 = (inp[9]) ? node5755 : node5716;
									assign node5716 = (inp[1]) ? node5738 : node5717;
										assign node5717 = (inp[15]) ? node5725 : node5718;
											assign node5718 = (inp[0]) ? 4'b1011 : node5719;
												assign node5719 = (inp[2]) ? 4'b1100 : node5720;
													assign node5720 = (inp[12]) ? 4'b1111 : 4'b1101;
											assign node5725 = (inp[12]) ? node5731 : node5726;
												assign node5726 = (inp[2]) ? node5728 : 4'b1000;
													assign node5728 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node5731 = (inp[7]) ? node5735 : node5732;
													assign node5732 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node5735 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node5738 = (inp[7]) ? node5748 : node5739;
											assign node5739 = (inp[2]) ? 4'b1111 : node5740;
												assign node5740 = (inp[11]) ? node5742 : 4'b1000;
													assign node5742 = (inp[4]) ? 4'b1011 : node5743;
														assign node5743 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node5748 = (inp[12]) ? 4'b1110 : node5749;
												assign node5749 = (inp[4]) ? 4'b1010 : node5750;
													assign node5750 = (inp[11]) ? 4'b1010 : 4'b1110;
									assign node5755 = (inp[11]) ? node5781 : node5756;
										assign node5756 = (inp[12]) ? node5768 : node5757;
											assign node5757 = (inp[7]) ? node5763 : node5758;
												assign node5758 = (inp[0]) ? node5760 : 4'b1001;
													assign node5760 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node5763 = (inp[0]) ? node5765 : 4'b1011;
													assign node5765 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node5768 = (inp[7]) ? node5776 : node5769;
												assign node5769 = (inp[15]) ? node5773 : node5770;
													assign node5770 = (inp[0]) ? 4'b1001 : 4'b1111;
													assign node5773 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5776 = (inp[1]) ? node5778 : 4'b1001;
													assign node5778 = (inp[0]) ? 4'b1110 : 4'b1000;
										assign node5781 = (inp[0]) ? node5797 : node5782;
											assign node5782 = (inp[2]) ? node5788 : node5783;
												assign node5783 = (inp[4]) ? 4'b1010 : node5784;
													assign node5784 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node5788 = (inp[1]) ? node5790 : 4'b1001;
													assign node5790 = (inp[4]) ? node5794 : node5791;
														assign node5791 = (inp[12]) ? 4'b1100 : 4'b1100;
														assign node5794 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node5797 = (inp[7]) ? 4'b1001 : node5798;
												assign node5798 = (inp[12]) ? node5802 : node5799;
													assign node5799 = (inp[4]) ? 4'b1011 : 4'b1100;
													assign node5802 = (inp[2]) ? node5806 : node5803;
														assign node5803 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node5806 = (inp[15]) ? 4'b1011 : 4'b1010;
								assign node5810 = (inp[1]) ? node5856 : node5811;
									assign node5811 = (inp[2]) ? node5841 : node5812;
										assign node5812 = (inp[4]) ? node5824 : node5813;
											assign node5813 = (inp[9]) ? node5819 : node5814;
												assign node5814 = (inp[7]) ? node5816 : 4'b1110;
													assign node5816 = (inp[11]) ? 4'b1101 : 4'b1111;
												assign node5819 = (inp[11]) ? node5821 : 4'b1100;
													assign node5821 = (inp[0]) ? 4'b1001 : 4'b1101;
											assign node5824 = (inp[12]) ? node5834 : node5825;
												assign node5825 = (inp[0]) ? 4'b1000 : node5826;
													assign node5826 = (inp[15]) ? node5830 : node5827;
														assign node5827 = (inp[11]) ? 4'b1001 : 4'b1110;
														assign node5830 = (inp[7]) ? 4'b1111 : 4'b1001;
												assign node5834 = (inp[11]) ? node5836 : 4'b1110;
													assign node5836 = (inp[15]) ? node5838 : 4'b1000;
														assign node5838 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node5841 = (inp[7]) ? node5849 : node5842;
											assign node5842 = (inp[12]) ? 4'b1011 : node5843;
												assign node5843 = (inp[15]) ? node5845 : 4'b1011;
													assign node5845 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node5849 = (inp[15]) ? node5851 : 4'b1101;
												assign node5851 = (inp[12]) ? node5853 : 4'b1010;
													assign node5853 = (inp[4]) ? 4'b1000 : 4'b1001;
									assign node5856 = (inp[2]) ? node5880 : node5857;
										assign node5857 = (inp[0]) ? node5867 : node5858;
											assign node5858 = (inp[9]) ? node5864 : node5859;
												assign node5859 = (inp[11]) ? 4'b1100 : node5860;
													assign node5860 = (inp[12]) ? 4'b1101 : 4'b1110;
												assign node5864 = (inp[15]) ? 4'b1001 : 4'b1101;
											assign node5867 = (inp[7]) ? node5871 : node5868;
												assign node5868 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node5871 = (inp[12]) ? node5877 : node5872;
													assign node5872 = (inp[11]) ? node5874 : 4'b1011;
														assign node5874 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node5877 = (inp[4]) ? 4'b1011 : 4'b1001;
										assign node5880 = (inp[4]) ? node5898 : node5881;
											assign node5881 = (inp[12]) ? node5891 : node5882;
												assign node5882 = (inp[7]) ? node5888 : node5883;
													assign node5883 = (inp[15]) ? 4'b1100 : node5884;
														assign node5884 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node5888 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node5891 = (inp[7]) ? 4'b1101 : node5892;
													assign node5892 = (inp[11]) ? node5894 : 4'b1110;
														assign node5894 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5898 = (inp[15]) ? node5906 : node5899;
												assign node5899 = (inp[7]) ? node5903 : node5900;
													assign node5900 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node5903 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node5906 = (inp[9]) ? 4'b1111 : node5907;
													assign node5907 = (inp[0]) ? 4'b1111 : 4'b1110;
							assign node5911 = (inp[12]) ? node5997 : node5912;
								assign node5912 = (inp[15]) ? node5956 : node5913;
									assign node5913 = (inp[7]) ? node5931 : node5914;
										assign node5914 = (inp[1]) ? node5922 : node5915;
											assign node5915 = (inp[2]) ? 4'b1100 : node5916;
												assign node5916 = (inp[0]) ? node5918 : 4'b1101;
													assign node5918 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node5922 = (inp[4]) ? node5926 : node5923;
												assign node5923 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node5926 = (inp[2]) ? node5928 : 4'b1101;
													assign node5928 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node5931 = (inp[4]) ? node5945 : node5932;
											assign node5932 = (inp[2]) ? node5940 : node5933;
												assign node5933 = (inp[0]) ? 4'b1110 : node5934;
													assign node5934 = (inp[10]) ? node5936 : 4'b1111;
														assign node5936 = (inp[11]) ? 4'b1110 : 4'b1110;
												assign node5940 = (inp[11]) ? 4'b1111 : node5941;
													assign node5941 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node5945 = (inp[1]) ? node5949 : node5946;
												assign node5946 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node5949 = (inp[10]) ? node5951 : 4'b1110;
													assign node5951 = (inp[9]) ? node5953 : 4'b1111;
														assign node5953 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node5956 = (inp[7]) ? node5976 : node5957;
										assign node5957 = (inp[0]) ? node5967 : node5958;
											assign node5958 = (inp[4]) ? 4'b1011 : node5959;
												assign node5959 = (inp[1]) ? 4'b1010 : node5960;
													assign node5960 = (inp[11]) ? 4'b1111 : node5961;
														assign node5961 = (inp[9]) ? 4'b1110 : 4'b1110;
											assign node5967 = (inp[4]) ? node5969 : 4'b1011;
												assign node5969 = (inp[1]) ? 4'b1110 : node5970;
													assign node5970 = (inp[9]) ? node5972 : 4'b1010;
														assign node5972 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node5976 = (inp[10]) ? node5986 : node5977;
											assign node5977 = (inp[11]) ? node5979 : 4'b1100;
												assign node5979 = (inp[9]) ? node5981 : 4'b1101;
													assign node5981 = (inp[1]) ? 4'b1000 : node5982;
														assign node5982 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node5986 = (inp[1]) ? node5992 : node5987;
												assign node5987 = (inp[4]) ? node5989 : 4'b1100;
													assign node5989 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node5992 = (inp[4]) ? 4'b1101 : node5993;
													assign node5993 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node5997 = (inp[15]) ? node6027 : node5998;
									assign node5998 = (inp[7]) ? node6012 : node5999;
										assign node5999 = (inp[4]) ? node6005 : node6000;
											assign node6000 = (inp[0]) ? node6002 : 4'b1101;
												assign node6002 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node6005 = (inp[0]) ? node6007 : 4'b1100;
												assign node6007 = (inp[11]) ? node6009 : 4'b1001;
													assign node6009 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node6012 = (inp[1]) ? node6020 : node6013;
											assign node6013 = (inp[4]) ? 4'b1111 : node6014;
												assign node6014 = (inp[9]) ? 4'b1011 : node6015;
													assign node6015 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node6020 = (inp[4]) ? node6022 : 4'b1110;
												assign node6022 = (inp[10]) ? 4'b1111 : node6023;
													assign node6023 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node6027 = (inp[7]) ? node6037 : node6028;
										assign node6028 = (inp[11]) ? 4'b1111 : node6029;
											assign node6029 = (inp[9]) ? 4'b1110 : node6030;
												assign node6030 = (inp[2]) ? 4'b1111 : node6031;
													assign node6031 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node6037 = (inp[10]) ? node6045 : node6038;
											assign node6038 = (inp[1]) ? 4'b1100 : node6039;
												assign node6039 = (inp[9]) ? 4'b1101 : node6040;
													assign node6040 = (inp[4]) ? 4'b1100 : 4'b1101;
											assign node6045 = (inp[2]) ? node6047 : 4'b1100;
												assign node6047 = (inp[9]) ? 4'b1100 : node6048;
													assign node6048 = (inp[1]) ? 4'b1101 : 4'b1100;
					assign node6052 = (inp[13]) ? node6390 : node6053;
						assign node6053 = (inp[2]) ? node6237 : node6054;
							assign node6054 = (inp[6]) ? node6158 : node6055;
								assign node6055 = (inp[9]) ? node6109 : node6056;
									assign node6056 = (inp[1]) ? node6086 : node6057;
										assign node6057 = (inp[15]) ? node6069 : node6058;
											assign node6058 = (inp[7]) ? node6066 : node6059;
												assign node6059 = (inp[11]) ? node6063 : node6060;
													assign node6060 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node6063 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node6066 = (inp[12]) ? 4'b1010 : 4'b1101;
											assign node6069 = (inp[10]) ? node6079 : node6070;
												assign node6070 = (inp[11]) ? 4'b1010 : node6071;
													assign node6071 = (inp[0]) ? node6075 : node6072;
														assign node6072 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node6075 = (inp[4]) ? 4'b1010 : 4'b1001;
												assign node6079 = (inp[4]) ? 4'b1000 : node6080;
													assign node6080 = (inp[0]) ? 4'b1001 : node6081;
														assign node6081 = (inp[7]) ? 4'b1010 : 4'b1001;
										assign node6086 = (inp[7]) ? node6098 : node6087;
											assign node6087 = (inp[12]) ? node6091 : node6088;
												assign node6088 = (inp[4]) ? 4'b1010 : 4'b1000;
												assign node6091 = (inp[4]) ? node6095 : node6092;
													assign node6092 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node6095 = (inp[11]) ? 4'b1011 : 4'b1101;
											assign node6098 = (inp[12]) ? node6106 : node6099;
												assign node6099 = (inp[15]) ? node6101 : 4'b1101;
													assign node6101 = (inp[11]) ? node6103 : 4'b1011;
														assign node6103 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node6106 = (inp[11]) ? 4'b1100 : 4'b1000;
									assign node6109 = (inp[12]) ? node6135 : node6110;
										assign node6110 = (inp[4]) ? node6122 : node6111;
											assign node6111 = (inp[7]) ? node6119 : node6112;
												assign node6112 = (inp[11]) ? 4'b1000 : node6113;
													assign node6113 = (inp[1]) ? 4'b1000 : node6114;
														assign node6114 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node6119 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node6122 = (inp[1]) ? node6130 : node6123;
												assign node6123 = (inp[0]) ? node6125 : 4'b1101;
													assign node6125 = (inp[7]) ? 4'b1100 : node6126;
														assign node6126 = (inp[10]) ? 4'b1100 : 4'b1011;
												assign node6130 = (inp[15]) ? node6132 : 4'b1011;
													assign node6132 = (inp[10]) ? 4'b1101 : 4'b1011;
										assign node6135 = (inp[0]) ? node6149 : node6136;
											assign node6136 = (inp[4]) ? node6144 : node6137;
												assign node6137 = (inp[7]) ? node6141 : node6138;
													assign node6138 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node6141 = (inp[1]) ? 4'b1000 : 4'b1101;
												assign node6144 = (inp[10]) ? 4'b1010 : node6145;
													assign node6145 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node6149 = (inp[7]) ? node6155 : node6150;
												assign node6150 = (inp[4]) ? node6152 : 4'b1010;
													assign node6152 = (inp[10]) ? 4'b1000 : 4'b1101;
												assign node6155 = (inp[11]) ? 4'b1000 : 4'b1100;
								assign node6158 = (inp[12]) ? node6202 : node6159;
									assign node6159 = (inp[15]) ? node6181 : node6160;
										assign node6160 = (inp[7]) ? node6172 : node6161;
											assign node6161 = (inp[1]) ? node6165 : node6162;
												assign node6162 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6165 = (inp[4]) ? node6167 : 4'b1000;
													assign node6167 = (inp[10]) ? 4'b1100 : node6168;
														assign node6168 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node6172 = (inp[0]) ? node6176 : node6173;
												assign node6173 = (inp[4]) ? 4'b1010 : 4'b1111;
												assign node6176 = (inp[1]) ? node6178 : 4'b1111;
													assign node6178 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node6181 = (inp[7]) ? node6187 : node6182;
											assign node6182 = (inp[1]) ? 4'b1010 : node6183;
												assign node6183 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node6187 = (inp[4]) ? node6193 : node6188;
												assign node6188 = (inp[0]) ? node6190 : 4'b1000;
													assign node6190 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node6193 = (inp[1]) ? 4'b1101 : node6194;
													assign node6194 = (inp[11]) ? node6198 : node6195;
														assign node6195 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node6198 = (inp[9]) ? 4'b1000 : 4'b1001;
									assign node6202 = (inp[10]) ? node6216 : node6203;
										assign node6203 = (inp[15]) ? node6207 : node6204;
											assign node6204 = (inp[7]) ? 4'b1110 : 4'b1100;
											assign node6207 = (inp[7]) ? node6211 : node6208;
												assign node6208 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node6211 = (inp[4]) ? node6213 : 4'b1100;
													assign node6213 = (inp[1]) ? 4'b1100 : 4'b1101;
										assign node6216 = (inp[7]) ? node6228 : node6217;
											assign node6217 = (inp[15]) ? node6225 : node6218;
												assign node6218 = (inp[11]) ? node6222 : node6219;
													assign node6219 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node6222 = (inp[0]) ? 4'b1000 : 4'b1100;
												assign node6225 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node6228 = (inp[15]) ? 4'b1101 : node6229;
												assign node6229 = (inp[0]) ? 4'b1110 : node6230;
													assign node6230 = (inp[1]) ? 4'b1111 : node6231;
														assign node6231 = (inp[9]) ? 4'b1010 : 4'b1011;
							assign node6237 = (inp[7]) ? node6311 : node6238;
								assign node6238 = (inp[15]) ? node6272 : node6239;
									assign node6239 = (inp[11]) ? node6257 : node6240;
										assign node6240 = (inp[6]) ? node6250 : node6241;
											assign node6241 = (inp[9]) ? node6245 : node6242;
												assign node6242 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node6245 = (inp[4]) ? node6247 : 4'b1111;
													assign node6247 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node6250 = (inp[9]) ? node6254 : node6251;
												assign node6251 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6254 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node6257 = (inp[1]) ? node6265 : node6258;
											assign node6258 = (inp[0]) ? 4'b1100 : node6259;
												assign node6259 = (inp[4]) ? 4'b1100 : node6260;
													assign node6260 = (inp[6]) ? 4'b1100 : 4'b1101;
											assign node6265 = (inp[6]) ? node6269 : node6266;
												assign node6266 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node6269 = (inp[12]) ? 4'b1101 : 4'b1001;
									assign node6272 = (inp[12]) ? node6296 : node6273;
										assign node6273 = (inp[6]) ? node6287 : node6274;
											assign node6274 = (inp[4]) ? 4'b1000 : node6275;
												assign node6275 = (inp[9]) ? node6281 : node6276;
													assign node6276 = (inp[10]) ? node6278 : 4'b1101;
														assign node6278 = (inp[1]) ? 4'b1100 : 4'b1100;
													assign node6281 = (inp[1]) ? node6283 : 4'b1100;
														assign node6283 = (inp[10]) ? 4'b1100 : 4'b1100;
											assign node6287 = (inp[4]) ? node6291 : node6288;
												assign node6288 = (inp[1]) ? 4'b1011 : 4'b1110;
												assign node6291 = (inp[1]) ? node6293 : 4'b1011;
													assign node6293 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node6296 = (inp[6]) ? node6302 : node6297;
											assign node6297 = (inp[0]) ? node6299 : 4'b1111;
												assign node6299 = (inp[4]) ? 4'b1110 : 4'b1111;
											assign node6302 = (inp[0]) ? 4'b1111 : node6303;
												assign node6303 = (inp[11]) ? node6307 : node6304;
													assign node6304 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6307 = (inp[9]) ? 4'b1110 : 4'b1111;
								assign node6311 = (inp[15]) ? node6359 : node6312;
									assign node6312 = (inp[6]) ? node6336 : node6313;
										assign node6313 = (inp[10]) ? node6327 : node6314;
											assign node6314 = (inp[9]) ? node6322 : node6315;
												assign node6315 = (inp[0]) ? node6319 : node6316;
													assign node6316 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node6319 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node6322 = (inp[4]) ? node6324 : 4'b1110;
													assign node6324 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node6327 = (inp[11]) ? node6333 : node6328;
												assign node6328 = (inp[9]) ? node6330 : 4'b1000;
													assign node6330 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node6333 = (inp[4]) ? 4'b1110 : 4'b1010;
										assign node6336 = (inp[1]) ? node6350 : node6337;
											assign node6337 = (inp[4]) ? node6343 : node6338;
												assign node6338 = (inp[12]) ? 4'b1011 : node6339;
													assign node6339 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node6343 = (inp[12]) ? node6345 : 4'b1010;
													assign node6345 = (inp[0]) ? node6347 : 4'b1110;
														assign node6347 = (inp[9]) ? 4'b1110 : 4'b1110;
											assign node6350 = (inp[4]) ? 4'b1111 : node6351;
												assign node6351 = (inp[9]) ? 4'b1110 : node6352;
													assign node6352 = (inp[12]) ? 4'b1111 : node6353;
														assign node6353 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node6359 = (inp[12]) ? node6377 : node6360;
										assign node6360 = (inp[6]) ? node6374 : node6361;
											assign node6361 = (inp[10]) ? node6371 : node6362;
												assign node6362 = (inp[1]) ? node6368 : node6363;
													assign node6363 = (inp[0]) ? node6365 : 4'b1111;
														assign node6365 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node6368 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node6371 = (inp[11]) ? 4'b1010 : 4'b1111;
											assign node6374 = (inp[9]) ? 4'b1000 : 4'b1101;
										assign node6377 = (inp[1]) ? node6385 : node6378;
											assign node6378 = (inp[0]) ? node6382 : node6379;
												assign node6379 = (inp[4]) ? 4'b1100 : 4'b1101;
												assign node6382 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node6385 = (inp[0]) ? node6387 : 4'b1100;
												assign node6387 = (inp[11]) ? 4'b1100 : 4'b1101;
						assign node6390 = (inp[12]) ? node6562 : node6391;
							assign node6391 = (inp[1]) ? node6471 : node6392;
								assign node6392 = (inp[4]) ? node6428 : node6393;
									assign node6393 = (inp[7]) ? node6407 : node6394;
										assign node6394 = (inp[15]) ? node6402 : node6395;
											assign node6395 = (inp[11]) ? node6397 : 4'b1001;
												assign node6397 = (inp[9]) ? 4'b1001 : node6398;
													assign node6398 = (inp[6]) ? 4'b1000 : 4'b1100;
											assign node6402 = (inp[6]) ? node6404 : 4'b1100;
												assign node6404 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node6407 = (inp[0]) ? node6417 : node6408;
											assign node6408 = (inp[10]) ? node6412 : node6409;
												assign node6409 = (inp[6]) ? 4'b1010 : 4'b1110;
												assign node6412 = (inp[9]) ? 4'b1010 : node6413;
													assign node6413 = (inp[15]) ? 4'b1010 : 4'b1011;
											assign node6417 = (inp[10]) ? 4'b1000 : node6418;
												assign node6418 = (inp[2]) ? node6422 : node6419;
													assign node6419 = (inp[6]) ? 4'b1010 : 4'b1011;
													assign node6422 = (inp[6]) ? 4'b1011 : node6423;
														assign node6423 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node6428 = (inp[2]) ? node6456 : node6429;
										assign node6429 = (inp[6]) ? node6451 : node6430;
											assign node6430 = (inp[15]) ? node6440 : node6431;
												assign node6431 = (inp[7]) ? node6437 : node6432;
													assign node6432 = (inp[10]) ? node6434 : 4'b1111;
														assign node6434 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6437 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6440 = (inp[7]) ? node6446 : node6441;
													assign node6441 = (inp[11]) ? 4'b1001 : node6442;
														assign node6442 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node6446 = (inp[11]) ? 4'b1010 : node6447;
														assign node6447 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node6451 = (inp[10]) ? node6453 : 4'b1111;
												assign node6453 = (inp[7]) ? 4'b1111 : 4'b1000;
										assign node6456 = (inp[15]) ? node6462 : node6457;
											assign node6457 = (inp[10]) ? 4'b1001 : node6458;
												assign node6458 = (inp[6]) ? 4'b1111 : 4'b1100;
											assign node6462 = (inp[6]) ? 4'b1110 : node6463;
												assign node6463 = (inp[7]) ? node6467 : node6464;
													assign node6464 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node6467 = (inp[9]) ? 4'b1111 : 4'b1110;
								assign node6471 = (inp[4]) ? node6521 : node6472;
									assign node6472 = (inp[15]) ? node6496 : node6473;
										assign node6473 = (inp[7]) ? node6483 : node6474;
											assign node6474 = (inp[10]) ? node6476 : 4'b1100;
												assign node6476 = (inp[9]) ? 4'b1101 : node6477;
													assign node6477 = (inp[0]) ? 4'b1101 : node6478;
														assign node6478 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node6483 = (inp[0]) ? node6485 : 4'b1110;
												assign node6485 = (inp[6]) ? node6489 : node6486;
													assign node6486 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node6489 = (inp[10]) ? node6493 : node6490;
														assign node6490 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node6493 = (inp[9]) ? 4'b1011 : 4'b1010;
										assign node6496 = (inp[7]) ? node6508 : node6497;
											assign node6497 = (inp[6]) ? node6501 : node6498;
												assign node6498 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node6501 = (inp[10]) ? node6503 : 4'b1111;
													assign node6503 = (inp[9]) ? node6505 : 4'b1110;
														assign node6505 = (inp[11]) ? 4'b1110 : 4'b1110;
											assign node6508 = (inp[6]) ? node6510 : 4'b1111;
												assign node6510 = (inp[0]) ? node6516 : node6511;
													assign node6511 = (inp[10]) ? node6513 : 4'b1101;
														assign node6513 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node6516 = (inp[9]) ? node6518 : 4'b1100;
														assign node6518 = (inp[11]) ? 4'b1100 : 4'b1101;
									assign node6521 = (inp[6]) ? node6545 : node6522;
										assign node6522 = (inp[15]) ? node6536 : node6523;
											assign node6523 = (inp[7]) ? 4'b1101 : node6524;
												assign node6524 = (inp[2]) ? node6530 : node6525;
													assign node6525 = (inp[0]) ? node6527 : 4'b1111;
														assign node6527 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6530 = (inp[0]) ? 4'b1011 : node6531;
														assign node6531 = (inp[9]) ? 4'b1010 : 4'b1010;
											assign node6536 = (inp[7]) ? node6542 : node6537;
												assign node6537 = (inp[9]) ? 4'b1001 : node6538;
													assign node6538 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node6542 = (inp[2]) ? 4'b1010 : 4'b1111;
										assign node6545 = (inp[0]) ? node6553 : node6546;
											assign node6546 = (inp[11]) ? 4'b1010 : node6547;
												assign node6547 = (inp[7]) ? 4'b1000 : node6548;
													assign node6548 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node6553 = (inp[11]) ? node6559 : node6554;
												assign node6554 = (inp[2]) ? 4'b1001 : node6555;
													assign node6555 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node6559 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node6562 = (inp[6]) ? node6626 : node6563;
								assign node6563 = (inp[2]) ? node6599 : node6564;
									assign node6564 = (inp[7]) ? node6580 : node6565;
										assign node6565 = (inp[4]) ? node6571 : node6566;
											assign node6566 = (inp[11]) ? node6568 : 4'b1111;
												assign node6568 = (inp[15]) ? 4'b1111 : 4'b1110;
											assign node6571 = (inp[10]) ? node6573 : 4'b1000;
												assign node6573 = (inp[15]) ? node6575 : 4'b1101;
													assign node6575 = (inp[0]) ? 4'b1110 : node6576;
														assign node6576 = (inp[1]) ? 4'b1110 : 4'b1111;
										assign node6580 = (inp[15]) ? node6592 : node6581;
											assign node6581 = (inp[4]) ? node6589 : node6582;
												assign node6582 = (inp[0]) ? 4'b1001 : node6583;
													assign node6583 = (inp[1]) ? node6585 : 4'b1000;
														assign node6585 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6589 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node6592 = (inp[11]) ? node6594 : 4'b1100;
												assign node6594 = (inp[9]) ? 4'b1101 : node6595;
													assign node6595 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node6599 = (inp[7]) ? node6615 : node6600;
										assign node6600 = (inp[15]) ? node6610 : node6601;
											assign node6601 = (inp[4]) ? node6603 : 4'b1010;
												assign node6603 = (inp[1]) ? 4'b1100 : node6604;
													assign node6604 = (inp[11]) ? node6606 : 4'b1000;
														assign node6606 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node6610 = (inp[11]) ? node6612 : 4'b1011;
												assign node6612 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node6615 = (inp[15]) ? node6619 : node6616;
											assign node6616 = (inp[4]) ? 4'b1011 : 4'b1100;
											assign node6619 = (inp[9]) ? 4'b1001 : node6620;
												assign node6620 = (inp[0]) ? node6622 : 4'b1000;
													assign node6622 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node6626 = (inp[15]) ? node6666 : node6627;
									assign node6627 = (inp[7]) ? node6649 : node6628;
										assign node6628 = (inp[1]) ? node6640 : node6629;
											assign node6629 = (inp[4]) ? node6635 : node6630;
												assign node6630 = (inp[0]) ? node6632 : 4'b1000;
													assign node6632 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6635 = (inp[11]) ? 4'b1001 : node6636;
													assign node6636 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node6640 = (inp[4]) ? node6644 : node6641;
												assign node6641 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node6644 = (inp[11]) ? node6646 : 4'b1101;
													assign node6646 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node6649 = (inp[1]) ? node6659 : node6650;
											assign node6650 = (inp[4]) ? node6656 : node6651;
												assign node6651 = (inp[2]) ? 4'b1111 : node6652;
													assign node6652 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node6656 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node6659 = (inp[2]) ? node6661 : 4'b1011;
												assign node6661 = (inp[9]) ? 4'b1010 : node6662;
													assign node6662 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node6666 = (inp[7]) ? node6682 : node6667;
										assign node6667 = (inp[10]) ? node6673 : node6668;
											assign node6668 = (inp[0]) ? 4'b1010 : node6669;
												assign node6669 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node6673 = (inp[9]) ? node6677 : node6674;
												assign node6674 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node6677 = (inp[11]) ? node6679 : 4'b1011;
													assign node6679 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node6682 = (inp[0]) ? node6696 : node6683;
											assign node6683 = (inp[11]) ? node6689 : node6684;
												assign node6684 = (inp[9]) ? node6686 : 4'b1000;
													assign node6686 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node6689 = (inp[9]) ? node6691 : 4'b1001;
													assign node6691 = (inp[1]) ? node6693 : 4'b1000;
														assign node6693 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node6696 = (inp[1]) ? node6702 : node6697;
												assign node6697 = (inp[11]) ? node6699 : 4'b1001;
													assign node6699 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6702 = (inp[10]) ? 4'b1000 : 4'b1001;
				assign node6705 = (inp[15]) ? node7311 : node6706;
					assign node6706 = (inp[12]) ? node7016 : node6707;
						assign node6707 = (inp[6]) ? node6865 : node6708;
							assign node6708 = (inp[11]) ? node6790 : node6709;
								assign node6709 = (inp[2]) ? node6747 : node6710;
									assign node6710 = (inp[7]) ? node6724 : node6711;
										assign node6711 = (inp[4]) ? node6721 : node6712;
											assign node6712 = (inp[0]) ? node6718 : node6713;
												assign node6713 = (inp[13]) ? 4'b0000 : node6714;
													assign node6714 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node6718 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node6721 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node6724 = (inp[1]) ? node6738 : node6725;
											assign node6725 = (inp[4]) ? node6733 : node6726;
												assign node6726 = (inp[10]) ? node6728 : 4'b0100;
													assign node6728 = (inp[9]) ? 4'b0100 : node6729;
														assign node6729 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node6733 = (inp[5]) ? node6735 : 4'b0100;
													assign node6735 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node6738 = (inp[0]) ? 4'b0101 : node6739;
												assign node6739 = (inp[10]) ? 4'b0100 : node6740;
													assign node6740 = (inp[13]) ? node6742 : 4'b0101;
														assign node6742 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node6747 = (inp[9]) ? node6777 : node6748;
										assign node6748 = (inp[13]) ? node6762 : node6749;
											assign node6749 = (inp[10]) ? node6757 : node6750;
												assign node6750 = (inp[7]) ? node6752 : 4'b0000;
													assign node6752 = (inp[4]) ? 4'b0101 : node6753;
														assign node6753 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node6757 = (inp[1]) ? 4'b0001 : node6758;
													assign node6758 = (inp[7]) ? 4'b0000 : 4'b0101;
											assign node6762 = (inp[10]) ? node6770 : node6763;
												assign node6763 = (inp[7]) ? node6767 : node6764;
													assign node6764 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node6767 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node6770 = (inp[4]) ? node6772 : 4'b0100;
													assign node6772 = (inp[0]) ? 4'b0001 : node6773;
														assign node6773 = (inp[7]) ? 4'b0101 : 4'b0000;
										assign node6777 = (inp[7]) ? node6783 : node6778;
											assign node6778 = (inp[10]) ? node6780 : 4'b0100;
												assign node6780 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node6783 = (inp[0]) ? 4'b0100 : node6784;
												assign node6784 = (inp[1]) ? node6786 : 4'b0000;
													assign node6786 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node6790 = (inp[2]) ? node6828 : node6791;
									assign node6791 = (inp[7]) ? node6807 : node6792;
										assign node6792 = (inp[5]) ? node6798 : node6793;
											assign node6793 = (inp[4]) ? node6795 : 4'b0001;
												assign node6795 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node6798 = (inp[4]) ? 4'b0101 : node6799;
												assign node6799 = (inp[13]) ? node6801 : 4'b0001;
													assign node6801 = (inp[1]) ? node6803 : 4'b0000;
														assign node6803 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node6807 = (inp[4]) ? node6815 : node6808;
											assign node6808 = (inp[0]) ? node6810 : 4'b0101;
												assign node6810 = (inp[13]) ? node6812 : 4'b0100;
													assign node6812 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node6815 = (inp[5]) ? node6821 : node6816;
												assign node6816 = (inp[9]) ? node6818 : 4'b0100;
													assign node6818 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node6821 = (inp[0]) ? node6823 : 4'b0000;
													assign node6823 = (inp[1]) ? node6825 : 4'b0001;
														assign node6825 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node6828 = (inp[7]) ? node6850 : node6829;
										assign node6829 = (inp[13]) ? node6841 : node6830;
											assign node6830 = (inp[5]) ? node6838 : node6831;
												assign node6831 = (inp[9]) ? 4'b0101 : node6832;
													assign node6832 = (inp[1]) ? 4'b0100 : node6833;
														assign node6833 = (inp[10]) ? 4'b0100 : 4'b0100;
												assign node6838 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node6841 = (inp[0]) ? node6847 : node6842;
												assign node6842 = (inp[5]) ? node6844 : 4'b0101;
													assign node6844 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node6847 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node6850 = (inp[13]) ? node6860 : node6851;
											assign node6851 = (inp[0]) ? node6857 : node6852;
												assign node6852 = (inp[4]) ? node6854 : 4'b0001;
													assign node6854 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node6857 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node6860 = (inp[9]) ? 4'b0000 : node6861;
												assign node6861 = (inp[10]) ? 4'b0000 : 4'b0100;
							assign node6865 = (inp[10]) ? node6951 : node6866;
								assign node6866 = (inp[0]) ? node6916 : node6867;
									assign node6867 = (inp[4]) ? node6891 : node6868;
										assign node6868 = (inp[9]) ? node6886 : node6869;
											assign node6869 = (inp[11]) ? node6875 : node6870;
												assign node6870 = (inp[7]) ? node6872 : 4'b0110;
													assign node6872 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node6875 = (inp[13]) ? node6881 : node6876;
													assign node6876 = (inp[2]) ? 4'b0011 : node6877;
														assign node6877 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node6881 = (inp[7]) ? node6883 : 4'b0011;
														assign node6883 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node6886 = (inp[5]) ? 4'b0110 : node6887;
												assign node6887 = (inp[7]) ? 4'b0110 : 4'b0010;
										assign node6891 = (inp[13]) ? node6909 : node6892;
											assign node6892 = (inp[1]) ? node6902 : node6893;
												assign node6893 = (inp[9]) ? node6899 : node6894;
													assign node6894 = (inp[11]) ? 4'b0011 : node6895;
														assign node6895 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node6899 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node6902 = (inp[2]) ? 4'b0111 : node6903;
													assign node6903 = (inp[5]) ? node6905 : 4'b0010;
														assign node6905 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node6909 = (inp[5]) ? node6913 : node6910;
												assign node6910 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node6913 = (inp[7]) ? 4'b0011 : 4'b0110;
									assign node6916 = (inp[1]) ? node6942 : node6917;
										assign node6917 = (inp[13]) ? node6925 : node6918;
											assign node6918 = (inp[11]) ? 4'b0111 : node6919;
												assign node6919 = (inp[9]) ? 4'b0110 : node6920;
													assign node6920 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node6925 = (inp[11]) ? node6933 : node6926;
												assign node6926 = (inp[2]) ? node6928 : 4'b0111;
													assign node6928 = (inp[4]) ? node6930 : 4'b0011;
														assign node6930 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node6933 = (inp[2]) ? 4'b0010 : node6934;
													assign node6934 = (inp[7]) ? node6938 : node6935;
														assign node6935 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node6938 = (inp[4]) ? 4'b0110 : 4'b0011;
										assign node6942 = (inp[13]) ? 4'b0111 : node6943;
											assign node6943 = (inp[11]) ? node6945 : 4'b0010;
												assign node6945 = (inp[2]) ? node6947 : 4'b0011;
													assign node6947 = (inp[7]) ? 4'b0011 : 4'b0111;
								assign node6951 = (inp[5]) ? node6985 : node6952;
									assign node6952 = (inp[7]) ? node6964 : node6953;
										assign node6953 = (inp[4]) ? node6955 : 4'b0010;
											assign node6955 = (inp[1]) ? node6961 : node6956;
												assign node6956 = (inp[13]) ? node6958 : 4'b0011;
													assign node6958 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node6961 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node6964 = (inp[2]) ? node6974 : node6965;
											assign node6965 = (inp[9]) ? node6967 : 4'b0110;
												assign node6967 = (inp[1]) ? node6969 : 4'b0111;
													assign node6969 = (inp[11]) ? node6971 : 4'b0110;
														assign node6971 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node6974 = (inp[1]) ? node6980 : node6975;
												assign node6975 = (inp[11]) ? node6977 : 4'b0110;
													assign node6977 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node6980 = (inp[11]) ? node6982 : 4'b0111;
													assign node6982 = (inp[13]) ? 4'b0111 : 4'b0110;
									assign node6985 = (inp[7]) ? node6997 : node6986;
										assign node6986 = (inp[2]) ? node6992 : node6987;
											assign node6987 = (inp[1]) ? node6989 : 4'b0111;
												assign node6989 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node6992 = (inp[1]) ? node6994 : 4'b0110;
												assign node6994 = (inp[4]) ? 4'b0110 : 4'b0111;
										assign node6997 = (inp[9]) ? node7003 : node6998;
											assign node6998 = (inp[0]) ? 4'b0010 : node6999;
												assign node6999 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node7003 = (inp[13]) ? node7007 : node7004;
												assign node7004 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node7007 = (inp[0]) ? node7009 : 4'b0011;
													assign node7009 = (inp[4]) ? node7013 : node7010;
														assign node7010 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node7013 = (inp[1]) ? 4'b0011 : 4'b0010;
						assign node7016 = (inp[4]) ? node7164 : node7017;
							assign node7017 = (inp[7]) ? node7097 : node7018;
								assign node7018 = (inp[2]) ? node7062 : node7019;
									assign node7019 = (inp[6]) ? node7041 : node7020;
										assign node7020 = (inp[10]) ? node7024 : node7021;
											assign node7021 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node7024 = (inp[5]) ? node7034 : node7025;
												assign node7025 = (inp[9]) ? node7027 : 4'b0011;
													assign node7027 = (inp[0]) ? node7031 : node7028;
														assign node7028 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node7031 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node7034 = (inp[1]) ? node7036 : 4'b0010;
													assign node7036 = (inp[11]) ? 4'b0011 : node7037;
														assign node7037 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node7041 = (inp[5]) ? node7051 : node7042;
											assign node7042 = (inp[10]) ? node7044 : 4'b0011;
												assign node7044 = (inp[13]) ? node7048 : node7045;
													assign node7045 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node7048 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node7051 = (inp[10]) ? 4'b0111 : node7052;
												assign node7052 = (inp[0]) ? node7058 : node7053;
													assign node7053 = (inp[1]) ? node7055 : 4'b0111;
														assign node7055 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node7058 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node7062 = (inp[6]) ? node7084 : node7063;
										assign node7063 = (inp[9]) ? node7071 : node7064;
											assign node7064 = (inp[5]) ? node7066 : 4'b0111;
												assign node7066 = (inp[10]) ? node7068 : 4'b0111;
													assign node7068 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node7071 = (inp[1]) ? node7077 : node7072;
												assign node7072 = (inp[13]) ? node7074 : 4'b0110;
													assign node7074 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node7077 = (inp[11]) ? 4'b0111 : node7078;
													assign node7078 = (inp[5]) ? node7080 : 4'b0110;
														assign node7080 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node7084 = (inp[5]) ? node7088 : node7085;
											assign node7085 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node7088 = (inp[1]) ? 4'b0110 : node7089;
												assign node7089 = (inp[9]) ? 4'b0111 : node7090;
													assign node7090 = (inp[13]) ? 4'b0110 : node7091;
														assign node7091 = (inp[11]) ? 4'b0111 : 4'b0110;
								assign node7097 = (inp[2]) ? node7137 : node7098;
									assign node7098 = (inp[0]) ? node7126 : node7099;
										assign node7099 = (inp[5]) ? node7113 : node7100;
											assign node7100 = (inp[1]) ? node7106 : node7101;
												assign node7101 = (inp[9]) ? 4'b0110 : node7102;
													assign node7102 = (inp[6]) ? 4'b0111 : 4'b0110;
												assign node7106 = (inp[10]) ? node7108 : 4'b0111;
													assign node7108 = (inp[11]) ? 4'b0111 : node7109;
														assign node7109 = (inp[6]) ? 4'b0110 : 4'b0111;
											assign node7113 = (inp[6]) ? node7123 : node7114;
												assign node7114 = (inp[9]) ? node7116 : 4'b0111;
													assign node7116 = (inp[10]) ? node7120 : node7117;
														assign node7117 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node7120 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node7123 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node7126 = (inp[10]) ? node7128 : 4'b0110;
											assign node7128 = (inp[6]) ? node7134 : node7129;
												assign node7129 = (inp[13]) ? node7131 : 4'b0110;
													assign node7131 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node7134 = (inp[5]) ? 4'b0011 : 4'b0111;
									assign node7137 = (inp[5]) ? node7153 : node7138;
										assign node7138 = (inp[6]) ? node7142 : node7139;
											assign node7139 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node7142 = (inp[0]) ? node7148 : node7143;
												assign node7143 = (inp[10]) ? 4'b0110 : node7144;
													assign node7144 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node7148 = (inp[11]) ? 4'b0111 : node7149;
													assign node7149 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node7153 = (inp[13]) ? 4'b0010 : node7154;
											assign node7154 = (inp[0]) ? node7156 : 4'b0011;
												assign node7156 = (inp[11]) ? node7158 : 4'b0010;
													assign node7158 = (inp[9]) ? 4'b0011 : node7159;
														assign node7159 = (inp[1]) ? 4'b0011 : 4'b0010;
							assign node7164 = (inp[6]) ? node7248 : node7165;
								assign node7165 = (inp[2]) ? node7211 : node7166;
									assign node7166 = (inp[5]) ? node7194 : node7167;
										assign node7167 = (inp[7]) ? node7179 : node7168;
											assign node7168 = (inp[1]) ? node7174 : node7169;
												assign node7169 = (inp[10]) ? 4'b0110 : node7170;
													assign node7170 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node7174 = (inp[10]) ? node7176 : 4'b0111;
													assign node7176 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node7179 = (inp[1]) ? node7185 : node7180;
												assign node7180 = (inp[0]) ? 4'b0011 : node7181;
													assign node7181 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node7185 = (inp[10]) ? 4'b0011 : node7186;
													assign node7186 = (inp[11]) ? node7190 : node7187;
														assign node7187 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node7190 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node7194 = (inp[7]) ? node7206 : node7195;
											assign node7195 = (inp[1]) ? node7199 : node7196;
												assign node7196 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node7199 = (inp[0]) ? 4'b0010 : node7200;
													assign node7200 = (inp[10]) ? 4'b0010 : node7201;
														assign node7201 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node7206 = (inp[13]) ? 4'b0110 : node7207;
												assign node7207 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node7211 = (inp[10]) ? node7239 : node7212;
										assign node7212 = (inp[13]) ? node7226 : node7213;
											assign node7213 = (inp[9]) ? node7219 : node7214;
												assign node7214 = (inp[5]) ? node7216 : 4'b0110;
													assign node7216 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node7219 = (inp[7]) ? 4'b0010 : node7220;
													assign node7220 = (inp[5]) ? 4'b0110 : node7221;
														assign node7221 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node7226 = (inp[9]) ? 4'b0110 : node7227;
												assign node7227 = (inp[5]) ? node7235 : node7228;
													assign node7228 = (inp[7]) ? node7232 : node7229;
														assign node7229 = (inp[0]) ? 4'b0010 : 4'b0010;
														assign node7232 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node7235 = (inp[7]) ? 4'b0011 : 4'b0111;
										assign node7239 = (inp[7]) ? node7243 : node7240;
											assign node7240 = (inp[5]) ? 4'b0111 : 4'b0011;
											assign node7243 = (inp[5]) ? node7245 : 4'b0110;
												assign node7245 = (inp[13]) ? 4'b0010 : 4'b0011;
								assign node7248 = (inp[13]) ? node7288 : node7249;
									assign node7249 = (inp[11]) ? node7267 : node7250;
										assign node7250 = (inp[0]) ? node7260 : node7251;
											assign node7251 = (inp[7]) ? node7257 : node7252;
												assign node7252 = (inp[2]) ? node7254 : 4'b0010;
													assign node7254 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node7257 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node7260 = (inp[5]) ? node7264 : node7261;
												assign node7261 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node7264 = (inp[7]) ? 4'b0010 : 4'b0110;
										assign node7267 = (inp[9]) ? node7281 : node7268;
											assign node7268 = (inp[2]) ? node7272 : node7269;
												assign node7269 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node7272 = (inp[1]) ? node7278 : node7273;
													assign node7273 = (inp[10]) ? node7275 : 4'b0111;
														assign node7275 = (inp[7]) ? 4'b0011 : 4'b0011;
													assign node7278 = (inp[5]) ? 4'b0111 : 4'b0010;
											assign node7281 = (inp[1]) ? 4'b0111 : node7282;
												assign node7282 = (inp[0]) ? node7284 : 4'b0110;
													assign node7284 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node7288 = (inp[11]) ? node7296 : node7289;
										assign node7289 = (inp[7]) ? node7293 : node7290;
											assign node7290 = (inp[5]) ? 4'b0111 : 4'b0011;
											assign node7293 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node7296 = (inp[7]) ? node7304 : node7297;
											assign node7297 = (inp[5]) ? 4'b0110 : node7298;
												assign node7298 = (inp[2]) ? node7300 : 4'b0010;
													assign node7300 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node7304 = (inp[2]) ? node7308 : node7305;
												assign node7305 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node7308 = (inp[5]) ? 4'b0010 : 4'b0110;
					assign node7311 = (inp[6]) ? node7497 : node7312;
						assign node7312 = (inp[12]) ? node7406 : node7313;
							assign node7313 = (inp[2]) ? node7365 : node7314;
								assign node7314 = (inp[4]) ? node7344 : node7315;
									assign node7315 = (inp[13]) ? node7333 : node7316;
										assign node7316 = (inp[10]) ? node7326 : node7317;
											assign node7317 = (inp[11]) ? node7319 : 4'b0010;
												assign node7319 = (inp[7]) ? node7321 : 4'b0010;
													assign node7321 = (inp[0]) ? 4'b0011 : node7322;
														assign node7322 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node7326 = (inp[1]) ? node7328 : 4'b0011;
												assign node7328 = (inp[5]) ? node7330 : 4'b0010;
													assign node7330 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node7333 = (inp[0]) ? node7335 : 4'b0011;
											assign node7335 = (inp[10]) ? node7339 : node7336;
												assign node7336 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node7339 = (inp[9]) ? node7341 : 4'b0011;
													assign node7341 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node7344 = (inp[1]) ? node7352 : node7345;
										assign node7345 = (inp[10]) ? 4'b0111 : node7346;
											assign node7346 = (inp[11]) ? node7348 : 4'b0110;
												assign node7348 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node7352 = (inp[10]) ? node7362 : node7353;
											assign node7353 = (inp[11]) ? node7355 : 4'b0111;
												assign node7355 = (inp[9]) ? node7357 : 4'b0111;
													assign node7357 = (inp[0]) ? node7359 : 4'b0110;
														assign node7359 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node7362 = (inp[11]) ? 4'b0111 : 4'b0110;
								assign node7365 = (inp[4]) ? node7387 : node7366;
									assign node7366 = (inp[5]) ? node7376 : node7367;
										assign node7367 = (inp[9]) ? 4'b0111 : node7368;
											assign node7368 = (inp[13]) ? 4'b0110 : node7369;
												assign node7369 = (inp[11]) ? node7371 : 4'b0111;
													assign node7371 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node7376 = (inp[10]) ? 4'b0110 : node7377;
											assign node7377 = (inp[11]) ? node7383 : node7378;
												assign node7378 = (inp[0]) ? 4'b0110 : node7379;
													assign node7379 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node7383 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node7387 = (inp[7]) ? node7393 : node7388;
										assign node7388 = (inp[10]) ? node7390 : 4'b0010;
											assign node7390 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node7393 = (inp[0]) ? node7399 : node7394;
											assign node7394 = (inp[5]) ? 4'b0010 : node7395;
												assign node7395 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node7399 = (inp[5]) ? 4'b0011 : node7400;
												assign node7400 = (inp[9]) ? 4'b0010 : node7401;
													assign node7401 = (inp[13]) ? 4'b0011 : 4'b0010;
							assign node7406 = (inp[4]) ? node7434 : node7407;
								assign node7407 = (inp[10]) ? node7417 : node7408;
									assign node7408 = (inp[2]) ? node7412 : node7409;
										assign node7409 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node7412 = (inp[5]) ? 4'b0001 : node7413;
											assign node7413 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node7417 = (inp[7]) ? node7425 : node7418;
										assign node7418 = (inp[2]) ? node7422 : node7419;
											assign node7419 = (inp[5]) ? 4'b0101 : 4'b0001;
											assign node7422 = (inp[5]) ? 4'b0000 : 4'b0101;
										assign node7425 = (inp[5]) ? node7429 : node7426;
											assign node7426 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node7429 = (inp[2]) ? node7431 : 4'b0101;
												assign node7431 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node7434 = (inp[7]) ? node7470 : node7435;
									assign node7435 = (inp[13]) ? node7465 : node7436;
										assign node7436 = (inp[0]) ? node7452 : node7437;
											assign node7437 = (inp[1]) ? node7445 : node7438;
												assign node7438 = (inp[2]) ? node7442 : node7439;
													assign node7439 = (inp[5]) ? 4'b0101 : 4'b0001;
													assign node7442 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node7445 = (inp[11]) ? node7447 : 4'b0100;
													assign node7447 = (inp[2]) ? 4'b0000 : node7448;
														assign node7448 = (inp[5]) ? 4'b0100 : 4'b0000;
											assign node7452 = (inp[10]) ? 4'b0001 : node7453;
												assign node7453 = (inp[5]) ? node7459 : node7454;
													assign node7454 = (inp[2]) ? node7456 : 4'b0000;
														assign node7456 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node7459 = (inp[2]) ? node7461 : 4'b0101;
														assign node7461 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node7465 = (inp[0]) ? node7467 : 4'b0000;
											assign node7467 = (inp[2]) ? 4'b0000 : 4'b0100;
									assign node7470 = (inp[0]) ? node7482 : node7471;
										assign node7471 = (inp[13]) ? 4'b0001 : node7472;
											assign node7472 = (inp[11]) ? node7474 : 4'b0101;
												assign node7474 = (inp[9]) ? node7476 : 4'b0000;
													assign node7476 = (inp[1]) ? node7478 : 4'b0001;
														assign node7478 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node7482 = (inp[2]) ? node7490 : node7483;
											assign node7483 = (inp[5]) ? node7487 : node7484;
												assign node7484 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node7487 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node7490 = (inp[5]) ? node7494 : node7491;
												assign node7491 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node7494 = (inp[9]) ? 4'b0001 : 4'b0000;
						assign node7497 = (inp[5]) ? node7557 : node7498;
							assign node7498 = (inp[12]) ? node7550 : node7499;
								assign node7499 = (inp[4]) ? node7521 : node7500;
									assign node7500 = (inp[1]) ? node7508 : node7501;
										assign node7501 = (inp[7]) ? node7505 : node7502;
											assign node7502 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node7505 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node7508 = (inp[7]) ? node7512 : node7509;
											assign node7509 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node7512 = (inp[10]) ? node7514 : 4'b0001;
												assign node7514 = (inp[11]) ? node7518 : node7515;
													assign node7515 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node7518 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node7521 = (inp[2]) ? node7539 : node7522;
										assign node7522 = (inp[9]) ? node7528 : node7523;
											assign node7523 = (inp[7]) ? 4'b0100 : node7524;
												assign node7524 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node7528 = (inp[10]) ? node7534 : node7529;
												assign node7529 = (inp[11]) ? 4'b0101 : node7530;
													assign node7530 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node7534 = (inp[1]) ? node7536 : 4'b0100;
													assign node7536 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node7539 = (inp[7]) ? 4'b0101 : node7540;
											assign node7540 = (inp[9]) ? node7542 : 4'b0101;
												assign node7542 = (inp[0]) ? 4'b0100 : node7543;
													assign node7543 = (inp[13]) ? 4'b0101 : node7544;
														assign node7544 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node7550 = (inp[11]) ? node7554 : node7551;
									assign node7551 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node7554 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node7557 = (inp[12]) ? node7607 : node7558;
								assign node7558 = (inp[4]) ? node7586 : node7559;
									assign node7559 = (inp[0]) ? node7573 : node7560;
										assign node7560 = (inp[1]) ? node7566 : node7561;
											assign node7561 = (inp[11]) ? 4'b0101 : node7562;
												assign node7562 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node7566 = (inp[11]) ? 4'b0100 : node7567;
												assign node7567 = (inp[2]) ? 4'b0101 : node7568;
													assign node7568 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node7573 = (inp[2]) ? node7579 : node7574;
											assign node7574 = (inp[7]) ? node7576 : 4'b0100;
												assign node7576 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node7579 = (inp[11]) ? node7583 : node7580;
												assign node7580 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node7583 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node7586 = (inp[2]) ? node7592 : node7587;
										assign node7587 = (inp[7]) ? node7589 : 4'b0001;
											assign node7589 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node7592 = (inp[9]) ? node7598 : node7593;
											assign node7593 = (inp[7]) ? node7595 : 4'b0001;
												assign node7595 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node7598 = (inp[10]) ? 4'b0000 : node7599;
												assign node7599 = (inp[11]) ? node7603 : node7600;
													assign node7600 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node7603 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node7607 = (inp[11]) ? node7613 : node7608;
									assign node7608 = (inp[2]) ? 4'b0001 : node7609;
										assign node7609 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node7613 = (inp[2]) ? 4'b0000 : node7614;
										assign node7614 = (inp[4]) ? 4'b0000 : 4'b0001;
			assign node7618 = (inp[6]) ? node8968 : node7619;
				assign node7619 = (inp[12]) ? node8367 : node7620;
					assign node7620 = (inp[8]) ? node7994 : node7621;
						assign node7621 = (inp[7]) ? node7811 : node7622;
							assign node7622 = (inp[4]) ? node7702 : node7623;
								assign node7623 = (inp[15]) ? node7667 : node7624;
									assign node7624 = (inp[1]) ? node7656 : node7625;
										assign node7625 = (inp[0]) ? node7639 : node7626;
											assign node7626 = (inp[9]) ? node7634 : node7627;
												assign node7627 = (inp[13]) ? node7631 : node7628;
													assign node7628 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node7631 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node7634 = (inp[10]) ? node7636 : 4'b0111;
													assign node7636 = (inp[13]) ? 4'b0111 : 4'b0010;
											assign node7639 = (inp[9]) ? node7647 : node7640;
												assign node7640 = (inp[13]) ? node7644 : node7641;
													assign node7641 = (inp[11]) ? 4'b0011 : 4'b0110;
													assign node7644 = (inp[11]) ? 4'b0110 : 4'b0011;
												assign node7647 = (inp[5]) ? node7649 : 4'b0011;
													assign node7649 = (inp[13]) ? node7653 : node7650;
														assign node7650 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node7653 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node7656 = (inp[2]) ? node7664 : node7657;
											assign node7657 = (inp[13]) ? 4'b0010 : node7658;
												assign node7658 = (inp[11]) ? 4'b0110 : node7659;
													assign node7659 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node7664 = (inp[11]) ? 4'b0011 : 4'b0010;
									assign node7667 = (inp[9]) ? node7687 : node7668;
										assign node7668 = (inp[11]) ? node7678 : node7669;
											assign node7669 = (inp[10]) ? 4'b0100 : node7670;
												assign node7670 = (inp[5]) ? 4'b0101 : node7671;
													assign node7671 = (inp[1]) ? node7673 : 4'b0100;
														assign node7673 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node7678 = (inp[10]) ? node7680 : 4'b0000;
												assign node7680 = (inp[2]) ? 4'b0100 : node7681;
													assign node7681 = (inp[13]) ? node7683 : 4'b0101;
														assign node7683 = (inp[0]) ? 4'b0101 : 4'b0001;
										assign node7687 = (inp[2]) ? node7695 : node7688;
											assign node7688 = (inp[10]) ? node7690 : 4'b0001;
												assign node7690 = (inp[0]) ? node7692 : 4'b0000;
													assign node7692 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node7695 = (inp[10]) ? node7697 : 4'b0000;
												assign node7697 = (inp[11]) ? node7699 : 4'b0101;
													assign node7699 = (inp[5]) ? 4'b0100 : 4'b0000;
								assign node7702 = (inp[11]) ? node7754 : node7703;
									assign node7703 = (inp[15]) ? node7729 : node7704;
										assign node7704 = (inp[9]) ? node7722 : node7705;
											assign node7705 = (inp[0]) ? node7713 : node7706;
												assign node7706 = (inp[5]) ? node7708 : 4'b0100;
													assign node7708 = (inp[2]) ? node7710 : 4'b0101;
														assign node7710 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node7713 = (inp[5]) ? 4'b0100 : node7714;
													assign node7714 = (inp[10]) ? node7718 : node7715;
														assign node7715 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node7718 = (inp[13]) ? 4'b0001 : 4'b0100;
											assign node7722 = (inp[13]) ? 4'b0000 : node7723;
												assign node7723 = (inp[1]) ? 4'b0001 : node7724;
													assign node7724 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node7729 = (inp[9]) ? node7743 : node7730;
											assign node7730 = (inp[0]) ? node7738 : node7731;
												assign node7731 = (inp[13]) ? node7733 : 4'b0001;
													assign node7733 = (inp[2]) ? node7735 : 4'b0000;
														assign node7735 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node7738 = (inp[2]) ? 4'b0000 : node7739;
													assign node7739 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node7743 = (inp[1]) ? 4'b0100 : node7744;
												assign node7744 = (inp[5]) ? node7746 : 4'b0100;
													assign node7746 = (inp[0]) ? node7750 : node7747;
														assign node7747 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node7750 = (inp[2]) ? 4'b0100 : 4'b0000;
									assign node7754 = (inp[9]) ? node7780 : node7755;
										assign node7755 = (inp[1]) ? node7763 : node7756;
											assign node7756 = (inp[13]) ? 4'b0101 : node7757;
												assign node7757 = (inp[5]) ? 4'b0001 : node7758;
													assign node7758 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node7763 = (inp[0]) ? node7773 : node7764;
												assign node7764 = (inp[5]) ? node7768 : node7765;
													assign node7765 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node7768 = (inp[2]) ? node7770 : 4'b0000;
														assign node7770 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node7773 = (inp[10]) ? node7777 : node7774;
													assign node7774 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node7777 = (inp[15]) ? 4'b0101 : 4'b0001;
										assign node7780 = (inp[13]) ? node7798 : node7781;
											assign node7781 = (inp[2]) ? node7791 : node7782;
												assign node7782 = (inp[0]) ? node7784 : 4'b0000;
													assign node7784 = (inp[1]) ? node7788 : node7785;
														assign node7785 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node7788 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node7791 = (inp[15]) ? 4'b0001 : node7792;
													assign node7792 = (inp[1]) ? 4'b0101 : node7793;
														assign node7793 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node7798 = (inp[15]) ? node7804 : node7799;
												assign node7799 = (inp[1]) ? 4'b0000 : node7800;
													assign node7800 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node7804 = (inp[5]) ? 4'b0001 : node7805;
													assign node7805 = (inp[1]) ? 4'b0001 : node7806;
														assign node7806 = (inp[0]) ? 4'b0000 : 4'b0001;
							assign node7811 = (inp[4]) ? node7917 : node7812;
								assign node7812 = (inp[15]) ? node7868 : node7813;
									assign node7813 = (inp[11]) ? node7845 : node7814;
										assign node7814 = (inp[1]) ? node7834 : node7815;
											assign node7815 = (inp[0]) ? node7825 : node7816;
												assign node7816 = (inp[5]) ? node7822 : node7817;
													assign node7817 = (inp[10]) ? 4'b0100 : node7818;
														assign node7818 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node7822 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node7825 = (inp[5]) ? node7829 : node7826;
													assign node7826 = (inp[2]) ? 4'b0100 : 4'b0001;
													assign node7829 = (inp[10]) ? 4'b0001 : node7830;
														assign node7830 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node7834 = (inp[5]) ? node7836 : 4'b0000;
												assign node7836 = (inp[10]) ? 4'b0100 : node7837;
													assign node7837 = (inp[9]) ? node7841 : node7838;
														assign node7838 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node7841 = (inp[2]) ? 4'b0000 : 4'b0101;
										assign node7845 = (inp[0]) ? node7861 : node7846;
											assign node7846 = (inp[1]) ? node7854 : node7847;
												assign node7847 = (inp[2]) ? node7849 : 4'b0100;
													assign node7849 = (inp[5]) ? node7851 : 4'b0100;
														assign node7851 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node7854 = (inp[5]) ? 4'b0000 : node7855;
													assign node7855 = (inp[10]) ? 4'b0101 : node7856;
														assign node7856 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node7861 = (inp[10]) ? node7865 : node7862;
												assign node7862 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node7865 = (inp[1]) ? 4'b0101 : 4'b0001;
									assign node7868 = (inp[10]) ? node7896 : node7869;
										assign node7869 = (inp[2]) ? node7883 : node7870;
											assign node7870 = (inp[5]) ? node7876 : node7871;
												assign node7871 = (inp[1]) ? node7873 : 4'b0110;
													assign node7873 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node7876 = (inp[13]) ? 4'b0011 : node7877;
													assign node7877 = (inp[1]) ? node7879 : 4'b0111;
														assign node7879 = (inp[9]) ? 4'b0110 : 4'b0110;
											assign node7883 = (inp[13]) ? node7887 : node7884;
												assign node7884 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node7887 = (inp[1]) ? 4'b0111 : node7888;
													assign node7888 = (inp[5]) ? node7892 : node7889;
														assign node7889 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node7892 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node7896 = (inp[1]) ? node7910 : node7897;
											assign node7897 = (inp[5]) ? 4'b0011 : node7898;
												assign node7898 = (inp[13]) ? node7904 : node7899;
													assign node7899 = (inp[2]) ? 4'b0111 : node7900;
														assign node7900 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node7904 = (inp[2]) ? 4'b0011 : node7905;
														assign node7905 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node7910 = (inp[2]) ? node7914 : node7911;
												assign node7911 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node7914 = (inp[5]) ? 4'b0011 : 4'b0010;
								assign node7917 = (inp[9]) ? node7947 : node7918;
									assign node7918 = (inp[13]) ? node7928 : node7919;
										assign node7919 = (inp[2]) ? node7925 : node7920;
											assign node7920 = (inp[10]) ? 4'b0011 : node7921;
												assign node7921 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node7925 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node7928 = (inp[2]) ? node7938 : node7929;
											assign node7929 = (inp[1]) ? node7933 : node7930;
												assign node7930 = (inp[0]) ? 4'b0110 : 4'b0010;
												assign node7933 = (inp[10]) ? node7935 : 4'b0110;
													assign node7935 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node7938 = (inp[10]) ? node7942 : node7939;
												assign node7939 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node7942 = (inp[1]) ? 4'b0011 : node7943;
													assign node7943 = (inp[15]) ? 4'b0010 : 4'b0011;
									assign node7947 = (inp[0]) ? node7969 : node7948;
										assign node7948 = (inp[5]) ? node7962 : node7949;
											assign node7949 = (inp[1]) ? node7955 : node7950;
												assign node7950 = (inp[11]) ? 4'b0011 : node7951;
													assign node7951 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node7955 = (inp[13]) ? 4'b0111 : node7956;
													assign node7956 = (inp[11]) ? node7958 : 4'b0010;
														assign node7958 = (inp[15]) ? 4'b0111 : 4'b0110;
											assign node7962 = (inp[10]) ? node7966 : node7963;
												assign node7963 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node7966 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node7969 = (inp[2]) ? node7983 : node7970;
											assign node7970 = (inp[13]) ? node7976 : node7971;
												assign node7971 = (inp[5]) ? 4'b0010 : node7972;
													assign node7972 = (inp[15]) ? 4'b0011 : 4'b0111;
												assign node7976 = (inp[5]) ? node7978 : 4'b0110;
													assign node7978 = (inp[1]) ? 4'b0111 : node7979;
														assign node7979 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node7983 = (inp[13]) ? node7989 : node7984;
												assign node7984 = (inp[5]) ? node7986 : 4'b0010;
													assign node7986 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node7989 = (inp[1]) ? node7991 : 4'b0010;
													assign node7991 = (inp[10]) ? 4'b0010 : 4'b0011;
						assign node7994 = (inp[0]) ? node8190 : node7995;
							assign node7995 = (inp[10]) ? node8083 : node7996;
								assign node7996 = (inp[1]) ? node8040 : node7997;
									assign node7997 = (inp[15]) ? node8015 : node7998;
										assign node7998 = (inp[9]) ? node8006 : node7999;
											assign node7999 = (inp[5]) ? 4'b0110 : node8000;
												assign node8000 = (inp[4]) ? node8002 : 4'b0011;
													assign node8002 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node8006 = (inp[7]) ? node8008 : 4'b0011;
												assign node8008 = (inp[5]) ? node8010 : 4'b0110;
													assign node8010 = (inp[2]) ? node8012 : 4'b0011;
														assign node8012 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node8015 = (inp[5]) ? node8023 : node8016;
											assign node8016 = (inp[2]) ? node8020 : node8017;
												assign node8017 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node8020 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node8023 = (inp[7]) ? node8031 : node8024;
												assign node8024 = (inp[11]) ? 4'b0010 : node8025;
													assign node8025 = (inp[2]) ? node8027 : 4'b0111;
														assign node8027 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node8031 = (inp[2]) ? node8037 : node8032;
													assign node8032 = (inp[4]) ? 4'b0110 : node8033;
														assign node8033 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node8037 = (inp[4]) ? 4'b0010 : 4'b0110;
									assign node8040 = (inp[13]) ? node8066 : node8041;
										assign node8041 = (inp[9]) ? node8051 : node8042;
											assign node8042 = (inp[4]) ? 4'b0011 : node8043;
												assign node8043 = (inp[2]) ? node8045 : 4'b0010;
													assign node8045 = (inp[5]) ? 4'b0110 : node8046;
														assign node8046 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node8051 = (inp[7]) ? node8063 : node8052;
												assign node8052 = (inp[15]) ? node8058 : node8053;
													assign node8053 = (inp[11]) ? 4'b0011 : node8054;
														assign node8054 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node8058 = (inp[2]) ? node8060 : 4'b0111;
														assign node8060 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node8063 = (inp[4]) ? 4'b0110 : 4'b0111;
										assign node8066 = (inp[11]) ? node8072 : node8067;
											assign node8067 = (inp[5]) ? 4'b0011 : node8068;
												assign node8068 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node8072 = (inp[15]) ? node8074 : 4'b0011;
												assign node8074 = (inp[5]) ? node8076 : 4'b0010;
													assign node8076 = (inp[4]) ? node8080 : node8077;
														assign node8077 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node8080 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node8083 = (inp[7]) ? node8145 : node8084;
									assign node8084 = (inp[5]) ? node8114 : node8085;
										assign node8085 = (inp[9]) ? node8099 : node8086;
											assign node8086 = (inp[11]) ? node8092 : node8087;
												assign node8087 = (inp[2]) ? 4'b0110 : node8088;
													assign node8088 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node8092 = (inp[1]) ? node8096 : node8093;
													assign node8093 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node8096 = (inp[2]) ? 4'b0011 : 4'b0111;
											assign node8099 = (inp[4]) ? node8103 : node8100;
												assign node8100 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node8103 = (inp[1]) ? node8111 : node8104;
													assign node8104 = (inp[11]) ? node8108 : node8105;
														assign node8105 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node8108 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node8111 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node8114 = (inp[1]) ? node8134 : node8115;
											assign node8115 = (inp[2]) ? node8125 : node8116;
												assign node8116 = (inp[13]) ? node8122 : node8117;
													assign node8117 = (inp[15]) ? 4'b0011 : node8118;
														assign node8118 = (inp[4]) ? 4'b0011 : 4'b0110;
													assign node8122 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node8125 = (inp[15]) ? node8131 : node8126;
													assign node8126 = (inp[4]) ? node8128 : 4'b0011;
														assign node8128 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node8131 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node8134 = (inp[2]) ? node8140 : node8135;
												assign node8135 = (inp[4]) ? node8137 : 4'b0110;
													assign node8137 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node8140 = (inp[9]) ? node8142 : 4'b0111;
													assign node8142 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node8145 = (inp[1]) ? node8171 : node8146;
										assign node8146 = (inp[9]) ? node8158 : node8147;
											assign node8147 = (inp[13]) ? node8151 : node8148;
												assign node8148 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node8151 = (inp[2]) ? node8153 : 4'b0010;
													assign node8153 = (inp[15]) ? node8155 : 4'b0010;
														assign node8155 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node8158 = (inp[4]) ? node8164 : node8159;
												assign node8159 = (inp[11]) ? node8161 : 4'b0111;
													assign node8161 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node8164 = (inp[2]) ? 4'b0011 : node8165;
													assign node8165 = (inp[15]) ? 4'b0111 : node8166;
														assign node8166 = (inp[13]) ? 4'b0111 : 4'b0110;
										assign node8171 = (inp[15]) ? node8185 : node8172;
											assign node8172 = (inp[13]) ? node8178 : node8173;
												assign node8173 = (inp[2]) ? node8175 : 4'b0111;
													assign node8175 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node8178 = (inp[2]) ? node8180 : 4'b0110;
													assign node8180 = (inp[5]) ? node8182 : 4'b0011;
														assign node8182 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node8185 = (inp[11]) ? 4'b0110 : node8186;
												assign node8186 = (inp[4]) ? 4'b0110 : 4'b0010;
							assign node8190 = (inp[1]) ? node8294 : node8191;
								assign node8191 = (inp[10]) ? node8231 : node8192;
									assign node8192 = (inp[5]) ? node8218 : node8193;
										assign node8193 = (inp[7]) ? node8209 : node8194;
											assign node8194 = (inp[2]) ? node8202 : node8195;
												assign node8195 = (inp[9]) ? node8197 : 4'b0010;
													assign node8197 = (inp[13]) ? node8199 : 4'b0011;
														assign node8199 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node8202 = (inp[4]) ? 4'b0011 : node8203;
													assign node8203 = (inp[15]) ? 4'b0110 : node8204;
														assign node8204 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node8209 = (inp[15]) ? node8215 : node8210;
												assign node8210 = (inp[13]) ? 4'b0111 : node8211;
													assign node8211 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node8215 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node8218 = (inp[4]) ? node8224 : node8219;
											assign node8219 = (inp[9]) ? node8221 : 4'b0010;
												assign node8221 = (inp[15]) ? 4'b0110 : 4'b0010;
											assign node8224 = (inp[7]) ? 4'b0010 : node8225;
												assign node8225 = (inp[13]) ? node8227 : 4'b0110;
													assign node8227 = (inp[2]) ? 4'b0011 : 4'b0111;
									assign node8231 = (inp[15]) ? node8273 : node8232;
										assign node8232 = (inp[5]) ? node8254 : node8233;
											assign node8233 = (inp[13]) ? node8243 : node8234;
												assign node8234 = (inp[11]) ? node8236 : 4'b0111;
													assign node8236 = (inp[2]) ? node8240 : node8237;
														assign node8237 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node8240 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node8243 = (inp[11]) ? node8249 : node8244;
													assign node8244 = (inp[2]) ? node8246 : 4'b0010;
														assign node8246 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node8249 = (inp[9]) ? 4'b0011 : node8250;
														assign node8250 = (inp[7]) ? 4'b0010 : 4'b0111;
											assign node8254 = (inp[9]) ? node8262 : node8255;
												assign node8255 = (inp[4]) ? node8259 : node8256;
													assign node8256 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node8259 = (inp[11]) ? 4'b0010 : 4'b0110;
												assign node8262 = (inp[2]) ? node8270 : node8263;
													assign node8263 = (inp[7]) ? node8267 : node8264;
														assign node8264 = (inp[4]) ? 4'b0011 : 4'b0110;
														assign node8267 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node8270 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node8273 = (inp[7]) ? node8281 : node8274;
											assign node8274 = (inp[9]) ? 4'b0010 : node8275;
												assign node8275 = (inp[5]) ? 4'b0011 : node8276;
													assign node8276 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node8281 = (inp[13]) ? node8285 : node8282;
												assign node8282 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node8285 = (inp[4]) ? node8291 : node8286;
													assign node8286 = (inp[2]) ? node8288 : 4'b0011;
														assign node8288 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node8291 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node8294 = (inp[4]) ? node8334 : node8295;
									assign node8295 = (inp[2]) ? node8319 : node8296;
										assign node8296 = (inp[15]) ? node8312 : node8297;
											assign node8297 = (inp[11]) ? node8309 : node8298;
												assign node8298 = (inp[13]) ? node8304 : node8299;
													assign node8299 = (inp[10]) ? 4'b0011 : node8300;
														assign node8300 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node8304 = (inp[9]) ? 4'b0011 : node8305;
														assign node8305 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node8309 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node8312 = (inp[7]) ? node8314 : 4'b0010;
												assign node8314 = (inp[13]) ? 4'b0011 : node8315;
													assign node8315 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node8319 = (inp[15]) ? node8329 : node8320;
											assign node8320 = (inp[5]) ? node8326 : node8321;
												assign node8321 = (inp[7]) ? 4'b0011 : node8322;
													assign node8322 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node8326 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node8329 = (inp[13]) ? 4'b0111 : node8330;
												assign node8330 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node8334 = (inp[2]) ? node8346 : node8335;
										assign node8335 = (inp[7]) ? node8341 : node8336;
											assign node8336 = (inp[15]) ? 4'b0110 : node8337;
												assign node8337 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node8341 = (inp[10]) ? 4'b0110 : node8342;
												assign node8342 = (inp[15]) ? 4'b0111 : 4'b0110;
										assign node8346 = (inp[15]) ? node8356 : node8347;
											assign node8347 = (inp[7]) ? 4'b0010 : node8348;
												assign node8348 = (inp[10]) ? 4'b0110 : node8349;
													assign node8349 = (inp[13]) ? node8351 : 4'b0111;
														assign node8351 = (inp[11]) ? 4'b0110 : 4'b0110;
											assign node8356 = (inp[9]) ? node8358 : 4'b0010;
												assign node8358 = (inp[7]) ? node8364 : node8359;
													assign node8359 = (inp[13]) ? node8361 : 4'b0010;
														assign node8361 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node8364 = (inp[10]) ? 4'b0010 : 4'b0011;
					assign node8367 = (inp[8]) ? node8711 : node8368;
						assign node8368 = (inp[7]) ? node8550 : node8369;
							assign node8369 = (inp[15]) ? node8445 : node8370;
								assign node8370 = (inp[4]) ? node8402 : node8371;
									assign node8371 = (inp[2]) ? node8391 : node8372;
										assign node8372 = (inp[13]) ? node8384 : node8373;
											assign node8373 = (inp[1]) ? node8377 : node8374;
												assign node8374 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node8377 = (inp[9]) ? node8381 : node8378;
													assign node8378 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node8381 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node8384 = (inp[5]) ? node8388 : node8385;
												assign node8385 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node8388 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node8391 = (inp[10]) ? node8395 : node8392;
											assign node8392 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node8395 = (inp[5]) ? 4'b0101 : node8396;
												assign node8396 = (inp[9]) ? node8398 : 4'b0001;
													assign node8398 = (inp[1]) ? 4'b0101 : 4'b0001;
									assign node8402 = (inp[0]) ? node8426 : node8403;
										assign node8403 = (inp[13]) ? node8411 : node8404;
											assign node8404 = (inp[2]) ? node8406 : 4'b0110;
												assign node8406 = (inp[1]) ? node8408 : 4'b0010;
													assign node8408 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node8411 = (inp[5]) ? node8423 : node8412;
												assign node8412 = (inp[9]) ? node8418 : node8413;
													assign node8413 = (inp[1]) ? node8415 : 4'b0011;
														assign node8415 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node8418 = (inp[2]) ? 4'b0011 : node8419;
														assign node8419 = (inp[1]) ? 4'b0011 : 4'b0110;
												assign node8423 = (inp[2]) ? 4'b0111 : 4'b0011;
										assign node8426 = (inp[5]) ? node8430 : node8427;
											assign node8427 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node8430 = (inp[13]) ? node8438 : node8431;
												assign node8431 = (inp[2]) ? 4'b0010 : node8432;
													assign node8432 = (inp[10]) ? 4'b0110 : node8433;
														assign node8433 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node8438 = (inp[2]) ? node8440 : 4'b0011;
													assign node8440 = (inp[1]) ? 4'b0111 : node8441;
														assign node8441 = (inp[11]) ? 4'b0110 : 4'b0110;
								assign node8445 = (inp[0]) ? node8497 : node8446;
									assign node8446 = (inp[9]) ? node8472 : node8447;
										assign node8447 = (inp[11]) ? node8459 : node8448;
											assign node8448 = (inp[1]) ? node8456 : node8449;
												assign node8449 = (inp[5]) ? node8451 : 4'b0010;
													assign node8451 = (inp[4]) ? 4'b0010 : node8452;
														assign node8452 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node8456 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node8459 = (inp[4]) ? node8463 : node8460;
												assign node8460 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node8463 = (inp[10]) ? node8467 : node8464;
													assign node8464 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node8467 = (inp[2]) ? node8469 : 4'b0011;
														assign node8469 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node8472 = (inp[5]) ? node8482 : node8473;
											assign node8473 = (inp[2]) ? node8477 : node8474;
												assign node8474 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node8477 = (inp[13]) ? node8479 : 4'b0110;
													assign node8479 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node8482 = (inp[2]) ? node8490 : node8483;
												assign node8483 = (inp[13]) ? 4'b0110 : node8484;
													assign node8484 = (inp[10]) ? node8486 : 4'b0010;
														assign node8486 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node8490 = (inp[13]) ? node8494 : node8491;
													assign node8491 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node8494 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node8497 = (inp[4]) ? node8519 : node8498;
										assign node8498 = (inp[2]) ? node8512 : node8499;
											assign node8499 = (inp[13]) ? node8503 : node8500;
												assign node8500 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node8503 = (inp[10]) ? node8507 : node8504;
													assign node8504 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node8507 = (inp[11]) ? 4'b0110 : node8508;
														assign node8508 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node8512 = (inp[5]) ? node8516 : node8513;
												assign node8513 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node8516 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node8519 = (inp[11]) ? node8531 : node8520;
											assign node8520 = (inp[10]) ? node8528 : node8521;
												assign node8521 = (inp[1]) ? 4'b0111 : node8522;
													assign node8522 = (inp[5]) ? 4'b0110 : node8523;
														assign node8523 = (inp[9]) ? 4'b0010 : 4'b0010;
												assign node8528 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node8531 = (inp[9]) ? node8539 : node8532;
												assign node8532 = (inp[5]) ? node8536 : node8533;
													assign node8533 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node8536 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node8539 = (inp[13]) ? node8545 : node8540;
													assign node8540 = (inp[5]) ? node8542 : 4'b0111;
														assign node8542 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node8545 = (inp[10]) ? node8547 : 4'b0011;
														assign node8547 = (inp[1]) ? 4'b0011 : 4'b0111;
							assign node8550 = (inp[15]) ? node8642 : node8551;
								assign node8551 = (inp[4]) ? node8597 : node8552;
									assign node8552 = (inp[11]) ? node8576 : node8553;
										assign node8553 = (inp[10]) ? node8565 : node8554;
											assign node8554 = (inp[0]) ? node8562 : node8555;
												assign node8555 = (inp[13]) ? node8559 : node8556;
													assign node8556 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node8559 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node8562 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node8565 = (inp[5]) ? node8569 : node8566;
												assign node8566 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node8569 = (inp[13]) ? node8571 : 4'b0010;
													assign node8571 = (inp[0]) ? node8573 : 4'b0011;
														assign node8573 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node8576 = (inp[0]) ? node8584 : node8577;
											assign node8577 = (inp[2]) ? node8581 : node8578;
												assign node8578 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node8581 = (inp[1]) ? 4'b0111 : 4'b0011;
											assign node8584 = (inp[9]) ? node8588 : node8585;
												assign node8585 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node8588 = (inp[2]) ? node8592 : node8589;
													assign node8589 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node8592 = (inp[5]) ? node8594 : 4'b0010;
														assign node8594 = (inp[10]) ? 4'b0111 : 4'b0011;
									assign node8597 = (inp[0]) ? node8619 : node8598;
										assign node8598 = (inp[10]) ? node8604 : node8599;
											assign node8599 = (inp[2]) ? node8601 : 4'b0000;
												assign node8601 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node8604 = (inp[1]) ? node8614 : node8605;
												assign node8605 = (inp[9]) ? node8609 : node8606;
													assign node8606 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node8609 = (inp[13]) ? node8611 : 4'b0001;
														assign node8611 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node8614 = (inp[2]) ? 4'b0101 : node8615;
													assign node8615 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node8619 = (inp[11]) ? node8633 : node8620;
											assign node8620 = (inp[10]) ? 4'b0101 : node8621;
												assign node8621 = (inp[5]) ? node8625 : node8622;
													assign node8622 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node8625 = (inp[9]) ? node8629 : node8626;
														assign node8626 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node8629 = (inp[13]) ? 4'b0001 : 4'b0100;
											assign node8633 = (inp[13]) ? node8637 : node8634;
												assign node8634 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node8637 = (inp[5]) ? node8639 : 4'b0100;
													assign node8639 = (inp[1]) ? 4'b0000 : 4'b0100;
								assign node8642 = (inp[2]) ? node8686 : node8643;
									assign node8643 = (inp[13]) ? node8661 : node8644;
										assign node8644 = (inp[11]) ? node8646 : 4'b0001;
											assign node8646 = (inp[1]) ? node8654 : node8647;
												assign node8647 = (inp[5]) ? node8649 : 4'b0101;
													assign node8649 = (inp[4]) ? node8651 : 4'b0000;
														assign node8651 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node8654 = (inp[0]) ? 4'b0000 : node8655;
													assign node8655 = (inp[4]) ? 4'b0000 : node8656;
														assign node8656 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node8661 = (inp[5]) ? node8673 : node8662;
											assign node8662 = (inp[1]) ? node8664 : 4'b0000;
												assign node8664 = (inp[9]) ? node8668 : node8665;
													assign node8665 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node8668 = (inp[10]) ? 4'b0100 : node8669;
														assign node8669 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node8673 = (inp[11]) ? node8677 : node8674;
												assign node8674 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node8677 = (inp[4]) ? node8681 : node8678;
													assign node8678 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node8681 = (inp[10]) ? 4'b0101 : node8682;
														assign node8682 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node8686 = (inp[13]) ? node8702 : node8687;
										assign node8687 = (inp[1]) ? node8693 : node8688;
											assign node8688 = (inp[5]) ? 4'b0101 : node8689;
												assign node8689 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node8693 = (inp[5]) ? node8697 : node8694;
												assign node8694 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node8697 = (inp[10]) ? 4'b0100 : node8698;
													assign node8698 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node8702 = (inp[1]) ? node8706 : node8703;
											assign node8703 = (inp[5]) ? 4'b0001 : 4'b0101;
											assign node8706 = (inp[4]) ? node8708 : 4'b0001;
												assign node8708 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node8711 = (inp[2]) ? node8851 : node8712;
							assign node8712 = (inp[15]) ? node8792 : node8713;
								assign node8713 = (inp[7]) ? node8757 : node8714;
									assign node8714 = (inp[5]) ? node8730 : node8715;
										assign node8715 = (inp[4]) ? node8723 : node8716;
											assign node8716 = (inp[10]) ? node8718 : 4'b0101;
												assign node8718 = (inp[0]) ? 4'b0101 : node8719;
													assign node8719 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node8723 = (inp[11]) ? node8725 : 4'b0000;
												assign node8725 = (inp[9]) ? 4'b0001 : node8726;
													assign node8726 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node8730 = (inp[0]) ? node8744 : node8731;
											assign node8731 = (inp[4]) ? node8737 : node8732;
												assign node8732 = (inp[11]) ? node8734 : 4'b0000;
													assign node8734 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node8737 = (inp[1]) ? node8739 : 4'b0001;
													assign node8739 = (inp[11]) ? 4'b0001 : node8740;
														assign node8740 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node8744 = (inp[11]) ? 4'b0000 : node8745;
												assign node8745 = (inp[10]) ? node8751 : node8746;
													assign node8746 = (inp[13]) ? node8748 : 4'b0000;
														assign node8748 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node8751 = (inp[1]) ? node8753 : 4'b0001;
														assign node8753 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node8757 = (inp[4]) ? node8777 : node8758;
										assign node8758 = (inp[5]) ? node8764 : node8759;
											assign node8759 = (inp[0]) ? node8761 : 4'b0000;
												assign node8761 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node8764 = (inp[1]) ? node8772 : node8765;
												assign node8765 = (inp[11]) ? node8767 : 4'b0100;
													assign node8767 = (inp[9]) ? 4'b0101 : node8768;
														assign node8768 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node8772 = (inp[11]) ? node8774 : 4'b0101;
													assign node8774 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node8777 = (inp[13]) ? node8783 : node8778;
											assign node8778 = (inp[5]) ? node8780 : 4'b0101;
												assign node8780 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node8783 = (inp[10]) ? node8787 : node8784;
												assign node8784 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node8787 = (inp[11]) ? 4'b0100 : node8788;
													assign node8788 = (inp[1]) ? 4'b0100 : 4'b0101;
								assign node8792 = (inp[13]) ? node8816 : node8793;
									assign node8793 = (inp[5]) ? node8809 : node8794;
										assign node8794 = (inp[7]) ? node8802 : node8795;
											assign node8795 = (inp[10]) ? 4'b0101 : node8796;
												assign node8796 = (inp[1]) ? node8798 : 4'b0100;
													assign node8798 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node8802 = (inp[4]) ? 4'b0100 : node8803;
												assign node8803 = (inp[9]) ? 4'b0101 : node8804;
													assign node8804 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node8809 = (inp[10]) ? node8813 : node8810;
											assign node8810 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node8813 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node8816 = (inp[11]) ? node8834 : node8817;
										assign node8817 = (inp[7]) ? node8825 : node8818;
											assign node8818 = (inp[10]) ? 4'b0101 : node8819;
												assign node8819 = (inp[9]) ? node8821 : 4'b0100;
													assign node8821 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node8825 = (inp[0]) ? node8827 : 4'b0100;
												assign node8827 = (inp[1]) ? 4'b0101 : node8828;
													assign node8828 = (inp[5]) ? node8830 : 4'b0100;
														assign node8830 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node8834 = (inp[7]) ? node8842 : node8835;
											assign node8835 = (inp[10]) ? node8837 : 4'b0101;
												assign node8837 = (inp[9]) ? 4'b0100 : node8838;
													assign node8838 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node8842 = (inp[0]) ? node8844 : 4'b0101;
												assign node8844 = (inp[4]) ? node8848 : node8845;
													assign node8845 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node8848 = (inp[10]) ? 4'b0100 : 4'b0101;
							assign node8851 = (inp[15]) ? node8935 : node8852;
								assign node8852 = (inp[7]) ? node8890 : node8853;
									assign node8853 = (inp[5]) ? node8871 : node8854;
										assign node8854 = (inp[4]) ? node8862 : node8855;
											assign node8855 = (inp[13]) ? 4'b0001 : node8856;
												assign node8856 = (inp[11]) ? node8858 : 4'b0000;
													assign node8858 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node8862 = (inp[13]) ? 4'b0101 : node8863;
												assign node8863 = (inp[0]) ? node8865 : 4'b0100;
													assign node8865 = (inp[10]) ? node8867 : 4'b0101;
														assign node8867 = (inp[1]) ? 4'b0100 : 4'b0100;
										assign node8871 = (inp[0]) ? node8883 : node8872;
											assign node8872 = (inp[9]) ? node8876 : node8873;
												assign node8873 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node8876 = (inp[4]) ? node8878 : 4'b0101;
													assign node8878 = (inp[11]) ? 4'b0101 : node8879;
														assign node8879 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node8883 = (inp[4]) ? 4'b0100 : node8884;
												assign node8884 = (inp[10]) ? node8886 : 4'b0101;
													assign node8886 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node8890 = (inp[5]) ? node8912 : node8891;
										assign node8891 = (inp[4]) ? node8901 : node8892;
											assign node8892 = (inp[13]) ? node8894 : 4'b0101;
												assign node8894 = (inp[0]) ? 4'b0100 : node8895;
													assign node8895 = (inp[9]) ? 4'b0101 : node8896;
														assign node8896 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node8901 = (inp[9]) ? 4'b0001 : node8902;
												assign node8902 = (inp[10]) ? node8908 : node8903;
													assign node8903 = (inp[1]) ? 4'b0000 : node8904;
														assign node8904 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node8908 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node8912 = (inp[9]) ? node8924 : node8913;
											assign node8913 = (inp[4]) ? 4'b0001 : node8914;
												assign node8914 = (inp[10]) ? node8918 : node8915;
													assign node8915 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node8918 = (inp[13]) ? node8920 : 4'b0001;
														assign node8920 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node8924 = (inp[1]) ? node8930 : node8925;
												assign node8925 = (inp[4]) ? 4'b0000 : node8926;
													assign node8926 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node8930 = (inp[10]) ? node8932 : 4'b0001;
													assign node8932 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node8935 = (inp[1]) ? node8947 : node8936;
									assign node8936 = (inp[7]) ? node8938 : 4'b0000;
										assign node8938 = (inp[10]) ? node8942 : node8939;
											assign node8939 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node8942 = (inp[11]) ? 4'b0000 : node8943;
												assign node8943 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node8947 = (inp[10]) ? node8961 : node8948;
										assign node8948 = (inp[5]) ? 4'b0001 : node8949;
											assign node8949 = (inp[7]) ? node8955 : node8950;
												assign node8950 = (inp[11]) ? 4'b0000 : node8951;
													assign node8951 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node8955 = (inp[11]) ? 4'b0001 : node8956;
													assign node8956 = (inp[4]) ? 4'b0001 : 4'b0000;
										assign node8961 = (inp[5]) ? 4'b0000 : node8962;
											assign node8962 = (inp[4]) ? node8964 : 4'b0001;
												assign node8964 = (inp[7]) ? 4'b0000 : 4'b0001;
				assign node8968 = (inp[8]) ? node9450 : node8969;
					assign node8969 = (inp[7]) ? node9235 : node8970;
						assign node8970 = (inp[15]) ? node9100 : node8971;
							assign node8971 = (inp[13]) ? node9047 : node8972;
								assign node8972 = (inp[4]) ? node9024 : node8973;
									assign node8973 = (inp[11]) ? node8997 : node8974;
										assign node8974 = (inp[12]) ? node8986 : node8975;
											assign node8975 = (inp[1]) ? node8983 : node8976;
												assign node8976 = (inp[5]) ? node8978 : 4'b0010;
													assign node8978 = (inp[10]) ? 4'b0011 : node8979;
														assign node8979 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node8983 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node8986 = (inp[1]) ? 4'b0011 : node8987;
												assign node8987 = (inp[9]) ? node8991 : node8988;
													assign node8988 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node8991 = (inp[2]) ? 4'b0110 : node8992;
														assign node8992 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node8997 = (inp[1]) ? node9011 : node8998;
											assign node8998 = (inp[2]) ? 4'b0011 : node8999;
												assign node8999 = (inp[0]) ? node9003 : node9000;
													assign node9000 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node9003 = (inp[9]) ? node9007 : node9004;
														assign node9004 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node9007 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node9011 = (inp[12]) ? node9017 : node9012;
												assign node9012 = (inp[0]) ? 4'b0111 : node9013;
													assign node9013 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node9017 = (inp[2]) ? node9019 : 4'b0011;
													assign node9019 = (inp[10]) ? node9021 : 4'b0010;
														assign node9021 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node9024 = (inp[5]) ? node9030 : node9025;
										assign node9025 = (inp[0]) ? node9027 : 4'b0011;
											assign node9027 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node9030 = (inp[9]) ? 4'b0010 : node9031;
											assign node9031 = (inp[0]) ? node9033 : 4'b0011;
												assign node9033 = (inp[10]) ? node9041 : node9034;
													assign node9034 = (inp[11]) ? node9038 : node9035;
														assign node9035 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node9038 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node9041 = (inp[11]) ? node9043 : 4'b0010;
														assign node9043 = (inp[1]) ? 4'b0010 : 4'b0010;
								assign node9047 = (inp[4]) ? node9081 : node9048;
									assign node9048 = (inp[12]) ? node9062 : node9049;
										assign node9049 = (inp[1]) ? node9055 : node9050;
											assign node9050 = (inp[0]) ? node9052 : 4'b0110;
												assign node9052 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node9055 = (inp[9]) ? node9057 : 4'b0010;
												assign node9057 = (inp[11]) ? 4'b0011 : node9058;
													assign node9058 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node9062 = (inp[1]) ? node9066 : node9063;
											assign node9063 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node9066 = (inp[5]) ? node9076 : node9067;
												assign node9067 = (inp[2]) ? 4'b0111 : node9068;
													assign node9068 = (inp[11]) ? node9072 : node9069;
														assign node9069 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node9072 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node9076 = (inp[11]) ? node9078 : 4'b0110;
													assign node9078 = (inp[2]) ? 4'b0111 : 4'b0110;
									assign node9081 = (inp[2]) ? node9087 : node9082;
										assign node9082 = (inp[5]) ? node9084 : 4'b0110;
											assign node9084 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node9087 = (inp[11]) ? node9095 : node9088;
											assign node9088 = (inp[10]) ? node9090 : 4'b0110;
												assign node9090 = (inp[9]) ? node9092 : 4'b0111;
													assign node9092 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node9095 = (inp[12]) ? 4'b0111 : node9096;
												assign node9096 = (inp[1]) ? 4'b0110 : 4'b0111;
							assign node9100 = (inp[13]) ? node9168 : node9101;
								assign node9101 = (inp[12]) ? node9129 : node9102;
									assign node9102 = (inp[4]) ? node9116 : node9103;
										assign node9103 = (inp[5]) ? node9111 : node9104;
											assign node9104 = (inp[11]) ? 4'b0010 : node9105;
												assign node9105 = (inp[2]) ? 4'b0011 : node9106;
													assign node9106 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node9111 = (inp[2]) ? node9113 : 4'b0011;
												assign node9113 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node9116 = (inp[9]) ? node9122 : node9117;
											assign node9117 = (inp[1]) ? node9119 : 4'b0111;
												assign node9119 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node9122 = (inp[10]) ? 4'b0110 : node9123;
												assign node9123 = (inp[5]) ? node9125 : 4'b0110;
													assign node9125 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node9129 = (inp[11]) ? node9141 : node9130;
										assign node9130 = (inp[0]) ? 4'b0110 : node9131;
											assign node9131 = (inp[2]) ? 4'b0111 : node9132;
												assign node9132 = (inp[9]) ? 4'b0111 : node9133;
													assign node9133 = (inp[10]) ? node9135 : 4'b0110;
														assign node9135 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node9141 = (inp[2]) ? node9157 : node9142;
											assign node9142 = (inp[0]) ? node9150 : node9143;
												assign node9143 = (inp[9]) ? node9147 : node9144;
													assign node9144 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node9147 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node9150 = (inp[1]) ? 4'b0111 : node9151;
													assign node9151 = (inp[9]) ? node9153 : 4'b0111;
														assign node9153 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node9157 = (inp[4]) ? node9163 : node9158;
												assign node9158 = (inp[0]) ? node9160 : 4'b0111;
													assign node9160 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node9163 = (inp[0]) ? node9165 : 4'b0110;
													assign node9165 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node9168 = (inp[12]) ? node9214 : node9169;
									assign node9169 = (inp[4]) ? node9197 : node9170;
										assign node9170 = (inp[10]) ? node9184 : node9171;
											assign node9171 = (inp[11]) ? node9173 : 4'b0111;
												assign node9173 = (inp[1]) ? node9179 : node9174;
													assign node9174 = (inp[5]) ? node9176 : 4'b0111;
														assign node9176 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node9179 = (inp[0]) ? 4'b0110 : node9180;
														assign node9180 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node9184 = (inp[9]) ? node9190 : node9185;
												assign node9185 = (inp[5]) ? node9187 : 4'b0111;
													assign node9187 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node9190 = (inp[5]) ? 4'b0111 : node9191;
													assign node9191 = (inp[11]) ? node9193 : 4'b0110;
														assign node9193 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node9197 = (inp[1]) ? node9205 : node9198;
											assign node9198 = (inp[9]) ? node9200 : 4'b0010;
												assign node9200 = (inp[5]) ? node9202 : 4'b0011;
													assign node9202 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node9205 = (inp[11]) ? 4'b0011 : node9206;
												assign node9206 = (inp[9]) ? node9210 : node9207;
													assign node9207 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node9210 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node9214 = (inp[4]) ? node9226 : node9215;
										assign node9215 = (inp[2]) ? node9219 : node9216;
											assign node9216 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node9219 = (inp[11]) ? node9221 : 4'b0010;
												assign node9221 = (inp[0]) ? 4'b0011 : node9222;
													assign node9222 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node9226 = (inp[1]) ? 4'b0010 : node9227;
											assign node9227 = (inp[0]) ? 4'b0010 : node9228;
												assign node9228 = (inp[10]) ? 4'b0010 : node9229;
													assign node9229 = (inp[5]) ? 4'b0011 : 4'b0010;
						assign node9235 = (inp[13]) ? node9365 : node9236;
							assign node9236 = (inp[4]) ? node9312 : node9237;
								assign node9237 = (inp[12]) ? node9269 : node9238;
									assign node9238 = (inp[15]) ? node9252 : node9239;
										assign node9239 = (inp[1]) ? node9249 : node9240;
											assign node9240 = (inp[2]) ? 4'b0101 : node9241;
												assign node9241 = (inp[0]) ? 4'b0100 : node9242;
													assign node9242 = (inp[9]) ? 4'b0101 : node9243;
														assign node9243 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node9249 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node9252 = (inp[1]) ? node9260 : node9253;
											assign node9253 = (inp[5]) ? node9255 : 4'b0000;
												assign node9255 = (inp[10]) ? 4'b0001 : node9256;
													assign node9256 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node9260 = (inp[2]) ? node9266 : node9261;
												assign node9261 = (inp[0]) ? 4'b0001 : node9262;
													assign node9262 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node9266 = (inp[9]) ? 4'b0001 : 4'b0000;
									assign node9269 = (inp[1]) ? node9281 : node9270;
										assign node9270 = (inp[15]) ? node9276 : node9271;
											assign node9271 = (inp[9]) ? 4'b0001 : node9272;
												assign node9272 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node9276 = (inp[9]) ? node9278 : 4'b0100;
												assign node9278 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node9281 = (inp[5]) ? node9289 : node9282;
											assign node9282 = (inp[15]) ? 4'b0100 : node9283;
												assign node9283 = (inp[9]) ? node9285 : 4'b0100;
													assign node9285 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node9289 = (inp[2]) ? node9297 : node9290;
												assign node9290 = (inp[0]) ? node9292 : 4'b0101;
													assign node9292 = (inp[15]) ? node9294 : 4'b0101;
														assign node9294 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node9297 = (inp[11]) ? node9305 : node9298;
													assign node9298 = (inp[10]) ? node9302 : node9299;
														assign node9299 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node9302 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node9305 = (inp[0]) ? node9309 : node9306;
														assign node9306 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node9309 = (inp[9]) ? 4'b0101 : 4'b0100;
								assign node9312 = (inp[2]) ? node9340 : node9313;
									assign node9313 = (inp[11]) ? node9331 : node9314;
										assign node9314 = (inp[0]) ? node9320 : node9315;
											assign node9315 = (inp[1]) ? node9317 : 4'b0101;
												assign node9317 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node9320 = (inp[9]) ? 4'b0100 : node9321;
												assign node9321 = (inp[5]) ? node9323 : 4'b0101;
													assign node9323 = (inp[12]) ? node9327 : node9324;
														assign node9324 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node9327 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node9331 = (inp[5]) ? node9337 : node9332;
											assign node9332 = (inp[12]) ? 4'b0100 : node9333;
												assign node9333 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node9337 = (inp[12]) ? 4'b0101 : 4'b0100;
									assign node9340 = (inp[0]) ? node9350 : node9341;
										assign node9341 = (inp[5]) ? 4'b0101 : node9342;
											assign node9342 = (inp[1]) ? 4'b0101 : node9343;
												assign node9343 = (inp[9]) ? node9345 : 4'b0100;
													assign node9345 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node9350 = (inp[10]) ? node9360 : node9351;
											assign node9351 = (inp[12]) ? 4'b0101 : node9352;
												assign node9352 = (inp[15]) ? node9354 : 4'b0100;
													assign node9354 = (inp[5]) ? 4'b0101 : node9355;
														assign node9355 = (inp[9]) ? 4'b0100 : 4'b0100;
											assign node9360 = (inp[12]) ? node9362 : 4'b0101;
												assign node9362 = (inp[9]) ? 4'b0100 : 4'b0101;
							assign node9365 = (inp[4]) ? node9427 : node9366;
								assign node9366 = (inp[12]) ? node9400 : node9367;
									assign node9367 = (inp[1]) ? node9381 : node9368;
										assign node9368 = (inp[15]) ? node9372 : node9369;
											assign node9369 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node9372 = (inp[9]) ? node9374 : 4'b0101;
												assign node9374 = (inp[2]) ? 4'b0101 : node9375;
													assign node9375 = (inp[11]) ? node9377 : 4'b0100;
														assign node9377 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node9381 = (inp[15]) ? node9393 : node9382;
											assign node9382 = (inp[5]) ? node9384 : 4'b0101;
												assign node9384 = (inp[11]) ? node9388 : node9385;
													assign node9385 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node9388 = (inp[10]) ? node9390 : 4'b0101;
														assign node9390 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node9393 = (inp[2]) ? 4'b0100 : node9394;
												assign node9394 = (inp[9]) ? 4'b0101 : node9395;
													assign node9395 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node9400 = (inp[1]) ? node9412 : node9401;
										assign node9401 = (inp[15]) ? 4'b0001 : node9402;
											assign node9402 = (inp[9]) ? 4'b0101 : node9403;
												assign node9403 = (inp[11]) ? node9405 : 4'b0100;
													assign node9405 = (inp[0]) ? node9407 : 4'b0101;
														assign node9407 = (inp[10]) ? 4'b0100 : 4'b0100;
										assign node9412 = (inp[15]) ? node9418 : node9413;
											assign node9413 = (inp[9]) ? node9415 : 4'b0001;
												assign node9415 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node9418 = (inp[10]) ? 4'b0000 : node9419;
												assign node9419 = (inp[9]) ? node9421 : 4'b0001;
													assign node9421 = (inp[2]) ? 4'b0000 : node9422;
														assign node9422 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node9427 = (inp[9]) ? node9439 : node9428;
									assign node9428 = (inp[1]) ? 4'b0001 : node9429;
										assign node9429 = (inp[12]) ? node9435 : node9430;
											assign node9430 = (inp[15]) ? 4'b0000 : node9431;
												assign node9431 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node9435 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node9439 = (inp[1]) ? 4'b0000 : node9440;
										assign node9440 = (inp[12]) ? node9444 : node9441;
											assign node9441 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node9444 = (inp[15]) ? 4'b0000 : node9445;
												assign node9445 = (inp[11]) ? 4'b0000 : 4'b0001;
					assign node9450 = (inp[15]) ? node9608 : node9451;
						assign node9451 = (inp[7]) ? node9537 : node9452;
							assign node9452 = (inp[12]) ? node9506 : node9453;
								assign node9453 = (inp[4]) ? node9485 : node9454;
									assign node9454 = (inp[10]) ? node9466 : node9455;
										assign node9455 = (inp[0]) ? 4'b0001 : node9456;
											assign node9456 = (inp[5]) ? node9460 : node9457;
												assign node9457 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node9460 = (inp[11]) ? node9462 : 4'b0001;
													assign node9462 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node9466 = (inp[2]) ? node9480 : node9467;
											assign node9467 = (inp[9]) ? node9475 : node9468;
												assign node9468 = (inp[1]) ? node9470 : 4'b0001;
													assign node9470 = (inp[11]) ? node9472 : 4'b0000;
														assign node9472 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node9475 = (inp[13]) ? 4'b0000 : node9476;
													assign node9476 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node9480 = (inp[1]) ? 4'b0000 : node9481;
												assign node9481 = (inp[13]) ? 4'b0000 : 4'b0001;
									assign node9485 = (inp[2]) ? node9493 : node9486;
										assign node9486 = (inp[5]) ? node9490 : node9487;
											assign node9487 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node9490 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node9493 = (inp[11]) ? node9501 : node9494;
											assign node9494 = (inp[13]) ? node9498 : node9495;
												assign node9495 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node9498 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node9501 = (inp[5]) ? 4'b0100 : node9502;
												assign node9502 = (inp[9]) ? 4'b0100 : 4'b0101;
								assign node9506 = (inp[5]) ? node9526 : node9507;
									assign node9507 = (inp[13]) ? node9515 : node9508;
										assign node9508 = (inp[4]) ? 4'b0100 : node9509;
											assign node9509 = (inp[2]) ? 4'b0101 : node9510;
												assign node9510 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node9515 = (inp[4]) ? 4'b0101 : node9516;
											assign node9516 = (inp[11]) ? node9518 : 4'b0100;
												assign node9518 = (inp[10]) ? 4'b0101 : node9519;
													assign node9519 = (inp[9]) ? node9521 : 4'b0101;
														assign node9521 = (inp[2]) ? 4'b0100 : 4'b0100;
									assign node9526 = (inp[13]) ? node9532 : node9527;
										assign node9527 = (inp[2]) ? 4'b0101 : node9528;
											assign node9528 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node9532 = (inp[4]) ? 4'b0100 : node9533;
											assign node9533 = (inp[2]) ? 4'b0100 : 4'b0101;
							assign node9537 = (inp[4]) ? node9597 : node9538;
								assign node9538 = (inp[12]) ? node9570 : node9539;
									assign node9539 = (inp[0]) ? node9555 : node9540;
										assign node9540 = (inp[11]) ? node9546 : node9541;
											assign node9541 = (inp[9]) ? node9543 : 4'b0100;
												assign node9543 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node9546 = (inp[10]) ? 4'b0101 : node9547;
												assign node9547 = (inp[2]) ? 4'b0101 : node9548;
													assign node9548 = (inp[9]) ? 4'b0100 : node9549;
														assign node9549 = (inp[1]) ? 4'b0100 : 4'b0100;
										assign node9555 = (inp[13]) ? node9563 : node9556;
											assign node9556 = (inp[2]) ? node9558 : 4'b0100;
												assign node9558 = (inp[9]) ? node9560 : 4'b0101;
													assign node9560 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node9563 = (inp[2]) ? node9565 : 4'b0101;
												assign node9565 = (inp[1]) ? 4'b0100 : node9566;
													assign node9566 = (inp[5]) ? 4'b0101 : 4'b0100;
									assign node9570 = (inp[11]) ? node9588 : node9571;
										assign node9571 = (inp[5]) ? node9581 : node9572;
											assign node9572 = (inp[1]) ? node9578 : node9573;
												assign node9573 = (inp[13]) ? 4'b0000 : node9574;
													assign node9574 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node9578 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node9581 = (inp[1]) ? 4'b0000 : node9582;
												assign node9582 = (inp[10]) ? 4'b0001 : node9583;
													assign node9583 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node9588 = (inp[10]) ? 4'b0000 : node9589;
											assign node9589 = (inp[5]) ? node9591 : 4'b0000;
												assign node9591 = (inp[2]) ? node9593 : 4'b0001;
													assign node9593 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node9597 = (inp[13]) ? node9603 : node9598;
									assign node9598 = (inp[12]) ? 4'b0001 : node9599;
										assign node9599 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node9603 = (inp[1]) ? 4'b0000 : node9604;
										assign node9604 = (inp[12]) ? 4'b0000 : 4'b0001;
						assign node9608 = (inp[4]) ? node9658 : node9609;
							assign node9609 = (inp[12]) ? node9647 : node9610;
								assign node9610 = (inp[10]) ? node9630 : node9611;
									assign node9611 = (inp[7]) ? node9619 : node9612;
										assign node9612 = (inp[2]) ? node9616 : node9613;
											assign node9613 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node9616 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node9619 = (inp[0]) ? 4'b0100 : node9620;
											assign node9620 = (inp[13]) ? node9622 : 4'b0100;
												assign node9622 = (inp[11]) ? node9624 : 4'b0101;
													assign node9624 = (inp[1]) ? node9626 : 4'b0100;
														assign node9626 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node9630 = (inp[7]) ? node9640 : node9631;
										assign node9631 = (inp[11]) ? node9633 : 4'b0100;
											assign node9633 = (inp[2]) ? node9637 : node9634;
												assign node9634 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node9637 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node9640 = (inp[1]) ? node9644 : node9641;
											assign node9641 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node9644 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node9647 = (inp[2]) ? node9653 : node9648;
									assign node9648 = (inp[7]) ? 4'b0001 : node9649;
										assign node9649 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node9653 = (inp[5]) ? 4'b0000 : node9654;
										assign node9654 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node9658 = (inp[7]) ? node9670 : node9659;
								assign node9659 = (inp[5]) ? node9665 : node9660;
									assign node9660 = (inp[1]) ? 4'b0001 : node9661;
										assign node9661 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node9665 = (inp[1]) ? 4'b0000 : node9666;
										assign node9666 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node9670 = (inp[12]) ? 4'b0000 : node9671;
									assign node9671 = (inp[1]) ? 4'b0000 : 4'b0001;

endmodule