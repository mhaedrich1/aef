module dtc_split125_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;

	assign outp = (inp[6]) ? node68 : node1;
		assign node1 = (inp[7]) ? node3 : 3'b000;
			assign node3 = (inp[0]) ? node49 : node4;
				assign node4 = (inp[9]) ? node30 : node5;
					assign node5 = (inp[10]) ? node23 : node6;
						assign node6 = (inp[1]) ? node10 : node7;
							assign node7 = (inp[11]) ? 3'b001 : 3'b101;
							assign node10 = (inp[5]) ? node16 : node11;
								assign node11 = (inp[2]) ? 3'b110 : node12;
									assign node12 = (inp[11]) ? 3'b110 : 3'b001;
								assign node16 = (inp[11]) ? node18 : 3'b110;
									assign node18 = (inp[8]) ? node20 : 3'b010;
										assign node20 = (inp[4]) ? 3'b110 : 3'b010;
						assign node23 = (inp[1]) ? node25 : 3'b110;
							assign node25 = (inp[4]) ? 3'b100 : node26;
								assign node26 = (inp[8]) ? 3'b010 : 3'b000;
					assign node30 = (inp[10]) ? 3'b000 : node31;
						assign node31 = (inp[4]) ? node43 : node32;
							assign node32 = (inp[2]) ? node38 : node33;
								assign node33 = (inp[11]) ? 3'b110 : node34;
									assign node34 = (inp[1]) ? 3'b000 : 3'b010;
								assign node38 = (inp[1]) ? 3'b000 : node39;
									assign node39 = (inp[11]) ? 3'b000 : 3'b100;
							assign node43 = (inp[2]) ? 3'b100 : node44;
								assign node44 = (inp[11]) ? 3'b100 : 3'b000;
				assign node49 = (inp[9]) ? 3'b000 : node50;
					assign node50 = (inp[10]) ? 3'b000 : node51;
						assign node51 = (inp[1]) ? node59 : node52;
							assign node52 = (inp[11]) ? node56 : node53;
								assign node53 = (inp[4]) ? 3'b010 : 3'b110;
								assign node56 = (inp[2]) ? 3'b100 : 3'b010;
							assign node59 = (inp[8]) ? node61 : 3'b000;
								assign node61 = (inp[11]) ? node63 : 3'b100;
									assign node63 = (inp[2]) ? 3'b000 : 3'b100;
		assign node68 = (inp[9]) ? node212 : node69;
			assign node69 = (inp[7]) ? node139 : node70;
				assign node70 = (inp[0]) ? node108 : node71;
					assign node71 = (inp[3]) ? node85 : node72;
						assign node72 = (inp[4]) ? node82 : node73;
							assign node73 = (inp[1]) ? node75 : 3'b001;
								assign node75 = (inp[11]) ? 3'b110 : node76;
									assign node76 = (inp[8]) ? 3'b101 : node77;
										assign node77 = (inp[10]) ? 3'b001 : 3'b101;
							assign node82 = (inp[11]) ? 3'b001 : 3'b011;
						assign node85 = (inp[1]) ? node97 : node86;
							assign node86 = (inp[8]) ? 3'b011 : node87;
								assign node87 = (inp[4]) ? 3'b101 : node88;
									assign node88 = (inp[10]) ? node90 : 3'b011;
										assign node90 = (inp[11]) ? node92 : 3'b001;
											assign node92 = (inp[2]) ? 3'b111 : 3'b001;
							assign node97 = (inp[8]) ? node103 : node98;
								assign node98 = (inp[11]) ? 3'b010 : node99;
									assign node99 = (inp[2]) ? 3'b010 : 3'b110;
								assign node103 = (inp[2]) ? node105 : 3'b011;
									assign node105 = (inp[4]) ? 3'b001 : 3'b101;
					assign node108 = (inp[8]) ? node124 : node109;
						assign node109 = (inp[10]) ? node115 : node110;
							assign node110 = (inp[3]) ? node112 : 3'b001;
								assign node112 = (inp[11]) ? 3'b010 : 3'b110;
							assign node115 = (inp[4]) ? node121 : node116;
								assign node116 = (inp[3]) ? node118 : 3'b100;
									assign node118 = (inp[2]) ? 3'b000 : 3'b100;
								assign node121 = (inp[2]) ? 3'b000 : 3'b010;
						assign node124 = (inp[11]) ? node132 : node125;
							assign node125 = (inp[2]) ? node129 : node126;
								assign node126 = (inp[10]) ? 3'b110 : 3'b101;
								assign node129 = (inp[10]) ? 3'b100 : 3'b110;
							assign node132 = (inp[4]) ? node134 : 3'b110;
								assign node134 = (inp[2]) ? node136 : 3'b010;
									assign node136 = (inp[3]) ? 3'b000 : 3'b001;
				assign node139 = (inp[0]) ? node161 : node140;
					assign node140 = (inp[10]) ? node142 : 3'b111;
						assign node142 = (inp[11]) ? node150 : node143;
							assign node143 = (inp[2]) ? node147 : node144;
								assign node144 = (inp[1]) ? 3'b101 : 3'b111;
								assign node147 = (inp[3]) ? 3'b011 : 3'b111;
							assign node150 = (inp[4]) ? node156 : node151;
								assign node151 = (inp[8]) ? node153 : 3'b001;
									assign node153 = (inp[2]) ? 3'b011 : 3'b111;
								assign node156 = (inp[2]) ? 3'b101 : node157;
									assign node157 = (inp[3]) ? 3'b101 : 3'b001;
					assign node161 = (inp[10]) ? node183 : node162;
						assign node162 = (inp[2]) ? node168 : node163;
							assign node163 = (inp[3]) ? node165 : 3'b011;
								assign node165 = (inp[1]) ? 3'b101 : 3'b011;
							assign node168 = (inp[11]) ? node176 : node169;
								assign node169 = (inp[1]) ? node173 : node170;
									assign node170 = (inp[8]) ? 3'b011 : 3'b101;
									assign node173 = (inp[8]) ? 3'b101 : 3'b001;
								assign node176 = (inp[8]) ? node180 : node177;
									assign node177 = (inp[1]) ? 3'b111 : 3'b101;
									assign node180 = (inp[1]) ? 3'b001 : 3'b011;
						assign node183 = (inp[1]) ? node201 : node184;
							assign node184 = (inp[4]) ? node194 : node185;
								assign node185 = (inp[11]) ? node191 : node186;
									assign node186 = (inp[3]) ? node188 : 3'b101;
										assign node188 = (inp[5]) ? 3'b001 : 3'b101;
									assign node191 = (inp[5]) ? 3'b101 : 3'b001;
								assign node194 = (inp[8]) ? node198 : node195;
									assign node195 = (inp[5]) ? 3'b110 : 3'b010;
									assign node198 = (inp[3]) ? 3'b001 : 3'b101;
							assign node201 = (inp[8]) ? node207 : node202;
								assign node202 = (inp[2]) ? 3'b010 : node203;
									assign node203 = (inp[11]) ? 3'b010 : 3'b110;
								assign node207 = (inp[11]) ? 3'b110 : node208;
									assign node208 = (inp[2]) ? 3'b111 : 3'b001;
			assign node212 = (inp[0]) ? node284 : node213;
				assign node213 = (inp[7]) ? node245 : node214;
					assign node214 = (inp[8]) ? node230 : node215;
						assign node215 = (inp[1]) ? node225 : node216;
							assign node216 = (inp[11]) ? node222 : node217;
								assign node217 = (inp[2]) ? node219 : 3'b100;
									assign node219 = (inp[4]) ? 3'b000 : 3'b010;
								assign node222 = (inp[2]) ? 3'b100 : 3'b000;
							assign node225 = (inp[11]) ? 3'b000 : node226;
								assign node226 = (inp[3]) ? 3'b000 : 3'b100;
						assign node230 = (inp[3]) ? node242 : node231;
							assign node231 = (inp[10]) ? node237 : node232;
								assign node232 = (inp[2]) ? 3'b010 : node233;
									assign node233 = (inp[4]) ? 3'b110 : 3'b001;
								assign node237 = (inp[4]) ? 3'b100 : node238;
									assign node238 = (inp[5]) ? 3'b010 : 3'b110;
							assign node242 = (inp[1]) ? 3'b000 : 3'b010;
					assign node245 = (inp[8]) ? node263 : node246;
						assign node246 = (inp[1]) ? node252 : node247;
							assign node247 = (inp[2]) ? node249 : 3'b101;
								assign node249 = (inp[11]) ? 3'b110 : 3'b101;
							assign node252 = (inp[10]) ? 3'b100 : node253;
								assign node253 = (inp[2]) ? node259 : node254;
									assign node254 = (inp[3]) ? node256 : 3'b110;
										assign node256 = (inp[4]) ? 3'b010 : 3'b110;
									assign node259 = (inp[11]) ? 3'b001 : 3'b110;
						assign node263 = (inp[10]) ? node275 : node264;
							assign node264 = (inp[11]) ? node270 : node265;
								assign node265 = (inp[3]) ? node267 : 3'b101;
									assign node267 = (inp[4]) ? 3'b001 : 3'b101;
								assign node270 = (inp[1]) ? 3'b010 : node271;
									assign node271 = (inp[2]) ? 3'b001 : 3'b101;
							assign node275 = (inp[4]) ? node279 : node276;
								assign node276 = (inp[11]) ? 3'b010 : 3'b001;
								assign node279 = (inp[3]) ? 3'b010 : node280;
									assign node280 = (inp[1]) ? 3'b100 : 3'b110;
				assign node284 = (inp[10]) ? node318 : node285;
					assign node285 = (inp[1]) ? node303 : node286;
						assign node286 = (inp[4]) ? node296 : node287;
							assign node287 = (inp[5]) ? 3'b010 : node288;
								assign node288 = (inp[11]) ? node290 : 3'b010;
									assign node290 = (inp[7]) ? 3'b100 : node291;
										assign node291 = (inp[2]) ? 3'b010 : 3'b100;
							assign node296 = (inp[7]) ? node298 : 3'b100;
								assign node298 = (inp[8]) ? 3'b010 : node299;
									assign node299 = (inp[11]) ? 3'b000 : 3'b100;
						assign node303 = (inp[7]) ? node305 : 3'b000;
							assign node305 = (inp[8]) ? node313 : node306;
								assign node306 = (inp[5]) ? 3'b000 : node307;
									assign node307 = (inp[4]) ? 3'b100 : node308;
										assign node308 = (inp[2]) ? 3'b100 : 3'b000;
								assign node313 = (inp[11]) ? node315 : 3'b010;
									assign node315 = (inp[4]) ? 3'b100 : 3'b110;
					assign node318 = (inp[1]) ? 3'b000 : node319;
						assign node319 = (inp[11]) ? 3'b000 : node320;
							assign node320 = (inp[3]) ? 3'b100 : 3'b000;

endmodule