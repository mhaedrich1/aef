module dtc_split875_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node443;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node870;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node896;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node909;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1057;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1152;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1159;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1200;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1277;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1302;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1311;
	wire [3-1:0] node1314;
	wire [3-1:0] node1315;
	wire [3-1:0] node1318;
	wire [3-1:0] node1321;
	wire [3-1:0] node1323;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1356;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1388;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1393;
	wire [3-1:0] node1396;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1417;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1425;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1444;
	wire [3-1:0] node1446;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1457;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1462;
	wire [3-1:0] node1464;
	wire [3-1:0] node1467;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1474;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1481;
	wire [3-1:0] node1483;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1494;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1501;
	wire [3-1:0] node1504;
	wire [3-1:0] node1507;
	wire [3-1:0] node1508;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1516;
	wire [3-1:0] node1518;
	wire [3-1:0] node1521;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1530;
	wire [3-1:0] node1532;
	wire [3-1:0] node1535;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1539;
	wire [3-1:0] node1542;
	wire [3-1:0] node1544;
	wire [3-1:0] node1547;
	wire [3-1:0] node1548;
	wire [3-1:0] node1551;
	wire [3-1:0] node1553;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1559;
	wire [3-1:0] node1561;
	wire [3-1:0] node1564;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1572;
	wire [3-1:0] node1575;
	wire [3-1:0] node1577;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1585;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1593;
	wire [3-1:0] node1596;
	wire [3-1:0] node1597;
	wire [3-1:0] node1600;
	wire [3-1:0] node1603;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1614;
	wire [3-1:0] node1615;
	wire [3-1:0] node1618;
	wire [3-1:0] node1621;
	wire [3-1:0] node1622;
	wire [3-1:0] node1623;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1639;
	wire [3-1:0] node1642;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1649;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1656;
	wire [3-1:0] node1659;
	wire [3-1:0] node1660;
	wire [3-1:0] node1661;
	wire [3-1:0] node1664;
	wire [3-1:0] node1667;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1677;
	wire [3-1:0] node1680;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1687;
	wire [3-1:0] node1690;
	wire [3-1:0] node1692;
	wire [3-1:0] node1694;
	wire [3-1:0] node1697;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1704;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1709;
	wire [3-1:0] node1712;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1719;
	wire [3-1:0] node1722;
	wire [3-1:0] node1723;
	wire [3-1:0] node1725;
	wire [3-1:0] node1726;
	wire [3-1:0] node1729;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1736;
	wire [3-1:0] node1739;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1742;
	wire [3-1:0] node1743;
	wire [3-1:0] node1746;
	wire [3-1:0] node1749;
	wire [3-1:0] node1751;
	wire [3-1:0] node1754;
	wire [3-1:0] node1755;
	wire [3-1:0] node1758;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1765;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1773;
	wire [3-1:0] node1776;
	wire [3-1:0] node1777;
	wire [3-1:0] node1778;
	wire [3-1:0] node1779;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1785;
	wire [3-1:0] node1788;
	wire [3-1:0] node1789;
	wire [3-1:0] node1790;
	wire [3-1:0] node1793;
	wire [3-1:0] node1796;
	wire [3-1:0] node1797;
	wire [3-1:0] node1800;
	wire [3-1:0] node1803;
	wire [3-1:0] node1804;
	wire [3-1:0] node1805;
	wire [3-1:0] node1808;
	wire [3-1:0] node1811;
	wire [3-1:0] node1812;
	wire [3-1:0] node1813;
	wire [3-1:0] node1816;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1828;
	wire [3-1:0] node1829;
	wire [3-1:0] node1833;
	wire [3-1:0] node1834;
	wire [3-1:0] node1835;
	wire [3-1:0] node1839;
	wire [3-1:0] node1840;
	wire [3-1:0] node1843;
	wire [3-1:0] node1846;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1852;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1865;
	wire [3-1:0] node1868;
	wire [3-1:0] node1869;
	wire [3-1:0] node1873;
	wire [3-1:0] node1874;
	wire [3-1:0] node1875;
	wire [3-1:0] node1876;
	wire [3-1:0] node1877;
	wire [3-1:0] node1878;
	wire [3-1:0] node1881;
	wire [3-1:0] node1884;
	wire [3-1:0] node1886;
	wire [3-1:0] node1889;
	wire [3-1:0] node1890;
	wire [3-1:0] node1891;
	wire [3-1:0] node1894;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1902;
	wire [3-1:0] node1903;
	wire [3-1:0] node1904;
	wire [3-1:0] node1905;
	wire [3-1:0] node1908;
	wire [3-1:0] node1911;
	wire [3-1:0] node1912;
	wire [3-1:0] node1915;
	wire [3-1:0] node1918;
	wire [3-1:0] node1919;
	wire [3-1:0] node1922;
	wire [3-1:0] node1925;
	wire [3-1:0] node1926;
	wire [3-1:0] node1927;
	wire [3-1:0] node1929;
	wire [3-1:0] node1930;
	wire [3-1:0] node1934;
	wire [3-1:0] node1935;
	wire [3-1:0] node1936;
	wire [3-1:0] node1940;
	wire [3-1:0] node1943;
	wire [3-1:0] node1944;
	wire [3-1:0] node1945;
	wire [3-1:0] node1946;
	wire [3-1:0] node1950;
	wire [3-1:0] node1953;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1959;
	wire [3-1:0] node1960;
	wire [3-1:0] node1964;
	wire [3-1:0] node1965;
	wire [3-1:0] node1966;
	wire [3-1:0] node1967;
	wire [3-1:0] node1968;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1974;
	wire [3-1:0] node1975;
	wire [3-1:0] node1979;
	wire [3-1:0] node1980;
	wire [3-1:0] node1981;
	wire [3-1:0] node1985;
	wire [3-1:0] node1986;
	wire [3-1:0] node1990;
	wire [3-1:0] node1991;
	wire [3-1:0] node1992;
	wire [3-1:0] node1995;
	wire [3-1:0] node1996;
	wire [3-1:0] node2000;
	wire [3-1:0] node2001;
	wire [3-1:0] node2002;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2011;
	wire [3-1:0] node2012;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2016;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2023;
	wire [3-1:0] node2026;
	wire [3-1:0] node2027;
	wire [3-1:0] node2030;
	wire [3-1:0] node2033;
	wire [3-1:0] node2034;
	wire [3-1:0] node2035;
	wire [3-1:0] node2036;
	wire [3-1:0] node2040;
	wire [3-1:0] node2041;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2050;
	wire [3-1:0] node2051;
	wire [3-1:0] node2052;
	wire [3-1:0] node2053;
	wire [3-1:0] node2054;
	wire [3-1:0] node2055;
	wire [3-1:0] node2058;
	wire [3-1:0] node2062;
	wire [3-1:0] node2063;
	wire [3-1:0] node2066;
	wire [3-1:0] node2069;
	wire [3-1:0] node2070;
	wire [3-1:0] node2071;
	wire [3-1:0] node2072;
	wire [3-1:0] node2076;
	wire [3-1:0] node2077;
	wire [3-1:0] node2080;
	wire [3-1:0] node2083;
	wire [3-1:0] node2084;
	wire [3-1:0] node2085;
	wire [3-1:0] node2088;
	wire [3-1:0] node2091;
	wire [3-1:0] node2092;
	wire [3-1:0] node2095;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2100;
	wire [3-1:0] node2101;
	wire [3-1:0] node2102;
	wire [3-1:0] node2105;
	wire [3-1:0] node2108;
	wire [3-1:0] node2109;
	wire [3-1:0] node2112;
	wire [3-1:0] node2115;
	wire [3-1:0] node2116;
	wire [3-1:0] node2119;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2125;
	wire [3-1:0] node2128;
	wire [3-1:0] node2129;
	wire [3-1:0] node2132;
	wire [3-1:0] node2133;
	wire [3-1:0] node2137;
	wire [3-1:0] node2138;
	wire [3-1:0] node2139;
	wire [3-1:0] node2140;
	wire [3-1:0] node2141;
	wire [3-1:0] node2142;
	wire [3-1:0] node2143;
	wire [3-1:0] node2144;
	wire [3-1:0] node2146;
	wire [3-1:0] node2149;
	wire [3-1:0] node2150;
	wire [3-1:0] node2153;
	wire [3-1:0] node2156;
	wire [3-1:0] node2157;
	wire [3-1:0] node2158;
	wire [3-1:0] node2161;
	wire [3-1:0] node2164;
	wire [3-1:0] node2166;
	wire [3-1:0] node2169;
	wire [3-1:0] node2170;
	wire [3-1:0] node2171;
	wire [3-1:0] node2172;
	wire [3-1:0] node2175;
	wire [3-1:0] node2178;
	wire [3-1:0] node2180;
	wire [3-1:0] node2183;
	wire [3-1:0] node2184;
	wire [3-1:0] node2185;
	wire [3-1:0] node2188;
	wire [3-1:0] node2191;
	wire [3-1:0] node2193;
	wire [3-1:0] node2196;
	wire [3-1:0] node2197;
	wire [3-1:0] node2198;
	wire [3-1:0] node2199;
	wire [3-1:0] node2201;
	wire [3-1:0] node2204;
	wire [3-1:0] node2206;
	wire [3-1:0] node2209;
	wire [3-1:0] node2210;
	wire [3-1:0] node2211;
	wire [3-1:0] node2214;
	wire [3-1:0] node2217;
	wire [3-1:0] node2218;
	wire [3-1:0] node2221;
	wire [3-1:0] node2224;
	wire [3-1:0] node2225;
	wire [3-1:0] node2226;
	wire [3-1:0] node2227;
	wire [3-1:0] node2230;
	wire [3-1:0] node2233;
	wire [3-1:0] node2234;
	wire [3-1:0] node2237;
	wire [3-1:0] node2240;
	wire [3-1:0] node2241;
	wire [3-1:0] node2242;
	wire [3-1:0] node2245;
	wire [3-1:0] node2248;
	wire [3-1:0] node2250;
	wire [3-1:0] node2253;
	wire [3-1:0] node2254;
	wire [3-1:0] node2255;
	wire [3-1:0] node2256;
	wire [3-1:0] node2257;
	wire [3-1:0] node2258;
	wire [3-1:0] node2261;
	wire [3-1:0] node2265;
	wire [3-1:0] node2266;
	wire [3-1:0] node2268;
	wire [3-1:0] node2271;
	wire [3-1:0] node2272;
	wire [3-1:0] node2275;
	wire [3-1:0] node2278;
	wire [3-1:0] node2279;
	wire [3-1:0] node2280;
	wire [3-1:0] node2281;
	wire [3-1:0] node2284;
	wire [3-1:0] node2287;
	wire [3-1:0] node2289;
	wire [3-1:0] node2292;
	wire [3-1:0] node2293;
	wire [3-1:0] node2294;
	wire [3-1:0] node2297;
	wire [3-1:0] node2300;
	wire [3-1:0] node2301;
	wire [3-1:0] node2304;
	wire [3-1:0] node2307;
	wire [3-1:0] node2308;
	wire [3-1:0] node2309;
	wire [3-1:0] node2310;
	wire [3-1:0] node2311;
	wire [3-1:0] node2314;
	wire [3-1:0] node2317;
	wire [3-1:0] node2318;
	wire [3-1:0] node2321;
	wire [3-1:0] node2324;
	wire [3-1:0] node2325;
	wire [3-1:0] node2326;
	wire [3-1:0] node2329;
	wire [3-1:0] node2332;
	wire [3-1:0] node2333;
	wire [3-1:0] node2336;
	wire [3-1:0] node2339;
	wire [3-1:0] node2340;
	wire [3-1:0] node2341;
	wire [3-1:0] node2342;
	wire [3-1:0] node2345;
	wire [3-1:0] node2348;
	wire [3-1:0] node2350;
	wire [3-1:0] node2353;
	wire [3-1:0] node2354;
	wire [3-1:0] node2355;
	wire [3-1:0] node2358;
	wire [3-1:0] node2361;
	wire [3-1:0] node2362;
	wire [3-1:0] node2365;
	wire [3-1:0] node2368;
	wire [3-1:0] node2369;
	wire [3-1:0] node2370;
	wire [3-1:0] node2371;
	wire [3-1:0] node2372;
	wire [3-1:0] node2373;
	wire [3-1:0] node2375;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2382;
	wire [3-1:0] node2385;
	wire [3-1:0] node2386;
	wire [3-1:0] node2387;
	wire [3-1:0] node2391;
	wire [3-1:0] node2392;
	wire [3-1:0] node2395;
	wire [3-1:0] node2398;
	wire [3-1:0] node2399;
	wire [3-1:0] node2400;
	wire [3-1:0] node2401;
	wire [3-1:0] node2404;
	wire [3-1:0] node2407;
	wire [3-1:0] node2408;
	wire [3-1:0] node2411;
	wire [3-1:0] node2414;
	wire [3-1:0] node2415;
	wire [3-1:0] node2416;
	wire [3-1:0] node2419;
	wire [3-1:0] node2422;
	wire [3-1:0] node2424;
	wire [3-1:0] node2427;
	wire [3-1:0] node2428;
	wire [3-1:0] node2429;
	wire [3-1:0] node2430;
	wire [3-1:0] node2431;
	wire [3-1:0] node2434;
	wire [3-1:0] node2437;
	wire [3-1:0] node2439;
	wire [3-1:0] node2442;
	wire [3-1:0] node2443;
	wire [3-1:0] node2444;
	wire [3-1:0] node2447;
	wire [3-1:0] node2450;
	wire [3-1:0] node2451;
	wire [3-1:0] node2454;
	wire [3-1:0] node2457;
	wire [3-1:0] node2458;
	wire [3-1:0] node2459;
	wire [3-1:0] node2460;
	wire [3-1:0] node2463;
	wire [3-1:0] node2466;
	wire [3-1:0] node2467;
	wire [3-1:0] node2470;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2476;
	wire [3-1:0] node2479;
	wire [3-1:0] node2480;
	wire [3-1:0] node2483;
	wire [3-1:0] node2486;
	wire [3-1:0] node2487;
	wire [3-1:0] node2488;
	wire [3-1:0] node2489;
	wire [3-1:0] node2490;
	wire [3-1:0] node2491;
	wire [3-1:0] node2494;
	wire [3-1:0] node2497;
	wire [3-1:0] node2498;
	wire [3-1:0] node2501;
	wire [3-1:0] node2504;
	wire [3-1:0] node2505;
	wire [3-1:0] node2506;
	wire [3-1:0] node2509;
	wire [3-1:0] node2512;
	wire [3-1:0] node2513;
	wire [3-1:0] node2516;
	wire [3-1:0] node2519;
	wire [3-1:0] node2520;
	wire [3-1:0] node2521;
	wire [3-1:0] node2522;
	wire [3-1:0] node2525;
	wire [3-1:0] node2528;
	wire [3-1:0] node2529;
	wire [3-1:0] node2532;
	wire [3-1:0] node2535;
	wire [3-1:0] node2536;
	wire [3-1:0] node2537;
	wire [3-1:0] node2540;
	wire [3-1:0] node2543;
	wire [3-1:0] node2545;
	wire [3-1:0] node2548;
	wire [3-1:0] node2549;
	wire [3-1:0] node2550;
	wire [3-1:0] node2551;
	wire [3-1:0] node2553;
	wire [3-1:0] node2556;
	wire [3-1:0] node2557;
	wire [3-1:0] node2560;
	wire [3-1:0] node2563;
	wire [3-1:0] node2564;
	wire [3-1:0] node2565;
	wire [3-1:0] node2568;
	wire [3-1:0] node2571;
	wire [3-1:0] node2572;
	wire [3-1:0] node2575;
	wire [3-1:0] node2578;
	wire [3-1:0] node2579;
	wire [3-1:0] node2580;
	wire [3-1:0] node2583;
	wire [3-1:0] node2586;
	wire [3-1:0] node2587;
	wire [3-1:0] node2588;
	wire [3-1:0] node2591;
	wire [3-1:0] node2594;
	wire [3-1:0] node2596;
	wire [3-1:0] node2599;
	wire [3-1:0] node2600;
	wire [3-1:0] node2601;
	wire [3-1:0] node2602;
	wire [3-1:0] node2603;
	wire [3-1:0] node2604;
	wire [3-1:0] node2605;
	wire [3-1:0] node2606;
	wire [3-1:0] node2609;
	wire [3-1:0] node2612;
	wire [3-1:0] node2615;
	wire [3-1:0] node2616;
	wire [3-1:0] node2617;
	wire [3-1:0] node2620;
	wire [3-1:0] node2623;
	wire [3-1:0] node2625;
	wire [3-1:0] node2628;
	wire [3-1:0] node2629;
	wire [3-1:0] node2630;
	wire [3-1:0] node2631;
	wire [3-1:0] node2634;
	wire [3-1:0] node2637;
	wire [3-1:0] node2639;
	wire [3-1:0] node2642;
	wire [3-1:0] node2643;
	wire [3-1:0] node2644;
	wire [3-1:0] node2647;
	wire [3-1:0] node2650;
	wire [3-1:0] node2652;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2657;
	wire [3-1:0] node2658;
	wire [3-1:0] node2659;
	wire [3-1:0] node2663;
	wire [3-1:0] node2664;
	wire [3-1:0] node2668;
	wire [3-1:0] node2669;
	wire [3-1:0] node2671;
	wire [3-1:0] node2674;
	wire [3-1:0] node2676;
	wire [3-1:0] node2679;
	wire [3-1:0] node2680;
	wire [3-1:0] node2681;
	wire [3-1:0] node2682;
	wire [3-1:0] node2685;
	wire [3-1:0] node2688;
	wire [3-1:0] node2689;
	wire [3-1:0] node2692;
	wire [3-1:0] node2695;
	wire [3-1:0] node2697;
	wire [3-1:0] node2698;
	wire [3-1:0] node2701;
	wire [3-1:0] node2704;
	wire [3-1:0] node2705;
	wire [3-1:0] node2706;
	wire [3-1:0] node2707;
	wire [3-1:0] node2708;
	wire [3-1:0] node2709;
	wire [3-1:0] node2712;
	wire [3-1:0] node2715;
	wire [3-1:0] node2716;
	wire [3-1:0] node2719;
	wire [3-1:0] node2722;
	wire [3-1:0] node2723;
	wire [3-1:0] node2724;
	wire [3-1:0] node2728;
	wire [3-1:0] node2729;
	wire [3-1:0] node2732;
	wire [3-1:0] node2735;
	wire [3-1:0] node2736;
	wire [3-1:0] node2737;
	wire [3-1:0] node2738;
	wire [3-1:0] node2743;
	wire [3-1:0] node2744;
	wire [3-1:0] node2745;
	wire [3-1:0] node2748;
	wire [3-1:0] node2751;
	wire [3-1:0] node2752;
	wire [3-1:0] node2756;
	wire [3-1:0] node2757;
	wire [3-1:0] node2758;
	wire [3-1:0] node2759;
	wire [3-1:0] node2760;
	wire [3-1:0] node2763;
	wire [3-1:0] node2766;
	wire [3-1:0] node2767;
	wire [3-1:0] node2770;
	wire [3-1:0] node2773;
	wire [3-1:0] node2774;
	wire [3-1:0] node2775;
	wire [3-1:0] node2778;
	wire [3-1:0] node2781;
	wire [3-1:0] node2783;
	wire [3-1:0] node2786;
	wire [3-1:0] node2787;
	wire [3-1:0] node2788;
	wire [3-1:0] node2791;
	wire [3-1:0] node2794;
	wire [3-1:0] node2795;
	wire [3-1:0] node2798;
	wire [3-1:0] node2801;
	wire [3-1:0] node2802;
	wire [3-1:0] node2803;
	wire [3-1:0] node2804;
	wire [3-1:0] node2805;
	wire [3-1:0] node2806;
	wire [3-1:0] node2808;
	wire [3-1:0] node2811;
	wire [3-1:0] node2812;
	wire [3-1:0] node2815;
	wire [3-1:0] node2818;
	wire [3-1:0] node2819;
	wire [3-1:0] node2820;
	wire [3-1:0] node2823;
	wire [3-1:0] node2826;
	wire [3-1:0] node2827;
	wire [3-1:0] node2830;
	wire [3-1:0] node2833;
	wire [3-1:0] node2834;
	wire [3-1:0] node2835;
	wire [3-1:0] node2836;
	wire [3-1:0] node2839;
	wire [3-1:0] node2842;
	wire [3-1:0] node2843;
	wire [3-1:0] node2846;
	wire [3-1:0] node2849;
	wire [3-1:0] node2850;
	wire [3-1:0] node2851;
	wire [3-1:0] node2854;
	wire [3-1:0] node2857;
	wire [3-1:0] node2858;
	wire [3-1:0] node2861;
	wire [3-1:0] node2864;
	wire [3-1:0] node2865;
	wire [3-1:0] node2866;
	wire [3-1:0] node2867;
	wire [3-1:0] node2868;
	wire [3-1:0] node2871;
	wire [3-1:0] node2874;
	wire [3-1:0] node2875;
	wire [3-1:0] node2878;
	wire [3-1:0] node2881;
	wire [3-1:0] node2882;
	wire [3-1:0] node2883;
	wire [3-1:0] node2886;
	wire [3-1:0] node2889;
	wire [3-1:0] node2890;
	wire [3-1:0] node2894;
	wire [3-1:0] node2895;
	wire [3-1:0] node2896;
	wire [3-1:0] node2897;
	wire [3-1:0] node2900;
	wire [3-1:0] node2903;
	wire [3-1:0] node2904;
	wire [3-1:0] node2907;
	wire [3-1:0] node2910;
	wire [3-1:0] node2911;
	wire [3-1:0] node2914;
	wire [3-1:0] node2917;
	wire [3-1:0] node2918;
	wire [3-1:0] node2919;
	wire [3-1:0] node2920;
	wire [3-1:0] node2921;
	wire [3-1:0] node2922;
	wire [3-1:0] node2925;
	wire [3-1:0] node2928;
	wire [3-1:0] node2929;
	wire [3-1:0] node2932;
	wire [3-1:0] node2935;
	wire [3-1:0] node2936;
	wire [3-1:0] node2937;
	wire [3-1:0] node2940;
	wire [3-1:0] node2944;
	wire [3-1:0] node2945;
	wire [3-1:0] node2946;
	wire [3-1:0] node2947;
	wire [3-1:0] node2950;
	wire [3-1:0] node2953;
	wire [3-1:0] node2955;
	wire [3-1:0] node2958;
	wire [3-1:0] node2959;
	wire [3-1:0] node2961;
	wire [3-1:0] node2964;
	wire [3-1:0] node2966;
	wire [3-1:0] node2969;
	wire [3-1:0] node2970;
	wire [3-1:0] node2971;
	wire [3-1:0] node2972;
	wire [3-1:0] node2973;
	wire [3-1:0] node2976;
	wire [3-1:0] node2980;
	wire [3-1:0] node2981;
	wire [3-1:0] node2982;
	wire [3-1:0] node2986;
	wire [3-1:0] node2988;
	wire [3-1:0] node2991;
	wire [3-1:0] node2992;
	wire [3-1:0] node2993;
	wire [3-1:0] node2994;
	wire [3-1:0] node2997;
	wire [3-1:0] node3000;
	wire [3-1:0] node3001;
	wire [3-1:0] node3004;
	wire [3-1:0] node3007;
	wire [3-1:0] node3008;
	wire [3-1:0] node3009;
	wire [3-1:0] node3012;
	wire [3-1:0] node3015;
	wire [3-1:0] node3017;
	wire [3-1:0] node3020;
	wire [3-1:0] node3021;
	wire [3-1:0] node3022;
	wire [3-1:0] node3023;
	wire [3-1:0] node3024;
	wire [3-1:0] node3025;
	wire [3-1:0] node3026;
	wire [3-1:0] node3027;
	wire [3-1:0] node3028;
	wire [3-1:0] node3031;
	wire [3-1:0] node3034;
	wire [3-1:0] node3035;
	wire [3-1:0] node3036;
	wire [3-1:0] node3039;
	wire [3-1:0] node3042;
	wire [3-1:0] node3044;
	wire [3-1:0] node3045;
	wire [3-1:0] node3048;
	wire [3-1:0] node3051;
	wire [3-1:0] node3052;
	wire [3-1:0] node3053;
	wire [3-1:0] node3056;
	wire [3-1:0] node3059;
	wire [3-1:0] node3060;
	wire [3-1:0] node3061;
	wire [3-1:0] node3064;
	wire [3-1:0] node3067;
	wire [3-1:0] node3068;
	wire [3-1:0] node3071;
	wire [3-1:0] node3074;
	wire [3-1:0] node3075;
	wire [3-1:0] node3076;
	wire [3-1:0] node3077;
	wire [3-1:0] node3080;
	wire [3-1:0] node3083;
	wire [3-1:0] node3084;
	wire [3-1:0] node3086;
	wire [3-1:0] node3087;
	wire [3-1:0] node3090;
	wire [3-1:0] node3093;
	wire [3-1:0] node3094;
	wire [3-1:0] node3097;
	wire [3-1:0] node3099;
	wire [3-1:0] node3102;
	wire [3-1:0] node3103;
	wire [3-1:0] node3104;
	wire [3-1:0] node3107;
	wire [3-1:0] node3110;
	wire [3-1:0] node3111;
	wire [3-1:0] node3112;
	wire [3-1:0] node3115;
	wire [3-1:0] node3118;
	wire [3-1:0] node3119;
	wire [3-1:0] node3120;
	wire [3-1:0] node3123;
	wire [3-1:0] node3126;
	wire [3-1:0] node3127;
	wire [3-1:0] node3130;
	wire [3-1:0] node3133;
	wire [3-1:0] node3134;
	wire [3-1:0] node3135;
	wire [3-1:0] node3136;
	wire [3-1:0] node3137;
	wire [3-1:0] node3138;
	wire [3-1:0] node3139;
	wire [3-1:0] node3142;
	wire [3-1:0] node3146;
	wire [3-1:0] node3147;
	wire [3-1:0] node3149;
	wire [3-1:0] node3152;
	wire [3-1:0] node3153;
	wire [3-1:0] node3156;
	wire [3-1:0] node3159;
	wire [3-1:0] node3160;
	wire [3-1:0] node3161;
	wire [3-1:0] node3164;
	wire [3-1:0] node3167;
	wire [3-1:0] node3168;
	wire [3-1:0] node3169;
	wire [3-1:0] node3172;
	wire [3-1:0] node3175;
	wire [3-1:0] node3176;
	wire [3-1:0] node3179;
	wire [3-1:0] node3182;
	wire [3-1:0] node3183;
	wire [3-1:0] node3184;
	wire [3-1:0] node3185;
	wire [3-1:0] node3188;
	wire [3-1:0] node3191;
	wire [3-1:0] node3192;
	wire [3-1:0] node3193;
	wire [3-1:0] node3197;
	wire [3-1:0] node3198;
	wire [3-1:0] node3201;
	wire [3-1:0] node3204;
	wire [3-1:0] node3205;
	wire [3-1:0] node3206;
	wire [3-1:0] node3207;
	wire [3-1:0] node3210;
	wire [3-1:0] node3213;
	wire [3-1:0] node3214;
	wire [3-1:0] node3218;
	wire [3-1:0] node3219;
	wire [3-1:0] node3222;
	wire [3-1:0] node3225;
	wire [3-1:0] node3226;
	wire [3-1:0] node3227;
	wire [3-1:0] node3228;
	wire [3-1:0] node3231;
	wire [3-1:0] node3234;
	wire [3-1:0] node3235;
	wire [3-1:0] node3236;
	wire [3-1:0] node3239;
	wire [3-1:0] node3242;
	wire [3-1:0] node3243;
	wire [3-1:0] node3246;
	wire [3-1:0] node3249;
	wire [3-1:0] node3250;
	wire [3-1:0] node3251;
	wire [3-1:0] node3254;
	wire [3-1:0] node3257;
	wire [3-1:0] node3258;
	wire [3-1:0] node3260;
	wire [3-1:0] node3261;
	wire [3-1:0] node3264;
	wire [3-1:0] node3267;
	wire [3-1:0] node3268;
	wire [3-1:0] node3271;
	wire [3-1:0] node3274;
	wire [3-1:0] node3275;
	wire [3-1:0] node3276;
	wire [3-1:0] node3277;
	wire [3-1:0] node3278;
	wire [3-1:0] node3279;
	wire [3-1:0] node3282;
	wire [3-1:0] node3285;
	wire [3-1:0] node3286;
	wire [3-1:0] node3287;
	wire [3-1:0] node3290;
	wire [3-1:0] node3293;
	wire [3-1:0] node3294;
	wire [3-1:0] node3297;
	wire [3-1:0] node3300;
	wire [3-1:0] node3301;
	wire [3-1:0] node3302;
	wire [3-1:0] node3304;
	wire [3-1:0] node3307;
	wire [3-1:0] node3310;
	wire [3-1:0] node3311;
	wire [3-1:0] node3313;
	wire [3-1:0] node3316;
	wire [3-1:0] node3318;
	wire [3-1:0] node3321;
	wire [3-1:0] node3322;
	wire [3-1:0] node3323;
	wire [3-1:0] node3324;
	wire [3-1:0] node3326;
	wire [3-1:0] node3329;
	wire [3-1:0] node3331;
	wire [3-1:0] node3334;
	wire [3-1:0] node3335;
	wire [3-1:0] node3337;
	wire [3-1:0] node3340;
	wire [3-1:0] node3342;
	wire [3-1:0] node3345;
	wire [3-1:0] node3346;
	wire [3-1:0] node3347;
	wire [3-1:0] node3348;
	wire [3-1:0] node3351;
	wire [3-1:0] node3354;
	wire [3-1:0] node3355;
	wire [3-1:0] node3357;
	wire [3-1:0] node3360;
	wire [3-1:0] node3362;
	wire [3-1:0] node3365;
	wire [3-1:0] node3366;
	wire [3-1:0] node3368;
	wire [3-1:0] node3371;
	wire [3-1:0] node3372;
	wire [3-1:0] node3375;
	wire [3-1:0] node3378;
	wire [3-1:0] node3379;
	wire [3-1:0] node3380;
	wire [3-1:0] node3381;
	wire [3-1:0] node3382;
	wire [3-1:0] node3384;
	wire [3-1:0] node3387;
	wire [3-1:0] node3389;
	wire [3-1:0] node3392;
	wire [3-1:0] node3393;
	wire [3-1:0] node3395;
	wire [3-1:0] node3398;
	wire [3-1:0] node3400;
	wire [3-1:0] node3403;
	wire [3-1:0] node3404;
	wire [3-1:0] node3405;
	wire [3-1:0] node3406;
	wire [3-1:0] node3410;
	wire [3-1:0] node3411;
	wire [3-1:0] node3415;
	wire [3-1:0] node3416;
	wire [3-1:0] node3417;
	wire [3-1:0] node3421;
	wire [3-1:0] node3422;
	wire [3-1:0] node3426;
	wire [3-1:0] node3427;
	wire [3-1:0] node3428;
	wire [3-1:0] node3429;
	wire [3-1:0] node3430;
	wire [3-1:0] node3434;
	wire [3-1:0] node3435;
	wire [3-1:0] node3439;
	wire [3-1:0] node3440;
	wire [3-1:0] node3441;
	wire [3-1:0] node3445;
	wire [3-1:0] node3446;
	wire [3-1:0] node3450;
	wire [3-1:0] node3451;
	wire [3-1:0] node3452;
	wire [3-1:0] node3453;
	wire [3-1:0] node3456;
	wire [3-1:0] node3459;
	wire [3-1:0] node3460;
	wire [3-1:0] node3461;
	wire [3-1:0] node3464;
	wire [3-1:0] node3467;
	wire [3-1:0] node3468;
	wire [3-1:0] node3471;
	wire [3-1:0] node3474;
	wire [3-1:0] node3475;
	wire [3-1:0] node3478;
	wire [3-1:0] node3481;
	wire [3-1:0] node3482;
	wire [3-1:0] node3483;
	wire [3-1:0] node3484;
	wire [3-1:0] node3485;
	wire [3-1:0] node3486;
	wire [3-1:0] node3487;
	wire [3-1:0] node3488;
	wire [3-1:0] node3491;
	wire [3-1:0] node3494;
	wire [3-1:0] node3495;
	wire [3-1:0] node3496;
	wire [3-1:0] node3500;
	wire [3-1:0] node3501;
	wire [3-1:0] node3504;
	wire [3-1:0] node3507;
	wire [3-1:0] node3508;
	wire [3-1:0] node3509;
	wire [3-1:0] node3512;
	wire [3-1:0] node3515;
	wire [3-1:0] node3516;
	wire [3-1:0] node3519;
	wire [3-1:0] node3522;
	wire [3-1:0] node3523;
	wire [3-1:0] node3524;
	wire [3-1:0] node3525;
	wire [3-1:0] node3527;
	wire [3-1:0] node3530;
	wire [3-1:0] node3533;
	wire [3-1:0] node3534;
	wire [3-1:0] node3536;
	wire [3-1:0] node3539;
	wire [3-1:0] node3542;
	wire [3-1:0] node3543;
	wire [3-1:0] node3545;
	wire [3-1:0] node3547;
	wire [3-1:0] node3550;
	wire [3-1:0] node3551;
	wire [3-1:0] node3553;
	wire [3-1:0] node3556;
	wire [3-1:0] node3558;
	wire [3-1:0] node3561;
	wire [3-1:0] node3562;
	wire [3-1:0] node3563;
	wire [3-1:0] node3564;
	wire [3-1:0] node3567;
	wire [3-1:0] node3570;
	wire [3-1:0] node3571;
	wire [3-1:0] node3572;
	wire [3-1:0] node3575;
	wire [3-1:0] node3578;
	wire [3-1:0] node3579;
	wire [3-1:0] node3580;
	wire [3-1:0] node3584;
	wire [3-1:0] node3585;
	wire [3-1:0] node3588;
	wire [3-1:0] node3591;
	wire [3-1:0] node3592;
	wire [3-1:0] node3593;
	wire [3-1:0] node3596;
	wire [3-1:0] node3599;
	wire [3-1:0] node3600;
	wire [3-1:0] node3601;
	wire [3-1:0] node3604;
	wire [3-1:0] node3607;
	wire [3-1:0] node3608;
	wire [3-1:0] node3611;
	wire [3-1:0] node3614;
	wire [3-1:0] node3615;
	wire [3-1:0] node3616;
	wire [3-1:0] node3617;
	wire [3-1:0] node3618;
	wire [3-1:0] node3621;
	wire [3-1:0] node3624;
	wire [3-1:0] node3625;
	wire [3-1:0] node3626;
	wire [3-1:0] node3627;
	wire [3-1:0] node3630;
	wire [3-1:0] node3633;
	wire [3-1:0] node3634;
	wire [3-1:0] node3637;
	wire [3-1:0] node3640;
	wire [3-1:0] node3641;
	wire [3-1:0] node3642;
	wire [3-1:0] node3645;
	wire [3-1:0] node3648;
	wire [3-1:0] node3649;
	wire [3-1:0] node3652;
	wire [3-1:0] node3655;
	wire [3-1:0] node3656;
	wire [3-1:0] node3657;
	wire [3-1:0] node3658;
	wire [3-1:0] node3662;
	wire [3-1:0] node3663;
	wire [3-1:0] node3667;
	wire [3-1:0] node3668;
	wire [3-1:0] node3669;
	wire [3-1:0] node3673;
	wire [3-1:0] node3674;
	wire [3-1:0] node3678;
	wire [3-1:0] node3679;
	wire [3-1:0] node3680;
	wire [3-1:0] node3681;
	wire [3-1:0] node3682;
	wire [3-1:0] node3683;
	wire [3-1:0] node3686;
	wire [3-1:0] node3689;
	wire [3-1:0] node3690;
	wire [3-1:0] node3693;
	wire [3-1:0] node3696;
	wire [3-1:0] node3697;
	wire [3-1:0] node3698;
	wire [3-1:0] node3701;
	wire [3-1:0] node3704;
	wire [3-1:0] node3705;
	wire [3-1:0] node3709;
	wire [3-1:0] node3710;
	wire [3-1:0] node3711;
	wire [3-1:0] node3714;
	wire [3-1:0] node3717;
	wire [3-1:0] node3718;
	wire [3-1:0] node3719;
	wire [3-1:0] node3722;
	wire [3-1:0] node3725;
	wire [3-1:0] node3726;
	wire [3-1:0] node3729;
	wire [3-1:0] node3732;
	wire [3-1:0] node3733;
	wire [3-1:0] node3734;
	wire [3-1:0] node3735;
	wire [3-1:0] node3736;
	wire [3-1:0] node3739;
	wire [3-1:0] node3742;
	wire [3-1:0] node3743;
	wire [3-1:0] node3746;
	wire [3-1:0] node3749;
	wire [3-1:0] node3750;
	wire [3-1:0] node3751;
	wire [3-1:0] node3754;
	wire [3-1:0] node3758;
	wire [3-1:0] node3759;
	wire [3-1:0] node3762;
	wire [3-1:0] node3765;
	wire [3-1:0] node3766;
	wire [3-1:0] node3767;
	wire [3-1:0] node3768;
	wire [3-1:0] node3769;
	wire [3-1:0] node3770;
	wire [3-1:0] node3771;
	wire [3-1:0] node3774;
	wire [3-1:0] node3777;
	wire [3-1:0] node3779;
	wire [3-1:0] node3782;
	wire [3-1:0] node3783;
	wire [3-1:0] node3784;
	wire [3-1:0] node3785;
	wire [3-1:0] node3788;
	wire [3-1:0] node3792;
	wire [3-1:0] node3793;
	wire [3-1:0] node3796;
	wire [3-1:0] node3799;
	wire [3-1:0] node3800;
	wire [3-1:0] node3801;
	wire [3-1:0] node3802;
	wire [3-1:0] node3805;
	wire [3-1:0] node3808;
	wire [3-1:0] node3809;
	wire [3-1:0] node3813;
	wire [3-1:0] node3814;
	wire [3-1:0] node3817;
	wire [3-1:0] node3820;
	wire [3-1:0] node3821;
	wire [3-1:0] node3822;
	wire [3-1:0] node3823;
	wire [3-1:0] node3824;
	wire [3-1:0] node3828;
	wire [3-1:0] node3829;
	wire [3-1:0] node3830;
	wire [3-1:0] node3833;
	wire [3-1:0] node3837;
	wire [3-1:0] node3838;
	wire [3-1:0] node3839;
	wire [3-1:0] node3842;
	wire [3-1:0] node3845;
	wire [3-1:0] node3846;
	wire [3-1:0] node3849;
	wire [3-1:0] node3852;
	wire [3-1:0] node3853;
	wire [3-1:0] node3854;
	wire [3-1:0] node3855;
	wire [3-1:0] node3858;
	wire [3-1:0] node3861;
	wire [3-1:0] node3862;
	wire [3-1:0] node3863;
	wire [3-1:0] node3866;
	wire [3-1:0] node3869;
	wire [3-1:0] node3871;
	wire [3-1:0] node3874;
	wire [3-1:0] node3875;
	wire [3-1:0] node3876;
	wire [3-1:0] node3879;
	wire [3-1:0] node3882;
	wire [3-1:0] node3883;
	wire [3-1:0] node3886;
	wire [3-1:0] node3888;
	wire [3-1:0] node3891;
	wire [3-1:0] node3892;
	wire [3-1:0] node3893;
	wire [3-1:0] node3894;
	wire [3-1:0] node3895;
	wire [3-1:0] node3897;
	wire [3-1:0] node3898;
	wire [3-1:0] node3901;
	wire [3-1:0] node3904;
	wire [3-1:0] node3905;
	wire [3-1:0] node3906;
	wire [3-1:0] node3909;
	wire [3-1:0] node3913;
	wire [3-1:0] node3914;
	wire [3-1:0] node3915;
	wire [3-1:0] node3916;
	wire [3-1:0] node3919;
	wire [3-1:0] node3922;
	wire [3-1:0] node3924;
	wire [3-1:0] node3927;
	wire [3-1:0] node3928;
	wire [3-1:0] node3931;
	wire [3-1:0] node3934;
	wire [3-1:0] node3935;
	wire [3-1:0] node3936;
	wire [3-1:0] node3937;
	wire [3-1:0] node3938;
	wire [3-1:0] node3943;
	wire [3-1:0] node3944;
	wire [3-1:0] node3945;
	wire [3-1:0] node3949;
	wire [3-1:0] node3950;
	wire [3-1:0] node3954;
	wire [3-1:0] node3955;
	wire [3-1:0] node3956;
	wire [3-1:0] node3957;
	wire [3-1:0] node3960;
	wire [3-1:0] node3963;
	wire [3-1:0] node3964;
	wire [3-1:0] node3967;
	wire [3-1:0] node3970;
	wire [3-1:0] node3971;
	wire [3-1:0] node3974;
	wire [3-1:0] node3977;
	wire [3-1:0] node3978;
	wire [3-1:0] node3979;
	wire [3-1:0] node3980;
	wire [3-1:0] node3981;
	wire [3-1:0] node3985;
	wire [3-1:0] node3986;
	wire [3-1:0] node3990;
	wire [3-1:0] node3991;
	wire [3-1:0] node3992;
	wire [3-1:0] node3996;
	wire [3-1:0] node3997;
	wire [3-1:0] node4001;
	wire [3-1:0] node4002;
	wire [3-1:0] node4003;
	wire [3-1:0] node4004;
	wire [3-1:0] node4008;
	wire [3-1:0] node4009;
	wire [3-1:0] node4013;
	wire [3-1:0] node4014;
	wire [3-1:0] node4015;
	wire [3-1:0] node4019;
	wire [3-1:0] node4020;
	wire [3-1:0] node4024;
	wire [3-1:0] node4025;
	wire [3-1:0] node4026;
	wire [3-1:0] node4027;
	wire [3-1:0] node4028;
	wire [3-1:0] node4029;
	wire [3-1:0] node4030;
	wire [3-1:0] node4031;
	wire [3-1:0] node4034;
	wire [3-1:0] node4036;
	wire [3-1:0] node4039;
	wire [3-1:0] node4040;
	wire [3-1:0] node4041;
	wire [3-1:0] node4044;
	wire [3-1:0] node4047;
	wire [3-1:0] node4049;
	wire [3-1:0] node4052;
	wire [3-1:0] node4053;
	wire [3-1:0] node4054;
	wire [3-1:0] node4057;
	wire [3-1:0] node4059;
	wire [3-1:0] node4062;
	wire [3-1:0] node4063;
	wire [3-1:0] node4066;
	wire [3-1:0] node4067;
	wire [3-1:0] node4071;
	wire [3-1:0] node4072;
	wire [3-1:0] node4073;
	wire [3-1:0] node4074;
	wire [3-1:0] node4075;
	wire [3-1:0] node4078;
	wire [3-1:0] node4081;
	wire [3-1:0] node4082;
	wire [3-1:0] node4085;
	wire [3-1:0] node4088;
	wire [3-1:0] node4089;
	wire [3-1:0] node4090;
	wire [3-1:0] node4093;
	wire [3-1:0] node4096;
	wire [3-1:0] node4097;
	wire [3-1:0] node4099;
	wire [3-1:0] node4102;
	wire [3-1:0] node4103;
	wire [3-1:0] node4106;
	wire [3-1:0] node4109;
	wire [3-1:0] node4110;
	wire [3-1:0] node4111;
	wire [3-1:0] node4112;
	wire [3-1:0] node4115;
	wire [3-1:0] node4118;
	wire [3-1:0] node4119;
	wire [3-1:0] node4120;
	wire [3-1:0] node4123;
	wire [3-1:0] node4126;
	wire [3-1:0] node4127;
	wire [3-1:0] node4130;
	wire [3-1:0] node4133;
	wire [3-1:0] node4134;
	wire [3-1:0] node4135;
	wire [3-1:0] node4138;
	wire [3-1:0] node4141;
	wire [3-1:0] node4142;
	wire [3-1:0] node4144;
	wire [3-1:0] node4147;
	wire [3-1:0] node4149;
	wire [3-1:0] node4152;
	wire [3-1:0] node4153;
	wire [3-1:0] node4154;
	wire [3-1:0] node4155;
	wire [3-1:0] node4156;
	wire [3-1:0] node4158;
	wire [3-1:0] node4161;
	wire [3-1:0] node4163;
	wire [3-1:0] node4166;
	wire [3-1:0] node4167;
	wire [3-1:0] node4169;
	wire [3-1:0] node4172;
	wire [3-1:0] node4174;
	wire [3-1:0] node4177;
	wire [3-1:0] node4178;
	wire [3-1:0] node4179;
	wire [3-1:0] node4180;
	wire [3-1:0] node4183;
	wire [3-1:0] node4186;
	wire [3-1:0] node4187;
	wire [3-1:0] node4190;
	wire [3-1:0] node4193;
	wire [3-1:0] node4194;
	wire [3-1:0] node4195;
	wire [3-1:0] node4196;
	wire [3-1:0] node4199;
	wire [3-1:0] node4202;
	wire [3-1:0] node4203;
	wire [3-1:0] node4207;
	wire [3-1:0] node4208;
	wire [3-1:0] node4211;
	wire [3-1:0] node4214;
	wire [3-1:0] node4215;
	wire [3-1:0] node4216;
	wire [3-1:0] node4217;
	wire [3-1:0] node4218;
	wire [3-1:0] node4219;
	wire [3-1:0] node4222;
	wire [3-1:0] node4225;
	wire [3-1:0] node4226;
	wire [3-1:0] node4229;
	wire [3-1:0] node4232;
	wire [3-1:0] node4233;
	wire [3-1:0] node4234;
	wire [3-1:0] node4237;
	wire [3-1:0] node4240;
	wire [3-1:0] node4241;
	wire [3-1:0] node4244;
	wire [3-1:0] node4247;
	wire [3-1:0] node4248;
	wire [3-1:0] node4249;
	wire [3-1:0] node4252;
	wire [3-1:0] node4255;
	wire [3-1:0] node4256;
	wire [3-1:0] node4257;
	wire [3-1:0] node4260;
	wire [3-1:0] node4263;
	wire [3-1:0] node4264;
	wire [3-1:0] node4268;
	wire [3-1:0] node4269;
	wire [3-1:0] node4270;
	wire [3-1:0] node4271;
	wire [3-1:0] node4274;
	wire [3-1:0] node4277;
	wire [3-1:0] node4278;
	wire [3-1:0] node4281;
	wire [3-1:0] node4284;
	wire [3-1:0] node4285;
	wire [3-1:0] node4286;
	wire [3-1:0] node4289;
	wire [3-1:0] node4292;
	wire [3-1:0] node4293;
	wire [3-1:0] node4296;
	wire [3-1:0] node4299;
	wire [3-1:0] node4300;
	wire [3-1:0] node4301;
	wire [3-1:0] node4302;
	wire [3-1:0] node4303;
	wire [3-1:0] node4304;
	wire [3-1:0] node4305;
	wire [3-1:0] node4308;
	wire [3-1:0] node4311;
	wire [3-1:0] node4312;
	wire [3-1:0] node4314;
	wire [3-1:0] node4317;
	wire [3-1:0] node4319;
	wire [3-1:0] node4322;
	wire [3-1:0] node4323;
	wire [3-1:0] node4326;
	wire [3-1:0] node4329;
	wire [3-1:0] node4330;
	wire [3-1:0] node4331;
	wire [3-1:0] node4332;
	wire [3-1:0] node4335;
	wire [3-1:0] node4338;
	wire [3-1:0] node4340;
	wire [3-1:0] node4343;
	wire [3-1:0] node4344;
	wire [3-1:0] node4347;
	wire [3-1:0] node4350;
	wire [3-1:0] node4351;
	wire [3-1:0] node4352;
	wire [3-1:0] node4353;
	wire [3-1:0] node4356;
	wire [3-1:0] node4359;
	wire [3-1:0] node4360;
	wire [3-1:0] node4363;
	wire [3-1:0] node4366;
	wire [3-1:0] node4367;
	wire [3-1:0] node4368;
	wire [3-1:0] node4371;
	wire [3-1:0] node4374;
	wire [3-1:0] node4375;
	wire [3-1:0] node4378;
	wire [3-1:0] node4381;
	wire [3-1:0] node4382;
	wire [3-1:0] node4383;
	wire [3-1:0] node4384;
	wire [3-1:0] node4385;
	wire [3-1:0] node4386;
	wire [3-1:0] node4387;
	wire [3-1:0] node4391;
	wire [3-1:0] node4393;
	wire [3-1:0] node4396;
	wire [3-1:0] node4398;
	wire [3-1:0] node4401;
	wire [3-1:0] node4402;
	wire [3-1:0] node4403;
	wire [3-1:0] node4404;
	wire [3-1:0] node4407;
	wire [3-1:0] node4410;
	wire [3-1:0] node4412;
	wire [3-1:0] node4415;
	wire [3-1:0] node4416;
	wire [3-1:0] node4419;
	wire [3-1:0] node4422;
	wire [3-1:0] node4423;
	wire [3-1:0] node4424;
	wire [3-1:0] node4427;
	wire [3-1:0] node4430;
	wire [3-1:0] node4431;
	wire [3-1:0] node4434;
	wire [3-1:0] node4437;
	wire [3-1:0] node4438;
	wire [3-1:0] node4439;
	wire [3-1:0] node4440;
	wire [3-1:0] node4441;
	wire [3-1:0] node4444;
	wire [3-1:0] node4447;
	wire [3-1:0] node4448;
	wire [3-1:0] node4451;
	wire [3-1:0] node4454;
	wire [3-1:0] node4455;
	wire [3-1:0] node4458;
	wire [3-1:0] node4461;
	wire [3-1:0] node4462;
	wire [3-1:0] node4463;
	wire [3-1:0] node4464;
	wire [3-1:0] node4465;
	wire [3-1:0] node4468;
	wire [3-1:0] node4471;
	wire [3-1:0] node4473;
	wire [3-1:0] node4476;
	wire [3-1:0] node4477;
	wire [3-1:0] node4480;
	wire [3-1:0] node4483;
	wire [3-1:0] node4484;
	wire [3-1:0] node4487;
	wire [3-1:0] node4490;
	wire [3-1:0] node4491;
	wire [3-1:0] node4492;
	wire [3-1:0] node4493;
	wire [3-1:0] node4494;
	wire [3-1:0] node4495;
	wire [3-1:0] node4496;
	wire [3-1:0] node4499;
	wire [3-1:0] node4502;
	wire [3-1:0] node4503;
	wire [3-1:0] node4506;
	wire [3-1:0] node4509;
	wire [3-1:0] node4510;
	wire [3-1:0] node4511;
	wire [3-1:0] node4514;
	wire [3-1:0] node4517;
	wire [3-1:0] node4518;
	wire [3-1:0] node4521;
	wire [3-1:0] node4524;
	wire [3-1:0] node4525;
	wire [3-1:0] node4526;
	wire [3-1:0] node4527;
	wire [3-1:0] node4528;
	wire [3-1:0] node4531;
	wire [3-1:0] node4534;
	wire [3-1:0] node4535;
	wire [3-1:0] node4536;
	wire [3-1:0] node4539;
	wire [3-1:0] node4542;
	wire [3-1:0] node4543;
	wire [3-1:0] node4546;
	wire [3-1:0] node4549;
	wire [3-1:0] node4550;
	wire [3-1:0] node4553;
	wire [3-1:0] node4556;
	wire [3-1:0] node4557;
	wire [3-1:0] node4558;
	wire [3-1:0] node4562;
	wire [3-1:0] node4565;
	wire [3-1:0] node4566;
	wire [3-1:0] node4567;
	wire [3-1:0] node4568;
	wire [3-1:0] node4569;
	wire [3-1:0] node4570;
	wire [3-1:0] node4574;
	wire [3-1:0] node4575;
	wire [3-1:0] node4578;
	wire [3-1:0] node4581;
	wire [3-1:0] node4582;
	wire [3-1:0] node4585;
	wire [3-1:0] node4588;
	wire [3-1:0] node4589;
	wire [3-1:0] node4590;
	wire [3-1:0] node4593;
	wire [3-1:0] node4596;
	wire [3-1:0] node4597;
	wire [3-1:0] node4600;
	wire [3-1:0] node4603;
	wire [3-1:0] node4604;
	wire [3-1:0] node4605;
	wire [3-1:0] node4606;
	wire [3-1:0] node4607;
	wire [3-1:0] node4608;
	wire [3-1:0] node4611;
	wire [3-1:0] node4614;
	wire [3-1:0] node4616;
	wire [3-1:0] node4619;
	wire [3-1:0] node4620;
	wire [3-1:0] node4623;
	wire [3-1:0] node4626;
	wire [3-1:0] node4627;
	wire [3-1:0] node4630;
	wire [3-1:0] node4633;
	wire [3-1:0] node4634;
	wire [3-1:0] node4635;
	wire [3-1:0] node4639;
	wire [3-1:0] node4642;
	wire [3-1:0] node4643;
	wire [3-1:0] node4644;
	wire [3-1:0] node4645;
	wire [3-1:0] node4646;
	wire [3-1:0] node4647;
	wire [3-1:0] node4650;
	wire [3-1:0] node4653;
	wire [3-1:0] node4654;
	wire [3-1:0] node4657;
	wire [3-1:0] node4660;
	wire [3-1:0] node4661;
	wire [3-1:0] node4662;
	wire [3-1:0] node4663;
	wire [3-1:0] node4666;
	wire [3-1:0] node4669;
	wire [3-1:0] node4670;
	wire [3-1:0] node4673;
	wire [3-1:0] node4676;
	wire [3-1:0] node4677;
	wire [3-1:0] node4680;
	wire [3-1:0] node4683;
	wire [3-1:0] node4684;
	wire [3-1:0] node4685;
	wire [3-1:0] node4686;
	wire [3-1:0] node4689;
	wire [3-1:0] node4692;
	wire [3-1:0] node4693;
	wire [3-1:0] node4696;
	wire [3-1:0] node4699;
	wire [3-1:0] node4700;
	wire [3-1:0] node4701;
	wire [3-1:0] node4702;
	wire [3-1:0] node4705;
	wire [3-1:0] node4708;
	wire [3-1:0] node4709;
	wire [3-1:0] node4712;
	wire [3-1:0] node4715;
	wire [3-1:0] node4716;
	wire [3-1:0] node4719;
	wire [3-1:0] node4722;
	wire [3-1:0] node4723;
	wire [3-1:0] node4724;
	wire [3-1:0] node4725;
	wire [3-1:0] node4726;
	wire [3-1:0] node4727;
	wire [3-1:0] node4730;
	wire [3-1:0] node4733;
	wire [3-1:0] node4734;
	wire [3-1:0] node4737;
	wire [3-1:0] node4740;
	wire [3-1:0] node4741;
	wire [3-1:0] node4744;
	wire [3-1:0] node4747;
	wire [3-1:0] node4748;
	wire [3-1:0] node4749;
	wire [3-1:0] node4750;
	wire [3-1:0] node4753;
	wire [3-1:0] node4756;
	wire [3-1:0] node4757;
	wire [3-1:0] node4760;
	wire [3-1:0] node4763;
	wire [3-1:0] node4764;
	wire [3-1:0] node4767;
	wire [3-1:0] node4770;
	wire [3-1:0] node4771;
	wire [3-1:0] node4772;
	wire [3-1:0] node4773;
	wire [3-1:0] node4774;
	wire [3-1:0] node4776;
	wire [3-1:0] node4779;
	wire [3-1:0] node4780;
	wire [3-1:0] node4784;
	wire [3-1:0] node4785;
	wire [3-1:0] node4788;
	wire [3-1:0] node4791;
	wire [3-1:0] node4792;
	wire [3-1:0] node4794;
	wire [3-1:0] node4797;
	wire [3-1:0] node4798;
	wire [3-1:0] node4801;
	wire [3-1:0] node4804;
	wire [3-1:0] node4805;
	wire [3-1:0] node4806;
	wire [3-1:0] node4807;
	wire [3-1:0] node4810;
	wire [3-1:0] node4813;
	wire [3-1:0] node4814;
	wire [3-1:0] node4817;
	wire [3-1:0] node4820;
	wire [3-1:0] node4821;
	wire [3-1:0] node4822;
	wire [3-1:0] node4825;
	wire [3-1:0] node4828;
	wire [3-1:0] node4829;
	wire [3-1:0] node4832;

	assign outp = (inp[11]) ? node3020 : node1;
		assign node1 = (inp[6]) ? node1435 : node2;
			assign node2 = (inp[0]) ? node684 : node3;
				assign node3 = (inp[1]) ? node349 : node4;
					assign node4 = (inp[10]) ? node186 : node5;
						assign node5 = (inp[9]) ? node89 : node6;
							assign node6 = (inp[7]) ? node48 : node7;
								assign node7 = (inp[2]) ? node31 : node8;
									assign node8 = (inp[4]) ? node20 : node9;
										assign node9 = (inp[8]) ? node15 : node10;
											assign node10 = (inp[3]) ? node12 : 3'b111;
												assign node12 = (inp[5]) ? 3'b101 : 3'b111;
											assign node15 = (inp[3]) ? node17 : 3'b101;
												assign node17 = (inp[5]) ? 3'b111 : 3'b101;
										assign node20 = (inp[8]) ? node26 : node21;
											assign node21 = (inp[5]) ? node23 : 3'b101;
												assign node23 = (inp[3]) ? 3'b111 : 3'b101;
											assign node26 = (inp[3]) ? node28 : 3'b111;
												assign node28 = (inp[5]) ? 3'b101 : 3'b111;
									assign node31 = (inp[4]) ? node37 : node32;
										assign node32 = (inp[8]) ? 3'b101 : node33;
											assign node33 = (inp[3]) ? 3'b101 : 3'b111;
										assign node37 = (inp[8]) ? node43 : node38;
											assign node38 = (inp[5]) ? node40 : 3'b101;
												assign node40 = (inp[3]) ? 3'b110 : 3'b101;
											assign node43 = (inp[3]) ? node45 : 3'b110;
												assign node45 = (inp[5]) ? 3'b100 : 3'b110;
								assign node48 = (inp[2]) ? node70 : node49;
									assign node49 = (inp[5]) ? node57 : node50;
										assign node50 = (inp[8]) ? node54 : node51;
											assign node51 = (inp[4]) ? 3'b100 : 3'b110;
											assign node54 = (inp[4]) ? 3'b110 : 3'b100;
										assign node57 = (inp[4]) ? node63 : node58;
											assign node58 = (inp[8]) ? node60 : 3'b100;
												assign node60 = (inp[3]) ? 3'b110 : 3'b100;
											assign node63 = (inp[3]) ? node67 : node64;
												assign node64 = (inp[8]) ? 3'b110 : 3'b100;
												assign node67 = (inp[8]) ? 3'b100 : 3'b110;
									assign node70 = (inp[8]) ? node80 : node71;
										assign node71 = (inp[5]) ? node75 : node72;
											assign node72 = (inp[4]) ? 3'b100 : 3'b110;
											assign node75 = (inp[3]) ? node77 : 3'b100;
												assign node77 = (inp[4]) ? 3'b111 : 3'b100;
										assign node80 = (inp[4]) ? node84 : node81;
											assign node81 = (inp[5]) ? 3'b111 : 3'b100;
											assign node84 = (inp[3]) ? node86 : 3'b111;
												assign node86 = (inp[5]) ? 3'b101 : 3'b111;
							assign node89 = (inp[7]) ? node141 : node90;
								assign node90 = (inp[2]) ? node118 : node91;
									assign node91 = (inp[3]) ? node105 : node92;
										assign node92 = (inp[5]) ? node100 : node93;
											assign node93 = (inp[4]) ? node97 : node94;
												assign node94 = (inp[8]) ? 3'b100 : 3'b110;
												assign node97 = (inp[8]) ? 3'b110 : 3'b100;
											assign node100 = (inp[8]) ? 3'b100 : node101;
												assign node101 = (inp[4]) ? 3'b100 : 3'b110;
										assign node105 = (inp[4]) ? node113 : node106;
											assign node106 = (inp[8]) ? node110 : node107;
												assign node107 = (inp[5]) ? 3'b100 : 3'b110;
												assign node110 = (inp[5]) ? 3'b110 : 3'b100;
											assign node113 = (inp[8]) ? 3'b110 : node114;
												assign node114 = (inp[5]) ? 3'b110 : 3'b100;
									assign node118 = (inp[8]) ? node130 : node119;
										assign node119 = (inp[4]) ? node125 : node120;
											assign node120 = (inp[3]) ? node122 : 3'b110;
												assign node122 = (inp[5]) ? 3'b100 : 3'b110;
											assign node125 = (inp[3]) ? node127 : 3'b100;
												assign node127 = (inp[5]) ? 3'b111 : 3'b100;
										assign node130 = (inp[4]) ? node136 : node131;
											assign node131 = (inp[3]) ? node133 : 3'b100;
												assign node133 = (inp[5]) ? 3'b111 : 3'b100;
											assign node136 = (inp[3]) ? node138 : 3'b111;
												assign node138 = (inp[5]) ? 3'b101 : 3'b111;
								assign node141 = (inp[2]) ? node165 : node142;
									assign node142 = (inp[3]) ? node150 : node143;
										assign node143 = (inp[4]) ? node147 : node144;
											assign node144 = (inp[8]) ? 3'b101 : 3'b111;
											assign node147 = (inp[8]) ? 3'b111 : 3'b101;
										assign node150 = (inp[4]) ? node158 : node151;
											assign node151 = (inp[5]) ? node155 : node152;
												assign node152 = (inp[8]) ? 3'b101 : 3'b111;
												assign node155 = (inp[8]) ? 3'b111 : 3'b101;
											assign node158 = (inp[5]) ? node162 : node159;
												assign node159 = (inp[8]) ? 3'b111 : 3'b101;
												assign node162 = (inp[8]) ? 3'b101 : 3'b111;
									assign node165 = (inp[8]) ? node177 : node166;
										assign node166 = (inp[4]) ? node172 : node167;
											assign node167 = (inp[5]) ? node169 : 3'b111;
												assign node169 = (inp[3]) ? 3'b101 : 3'b111;
											assign node172 = (inp[5]) ? node174 : 3'b101;
												assign node174 = (inp[3]) ? 3'b110 : 3'b101;
										assign node177 = (inp[4]) ? node181 : node178;
											assign node178 = (inp[5]) ? 3'b110 : 3'b101;
											assign node181 = (inp[3]) ? node183 : 3'b110;
												assign node183 = (inp[5]) ? 3'b100 : 3'b110;
						assign node186 = (inp[5]) ? node246 : node187;
							assign node187 = (inp[8]) ? node223 : node188;
								assign node188 = (inp[4]) ? node208 : node189;
									assign node189 = (inp[3]) ? node201 : node190;
										assign node190 = (inp[2]) ? node196 : node191;
											assign node191 = (inp[9]) ? 3'b010 : node192;
												assign node192 = (inp[7]) ? 3'b010 : 3'b011;
											assign node196 = (inp[9]) ? node198 : 3'b010;
												assign node198 = (inp[7]) ? 3'b011 : 3'b010;
										assign node201 = (inp[7]) ? node205 : node202;
											assign node202 = (inp[9]) ? 3'b010 : 3'b011;
											assign node205 = (inp[9]) ? 3'b011 : 3'b010;
									assign node208 = (inp[2]) ? node216 : node209;
										assign node209 = (inp[9]) ? node213 : node210;
											assign node210 = (inp[7]) ? 3'b000 : 3'b001;
											assign node213 = (inp[7]) ? 3'b001 : 3'b000;
										assign node216 = (inp[3]) ? node218 : 3'b000;
											assign node218 = (inp[7]) ? node220 : 3'b000;
												assign node220 = (inp[9]) ? 3'b001 : 3'b000;
								assign node223 = (inp[4]) ? node231 : node224;
									assign node224 = (inp[9]) ? node228 : node225;
										assign node225 = (inp[7]) ? 3'b000 : 3'b001;
										assign node228 = (inp[7]) ? 3'b001 : 3'b000;
									assign node231 = (inp[9]) ? node239 : node232;
										assign node232 = (inp[2]) ? node236 : node233;
											assign node233 = (inp[7]) ? 3'b010 : 3'b011;
											assign node236 = (inp[7]) ? 3'b011 : 3'b010;
										assign node239 = (inp[7]) ? node243 : node240;
											assign node240 = (inp[2]) ? 3'b011 : 3'b010;
											assign node243 = (inp[2]) ? 3'b010 : 3'b011;
							assign node246 = (inp[7]) ? node298 : node247;
								assign node247 = (inp[9]) ? node271 : node248;
									assign node248 = (inp[2]) ? node258 : node249;
										assign node249 = (inp[8]) ? node251 : 3'b011;
											assign node251 = (inp[3]) ? node255 : node252;
												assign node252 = (inp[4]) ? 3'b011 : 3'b001;
												assign node255 = (inp[4]) ? 3'b001 : 3'b011;
										assign node258 = (inp[8]) ? node266 : node259;
											assign node259 = (inp[3]) ? node263 : node260;
												assign node260 = (inp[4]) ? 3'b001 : 3'b011;
												assign node263 = (inp[4]) ? 3'b010 : 3'b001;
											assign node266 = (inp[3]) ? node268 : 3'b010;
												assign node268 = (inp[4]) ? 3'b000 : 3'b010;
									assign node271 = (inp[2]) ? node285 : node272;
										assign node272 = (inp[3]) ? node280 : node273;
											assign node273 = (inp[8]) ? node277 : node274;
												assign node274 = (inp[4]) ? 3'b000 : 3'b010;
												assign node277 = (inp[4]) ? 3'b010 : 3'b000;
											assign node280 = (inp[4]) ? 3'b000 : node281;
												assign node281 = (inp[8]) ? 3'b010 : 3'b000;
										assign node285 = (inp[4]) ? node291 : node286;
											assign node286 = (inp[3]) ? 3'b000 : node287;
												assign node287 = (inp[8]) ? 3'b000 : 3'b010;
											assign node291 = (inp[3]) ? node295 : node292;
												assign node292 = (inp[8]) ? 3'b011 : 3'b000;
												assign node295 = (inp[8]) ? 3'b001 : 3'b011;
								assign node298 = (inp[9]) ? node326 : node299;
									assign node299 = (inp[2]) ? node313 : node300;
										assign node300 = (inp[3]) ? node306 : node301;
											assign node301 = (inp[4]) ? node303 : 3'b000;
												assign node303 = (inp[8]) ? 3'b010 : 3'b000;
											assign node306 = (inp[8]) ? node310 : node307;
												assign node307 = (inp[4]) ? 3'b010 : 3'b000;
												assign node310 = (inp[4]) ? 3'b000 : 3'b010;
										assign node313 = (inp[3]) ? node321 : node314;
											assign node314 = (inp[4]) ? node318 : node315;
												assign node315 = (inp[8]) ? 3'b000 : 3'b010;
												assign node318 = (inp[8]) ? 3'b011 : 3'b000;
											assign node321 = (inp[4]) ? node323 : 3'b011;
												assign node323 = (inp[8]) ? 3'b001 : 3'b011;
									assign node326 = (inp[2]) ? node334 : node327;
										assign node327 = (inp[4]) ? node329 : 3'b011;
											assign node329 = (inp[3]) ? 3'b011 : node330;
												assign node330 = (inp[8]) ? 3'b011 : 3'b001;
										assign node334 = (inp[4]) ? node342 : node335;
											assign node335 = (inp[3]) ? node339 : node336;
												assign node336 = (inp[8]) ? 3'b001 : 3'b011;
												assign node339 = (inp[8]) ? 3'b010 : 3'b001;
											assign node342 = (inp[8]) ? node346 : node343;
												assign node343 = (inp[3]) ? 3'b010 : 3'b001;
												assign node346 = (inp[3]) ? 3'b000 : 3'b010;
					assign node349 = (inp[10]) ? node511 : node350;
						assign node350 = (inp[9]) ? node428 : node351;
							assign node351 = (inp[7]) ? node389 : node352;
								assign node352 = (inp[2]) ? node372 : node353;
									assign node353 = (inp[4]) ? node363 : node354;
										assign node354 = (inp[8]) ? node358 : node355;
											assign node355 = (inp[5]) ? 3'b001 : 3'b011;
											assign node358 = (inp[5]) ? node360 : 3'b001;
												assign node360 = (inp[3]) ? 3'b011 : 3'b001;
										assign node363 = (inp[3]) ? node365 : 3'b011;
											assign node365 = (inp[8]) ? node369 : node366;
												assign node366 = (inp[5]) ? 3'b011 : 3'b001;
												assign node369 = (inp[5]) ? 3'b001 : 3'b011;
									assign node372 = (inp[8]) ? node378 : node373;
										assign node373 = (inp[4]) ? node375 : 3'b011;
											assign node375 = (inp[3]) ? 3'b010 : 3'b001;
										assign node378 = (inp[4]) ? node384 : node379;
											assign node379 = (inp[5]) ? node381 : 3'b001;
												assign node381 = (inp[3]) ? 3'b010 : 3'b001;
											assign node384 = (inp[5]) ? node386 : 3'b010;
												assign node386 = (inp[3]) ? 3'b000 : 3'b010;
								assign node389 = (inp[2]) ? node413 : node390;
									assign node390 = (inp[8]) ? node402 : node391;
										assign node391 = (inp[4]) ? node397 : node392;
											assign node392 = (inp[5]) ? node394 : 3'b010;
												assign node394 = (inp[3]) ? 3'b000 : 3'b010;
											assign node397 = (inp[5]) ? node399 : 3'b000;
												assign node399 = (inp[3]) ? 3'b010 : 3'b000;
										assign node402 = (inp[4]) ? node408 : node403;
											assign node403 = (inp[5]) ? node405 : 3'b000;
												assign node405 = (inp[3]) ? 3'b010 : 3'b000;
											assign node408 = (inp[3]) ? node410 : 3'b010;
												assign node410 = (inp[5]) ? 3'b000 : 3'b010;
									assign node413 = (inp[8]) ? node421 : node414;
										assign node414 = (inp[4]) ? node416 : 3'b010;
											assign node416 = (inp[3]) ? node418 : 3'b000;
												assign node418 = (inp[5]) ? 3'b011 : 3'b000;
										assign node421 = (inp[4]) ? 3'b011 : node422;
											assign node422 = (inp[3]) ? node424 : 3'b000;
												assign node424 = (inp[5]) ? 3'b011 : 3'b000;
							assign node428 = (inp[7]) ? node466 : node429;
								assign node429 = (inp[2]) ? node447 : node430;
									assign node430 = (inp[8]) ? node440 : node431;
										assign node431 = (inp[4]) ? node435 : node432;
											assign node432 = (inp[3]) ? 3'b000 : 3'b010;
											assign node435 = (inp[3]) ? node437 : 3'b000;
												assign node437 = (inp[5]) ? 3'b010 : 3'b000;
										assign node440 = (inp[4]) ? 3'b010 : node441;
											assign node441 = (inp[5]) ? node443 : 3'b000;
												assign node443 = (inp[3]) ? 3'b010 : 3'b000;
									assign node447 = (inp[4]) ? node459 : node448;
										assign node448 = (inp[8]) ? node454 : node449;
											assign node449 = (inp[3]) ? node451 : 3'b010;
												assign node451 = (inp[5]) ? 3'b000 : 3'b010;
											assign node454 = (inp[3]) ? node456 : 3'b000;
												assign node456 = (inp[5]) ? 3'b011 : 3'b000;
										assign node459 = (inp[8]) ? node463 : node460;
											assign node460 = (inp[3]) ? 3'b011 : 3'b000;
											assign node463 = (inp[5]) ? 3'b001 : 3'b011;
								assign node466 = (inp[2]) ? node490 : node467;
									assign node467 = (inp[5]) ? node481 : node468;
										assign node468 = (inp[3]) ? node476 : node469;
											assign node469 = (inp[8]) ? node473 : node470;
												assign node470 = (inp[4]) ? 3'b001 : 3'b011;
												assign node473 = (inp[4]) ? 3'b011 : 3'b001;
											assign node476 = (inp[4]) ? 3'b011 : node477;
												assign node477 = (inp[8]) ? 3'b001 : 3'b011;
										assign node481 = (inp[4]) ? node483 : 3'b001;
											assign node483 = (inp[8]) ? node487 : node484;
												assign node484 = (inp[3]) ? 3'b011 : 3'b001;
												assign node487 = (inp[3]) ? 3'b001 : 3'b011;
									assign node490 = (inp[4]) ? node502 : node491;
										assign node491 = (inp[8]) ? node497 : node492;
											assign node492 = (inp[5]) ? node494 : 3'b011;
												assign node494 = (inp[3]) ? 3'b001 : 3'b011;
											assign node497 = (inp[5]) ? node499 : 3'b001;
												assign node499 = (inp[3]) ? 3'b010 : 3'b001;
										assign node502 = (inp[8]) ? node508 : node503;
											assign node503 = (inp[3]) ? node505 : 3'b001;
												assign node505 = (inp[5]) ? 3'b010 : 3'b001;
											assign node508 = (inp[5]) ? 3'b000 : 3'b010;
						assign node511 = (inp[9]) ? node605 : node512;
							assign node512 = (inp[7]) ? node558 : node513;
								assign node513 = (inp[2]) ? node535 : node514;
									assign node514 = (inp[5]) ? node528 : node515;
										assign node515 = (inp[4]) ? node523 : node516;
											assign node516 = (inp[8]) ? node520 : node517;
												assign node517 = (inp[3]) ? 3'b101 : 3'b111;
												assign node520 = (inp[3]) ? 3'b111 : 3'b101;
											assign node523 = (inp[8]) ? node525 : 3'b111;
												assign node525 = (inp[3]) ? 3'b101 : 3'b111;
										assign node528 = (inp[8]) ? node532 : node529;
											assign node529 = (inp[4]) ? 3'b111 : 3'b101;
											assign node532 = (inp[4]) ? 3'b101 : 3'b111;
									assign node535 = (inp[8]) ? node547 : node536;
										assign node536 = (inp[4]) ? node542 : node537;
											assign node537 = (inp[3]) ? 3'b101 : node538;
												assign node538 = (inp[5]) ? 3'b101 : 3'b111;
											assign node542 = (inp[5]) ? 3'b110 : node543;
												assign node543 = (inp[3]) ? 3'b110 : 3'b101;
										assign node547 = (inp[4]) ? node553 : node548;
											assign node548 = (inp[3]) ? 3'b110 : node549;
												assign node549 = (inp[5]) ? 3'b110 : 3'b101;
											assign node553 = (inp[5]) ? 3'b100 : node554;
												assign node554 = (inp[3]) ? 3'b100 : 3'b110;
								assign node558 = (inp[2]) ? node582 : node559;
									assign node559 = (inp[4]) ? node571 : node560;
										assign node560 = (inp[8]) ? node566 : node561;
											assign node561 = (inp[5]) ? 3'b100 : node562;
												assign node562 = (inp[3]) ? 3'b100 : 3'b110;
											assign node566 = (inp[3]) ? 3'b110 : node567;
												assign node567 = (inp[5]) ? 3'b110 : 3'b100;
										assign node571 = (inp[8]) ? node577 : node572;
											assign node572 = (inp[5]) ? 3'b110 : node573;
												assign node573 = (inp[3]) ? 3'b110 : 3'b100;
											assign node577 = (inp[3]) ? 3'b100 : node578;
												assign node578 = (inp[5]) ? 3'b100 : 3'b110;
									assign node582 = (inp[4]) ? node594 : node583;
										assign node583 = (inp[8]) ? node589 : node584;
											assign node584 = (inp[5]) ? 3'b100 : node585;
												assign node585 = (inp[3]) ? 3'b100 : 3'b110;
											assign node589 = (inp[5]) ? 3'b111 : node590;
												assign node590 = (inp[3]) ? 3'b111 : 3'b100;
										assign node594 = (inp[8]) ? node600 : node595;
											assign node595 = (inp[5]) ? 3'b111 : node596;
												assign node596 = (inp[3]) ? 3'b111 : 3'b100;
											assign node600 = (inp[3]) ? 3'b101 : node601;
												assign node601 = (inp[5]) ? 3'b101 : 3'b111;
							assign node605 = (inp[7]) ? node649 : node606;
								assign node606 = (inp[2]) ? node630 : node607;
									assign node607 = (inp[4]) ? node619 : node608;
										assign node608 = (inp[8]) ? node614 : node609;
											assign node609 = (inp[3]) ? 3'b100 : node610;
												assign node610 = (inp[5]) ? 3'b100 : 3'b110;
											assign node614 = (inp[5]) ? 3'b110 : node615;
												assign node615 = (inp[3]) ? 3'b110 : 3'b100;
										assign node619 = (inp[8]) ? node625 : node620;
											assign node620 = (inp[3]) ? 3'b110 : node621;
												assign node621 = (inp[5]) ? 3'b110 : 3'b100;
											assign node625 = (inp[5]) ? 3'b100 : node626;
												assign node626 = (inp[3]) ? 3'b100 : 3'b110;
									assign node630 = (inp[4]) ? node642 : node631;
										assign node631 = (inp[8]) ? node637 : node632;
											assign node632 = (inp[5]) ? 3'b100 : node633;
												assign node633 = (inp[3]) ? 3'b100 : 3'b110;
											assign node637 = (inp[3]) ? 3'b111 : node638;
												assign node638 = (inp[5]) ? 3'b111 : 3'b100;
										assign node642 = (inp[8]) ? 3'b101 : node643;
											assign node643 = (inp[3]) ? 3'b111 : node644;
												assign node644 = (inp[5]) ? 3'b111 : 3'b100;
								assign node649 = (inp[2]) ? node667 : node650;
									assign node650 = (inp[5]) ? node660 : node651;
										assign node651 = (inp[4]) ? node653 : 3'b111;
											assign node653 = (inp[3]) ? node657 : node654;
												assign node654 = (inp[8]) ? 3'b111 : 3'b101;
												assign node657 = (inp[8]) ? 3'b101 : 3'b111;
										assign node660 = (inp[4]) ? node664 : node661;
											assign node661 = (inp[8]) ? 3'b111 : 3'b101;
											assign node664 = (inp[8]) ? 3'b101 : 3'b111;
									assign node667 = (inp[4]) ? node677 : node668;
										assign node668 = (inp[8]) ? node672 : node669;
											assign node669 = (inp[5]) ? 3'b101 : 3'b111;
											assign node672 = (inp[3]) ? 3'b110 : node673;
												assign node673 = (inp[5]) ? 3'b110 : 3'b101;
										assign node677 = (inp[8]) ? node679 : 3'b110;
											assign node679 = (inp[5]) ? 3'b100 : node680;
												assign node680 = (inp[3]) ? 3'b100 : 3'b110;
				assign node684 = (inp[10]) ? node1014 : node685;
					assign node685 = (inp[1]) ? node841 : node686;
						assign node686 = (inp[4]) ? node770 : node687;
							assign node687 = (inp[8]) ? node725 : node688;
								assign node688 = (inp[3]) ? node704 : node689;
									assign node689 = (inp[9]) ? node697 : node690;
										assign node690 = (inp[2]) ? node694 : node691;
											assign node691 = (inp[7]) ? 3'b110 : 3'b111;
											assign node694 = (inp[7]) ? 3'b111 : 3'b110;
										assign node697 = (inp[2]) ? node701 : node698;
											assign node698 = (inp[7]) ? 3'b111 : 3'b110;
											assign node701 = (inp[7]) ? 3'b110 : 3'b111;
									assign node704 = (inp[5]) ? node712 : node705;
										assign node705 = (inp[2]) ? 3'b110 : node706;
											assign node706 = (inp[7]) ? 3'b110 : node707;
												assign node707 = (inp[9]) ? 3'b110 : 3'b111;
										assign node712 = (inp[9]) ? node720 : node713;
											assign node713 = (inp[2]) ? node717 : node714;
												assign node714 = (inp[7]) ? 3'b100 : 3'b101;
												assign node717 = (inp[7]) ? 3'b101 : 3'b100;
											assign node720 = (inp[2]) ? 3'b100 : node721;
												assign node721 = (inp[7]) ? 3'b101 : 3'b100;
								assign node725 = (inp[3]) ? node753 : node726;
									assign node726 = (inp[5]) ? node740 : node727;
										assign node727 = (inp[9]) ? node735 : node728;
											assign node728 = (inp[2]) ? node732 : node729;
												assign node729 = (inp[7]) ? 3'b100 : 3'b101;
												assign node732 = (inp[7]) ? 3'b101 : 3'b100;
											assign node735 = (inp[7]) ? node737 : 3'b100;
												assign node737 = (inp[2]) ? 3'b100 : 3'b101;
										assign node740 = (inp[2]) ? node748 : node741;
											assign node741 = (inp[7]) ? node745 : node742;
												assign node742 = (inp[9]) ? 3'b100 : 3'b101;
												assign node745 = (inp[9]) ? 3'b101 : 3'b100;
											assign node748 = (inp[9]) ? 3'b101 : node749;
												assign node749 = (inp[7]) ? 3'b101 : 3'b100;
									assign node753 = (inp[5]) ? node765 : node754;
										assign node754 = (inp[9]) ? node760 : node755;
											assign node755 = (inp[2]) ? 3'b101 : node756;
												assign node756 = (inp[7]) ? 3'b100 : 3'b101;
											assign node760 = (inp[7]) ? node762 : 3'b100;
												assign node762 = (inp[2]) ? 3'b100 : 3'b101;
										assign node765 = (inp[9]) ? 3'b110 : node766;
											assign node766 = (inp[7]) ? 3'b111 : 3'b110;
							assign node770 = (inp[8]) ? node810 : node771;
								assign node771 = (inp[5]) ? node795 : node772;
									assign node772 = (inp[9]) ? node782 : node773;
										assign node773 = (inp[3]) ? 3'b101 : node774;
											assign node774 = (inp[2]) ? node778 : node775;
												assign node775 = (inp[7]) ? 3'b100 : 3'b101;
												assign node778 = (inp[7]) ? 3'b101 : 3'b100;
										assign node782 = (inp[3]) ? node790 : node783;
											assign node783 = (inp[7]) ? node787 : node784;
												assign node784 = (inp[2]) ? 3'b101 : 3'b100;
												assign node787 = (inp[2]) ? 3'b100 : 3'b101;
											assign node790 = (inp[7]) ? node792 : 3'b100;
												assign node792 = (inp[2]) ? 3'b100 : 3'b101;
									assign node795 = (inp[3]) ? node803 : node796;
										assign node796 = (inp[2]) ? 3'b101 : node797;
											assign node797 = (inp[9]) ? node799 : 3'b100;
												assign node799 = (inp[7]) ? 3'b101 : 3'b100;
										assign node803 = (inp[7]) ? node807 : node804;
											assign node804 = (inp[9]) ? 3'b111 : 3'b110;
											assign node807 = (inp[9]) ? 3'b110 : 3'b111;
								assign node810 = (inp[5]) ? node826 : node811;
									assign node811 = (inp[3]) ? node819 : node812;
										assign node812 = (inp[7]) ? node816 : node813;
											assign node813 = (inp[9]) ? 3'b111 : 3'b110;
											assign node816 = (inp[9]) ? 3'b110 : 3'b111;
										assign node819 = (inp[9]) ? node823 : node820;
											assign node820 = (inp[7]) ? 3'b111 : 3'b110;
											assign node823 = (inp[7]) ? 3'b110 : 3'b111;
									assign node826 = (inp[3]) ? node834 : node827;
										assign node827 = (inp[7]) ? node831 : node828;
											assign node828 = (inp[9]) ? 3'b111 : 3'b110;
											assign node831 = (inp[9]) ? 3'b110 : 3'b111;
										assign node834 = (inp[7]) ? node838 : node835;
											assign node835 = (inp[9]) ? 3'b101 : 3'b100;
											assign node838 = (inp[9]) ? 3'b100 : 3'b101;
						assign node841 = (inp[2]) ? node923 : node842;
							assign node842 = (inp[9]) ? node880 : node843;
								assign node843 = (inp[7]) ? node861 : node844;
									assign node844 = (inp[8]) ? node854 : node845;
										assign node845 = (inp[4]) ? node851 : node846;
											assign node846 = (inp[5]) ? node848 : 3'b011;
												assign node848 = (inp[3]) ? 3'b001 : 3'b011;
											assign node851 = (inp[5]) ? 3'b010 : 3'b001;
										assign node854 = (inp[3]) ? node856 : 3'b010;
											assign node856 = (inp[5]) ? node858 : 3'b010;
												assign node858 = (inp[4]) ? 3'b000 : 3'b010;
									assign node861 = (inp[8]) ? node873 : node862;
										assign node862 = (inp[4]) ? node868 : node863;
											assign node863 = (inp[3]) ? node865 : 3'b010;
												assign node865 = (inp[5]) ? 3'b000 : 3'b010;
											assign node868 = (inp[5]) ? node870 : 3'b000;
												assign node870 = (inp[3]) ? 3'b011 : 3'b000;
										assign node873 = (inp[4]) ? 3'b011 : node874;
											assign node874 = (inp[5]) ? node876 : 3'b000;
												assign node876 = (inp[3]) ? 3'b011 : 3'b000;
								assign node880 = (inp[7]) ? node900 : node881;
									assign node881 = (inp[8]) ? node893 : node882;
										assign node882 = (inp[4]) ? node888 : node883;
											assign node883 = (inp[3]) ? node885 : 3'b010;
												assign node885 = (inp[5]) ? 3'b000 : 3'b010;
											assign node888 = (inp[5]) ? node890 : 3'b000;
												assign node890 = (inp[3]) ? 3'b011 : 3'b000;
										assign node893 = (inp[4]) ? 3'b011 : node894;
											assign node894 = (inp[5]) ? node896 : 3'b000;
												assign node896 = (inp[3]) ? 3'b011 : 3'b000;
									assign node900 = (inp[8]) ? node912 : node901;
										assign node901 = (inp[4]) ? node907 : node902;
											assign node902 = (inp[3]) ? node904 : 3'b011;
												assign node904 = (inp[5]) ? 3'b001 : 3'b011;
											assign node907 = (inp[3]) ? node909 : 3'b001;
												assign node909 = (inp[5]) ? 3'b010 : 3'b001;
										assign node912 = (inp[4]) ? node918 : node913;
											assign node913 = (inp[3]) ? node915 : 3'b001;
												assign node915 = (inp[5]) ? 3'b010 : 3'b001;
											assign node918 = (inp[3]) ? node920 : 3'b010;
												assign node920 = (inp[5]) ? 3'b000 : 3'b010;
							assign node923 = (inp[8]) ? node963 : node924;
								assign node924 = (inp[4]) ? node942 : node925;
									assign node925 = (inp[5]) ? node933 : node926;
										assign node926 = (inp[9]) ? node930 : node927;
											assign node927 = (inp[7]) ? 3'b011 : 3'b010;
											assign node930 = (inp[7]) ? 3'b010 : 3'b011;
										assign node933 = (inp[3]) ? node939 : node934;
											assign node934 = (inp[9]) ? node936 : 3'b011;
												assign node936 = (inp[7]) ? 3'b010 : 3'b011;
											assign node939 = (inp[9]) ? 3'b000 : 3'b001;
									assign node942 = (inp[5]) ? node950 : node943;
										assign node943 = (inp[9]) ? node947 : node944;
											assign node944 = (inp[7]) ? 3'b001 : 3'b000;
											assign node947 = (inp[7]) ? 3'b000 : 3'b001;
										assign node950 = (inp[3]) ? node956 : node951;
											assign node951 = (inp[7]) ? 3'b000 : node952;
												assign node952 = (inp[9]) ? 3'b001 : 3'b000;
											assign node956 = (inp[9]) ? node960 : node957;
												assign node957 = (inp[7]) ? 3'b011 : 3'b010;
												assign node960 = (inp[7]) ? 3'b010 : 3'b011;
								assign node963 = (inp[4]) ? node991 : node964;
									assign node964 = (inp[5]) ? node978 : node965;
										assign node965 = (inp[3]) ? node971 : node966;
											assign node966 = (inp[9]) ? 3'b001 : node967;
												assign node967 = (inp[7]) ? 3'b001 : 3'b000;
											assign node971 = (inp[7]) ? node975 : node972;
												assign node972 = (inp[9]) ? 3'b001 : 3'b000;
												assign node975 = (inp[9]) ? 3'b000 : 3'b001;
										assign node978 = (inp[3]) ? node986 : node979;
											assign node979 = (inp[9]) ? node983 : node980;
												assign node980 = (inp[7]) ? 3'b001 : 3'b000;
												assign node983 = (inp[7]) ? 3'b000 : 3'b001;
											assign node986 = (inp[7]) ? 3'b011 : node987;
												assign node987 = (inp[9]) ? 3'b011 : 3'b010;
									assign node991 = (inp[5]) ? node1003 : node992;
										assign node992 = (inp[3]) ? node998 : node993;
											assign node993 = (inp[7]) ? node995 : 3'b010;
												assign node995 = (inp[9]) ? 3'b010 : 3'b011;
											assign node998 = (inp[7]) ? node1000 : 3'b011;
												assign node1000 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1003 = (inp[3]) ? node1009 : node1004;
											assign node1004 = (inp[9]) ? 3'b011 : node1005;
												assign node1005 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1009 = (inp[9]) ? 3'b000 : node1010;
												assign node1010 = (inp[7]) ? 3'b001 : 3'b000;
					assign node1014 = (inp[1]) ? node1228 : node1015;
						assign node1015 = (inp[3]) ? node1115 : node1016;
							assign node1016 = (inp[5]) ? node1062 : node1017;
								assign node1017 = (inp[7]) ? node1037 : node1018;
									assign node1018 = (inp[9]) ? node1026 : node1019;
										assign node1019 = (inp[8]) ? 3'b010 : node1020;
											assign node1020 = (inp[4]) ? node1022 : 3'b011;
												assign node1022 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1026 = (inp[2]) ? node1032 : node1027;
											assign node1027 = (inp[4]) ? 3'b011 : node1028;
												assign node1028 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1032 = (inp[4]) ? 3'b011 : node1033;
												assign node1033 = (inp[8]) ? 3'b001 : 3'b011;
									assign node1037 = (inp[9]) ? node1051 : node1038;
										assign node1038 = (inp[2]) ? node1044 : node1039;
											assign node1039 = (inp[8]) ? 3'b011 : node1040;
												assign node1040 = (inp[4]) ? 3'b000 : 3'b010;
											assign node1044 = (inp[4]) ? node1048 : node1045;
												assign node1045 = (inp[8]) ? 3'b001 : 3'b011;
												assign node1048 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1051 = (inp[2]) ? node1057 : node1052;
											assign node1052 = (inp[4]) ? 3'b001 : node1053;
												assign node1053 = (inp[8]) ? 3'b001 : 3'b011;
											assign node1057 = (inp[8]) ? node1059 : 3'b010;
												assign node1059 = (inp[4]) ? 3'b010 : 3'b000;
								assign node1062 = (inp[2]) ? node1088 : node1063;
									assign node1063 = (inp[9]) ? node1075 : node1064;
										assign node1064 = (inp[7]) ? node1070 : node1065;
											assign node1065 = (inp[8]) ? 3'b001 : node1066;
												assign node1066 = (inp[4]) ? 3'b001 : 3'b011;
											assign node1070 = (inp[4]) ? node1072 : 3'b000;
												assign node1072 = (inp[8]) ? 3'b011 : 3'b000;
										assign node1075 = (inp[7]) ? node1081 : node1076;
											assign node1076 = (inp[4]) ? 3'b011 : node1077;
												assign node1077 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1081 = (inp[8]) ? node1085 : node1082;
												assign node1082 = (inp[4]) ? 3'b001 : 3'b011;
												assign node1085 = (inp[4]) ? 3'b010 : 3'b001;
									assign node1088 = (inp[9]) ? node1102 : node1089;
										assign node1089 = (inp[7]) ? node1095 : node1090;
											assign node1090 = (inp[4]) ? node1092 : 3'b010;
												assign node1092 = (inp[8]) ? 3'b010 : 3'b000;
											assign node1095 = (inp[4]) ? node1099 : node1096;
												assign node1096 = (inp[8]) ? 3'b001 : 3'b011;
												assign node1099 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1102 = (inp[7]) ? node1108 : node1103;
											assign node1103 = (inp[8]) ? 3'b001 : node1104;
												assign node1104 = (inp[4]) ? 3'b001 : 3'b011;
											assign node1108 = (inp[8]) ? node1112 : node1109;
												assign node1109 = (inp[4]) ? 3'b000 : 3'b010;
												assign node1112 = (inp[4]) ? 3'b010 : 3'b000;
							assign node1115 = (inp[8]) ? node1177 : node1116;
								assign node1116 = (inp[4]) ? node1148 : node1117;
									assign node1117 = (inp[5]) ? node1133 : node1118;
										assign node1118 = (inp[2]) ? node1126 : node1119;
											assign node1119 = (inp[7]) ? node1123 : node1120;
												assign node1120 = (inp[9]) ? 3'b010 : 3'b011;
												assign node1123 = (inp[9]) ? 3'b011 : 3'b010;
											assign node1126 = (inp[9]) ? node1130 : node1127;
												assign node1127 = (inp[7]) ? 3'b011 : 3'b010;
												assign node1130 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1133 = (inp[9]) ? node1141 : node1134;
											assign node1134 = (inp[7]) ? node1138 : node1135;
												assign node1135 = (inp[2]) ? 3'b000 : 3'b001;
												assign node1138 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1141 = (inp[7]) ? node1145 : node1142;
												assign node1142 = (inp[2]) ? 3'b001 : 3'b000;
												assign node1145 = (inp[2]) ? 3'b000 : 3'b001;
									assign node1148 = (inp[5]) ? node1162 : node1149;
										assign node1149 = (inp[7]) ? node1155 : node1150;
											assign node1150 = (inp[2]) ? node1152 : 3'b000;
												assign node1152 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1155 = (inp[2]) ? node1159 : node1156;
												assign node1156 = (inp[9]) ? 3'b001 : 3'b000;
												assign node1159 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1162 = (inp[2]) ? node1170 : node1163;
											assign node1163 = (inp[7]) ? node1167 : node1164;
												assign node1164 = (inp[9]) ? 3'b011 : 3'b010;
												assign node1167 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1170 = (inp[7]) ? node1174 : node1171;
												assign node1171 = (inp[9]) ? 3'b011 : 3'b010;
												assign node1174 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1177 = (inp[2]) ? node1205 : node1178;
									assign node1178 = (inp[9]) ? node1194 : node1179;
										assign node1179 = (inp[7]) ? node1187 : node1180;
											assign node1180 = (inp[4]) ? node1184 : node1181;
												assign node1181 = (inp[5]) ? 3'b010 : 3'b001;
												assign node1184 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1187 = (inp[4]) ? node1191 : node1188;
												assign node1188 = (inp[5]) ? 3'b011 : 3'b000;
												assign node1191 = (inp[5]) ? 3'b001 : 3'b011;
										assign node1194 = (inp[4]) ? node1200 : node1195;
											assign node1195 = (inp[5]) ? 3'b011 : node1196;
												assign node1196 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1200 = (inp[7]) ? node1202 : 3'b001;
												assign node1202 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1205 = (inp[7]) ? node1215 : node1206;
										assign node1206 = (inp[9]) ? node1208 : 3'b010;
											assign node1208 = (inp[5]) ? node1212 : node1209;
												assign node1209 = (inp[4]) ? 3'b011 : 3'b001;
												assign node1212 = (inp[4]) ? 3'b001 : 3'b011;
										assign node1215 = (inp[9]) ? node1221 : node1216;
											assign node1216 = (inp[5]) ? 3'b001 : node1217;
												assign node1217 = (inp[4]) ? 3'b011 : 3'b001;
											assign node1221 = (inp[5]) ? node1225 : node1222;
												assign node1222 = (inp[4]) ? 3'b010 : 3'b000;
												assign node1225 = (inp[4]) ? 3'b000 : 3'b010;
						assign node1228 = (inp[5]) ? node1328 : node1229;
							assign node1229 = (inp[4]) ? node1287 : node1230;
								assign node1230 = (inp[7]) ? node1256 : node1231;
									assign node1231 = (inp[9]) ? node1245 : node1232;
										assign node1232 = (inp[2]) ? node1238 : node1233;
											assign node1233 = (inp[8]) ? node1235 : 3'b101;
												assign node1235 = (inp[3]) ? 3'b110 : 3'b101;
											assign node1238 = (inp[8]) ? node1242 : node1239;
												assign node1239 = (inp[3]) ? 3'b100 : 3'b110;
												assign node1242 = (inp[3]) ? 3'b110 : 3'b100;
										assign node1245 = (inp[2]) ? node1251 : node1246;
											assign node1246 = (inp[3]) ? 3'b111 : node1247;
												assign node1247 = (inp[8]) ? 3'b100 : 3'b110;
											assign node1251 = (inp[8]) ? 3'b101 : node1252;
												assign node1252 = (inp[3]) ? 3'b101 : 3'b111;
									assign node1256 = (inp[9]) ? node1272 : node1257;
										assign node1257 = (inp[2]) ? node1265 : node1258;
											assign node1258 = (inp[3]) ? node1262 : node1259;
												assign node1259 = (inp[8]) ? 3'b100 : 3'b110;
												assign node1262 = (inp[8]) ? 3'b111 : 3'b100;
											assign node1265 = (inp[3]) ? node1269 : node1266;
												assign node1266 = (inp[8]) ? 3'b101 : 3'b111;
												assign node1269 = (inp[8]) ? 3'b111 : 3'b101;
										assign node1272 = (inp[2]) ? node1280 : node1273;
											assign node1273 = (inp[3]) ? node1277 : node1274;
												assign node1274 = (inp[8]) ? 3'b101 : 3'b111;
												assign node1277 = (inp[8]) ? 3'b110 : 3'b101;
											assign node1280 = (inp[8]) ? node1284 : node1281;
												assign node1281 = (inp[3]) ? 3'b100 : 3'b110;
												assign node1284 = (inp[3]) ? 3'b110 : 3'b100;
								assign node1287 = (inp[8]) ? node1305 : node1288;
									assign node1288 = (inp[3]) ? node1298 : node1289;
										assign node1289 = (inp[9]) ? 3'b100 : node1290;
											assign node1290 = (inp[7]) ? node1294 : node1291;
												assign node1291 = (inp[2]) ? 3'b100 : 3'b101;
												assign node1294 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1298 = (inp[9]) ? node1302 : node1299;
											assign node1299 = (inp[7]) ? 3'b111 : 3'b110;
											assign node1302 = (inp[7]) ? 3'b110 : 3'b111;
									assign node1305 = (inp[3]) ? node1321 : node1306;
										assign node1306 = (inp[2]) ? node1314 : node1307;
											assign node1307 = (inp[9]) ? node1311 : node1308;
												assign node1308 = (inp[7]) ? 3'b111 : 3'b110;
												assign node1311 = (inp[7]) ? 3'b110 : 3'b111;
											assign node1314 = (inp[7]) ? node1318 : node1315;
												assign node1315 = (inp[9]) ? 3'b111 : 3'b110;
												assign node1318 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1321 = (inp[2]) ? node1323 : 3'b100;
											assign node1323 = (inp[9]) ? node1325 : 3'b100;
												assign node1325 = (inp[7]) ? 3'b100 : 3'b101;
							assign node1328 = (inp[3]) ? node1374 : node1329;
								assign node1329 = (inp[4]) ? node1353 : node1330;
									assign node1330 = (inp[8]) ? node1346 : node1331;
										assign node1331 = (inp[9]) ? node1339 : node1332;
											assign node1332 = (inp[2]) ? node1336 : node1333;
												assign node1333 = (inp[7]) ? 3'b100 : 3'b101;
												assign node1336 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1339 = (inp[7]) ? node1343 : node1340;
												assign node1340 = (inp[2]) ? 3'b101 : 3'b100;
												assign node1343 = (inp[2]) ? 3'b100 : 3'b101;
										assign node1346 = (inp[7]) ? node1350 : node1347;
											assign node1347 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1350 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1353 = (inp[8]) ? node1359 : node1354;
										assign node1354 = (inp[7]) ? node1356 : 3'b111;
											assign node1356 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1359 = (inp[2]) ? node1367 : node1360;
											assign node1360 = (inp[7]) ? node1364 : node1361;
												assign node1361 = (inp[9]) ? 3'b101 : 3'b100;
												assign node1364 = (inp[9]) ? 3'b100 : 3'b101;
											assign node1367 = (inp[9]) ? node1371 : node1368;
												assign node1368 = (inp[7]) ? 3'b101 : 3'b100;
												assign node1371 = (inp[7]) ? 3'b100 : 3'b101;
								assign node1374 = (inp[2]) ? node1406 : node1375;
									assign node1375 = (inp[7]) ? node1391 : node1376;
										assign node1376 = (inp[9]) ? node1384 : node1377;
											assign node1377 = (inp[4]) ? node1381 : node1378;
												assign node1378 = (inp[8]) ? 3'b110 : 3'b101;
												assign node1381 = (inp[8]) ? 3'b100 : 3'b110;
											assign node1384 = (inp[4]) ? node1388 : node1385;
												assign node1385 = (inp[8]) ? 3'b111 : 3'b100;
												assign node1388 = (inp[8]) ? 3'b101 : 3'b111;
										assign node1391 = (inp[9]) ? node1399 : node1392;
											assign node1392 = (inp[4]) ? node1396 : node1393;
												assign node1393 = (inp[8]) ? 3'b111 : 3'b100;
												assign node1396 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1399 = (inp[8]) ? node1403 : node1400;
												assign node1400 = (inp[4]) ? 3'b110 : 3'b101;
												assign node1403 = (inp[4]) ? 3'b100 : 3'b110;
									assign node1406 = (inp[8]) ? node1420 : node1407;
										assign node1407 = (inp[4]) ? node1415 : node1408;
											assign node1408 = (inp[7]) ? node1412 : node1409;
												assign node1409 = (inp[9]) ? 3'b101 : 3'b100;
												assign node1412 = (inp[9]) ? 3'b100 : 3'b101;
											assign node1415 = (inp[7]) ? node1417 : 3'b111;
												assign node1417 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1420 = (inp[4]) ? node1428 : node1421;
											assign node1421 = (inp[9]) ? node1425 : node1422;
												assign node1422 = (inp[7]) ? 3'b111 : 3'b110;
												assign node1425 = (inp[7]) ? 3'b110 : 3'b111;
											assign node1428 = (inp[7]) ? node1432 : node1429;
												assign node1429 = (inp[9]) ? 3'b101 : 3'b100;
												assign node1432 = (inp[9]) ? 3'b100 : 3'b101;
			assign node1435 = (inp[5]) ? node2137 : node1436;
				assign node1436 = (inp[4]) ? node1776 : node1437;
					assign node1437 = (inp[8]) ? node1603 : node1438;
						assign node1438 = (inp[3]) ? node1512 : node1439;
							assign node1439 = (inp[1]) ? node1477 : node1440;
								assign node1440 = (inp[10]) ? node1460 : node1441;
									assign node1441 = (inp[9]) ? node1449 : node1442;
										assign node1442 = (inp[7]) ? node1444 : 3'b011;
											assign node1444 = (inp[2]) ? node1446 : 3'b010;
												assign node1446 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1449 = (inp[7]) ? node1455 : node1450;
											assign node1450 = (inp[2]) ? node1452 : 3'b010;
												assign node1452 = (inp[0]) ? 3'b011 : 3'b010;
											assign node1455 = (inp[0]) ? node1457 : 3'b011;
												assign node1457 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1460 = (inp[7]) ? node1472 : node1461;
										assign node1461 = (inp[9]) ? node1467 : node1462;
											assign node1462 = (inp[2]) ? node1464 : 3'b111;
												assign node1464 = (inp[0]) ? 3'b110 : 3'b111;
											assign node1467 = (inp[0]) ? node1469 : 3'b110;
												assign node1469 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1472 = (inp[9]) ? node1474 : 3'b110;
											assign node1474 = (inp[2]) ? 3'b110 : 3'b111;
								assign node1477 = (inp[10]) ? node1497 : node1478;
									assign node1478 = (inp[7]) ? node1486 : node1479;
										assign node1479 = (inp[9]) ? node1481 : 3'b111;
											assign node1481 = (inp[0]) ? node1483 : 3'b110;
												assign node1483 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1486 = (inp[9]) ? node1492 : node1487;
											assign node1487 = (inp[2]) ? node1489 : 3'b110;
												assign node1489 = (inp[0]) ? 3'b111 : 3'b110;
											assign node1492 = (inp[2]) ? node1494 : 3'b111;
												assign node1494 = (inp[0]) ? 3'b110 : 3'b111;
									assign node1497 = (inp[9]) ? node1507 : node1498;
										assign node1498 = (inp[7]) ? node1504 : node1499;
											assign node1499 = (inp[0]) ? node1501 : 3'b011;
												assign node1501 = (inp[2]) ? 3'b010 : 3'b011;
											assign node1504 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1507 = (inp[7]) ? 3'b011 : node1508;
											assign node1508 = (inp[2]) ? 3'b011 : 3'b010;
							assign node1512 = (inp[10]) ? node1556 : node1513;
								assign node1513 = (inp[1]) ? node1535 : node1514;
									assign node1514 = (inp[7]) ? node1526 : node1515;
										assign node1515 = (inp[9]) ? node1521 : node1516;
											assign node1516 = (inp[0]) ? node1518 : 3'b011;
												assign node1518 = (inp[2]) ? 3'b010 : 3'b011;
											assign node1521 = (inp[2]) ? node1523 : 3'b010;
												assign node1523 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1526 = (inp[9]) ? node1530 : node1527;
											assign node1527 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1530 = (inp[0]) ? node1532 : 3'b011;
												assign node1532 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1535 = (inp[7]) ? node1547 : node1536;
										assign node1536 = (inp[9]) ? node1542 : node1537;
											assign node1537 = (inp[2]) ? node1539 : 3'b101;
												assign node1539 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1542 = (inp[2]) ? node1544 : 3'b100;
												assign node1544 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1547 = (inp[9]) ? node1551 : node1548;
											assign node1548 = (inp[2]) ? 3'b101 : 3'b100;
											assign node1551 = (inp[2]) ? node1553 : 3'b101;
												assign node1553 = (inp[0]) ? 3'b100 : 3'b101;
								assign node1556 = (inp[1]) ? node1580 : node1557;
									assign node1557 = (inp[7]) ? node1569 : node1558;
										assign node1558 = (inp[9]) ? node1564 : node1559;
											assign node1559 = (inp[2]) ? node1561 : 3'b101;
												assign node1561 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1564 = (inp[2]) ? node1566 : 3'b100;
												assign node1566 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1569 = (inp[9]) ? node1575 : node1570;
											assign node1570 = (inp[2]) ? node1572 : 3'b100;
												assign node1572 = (inp[0]) ? 3'b101 : 3'b100;
											assign node1575 = (inp[0]) ? node1577 : 3'b101;
												assign node1577 = (inp[2]) ? 3'b100 : 3'b101;
									assign node1580 = (inp[0]) ? node1588 : node1581;
										assign node1581 = (inp[7]) ? node1585 : node1582;
											assign node1582 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1585 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1588 = (inp[9]) ? node1596 : node1589;
											assign node1589 = (inp[7]) ? node1593 : node1590;
												assign node1590 = (inp[2]) ? 3'b000 : 3'b001;
												assign node1593 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1596 = (inp[7]) ? node1600 : node1597;
												assign node1597 = (inp[2]) ? 3'b001 : 3'b000;
												assign node1600 = (inp[2]) ? 3'b000 : 3'b001;
						assign node1603 = (inp[3]) ? node1697 : node1604;
							assign node1604 = (inp[0]) ? node1642 : node1605;
								assign node1605 = (inp[10]) ? node1621 : node1606;
									assign node1606 = (inp[1]) ? node1614 : node1607;
										assign node1607 = (inp[9]) ? node1611 : node1608;
											assign node1608 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1611 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1614 = (inp[7]) ? node1618 : node1615;
											assign node1615 = (inp[9]) ? 3'b100 : 3'b101;
											assign node1618 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1621 = (inp[1]) ? node1635 : node1622;
										assign node1622 = (inp[2]) ? node1630 : node1623;
											assign node1623 = (inp[7]) ? node1627 : node1624;
												assign node1624 = (inp[9]) ? 3'b100 : 3'b101;
												assign node1627 = (inp[9]) ? 3'b101 : 3'b100;
											assign node1630 = (inp[7]) ? 3'b101 : node1631;
												assign node1631 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1635 = (inp[7]) ? node1639 : node1636;
											assign node1636 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1639 = (inp[9]) ? 3'b001 : 3'b000;
								assign node1642 = (inp[10]) ? node1674 : node1643;
									assign node1643 = (inp[1]) ? node1659 : node1644;
										assign node1644 = (inp[2]) ? node1652 : node1645;
											assign node1645 = (inp[9]) ? node1649 : node1646;
												assign node1646 = (inp[7]) ? 3'b000 : 3'b001;
												assign node1649 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1652 = (inp[9]) ? node1656 : node1653;
												assign node1653 = (inp[7]) ? 3'b001 : 3'b000;
												assign node1656 = (inp[7]) ? 3'b000 : 3'b001;
										assign node1659 = (inp[2]) ? node1667 : node1660;
											assign node1660 = (inp[9]) ? node1664 : node1661;
												assign node1661 = (inp[7]) ? 3'b100 : 3'b101;
												assign node1664 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1667 = (inp[7]) ? node1671 : node1668;
												assign node1668 = (inp[9]) ? 3'b101 : 3'b100;
												assign node1671 = (inp[9]) ? 3'b100 : 3'b101;
									assign node1674 = (inp[1]) ? node1690 : node1675;
										assign node1675 = (inp[9]) ? node1683 : node1676;
											assign node1676 = (inp[2]) ? node1680 : node1677;
												assign node1677 = (inp[7]) ? 3'b100 : 3'b101;
												assign node1680 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1683 = (inp[2]) ? node1687 : node1684;
												assign node1684 = (inp[7]) ? 3'b101 : 3'b100;
												assign node1687 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1690 = (inp[9]) ? node1692 : 3'b000;
											assign node1692 = (inp[2]) ? node1694 : 3'b001;
												assign node1694 = (inp[7]) ? 3'b000 : 3'b001;
							assign node1697 = (inp[1]) ? node1739 : node1698;
								assign node1698 = (inp[10]) ? node1722 : node1699;
									assign node1699 = (inp[2]) ? node1707 : node1700;
										assign node1700 = (inp[9]) ? node1704 : node1701;
											assign node1701 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1704 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1707 = (inp[0]) ? node1715 : node1708;
											assign node1708 = (inp[9]) ? node1712 : node1709;
												assign node1709 = (inp[7]) ? 3'b000 : 3'b001;
												assign node1712 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1715 = (inp[7]) ? node1719 : node1716;
												assign node1716 = (inp[9]) ? 3'b001 : 3'b000;
												assign node1719 = (inp[9]) ? 3'b000 : 3'b001;
									assign node1722 = (inp[2]) ? node1732 : node1723;
										assign node1723 = (inp[9]) ? node1725 : 3'b110;
											assign node1725 = (inp[0]) ? node1729 : node1726;
												assign node1726 = (inp[7]) ? 3'b111 : 3'b110;
												assign node1729 = (inp[7]) ? 3'b110 : 3'b111;
										assign node1732 = (inp[7]) ? node1736 : node1733;
											assign node1733 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1736 = (inp[9]) ? 3'b110 : 3'b111;
								assign node1739 = (inp[10]) ? node1761 : node1740;
									assign node1740 = (inp[2]) ? node1754 : node1741;
										assign node1741 = (inp[9]) ? node1749 : node1742;
											assign node1742 = (inp[0]) ? node1746 : node1743;
												assign node1743 = (inp[7]) ? 3'b110 : 3'b111;
												assign node1746 = (inp[7]) ? 3'b111 : 3'b110;
											assign node1749 = (inp[0]) ? node1751 : 3'b110;
												assign node1751 = (inp[7]) ? 3'b110 : 3'b111;
										assign node1754 = (inp[9]) ? node1758 : node1755;
											assign node1755 = (inp[7]) ? 3'b111 : 3'b110;
											assign node1758 = (inp[7]) ? 3'b110 : 3'b111;
									assign node1761 = (inp[2]) ? node1769 : node1762;
										assign node1762 = (inp[9]) ? 3'b010 : node1763;
											assign node1763 = (inp[0]) ? node1765 : 3'b010;
												assign node1765 = (inp[7]) ? 3'b011 : 3'b010;
										assign node1769 = (inp[9]) ? node1773 : node1770;
											assign node1770 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1773 = (inp[7]) ? 3'b010 : 3'b011;
					assign node1776 = (inp[8]) ? node1964 : node1777;
						assign node1777 = (inp[3]) ? node1873 : node1778;
							assign node1778 = (inp[7]) ? node1826 : node1779;
								assign node1779 = (inp[9]) ? node1803 : node1780;
									assign node1780 = (inp[2]) ? node1788 : node1781;
										assign node1781 = (inp[1]) ? node1785 : node1782;
											assign node1782 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1785 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1788 = (inp[0]) ? node1796 : node1789;
											assign node1789 = (inp[1]) ? node1793 : node1790;
												assign node1790 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1793 = (inp[10]) ? 3'b001 : 3'b101;
											assign node1796 = (inp[10]) ? node1800 : node1797;
												assign node1797 = (inp[1]) ? 3'b100 : 3'b000;
												assign node1800 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1803 = (inp[0]) ? node1811 : node1804;
										assign node1804 = (inp[10]) ? node1808 : node1805;
											assign node1805 = (inp[1]) ? 3'b100 : 3'b000;
											assign node1808 = (inp[1]) ? 3'b000 : 3'b100;
										assign node1811 = (inp[2]) ? node1819 : node1812;
											assign node1812 = (inp[10]) ? node1816 : node1813;
												assign node1813 = (inp[1]) ? 3'b100 : 3'b000;
												assign node1816 = (inp[1]) ? 3'b000 : 3'b100;
											assign node1819 = (inp[10]) ? node1823 : node1820;
												assign node1820 = (inp[1]) ? 3'b101 : 3'b001;
												assign node1823 = (inp[1]) ? 3'b001 : 3'b101;
								assign node1826 = (inp[9]) ? node1846 : node1827;
									assign node1827 = (inp[2]) ? node1833 : node1828;
										assign node1828 = (inp[10]) ? 3'b100 : node1829;
											assign node1829 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1833 = (inp[0]) ? node1839 : node1834;
											assign node1834 = (inp[10]) ? 3'b100 : node1835;
												assign node1835 = (inp[1]) ? 3'b100 : 3'b000;
											assign node1839 = (inp[1]) ? node1843 : node1840;
												assign node1840 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1843 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1846 = (inp[0]) ? node1862 : node1847;
										assign node1847 = (inp[2]) ? node1855 : node1848;
											assign node1848 = (inp[1]) ? node1852 : node1849;
												assign node1849 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1852 = (inp[10]) ? 3'b001 : 3'b101;
											assign node1855 = (inp[1]) ? node1859 : node1856;
												assign node1856 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1859 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1862 = (inp[2]) ? node1868 : node1863;
											assign node1863 = (inp[1]) ? node1865 : 3'b101;
												assign node1865 = (inp[10]) ? 3'b001 : 3'b101;
											assign node1868 = (inp[1]) ? 3'b100 : node1869;
												assign node1869 = (inp[10]) ? 3'b100 : 3'b000;
							assign node1873 = (inp[10]) ? node1925 : node1874;
								assign node1874 = (inp[1]) ? node1902 : node1875;
									assign node1875 = (inp[2]) ? node1889 : node1876;
										assign node1876 = (inp[0]) ? node1884 : node1877;
											assign node1877 = (inp[7]) ? node1881 : node1878;
												assign node1878 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1881 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1884 = (inp[9]) ? node1886 : 3'b000;
												assign node1886 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1889 = (inp[7]) ? node1897 : node1890;
											assign node1890 = (inp[0]) ? node1894 : node1891;
												assign node1891 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1894 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1897 = (inp[9]) ? 3'b000 : node1898;
												assign node1898 = (inp[0]) ? 3'b001 : 3'b000;
									assign node1902 = (inp[2]) ? node1918 : node1903;
										assign node1903 = (inp[0]) ? node1911 : node1904;
											assign node1904 = (inp[9]) ? node1908 : node1905;
												assign node1905 = (inp[7]) ? 3'b110 : 3'b111;
												assign node1908 = (inp[7]) ? 3'b111 : 3'b110;
											assign node1911 = (inp[9]) ? node1915 : node1912;
												assign node1912 = (inp[7]) ? 3'b111 : 3'b110;
												assign node1915 = (inp[7]) ? 3'b110 : 3'b111;
										assign node1918 = (inp[7]) ? node1922 : node1919;
											assign node1919 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1922 = (inp[9]) ? 3'b110 : 3'b111;
								assign node1925 = (inp[1]) ? node1943 : node1926;
									assign node1926 = (inp[9]) ? node1934 : node1927;
										assign node1927 = (inp[7]) ? node1929 : 3'b110;
											assign node1929 = (inp[2]) ? 3'b111 : node1930;
												assign node1930 = (inp[0]) ? 3'b111 : 3'b110;
										assign node1934 = (inp[7]) ? node1940 : node1935;
											assign node1935 = (inp[2]) ? 3'b111 : node1936;
												assign node1936 = (inp[0]) ? 3'b111 : 3'b110;
											assign node1940 = (inp[0]) ? 3'b110 : 3'b111;
									assign node1943 = (inp[9]) ? node1953 : node1944;
										assign node1944 = (inp[7]) ? node1950 : node1945;
											assign node1945 = (inp[2]) ? 3'b010 : node1946;
												assign node1946 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1950 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1953 = (inp[7]) ? node1959 : node1954;
											assign node1954 = (inp[2]) ? 3'b011 : node1955;
												assign node1955 = (inp[0]) ? 3'b011 : 3'b010;
											assign node1959 = (inp[0]) ? 3'b010 : node1960;
												assign node1960 = (inp[2]) ? 3'b010 : 3'b011;
						assign node1964 = (inp[3]) ? node2050 : node1965;
							assign node1965 = (inp[10]) ? node2011 : node1966;
								assign node1966 = (inp[1]) ? node1990 : node1967;
									assign node1967 = (inp[9]) ? node1979 : node1968;
										assign node1968 = (inp[7]) ? node1974 : node1969;
											assign node1969 = (inp[2]) ? 3'b010 : node1970;
												assign node1970 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1974 = (inp[0]) ? 3'b011 : node1975;
												assign node1975 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1979 = (inp[7]) ? node1985 : node1980;
											assign node1980 = (inp[0]) ? 3'b011 : node1981;
												assign node1981 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1985 = (inp[0]) ? 3'b010 : node1986;
												assign node1986 = (inp[2]) ? 3'b010 : 3'b011;
									assign node1990 = (inp[7]) ? node2000 : node1991;
										assign node1991 = (inp[9]) ? node1995 : node1992;
											assign node1992 = (inp[0]) ? 3'b110 : 3'b111;
											assign node1995 = (inp[0]) ? 3'b111 : node1996;
												assign node1996 = (inp[2]) ? 3'b111 : 3'b110;
										assign node2000 = (inp[9]) ? node2006 : node2001;
											assign node2001 = (inp[0]) ? 3'b111 : node2002;
												assign node2002 = (inp[2]) ? 3'b111 : 3'b110;
											assign node2006 = (inp[2]) ? 3'b110 : node2007;
												assign node2007 = (inp[0]) ? 3'b110 : 3'b111;
								assign node2011 = (inp[1]) ? node2033 : node2012;
									assign node2012 = (inp[2]) ? node2026 : node2013;
										assign node2013 = (inp[0]) ? node2019 : node2014;
											assign node2014 = (inp[7]) ? node2016 : 3'b111;
												assign node2016 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2019 = (inp[7]) ? node2023 : node2020;
												assign node2020 = (inp[9]) ? 3'b111 : 3'b110;
												assign node2023 = (inp[9]) ? 3'b110 : 3'b111;
										assign node2026 = (inp[9]) ? node2030 : node2027;
											assign node2027 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2030 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2033 = (inp[9]) ? node2045 : node2034;
										assign node2034 = (inp[7]) ? node2040 : node2035;
											assign node2035 = (inp[2]) ? 3'b010 : node2036;
												assign node2036 = (inp[0]) ? 3'b010 : 3'b011;
											assign node2040 = (inp[2]) ? 3'b011 : node2041;
												assign node2041 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2045 = (inp[7]) ? 3'b010 : node2046;
											assign node2046 = (inp[0]) ? 3'b011 : 3'b010;
							assign node2050 = (inp[1]) ? node2098 : node2051;
								assign node2051 = (inp[10]) ? node2069 : node2052;
									assign node2052 = (inp[2]) ? node2062 : node2053;
										assign node2053 = (inp[9]) ? 3'b010 : node2054;
											assign node2054 = (inp[0]) ? node2058 : node2055;
												assign node2055 = (inp[7]) ? 3'b010 : 3'b011;
												assign node2058 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2062 = (inp[9]) ? node2066 : node2063;
											assign node2063 = (inp[7]) ? 3'b011 : 3'b010;
											assign node2066 = (inp[7]) ? 3'b010 : 3'b011;
									assign node2069 = (inp[2]) ? node2083 : node2070;
										assign node2070 = (inp[0]) ? node2076 : node2071;
											assign node2071 = (inp[9]) ? 3'b101 : node2072;
												assign node2072 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2076 = (inp[9]) ? node2080 : node2077;
												assign node2077 = (inp[7]) ? 3'b101 : 3'b100;
												assign node2080 = (inp[7]) ? 3'b100 : 3'b101;
										assign node2083 = (inp[0]) ? node2091 : node2084;
											assign node2084 = (inp[7]) ? node2088 : node2085;
												assign node2085 = (inp[9]) ? 3'b101 : 3'b100;
												assign node2088 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2091 = (inp[7]) ? node2095 : node2092;
												assign node2092 = (inp[9]) ? 3'b101 : 3'b100;
												assign node2095 = (inp[9]) ? 3'b100 : 3'b101;
								assign node2098 = (inp[10]) ? node2122 : node2099;
									assign node2099 = (inp[0]) ? node2115 : node2100;
										assign node2100 = (inp[7]) ? node2108 : node2101;
											assign node2101 = (inp[9]) ? node2105 : node2102;
												assign node2102 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2105 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2108 = (inp[2]) ? node2112 : node2109;
												assign node2109 = (inp[9]) ? 3'b101 : 3'b100;
												assign node2112 = (inp[9]) ? 3'b100 : 3'b101;
										assign node2115 = (inp[7]) ? node2119 : node2116;
											assign node2116 = (inp[9]) ? 3'b101 : 3'b100;
											assign node2119 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2122 = (inp[9]) ? node2128 : node2123;
										assign node2123 = (inp[7]) ? node2125 : 3'b000;
											assign node2125 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2128 = (inp[7]) ? node2132 : node2129;
											assign node2129 = (inp[2]) ? 3'b001 : 3'b000;
											assign node2132 = (inp[2]) ? 3'b000 : node2133;
												assign node2133 = (inp[0]) ? 3'b000 : 3'b001;
				assign node2137 = (inp[3]) ? node2599 : node2138;
					assign node2138 = (inp[7]) ? node2368 : node2139;
						assign node2139 = (inp[9]) ? node2253 : node2140;
							assign node2140 = (inp[2]) ? node2196 : node2141;
								assign node2141 = (inp[0]) ? node2169 : node2142;
									assign node2142 = (inp[4]) ? node2156 : node2143;
										assign node2143 = (inp[8]) ? node2149 : node2144;
											assign node2144 = (inp[10]) ? node2146 : 3'b101;
												assign node2146 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2149 = (inp[1]) ? node2153 : node2150;
												assign node2150 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2153 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2156 = (inp[8]) ? node2164 : node2157;
											assign node2157 = (inp[1]) ? node2161 : node2158;
												assign node2158 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2161 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2164 = (inp[1]) ? node2166 : 3'b011;
												assign node2166 = (inp[10]) ? 3'b001 : 3'b101;
									assign node2169 = (inp[8]) ? node2183 : node2170;
										assign node2170 = (inp[4]) ? node2178 : node2171;
											assign node2171 = (inp[1]) ? node2175 : node2172;
												assign node2172 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2175 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2178 = (inp[10]) ? node2180 : 3'b001;
												assign node2180 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2183 = (inp[4]) ? node2191 : node2184;
											assign node2184 = (inp[1]) ? node2188 : node2185;
												assign node2185 = (inp[10]) ? 3'b110 : 3'b001;
												assign node2188 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2191 = (inp[1]) ? node2193 : 3'b010;
												assign node2193 = (inp[10]) ? 3'b000 : 3'b100;
								assign node2196 = (inp[0]) ? node2224 : node2197;
									assign node2197 = (inp[8]) ? node2209 : node2198;
										assign node2198 = (inp[4]) ? node2204 : node2199;
											assign node2199 = (inp[1]) ? node2201 : 3'b101;
												assign node2201 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2204 = (inp[10]) ? node2206 : 3'b001;
												assign node2206 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2209 = (inp[4]) ? node2217 : node2210;
											assign node2210 = (inp[1]) ? node2214 : node2211;
												assign node2211 = (inp[10]) ? 3'b110 : 3'b001;
												assign node2214 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2217 = (inp[10]) ? node2221 : node2218;
												assign node2218 = (inp[1]) ? 3'b100 : 3'b010;
												assign node2221 = (inp[1]) ? 3'b000 : 3'b100;
									assign node2224 = (inp[4]) ? node2240 : node2225;
										assign node2225 = (inp[8]) ? node2233 : node2226;
											assign node2226 = (inp[1]) ? node2230 : node2227;
												assign node2227 = (inp[10]) ? 3'b100 : 3'b010;
												assign node2230 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2233 = (inp[1]) ? node2237 : node2234;
												assign node2234 = (inp[10]) ? 3'b110 : 3'b000;
												assign node2237 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2240 = (inp[8]) ? node2248 : node2241;
											assign node2241 = (inp[10]) ? node2245 : node2242;
												assign node2242 = (inp[1]) ? 3'b110 : 3'b000;
												assign node2245 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2248 = (inp[1]) ? node2250 : 3'b100;
												assign node2250 = (inp[10]) ? 3'b000 : 3'b100;
							assign node2253 = (inp[0]) ? node2307 : node2254;
								assign node2254 = (inp[2]) ? node2278 : node2255;
									assign node2255 = (inp[8]) ? node2265 : node2256;
										assign node2256 = (inp[4]) ? 3'b110 : node2257;
											assign node2257 = (inp[10]) ? node2261 : node2258;
												assign node2258 = (inp[1]) ? 3'b100 : 3'b010;
												assign node2261 = (inp[1]) ? 3'b000 : 3'b100;
										assign node2265 = (inp[4]) ? node2271 : node2266;
											assign node2266 = (inp[10]) ? node2268 : 3'b000;
												assign node2268 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2271 = (inp[10]) ? node2275 : node2272;
												assign node2272 = (inp[1]) ? 3'b100 : 3'b010;
												assign node2275 = (inp[1]) ? 3'b000 : 3'b100;
									assign node2278 = (inp[8]) ? node2292 : node2279;
										assign node2279 = (inp[4]) ? node2287 : node2280;
											assign node2280 = (inp[10]) ? node2284 : node2281;
												assign node2281 = (inp[1]) ? 3'b100 : 3'b010;
												assign node2284 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2287 = (inp[10]) ? node2289 : 3'b000;
												assign node2289 = (inp[1]) ? 3'b011 : 3'b111;
										assign node2292 = (inp[4]) ? node2300 : node2293;
											assign node2293 = (inp[1]) ? node2297 : node2294;
												assign node2294 = (inp[10]) ? 3'b111 : 3'b000;
												assign node2297 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2300 = (inp[1]) ? node2304 : node2301;
												assign node2301 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2304 = (inp[10]) ? 3'b001 : 3'b101;
								assign node2307 = (inp[2]) ? node2339 : node2308;
									assign node2308 = (inp[4]) ? node2324 : node2309;
										assign node2309 = (inp[8]) ? node2317 : node2310;
											assign node2310 = (inp[1]) ? node2314 : node2311;
												assign node2311 = (inp[10]) ? 3'b100 : 3'b010;
												assign node2314 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2317 = (inp[1]) ? node2321 : node2318;
												assign node2318 = (inp[10]) ? 3'b111 : 3'b000;
												assign node2321 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2324 = (inp[8]) ? node2332 : node2325;
											assign node2325 = (inp[10]) ? node2329 : node2326;
												assign node2326 = (inp[1]) ? 3'b111 : 3'b000;
												assign node2329 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2332 = (inp[10]) ? node2336 : node2333;
												assign node2333 = (inp[1]) ? 3'b101 : 3'b011;
												assign node2336 = (inp[1]) ? 3'b001 : 3'b101;
									assign node2339 = (inp[4]) ? node2353 : node2340;
										assign node2340 = (inp[8]) ? node2348 : node2341;
											assign node2341 = (inp[10]) ? node2345 : node2342;
												assign node2342 = (inp[1]) ? 3'b101 : 3'b011;
												assign node2345 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2348 = (inp[10]) ? node2350 : 3'b001;
												assign node2350 = (inp[1]) ? 3'b011 : 3'b111;
										assign node2353 = (inp[8]) ? node2361 : node2354;
											assign node2354 = (inp[1]) ? node2358 : node2355;
												assign node2355 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2358 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2361 = (inp[1]) ? node2365 : node2362;
												assign node2362 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2365 = (inp[10]) ? 3'b001 : 3'b101;
						assign node2368 = (inp[9]) ? node2486 : node2369;
							assign node2369 = (inp[2]) ? node2427 : node2370;
								assign node2370 = (inp[0]) ? node2398 : node2371;
									assign node2371 = (inp[8]) ? node2385 : node2372;
										assign node2372 = (inp[4]) ? node2378 : node2373;
											assign node2373 = (inp[10]) ? node2375 : 3'b010;
												assign node2375 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2378 = (inp[10]) ? node2382 : node2379;
												assign node2379 = (inp[1]) ? 3'b110 : 3'b000;
												assign node2382 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2385 = (inp[4]) ? node2391 : node2386;
											assign node2386 = (inp[10]) ? 3'b110 : node2387;
												assign node2387 = (inp[1]) ? 3'b110 : 3'b000;
											assign node2391 = (inp[10]) ? node2395 : node2392;
												assign node2392 = (inp[1]) ? 3'b100 : 3'b010;
												assign node2395 = (inp[1]) ? 3'b000 : 3'b100;
									assign node2398 = (inp[4]) ? node2414 : node2399;
										assign node2399 = (inp[8]) ? node2407 : node2400;
											assign node2400 = (inp[1]) ? node2404 : node2401;
												assign node2401 = (inp[10]) ? 3'b100 : 3'b010;
												assign node2404 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2407 = (inp[10]) ? node2411 : node2408;
												assign node2408 = (inp[1]) ? 3'b111 : 3'b000;
												assign node2411 = (inp[1]) ? 3'b011 : 3'b111;
										assign node2414 = (inp[8]) ? node2422 : node2415;
											assign node2415 = (inp[1]) ? node2419 : node2416;
												assign node2416 = (inp[10]) ? 3'b111 : 3'b000;
												assign node2419 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2422 = (inp[1]) ? node2424 : 3'b011;
												assign node2424 = (inp[10]) ? 3'b001 : 3'b101;
								assign node2427 = (inp[0]) ? node2457 : node2428;
									assign node2428 = (inp[8]) ? node2442 : node2429;
										assign node2429 = (inp[4]) ? node2437 : node2430;
											assign node2430 = (inp[1]) ? node2434 : node2431;
												assign node2431 = (inp[10]) ? 3'b100 : 3'b010;
												assign node2434 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2437 = (inp[1]) ? node2439 : 3'b000;
												assign node2439 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2442 = (inp[4]) ? node2450 : node2443;
											assign node2443 = (inp[10]) ? node2447 : node2444;
												assign node2444 = (inp[1]) ? 3'b111 : 3'b000;
												assign node2447 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2450 = (inp[1]) ? node2454 : node2451;
												assign node2451 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2454 = (inp[10]) ? 3'b001 : 3'b101;
									assign node2457 = (inp[4]) ? node2473 : node2458;
										assign node2458 = (inp[8]) ? node2466 : node2459;
											assign node2459 = (inp[1]) ? node2463 : node2460;
												assign node2460 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2463 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2466 = (inp[1]) ? node2470 : node2467;
												assign node2467 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2470 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2473 = (inp[8]) ? node2479 : node2474;
											assign node2474 = (inp[1]) ? node2476 : 3'b001;
												assign node2476 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2479 = (inp[10]) ? node2483 : node2480;
												assign node2480 = (inp[1]) ? 3'b101 : 3'b011;
												assign node2483 = (inp[1]) ? 3'b001 : 3'b101;
							assign node2486 = (inp[2]) ? node2548 : node2487;
								assign node2487 = (inp[0]) ? node2519 : node2488;
									assign node2488 = (inp[4]) ? node2504 : node2489;
										assign node2489 = (inp[8]) ? node2497 : node2490;
											assign node2490 = (inp[1]) ? node2494 : node2491;
												assign node2491 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2494 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2497 = (inp[1]) ? node2501 : node2498;
												assign node2498 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2501 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2504 = (inp[8]) ? node2512 : node2505;
											assign node2505 = (inp[1]) ? node2509 : node2506;
												assign node2506 = (inp[10]) ? 3'b111 : 3'b001;
												assign node2509 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2512 = (inp[10]) ? node2516 : node2513;
												assign node2513 = (inp[1]) ? 3'b101 : 3'b011;
												assign node2516 = (inp[1]) ? 3'b001 : 3'b101;
									assign node2519 = (inp[8]) ? node2535 : node2520;
										assign node2520 = (inp[4]) ? node2528 : node2521;
											assign node2521 = (inp[1]) ? node2525 : node2522;
												assign node2522 = (inp[10]) ? 3'b101 : 3'b011;
												assign node2525 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2528 = (inp[1]) ? node2532 : node2529;
												assign node2529 = (inp[10]) ? 3'b110 : 3'b001;
												assign node2532 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2535 = (inp[4]) ? node2543 : node2536;
											assign node2536 = (inp[10]) ? node2540 : node2537;
												assign node2537 = (inp[1]) ? 3'b110 : 3'b001;
												assign node2540 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2543 = (inp[1]) ? node2545 : 3'b010;
												assign node2545 = (inp[10]) ? 3'b000 : 3'b100;
								assign node2548 = (inp[0]) ? node2578 : node2549;
									assign node2549 = (inp[8]) ? node2563 : node2550;
										assign node2550 = (inp[4]) ? node2556 : node2551;
											assign node2551 = (inp[1]) ? node2553 : 3'b011;
												assign node2553 = (inp[10]) ? 3'b001 : 3'b101;
											assign node2556 = (inp[1]) ? node2560 : node2557;
												assign node2557 = (inp[10]) ? 3'b110 : 3'b001;
												assign node2560 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2563 = (inp[4]) ? node2571 : node2564;
											assign node2564 = (inp[10]) ? node2568 : node2565;
												assign node2565 = (inp[1]) ? 3'b110 : 3'b001;
												assign node2568 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2571 = (inp[1]) ? node2575 : node2572;
												assign node2572 = (inp[10]) ? 3'b100 : 3'b010;
												assign node2575 = (inp[10]) ? 3'b000 : 3'b100;
									assign node2578 = (inp[4]) ? node2586 : node2579;
										assign node2579 = (inp[1]) ? node2583 : node2580;
											assign node2580 = (inp[8]) ? 3'b000 : 3'b010;
											assign node2583 = (inp[8]) ? 3'b010 : 3'b000;
										assign node2586 = (inp[8]) ? node2594 : node2587;
											assign node2587 = (inp[10]) ? node2591 : node2588;
												assign node2588 = (inp[1]) ? 3'b110 : 3'b000;
												assign node2591 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2594 = (inp[10]) ? node2596 : 3'b010;
												assign node2596 = (inp[1]) ? 3'b000 : 3'b100;
					assign node2599 = (inp[7]) ? node2801 : node2600;
						assign node2600 = (inp[9]) ? node2704 : node2601;
							assign node2601 = (inp[0]) ? node2655 : node2602;
								assign node2602 = (inp[2]) ? node2628 : node2603;
									assign node2603 = (inp[4]) ? node2615 : node2604;
										assign node2604 = (inp[8]) ? node2612 : node2605;
											assign node2605 = (inp[10]) ? node2609 : node2606;
												assign node2606 = (inp[1]) ? 3'b101 : 3'b001;
												assign node2609 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2612 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2615 = (inp[8]) ? node2623 : node2616;
											assign node2616 = (inp[10]) ? node2620 : node2617;
												assign node2617 = (inp[1]) ? 3'b111 : 3'b011;
												assign node2620 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2623 = (inp[10]) ? node2625 : 3'b101;
												assign node2625 = (inp[1]) ? 3'b001 : 3'b101;
									assign node2628 = (inp[8]) ? node2642 : node2629;
										assign node2629 = (inp[4]) ? node2637 : node2630;
											assign node2630 = (inp[10]) ? node2634 : node2631;
												assign node2631 = (inp[1]) ? 3'b101 : 3'b001;
												assign node2634 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2637 = (inp[1]) ? node2639 : 3'b010;
												assign node2639 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2642 = (inp[4]) ? node2650 : node2643;
											assign node2643 = (inp[10]) ? node2647 : node2644;
												assign node2644 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2647 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2650 = (inp[10]) ? node2652 : 3'b100;
												assign node2652 = (inp[1]) ? 3'b000 : 3'b100;
								assign node2655 = (inp[2]) ? node2679 : node2656;
									assign node2656 = (inp[8]) ? node2668 : node2657;
										assign node2657 = (inp[4]) ? node2663 : node2658;
											assign node2658 = (inp[10]) ? 3'b101 : node2659;
												assign node2659 = (inp[1]) ? 3'b101 : 3'b001;
											assign node2663 = (inp[1]) ? 3'b110 : node2664;
												assign node2664 = (inp[10]) ? 3'b110 : 3'b010;
										assign node2668 = (inp[4]) ? node2674 : node2669;
											assign node2669 = (inp[10]) ? node2671 : 3'b010;
												assign node2671 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2674 = (inp[1]) ? node2676 : 3'b100;
												assign node2676 = (inp[10]) ? 3'b000 : 3'b100;
									assign node2679 = (inp[4]) ? node2695 : node2680;
										assign node2680 = (inp[8]) ? node2688 : node2681;
											assign node2681 = (inp[10]) ? node2685 : node2682;
												assign node2682 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2685 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2688 = (inp[10]) ? node2692 : node2689;
												assign node2689 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2692 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2695 = (inp[8]) ? node2697 : 3'b010;
											assign node2697 = (inp[1]) ? node2701 : node2698;
												assign node2698 = (inp[10]) ? 3'b100 : 3'b000;
												assign node2701 = (inp[10]) ? 3'b000 : 3'b100;
							assign node2704 = (inp[2]) ? node2756 : node2705;
								assign node2705 = (inp[0]) ? node2735 : node2706;
									assign node2706 = (inp[4]) ? node2722 : node2707;
										assign node2707 = (inp[8]) ? node2715 : node2708;
											assign node2708 = (inp[10]) ? node2712 : node2709;
												assign node2709 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2712 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2715 = (inp[10]) ? node2719 : node2716;
												assign node2716 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2719 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2722 = (inp[8]) ? node2728 : node2723;
											assign node2723 = (inp[1]) ? 3'b010 : node2724;
												assign node2724 = (inp[10]) ? 3'b110 : 3'b010;
											assign node2728 = (inp[10]) ? node2732 : node2729;
												assign node2729 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2732 = (inp[1]) ? 3'b000 : 3'b100;
									assign node2735 = (inp[4]) ? node2743 : node2736;
										assign node2736 = (inp[8]) ? 3'b011 : node2737;
											assign node2737 = (inp[1]) ? 3'b000 : node2738;
												assign node2738 = (inp[10]) ? 3'b100 : 3'b000;
										assign node2743 = (inp[8]) ? node2751 : node2744;
											assign node2744 = (inp[1]) ? node2748 : node2745;
												assign node2745 = (inp[10]) ? 3'b111 : 3'b011;
												assign node2748 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2751 = (inp[1]) ? 3'b101 : node2752;
												assign node2752 = (inp[10]) ? 3'b101 : 3'b001;
								assign node2756 = (inp[4]) ? node2786 : node2757;
									assign node2757 = (inp[8]) ? node2773 : node2758;
										assign node2758 = (inp[0]) ? node2766 : node2759;
											assign node2759 = (inp[10]) ? node2763 : node2760;
												assign node2760 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2763 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2766 = (inp[1]) ? node2770 : node2767;
												assign node2767 = (inp[10]) ? 3'b101 : 3'b001;
												assign node2770 = (inp[10]) ? 3'b001 : 3'b101;
										assign node2773 = (inp[0]) ? node2781 : node2774;
											assign node2774 = (inp[1]) ? node2778 : node2775;
												assign node2775 = (inp[10]) ? 3'b111 : 3'b011;
												assign node2778 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2781 = (inp[10]) ? node2783 : 3'b011;
												assign node2783 = (inp[1]) ? 3'b011 : 3'b111;
									assign node2786 = (inp[8]) ? node2794 : node2787;
										assign node2787 = (inp[10]) ? node2791 : node2788;
											assign node2788 = (inp[1]) ? 3'b111 : 3'b011;
											assign node2791 = (inp[1]) ? 3'b011 : 3'b111;
										assign node2794 = (inp[1]) ? node2798 : node2795;
											assign node2795 = (inp[10]) ? 3'b101 : 3'b001;
											assign node2798 = (inp[10]) ? 3'b001 : 3'b101;
						assign node2801 = (inp[9]) ? node2917 : node2802;
							assign node2802 = (inp[0]) ? node2864 : node2803;
								assign node2803 = (inp[2]) ? node2833 : node2804;
									assign node2804 = (inp[8]) ? node2818 : node2805;
										assign node2805 = (inp[4]) ? node2811 : node2806;
											assign node2806 = (inp[10]) ? node2808 : 3'b000;
												assign node2808 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2811 = (inp[10]) ? node2815 : node2812;
												assign node2812 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2815 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2818 = (inp[4]) ? node2826 : node2819;
											assign node2819 = (inp[10]) ? node2823 : node2820;
												assign node2820 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2823 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2826 = (inp[1]) ? node2830 : node2827;
												assign node2827 = (inp[10]) ? 3'b100 : 3'b000;
												assign node2830 = (inp[10]) ? 3'b000 : 3'b100;
									assign node2833 = (inp[4]) ? node2849 : node2834;
										assign node2834 = (inp[8]) ? node2842 : node2835;
											assign node2835 = (inp[10]) ? node2839 : node2836;
												assign node2836 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2839 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2842 = (inp[1]) ? node2846 : node2843;
												assign node2843 = (inp[10]) ? 3'b111 : 3'b011;
												assign node2846 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2849 = (inp[8]) ? node2857 : node2850;
											assign node2850 = (inp[10]) ? node2854 : node2851;
												assign node2851 = (inp[1]) ? 3'b111 : 3'b011;
												assign node2854 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2857 = (inp[10]) ? node2861 : node2858;
												assign node2858 = (inp[1]) ? 3'b101 : 3'b001;
												assign node2861 = (inp[1]) ? 3'b001 : 3'b101;
								assign node2864 = (inp[8]) ? node2894 : node2865;
									assign node2865 = (inp[4]) ? node2881 : node2866;
										assign node2866 = (inp[2]) ? node2874 : node2867;
											assign node2867 = (inp[10]) ? node2871 : node2868;
												assign node2868 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2871 = (inp[1]) ? 3'b000 : 3'b100;
											assign node2874 = (inp[1]) ? node2878 : node2875;
												assign node2875 = (inp[10]) ? 3'b101 : 3'b001;
												assign node2878 = (inp[10]) ? 3'b001 : 3'b101;
										assign node2881 = (inp[2]) ? node2889 : node2882;
											assign node2882 = (inp[1]) ? node2886 : node2883;
												assign node2883 = (inp[10]) ? 3'b111 : 3'b011;
												assign node2886 = (inp[10]) ? 3'b011 : 3'b111;
											assign node2889 = (inp[10]) ? 3'b111 : node2890;
												assign node2890 = (inp[1]) ? 3'b111 : 3'b011;
									assign node2894 = (inp[4]) ? node2910 : node2895;
										assign node2895 = (inp[2]) ? node2903 : node2896;
											assign node2896 = (inp[10]) ? node2900 : node2897;
												assign node2897 = (inp[1]) ? 3'b111 : 3'b011;
												assign node2900 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2903 = (inp[1]) ? node2907 : node2904;
												assign node2904 = (inp[10]) ? 3'b111 : 3'b011;
												assign node2907 = (inp[10]) ? 3'b011 : 3'b111;
										assign node2910 = (inp[10]) ? node2914 : node2911;
											assign node2911 = (inp[1]) ? 3'b101 : 3'b001;
											assign node2914 = (inp[1]) ? 3'b001 : 3'b101;
							assign node2917 = (inp[0]) ? node2969 : node2918;
								assign node2918 = (inp[2]) ? node2944 : node2919;
									assign node2919 = (inp[10]) ? node2935 : node2920;
										assign node2920 = (inp[1]) ? node2928 : node2921;
											assign node2921 = (inp[4]) ? node2925 : node2922;
												assign node2922 = (inp[8]) ? 3'b011 : 3'b001;
												assign node2925 = (inp[8]) ? 3'b001 : 3'b011;
											assign node2928 = (inp[8]) ? node2932 : node2929;
												assign node2929 = (inp[4]) ? 3'b111 : 3'b101;
												assign node2932 = (inp[4]) ? 3'b101 : 3'b111;
										assign node2935 = (inp[1]) ? 3'b011 : node2936;
											assign node2936 = (inp[8]) ? node2940 : node2937;
												assign node2937 = (inp[4]) ? 3'b111 : 3'b101;
												assign node2940 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2944 = (inp[8]) ? node2958 : node2945;
										assign node2945 = (inp[4]) ? node2953 : node2946;
											assign node2946 = (inp[10]) ? node2950 : node2947;
												assign node2947 = (inp[1]) ? 3'b101 : 3'b001;
												assign node2950 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2953 = (inp[1]) ? node2955 : 3'b110;
												assign node2955 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2958 = (inp[4]) ? node2964 : node2959;
											assign node2959 = (inp[10]) ? node2961 : 3'b110;
												assign node2961 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2964 = (inp[10]) ? node2966 : 3'b100;
												assign node2966 = (inp[1]) ? 3'b000 : 3'b100;
								assign node2969 = (inp[8]) ? node2991 : node2970;
									assign node2970 = (inp[4]) ? node2980 : node2971;
										assign node2971 = (inp[2]) ? 3'b100 : node2972;
											assign node2972 = (inp[1]) ? node2976 : node2973;
												assign node2973 = (inp[10]) ? 3'b101 : 3'b001;
												assign node2976 = (inp[10]) ? 3'b001 : 3'b101;
										assign node2980 = (inp[2]) ? node2986 : node2981;
											assign node2981 = (inp[10]) ? 3'b110 : node2982;
												assign node2982 = (inp[1]) ? 3'b110 : 3'b010;
											assign node2986 = (inp[1]) ? node2988 : 3'b010;
												assign node2988 = (inp[10]) ? 3'b010 : 3'b110;
									assign node2991 = (inp[4]) ? node3007 : node2992;
										assign node2992 = (inp[2]) ? node3000 : node2993;
											assign node2993 = (inp[10]) ? node2997 : node2994;
												assign node2994 = (inp[1]) ? 3'b110 : 3'b010;
												assign node2997 = (inp[1]) ? 3'b010 : 3'b110;
											assign node3000 = (inp[10]) ? node3004 : node3001;
												assign node3001 = (inp[1]) ? 3'b110 : 3'b010;
												assign node3004 = (inp[1]) ? 3'b010 : 3'b110;
										assign node3007 = (inp[2]) ? node3015 : node3008;
											assign node3008 = (inp[10]) ? node3012 : node3009;
												assign node3009 = (inp[1]) ? 3'b100 : 3'b000;
												assign node3012 = (inp[1]) ? 3'b000 : 3'b100;
											assign node3015 = (inp[1]) ? node3017 : 3'b100;
												assign node3017 = (inp[10]) ? 3'b000 : 3'b100;
		assign node3020 = (inp[3]) ? node4024 : node3021;
			assign node3021 = (inp[4]) ? node3481 : node3022;
				assign node3022 = (inp[8]) ? node3274 : node3023;
					assign node3023 = (inp[5]) ? node3133 : node3024;
						assign node3024 = (inp[9]) ? node3074 : node3025;
							assign node3025 = (inp[7]) ? node3051 : node3026;
								assign node3026 = (inp[0]) ? node3034 : node3027;
									assign node3027 = (inp[6]) ? node3031 : node3028;
										assign node3028 = (inp[10]) ? 3'b111 : 3'b011;
										assign node3031 = (inp[10]) ? 3'b011 : 3'b111;
									assign node3034 = (inp[2]) ? node3042 : node3035;
										assign node3035 = (inp[6]) ? node3039 : node3036;
											assign node3036 = (inp[10]) ? 3'b111 : 3'b011;
											assign node3039 = (inp[10]) ? 3'b011 : 3'b111;
										assign node3042 = (inp[1]) ? node3044 : 3'b010;
											assign node3044 = (inp[6]) ? node3048 : node3045;
												assign node3045 = (inp[10]) ? 3'b110 : 3'b010;
												assign node3048 = (inp[10]) ? 3'b010 : 3'b110;
								assign node3051 = (inp[0]) ? node3059 : node3052;
									assign node3052 = (inp[6]) ? node3056 : node3053;
										assign node3053 = (inp[10]) ? 3'b110 : 3'b010;
										assign node3056 = (inp[10]) ? 3'b010 : 3'b110;
									assign node3059 = (inp[2]) ? node3067 : node3060;
										assign node3060 = (inp[10]) ? node3064 : node3061;
											assign node3061 = (inp[6]) ? 3'b110 : 3'b010;
											assign node3064 = (inp[6]) ? 3'b010 : 3'b110;
										assign node3067 = (inp[6]) ? node3071 : node3068;
											assign node3068 = (inp[10]) ? 3'b111 : 3'b011;
											assign node3071 = (inp[10]) ? 3'b011 : 3'b111;
							assign node3074 = (inp[7]) ? node3102 : node3075;
								assign node3075 = (inp[2]) ? node3083 : node3076;
									assign node3076 = (inp[6]) ? node3080 : node3077;
										assign node3077 = (inp[10]) ? 3'b110 : 3'b010;
										assign node3080 = (inp[10]) ? 3'b010 : 3'b110;
									assign node3083 = (inp[0]) ? node3093 : node3084;
										assign node3084 = (inp[1]) ? node3086 : 3'b010;
											assign node3086 = (inp[10]) ? node3090 : node3087;
												assign node3087 = (inp[6]) ? 3'b110 : 3'b010;
												assign node3090 = (inp[6]) ? 3'b010 : 3'b110;
										assign node3093 = (inp[1]) ? node3097 : node3094;
											assign node3094 = (inp[6]) ? 3'b111 : 3'b011;
											assign node3097 = (inp[10]) ? node3099 : 3'b011;
												assign node3099 = (inp[6]) ? 3'b011 : 3'b111;
								assign node3102 = (inp[0]) ? node3110 : node3103;
									assign node3103 = (inp[10]) ? node3107 : node3104;
										assign node3104 = (inp[6]) ? 3'b111 : 3'b011;
										assign node3107 = (inp[6]) ? 3'b011 : 3'b111;
									assign node3110 = (inp[2]) ? node3118 : node3111;
										assign node3111 = (inp[6]) ? node3115 : node3112;
											assign node3112 = (inp[10]) ? 3'b111 : 3'b011;
											assign node3115 = (inp[10]) ? 3'b011 : 3'b111;
										assign node3118 = (inp[1]) ? node3126 : node3119;
											assign node3119 = (inp[6]) ? node3123 : node3120;
												assign node3120 = (inp[10]) ? 3'b110 : 3'b010;
												assign node3123 = (inp[10]) ? 3'b010 : 3'b110;
											assign node3126 = (inp[6]) ? node3130 : node3127;
												assign node3127 = (inp[10]) ? 3'b110 : 3'b010;
												assign node3130 = (inp[10]) ? 3'b010 : 3'b110;
						assign node3133 = (inp[6]) ? node3225 : node3134;
							assign node3134 = (inp[10]) ? node3182 : node3135;
								assign node3135 = (inp[1]) ? node3159 : node3136;
									assign node3136 = (inp[0]) ? node3146 : node3137;
										assign node3137 = (inp[2]) ? 3'b010 : node3138;
											assign node3138 = (inp[7]) ? node3142 : node3139;
												assign node3139 = (inp[9]) ? 3'b010 : 3'b011;
												assign node3142 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3146 = (inp[7]) ? node3152 : node3147;
											assign node3147 = (inp[9]) ? node3149 : 3'b010;
												assign node3149 = (inp[2]) ? 3'b011 : 3'b010;
											assign node3152 = (inp[9]) ? node3156 : node3153;
												assign node3153 = (inp[2]) ? 3'b011 : 3'b010;
												assign node3156 = (inp[2]) ? 3'b010 : 3'b011;
									assign node3159 = (inp[0]) ? node3167 : node3160;
										assign node3160 = (inp[9]) ? node3164 : node3161;
											assign node3161 = (inp[7]) ? 3'b010 : 3'b011;
											assign node3164 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3167 = (inp[2]) ? node3175 : node3168;
											assign node3168 = (inp[9]) ? node3172 : node3169;
												assign node3169 = (inp[7]) ? 3'b010 : 3'b011;
												assign node3172 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3175 = (inp[9]) ? node3179 : node3176;
												assign node3176 = (inp[7]) ? 3'b011 : 3'b010;
												assign node3179 = (inp[7]) ? 3'b010 : 3'b011;
								assign node3182 = (inp[2]) ? node3204 : node3183;
									assign node3183 = (inp[1]) ? node3191 : node3184;
										assign node3184 = (inp[7]) ? node3188 : node3185;
											assign node3185 = (inp[9]) ? 3'b100 : 3'b101;
											assign node3188 = (inp[9]) ? 3'b101 : 3'b100;
										assign node3191 = (inp[0]) ? node3197 : node3192;
											assign node3192 = (inp[9]) ? 3'b100 : node3193;
												assign node3193 = (inp[7]) ? 3'b100 : 3'b101;
											assign node3197 = (inp[9]) ? node3201 : node3198;
												assign node3198 = (inp[7]) ? 3'b100 : 3'b101;
												assign node3201 = (inp[7]) ? 3'b101 : 3'b100;
									assign node3204 = (inp[0]) ? node3218 : node3205;
										assign node3205 = (inp[1]) ? node3213 : node3206;
											assign node3206 = (inp[9]) ? node3210 : node3207;
												assign node3207 = (inp[7]) ? 3'b100 : 3'b101;
												assign node3210 = (inp[7]) ? 3'b101 : 3'b100;
											assign node3213 = (inp[7]) ? 3'b101 : node3214;
												assign node3214 = (inp[9]) ? 3'b100 : 3'b101;
										assign node3218 = (inp[7]) ? node3222 : node3219;
											assign node3219 = (inp[9]) ? 3'b101 : 3'b100;
											assign node3222 = (inp[9]) ? 3'b100 : 3'b101;
							assign node3225 = (inp[10]) ? node3249 : node3226;
								assign node3226 = (inp[0]) ? node3234 : node3227;
									assign node3227 = (inp[7]) ? node3231 : node3228;
										assign node3228 = (inp[9]) ? 3'b100 : 3'b101;
										assign node3231 = (inp[9]) ? 3'b101 : 3'b100;
									assign node3234 = (inp[9]) ? node3242 : node3235;
										assign node3235 = (inp[7]) ? node3239 : node3236;
											assign node3236 = (inp[2]) ? 3'b100 : 3'b101;
											assign node3239 = (inp[2]) ? 3'b101 : 3'b100;
										assign node3242 = (inp[7]) ? node3246 : node3243;
											assign node3243 = (inp[2]) ? 3'b101 : 3'b100;
											assign node3246 = (inp[2]) ? 3'b100 : 3'b101;
								assign node3249 = (inp[2]) ? node3257 : node3250;
									assign node3250 = (inp[7]) ? node3254 : node3251;
										assign node3251 = (inp[9]) ? 3'b000 : 3'b001;
										assign node3254 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3257 = (inp[0]) ? node3267 : node3258;
										assign node3258 = (inp[1]) ? node3260 : 3'b001;
											assign node3260 = (inp[7]) ? node3264 : node3261;
												assign node3261 = (inp[9]) ? 3'b000 : 3'b001;
												assign node3264 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3267 = (inp[9]) ? node3271 : node3268;
											assign node3268 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3271 = (inp[7]) ? 3'b000 : 3'b001;
					assign node3274 = (inp[5]) ? node3378 : node3275;
						assign node3275 = (inp[6]) ? node3321 : node3276;
							assign node3276 = (inp[10]) ? node3300 : node3277;
								assign node3277 = (inp[2]) ? node3285 : node3278;
									assign node3278 = (inp[7]) ? node3282 : node3279;
										assign node3279 = (inp[9]) ? 3'b000 : 3'b001;
										assign node3282 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3285 = (inp[7]) ? node3293 : node3286;
										assign node3286 = (inp[0]) ? node3290 : node3287;
											assign node3287 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3290 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3293 = (inp[9]) ? node3297 : node3294;
											assign node3294 = (inp[0]) ? 3'b001 : 3'b000;
											assign node3297 = (inp[0]) ? 3'b000 : 3'b001;
								assign node3300 = (inp[7]) ? node3310 : node3301;
									assign node3301 = (inp[9]) ? node3307 : node3302;
										assign node3302 = (inp[2]) ? node3304 : 3'b101;
											assign node3304 = (inp[0]) ? 3'b100 : 3'b101;
										assign node3307 = (inp[0]) ? 3'b101 : 3'b100;
									assign node3310 = (inp[9]) ? node3316 : node3311;
										assign node3311 = (inp[2]) ? node3313 : 3'b100;
											assign node3313 = (inp[0]) ? 3'b101 : 3'b100;
										assign node3316 = (inp[0]) ? node3318 : 3'b101;
											assign node3318 = (inp[2]) ? 3'b100 : 3'b101;
							assign node3321 = (inp[10]) ? node3345 : node3322;
								assign node3322 = (inp[7]) ? node3334 : node3323;
									assign node3323 = (inp[9]) ? node3329 : node3324;
										assign node3324 = (inp[0]) ? node3326 : 3'b101;
											assign node3326 = (inp[2]) ? 3'b100 : 3'b101;
										assign node3329 = (inp[0]) ? node3331 : 3'b100;
											assign node3331 = (inp[2]) ? 3'b101 : 3'b100;
									assign node3334 = (inp[9]) ? node3340 : node3335;
										assign node3335 = (inp[2]) ? node3337 : 3'b100;
											assign node3337 = (inp[0]) ? 3'b101 : 3'b100;
										assign node3340 = (inp[0]) ? node3342 : 3'b101;
											assign node3342 = (inp[2]) ? 3'b100 : 3'b101;
								assign node3345 = (inp[2]) ? node3365 : node3346;
									assign node3346 = (inp[0]) ? node3354 : node3347;
										assign node3347 = (inp[7]) ? node3351 : node3348;
											assign node3348 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3351 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3354 = (inp[1]) ? node3360 : node3355;
											assign node3355 = (inp[9]) ? node3357 : 3'b001;
												assign node3357 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3360 = (inp[7]) ? node3362 : 3'b001;
												assign node3362 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3365 = (inp[7]) ? node3371 : node3366;
										assign node3366 = (inp[0]) ? node3368 : 3'b000;
											assign node3368 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3371 = (inp[0]) ? node3375 : node3372;
											assign node3372 = (inp[9]) ? 3'b001 : 3'b000;
											assign node3375 = (inp[9]) ? 3'b000 : 3'b001;
						assign node3378 = (inp[6]) ? node3426 : node3379;
							assign node3379 = (inp[10]) ? node3403 : node3380;
								assign node3380 = (inp[9]) ? node3392 : node3381;
									assign node3381 = (inp[7]) ? node3387 : node3382;
										assign node3382 = (inp[2]) ? node3384 : 3'b001;
											assign node3384 = (inp[0]) ? 3'b000 : 3'b001;
										assign node3387 = (inp[0]) ? node3389 : 3'b000;
											assign node3389 = (inp[2]) ? 3'b001 : 3'b000;
									assign node3392 = (inp[7]) ? node3398 : node3393;
										assign node3393 = (inp[2]) ? node3395 : 3'b000;
											assign node3395 = (inp[0]) ? 3'b001 : 3'b000;
										assign node3398 = (inp[0]) ? node3400 : 3'b001;
											assign node3400 = (inp[2]) ? 3'b000 : 3'b001;
								assign node3403 = (inp[7]) ? node3415 : node3404;
									assign node3404 = (inp[9]) ? node3410 : node3405;
										assign node3405 = (inp[0]) ? 3'b110 : node3406;
											assign node3406 = (inp[2]) ? 3'b110 : 3'b111;
										assign node3410 = (inp[2]) ? 3'b111 : node3411;
											assign node3411 = (inp[0]) ? 3'b111 : 3'b110;
									assign node3415 = (inp[9]) ? node3421 : node3416;
										assign node3416 = (inp[0]) ? 3'b111 : node3417;
											assign node3417 = (inp[2]) ? 3'b111 : 3'b110;
										assign node3421 = (inp[2]) ? 3'b110 : node3422;
											assign node3422 = (inp[0]) ? 3'b110 : 3'b111;
							assign node3426 = (inp[10]) ? node3450 : node3427;
								assign node3427 = (inp[7]) ? node3439 : node3428;
									assign node3428 = (inp[9]) ? node3434 : node3429;
										assign node3429 = (inp[0]) ? 3'b110 : node3430;
											assign node3430 = (inp[2]) ? 3'b110 : 3'b111;
										assign node3434 = (inp[2]) ? 3'b111 : node3435;
											assign node3435 = (inp[0]) ? 3'b111 : 3'b110;
									assign node3439 = (inp[9]) ? node3445 : node3440;
										assign node3440 = (inp[2]) ? 3'b111 : node3441;
											assign node3441 = (inp[0]) ? 3'b111 : 3'b110;
										assign node3445 = (inp[0]) ? 3'b110 : node3446;
											assign node3446 = (inp[2]) ? 3'b110 : 3'b111;
								assign node3450 = (inp[0]) ? node3474 : node3451;
									assign node3451 = (inp[7]) ? node3459 : node3452;
										assign node3452 = (inp[9]) ? node3456 : node3453;
											assign node3453 = (inp[2]) ? 3'b010 : 3'b011;
											assign node3456 = (inp[2]) ? 3'b011 : 3'b010;
										assign node3459 = (inp[1]) ? node3467 : node3460;
											assign node3460 = (inp[9]) ? node3464 : node3461;
												assign node3461 = (inp[2]) ? 3'b011 : 3'b010;
												assign node3464 = (inp[2]) ? 3'b010 : 3'b011;
											assign node3467 = (inp[9]) ? node3471 : node3468;
												assign node3468 = (inp[2]) ? 3'b011 : 3'b010;
												assign node3471 = (inp[2]) ? 3'b010 : 3'b011;
									assign node3474 = (inp[7]) ? node3478 : node3475;
										assign node3475 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3478 = (inp[9]) ? 3'b010 : 3'b011;
				assign node3481 = (inp[8]) ? node3765 : node3482;
					assign node3482 = (inp[5]) ? node3614 : node3483;
						assign node3483 = (inp[10]) ? node3561 : node3484;
							assign node3484 = (inp[6]) ? node3522 : node3485;
								assign node3485 = (inp[0]) ? node3507 : node3486;
									assign node3486 = (inp[2]) ? node3494 : node3487;
										assign node3487 = (inp[7]) ? node3491 : node3488;
											assign node3488 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3491 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3494 = (inp[1]) ? node3500 : node3495;
											assign node3495 = (inp[9]) ? 3'b001 : node3496;
												assign node3496 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3500 = (inp[7]) ? node3504 : node3501;
												assign node3501 = (inp[9]) ? 3'b000 : 3'b001;
												assign node3504 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3507 = (inp[7]) ? node3515 : node3508;
										assign node3508 = (inp[2]) ? node3512 : node3509;
											assign node3509 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3512 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3515 = (inp[9]) ? node3519 : node3516;
											assign node3516 = (inp[2]) ? 3'b001 : 3'b000;
											assign node3519 = (inp[2]) ? 3'b000 : 3'b001;
								assign node3522 = (inp[1]) ? node3542 : node3523;
									assign node3523 = (inp[9]) ? node3533 : node3524;
										assign node3524 = (inp[7]) ? node3530 : node3525;
											assign node3525 = (inp[2]) ? node3527 : 3'b101;
												assign node3527 = (inp[0]) ? 3'b100 : 3'b101;
											assign node3530 = (inp[2]) ? 3'b101 : 3'b100;
										assign node3533 = (inp[7]) ? node3539 : node3534;
											assign node3534 = (inp[0]) ? node3536 : 3'b100;
												assign node3536 = (inp[2]) ? 3'b101 : 3'b100;
											assign node3539 = (inp[0]) ? 3'b100 : 3'b101;
									assign node3542 = (inp[7]) ? node3550 : node3543;
										assign node3543 = (inp[9]) ? node3545 : 3'b101;
											assign node3545 = (inp[0]) ? node3547 : 3'b100;
												assign node3547 = (inp[2]) ? 3'b101 : 3'b100;
										assign node3550 = (inp[9]) ? node3556 : node3551;
											assign node3551 = (inp[2]) ? node3553 : 3'b100;
												assign node3553 = (inp[0]) ? 3'b101 : 3'b100;
											assign node3556 = (inp[0]) ? node3558 : 3'b101;
												assign node3558 = (inp[2]) ? 3'b100 : 3'b101;
							assign node3561 = (inp[6]) ? node3591 : node3562;
								assign node3562 = (inp[2]) ? node3570 : node3563;
									assign node3563 = (inp[9]) ? node3567 : node3564;
										assign node3564 = (inp[7]) ? 3'b100 : 3'b101;
										assign node3567 = (inp[7]) ? 3'b101 : 3'b100;
									assign node3570 = (inp[0]) ? node3578 : node3571;
										assign node3571 = (inp[9]) ? node3575 : node3572;
											assign node3572 = (inp[7]) ? 3'b100 : 3'b101;
											assign node3575 = (inp[7]) ? 3'b101 : 3'b100;
										assign node3578 = (inp[1]) ? node3584 : node3579;
											assign node3579 = (inp[9]) ? 3'b100 : node3580;
												assign node3580 = (inp[7]) ? 3'b101 : 3'b100;
											assign node3584 = (inp[9]) ? node3588 : node3585;
												assign node3585 = (inp[7]) ? 3'b101 : 3'b100;
												assign node3588 = (inp[7]) ? 3'b100 : 3'b101;
								assign node3591 = (inp[0]) ? node3599 : node3592;
									assign node3592 = (inp[7]) ? node3596 : node3593;
										assign node3593 = (inp[9]) ? 3'b000 : 3'b001;
										assign node3596 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3599 = (inp[2]) ? node3607 : node3600;
										assign node3600 = (inp[7]) ? node3604 : node3601;
											assign node3601 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3604 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3607 = (inp[7]) ? node3611 : node3608;
											assign node3608 = (inp[9]) ? 3'b001 : 3'b000;
											assign node3611 = (inp[9]) ? 3'b000 : 3'b001;
						assign node3614 = (inp[10]) ? node3678 : node3615;
							assign node3615 = (inp[6]) ? node3655 : node3616;
								assign node3616 = (inp[0]) ? node3624 : node3617;
									assign node3617 = (inp[9]) ? node3621 : node3618;
										assign node3618 = (inp[7]) ? 3'b000 : 3'b001;
										assign node3621 = (inp[7]) ? 3'b001 : 3'b000;
									assign node3624 = (inp[9]) ? node3640 : node3625;
										assign node3625 = (inp[1]) ? node3633 : node3626;
											assign node3626 = (inp[2]) ? node3630 : node3627;
												assign node3627 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3630 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3633 = (inp[2]) ? node3637 : node3634;
												assign node3634 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3637 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3640 = (inp[1]) ? node3648 : node3641;
											assign node3641 = (inp[7]) ? node3645 : node3642;
												assign node3642 = (inp[2]) ? 3'b001 : 3'b000;
												assign node3645 = (inp[2]) ? 3'b000 : 3'b001;
											assign node3648 = (inp[2]) ? node3652 : node3649;
												assign node3649 = (inp[7]) ? 3'b001 : 3'b000;
												assign node3652 = (inp[7]) ? 3'b000 : 3'b001;
								assign node3655 = (inp[7]) ? node3667 : node3656;
									assign node3656 = (inp[9]) ? node3662 : node3657;
										assign node3657 = (inp[2]) ? 3'b110 : node3658;
											assign node3658 = (inp[0]) ? 3'b110 : 3'b111;
										assign node3662 = (inp[2]) ? 3'b111 : node3663;
											assign node3663 = (inp[0]) ? 3'b111 : 3'b110;
									assign node3667 = (inp[9]) ? node3673 : node3668;
										assign node3668 = (inp[0]) ? 3'b111 : node3669;
											assign node3669 = (inp[2]) ? 3'b111 : 3'b110;
										assign node3673 = (inp[0]) ? 3'b110 : node3674;
											assign node3674 = (inp[2]) ? 3'b110 : 3'b111;
							assign node3678 = (inp[6]) ? node3732 : node3679;
								assign node3679 = (inp[2]) ? node3709 : node3680;
									assign node3680 = (inp[1]) ? node3696 : node3681;
										assign node3681 = (inp[0]) ? node3689 : node3682;
											assign node3682 = (inp[9]) ? node3686 : node3683;
												assign node3683 = (inp[7]) ? 3'b110 : 3'b111;
												assign node3686 = (inp[7]) ? 3'b111 : 3'b110;
											assign node3689 = (inp[7]) ? node3693 : node3690;
												assign node3690 = (inp[9]) ? 3'b111 : 3'b110;
												assign node3693 = (inp[9]) ? 3'b110 : 3'b111;
										assign node3696 = (inp[9]) ? node3704 : node3697;
											assign node3697 = (inp[7]) ? node3701 : node3698;
												assign node3698 = (inp[0]) ? 3'b110 : 3'b111;
												assign node3701 = (inp[0]) ? 3'b111 : 3'b110;
											assign node3704 = (inp[0]) ? 3'b110 : node3705;
												assign node3705 = (inp[7]) ? 3'b111 : 3'b110;
									assign node3709 = (inp[0]) ? node3717 : node3710;
										assign node3710 = (inp[9]) ? node3714 : node3711;
											assign node3711 = (inp[7]) ? 3'b111 : 3'b110;
											assign node3714 = (inp[7]) ? 3'b110 : 3'b111;
										assign node3717 = (inp[1]) ? node3725 : node3718;
											assign node3718 = (inp[7]) ? node3722 : node3719;
												assign node3719 = (inp[9]) ? 3'b111 : 3'b110;
												assign node3722 = (inp[9]) ? 3'b110 : 3'b111;
											assign node3725 = (inp[9]) ? node3729 : node3726;
												assign node3726 = (inp[7]) ? 3'b111 : 3'b110;
												assign node3729 = (inp[7]) ? 3'b110 : 3'b111;
								assign node3732 = (inp[2]) ? node3758 : node3733;
									assign node3733 = (inp[1]) ? node3749 : node3734;
										assign node3734 = (inp[0]) ? node3742 : node3735;
											assign node3735 = (inp[7]) ? node3739 : node3736;
												assign node3736 = (inp[9]) ? 3'b010 : 3'b011;
												assign node3739 = (inp[9]) ? 3'b011 : 3'b010;
											assign node3742 = (inp[7]) ? node3746 : node3743;
												assign node3743 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3746 = (inp[9]) ? 3'b010 : 3'b011;
										assign node3749 = (inp[0]) ? 3'b011 : node3750;
											assign node3750 = (inp[9]) ? node3754 : node3751;
												assign node3751 = (inp[7]) ? 3'b010 : 3'b011;
												assign node3754 = (inp[7]) ? 3'b011 : 3'b010;
									assign node3758 = (inp[9]) ? node3762 : node3759;
										assign node3759 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3762 = (inp[7]) ? 3'b010 : 3'b011;
					assign node3765 = (inp[5]) ? node3891 : node3766;
						assign node3766 = (inp[7]) ? node3820 : node3767;
							assign node3767 = (inp[9]) ? node3799 : node3768;
								assign node3768 = (inp[0]) ? node3782 : node3769;
									assign node3769 = (inp[2]) ? node3777 : node3770;
										assign node3770 = (inp[6]) ? node3774 : node3771;
											assign node3771 = (inp[10]) ? 3'b111 : 3'b011;
											assign node3774 = (inp[10]) ? 3'b011 : 3'b111;
										assign node3777 = (inp[6]) ? node3779 : 3'b010;
											assign node3779 = (inp[10]) ? 3'b010 : 3'b110;
									assign node3782 = (inp[1]) ? node3792 : node3783;
										assign node3783 = (inp[2]) ? 3'b110 : node3784;
											assign node3784 = (inp[10]) ? node3788 : node3785;
												assign node3785 = (inp[6]) ? 3'b110 : 3'b010;
												assign node3788 = (inp[6]) ? 3'b010 : 3'b110;
										assign node3792 = (inp[6]) ? node3796 : node3793;
											assign node3793 = (inp[10]) ? 3'b110 : 3'b010;
											assign node3796 = (inp[10]) ? 3'b010 : 3'b110;
								assign node3799 = (inp[0]) ? node3813 : node3800;
									assign node3800 = (inp[2]) ? node3808 : node3801;
										assign node3801 = (inp[10]) ? node3805 : node3802;
											assign node3802 = (inp[6]) ? 3'b110 : 3'b010;
											assign node3805 = (inp[6]) ? 3'b010 : 3'b110;
										assign node3808 = (inp[10]) ? 3'b011 : node3809;
											assign node3809 = (inp[6]) ? 3'b111 : 3'b011;
									assign node3813 = (inp[6]) ? node3817 : node3814;
										assign node3814 = (inp[10]) ? 3'b111 : 3'b011;
										assign node3817 = (inp[10]) ? 3'b011 : 3'b111;
							assign node3820 = (inp[9]) ? node3852 : node3821;
								assign node3821 = (inp[2]) ? node3837 : node3822;
									assign node3822 = (inp[0]) ? node3828 : node3823;
										assign node3823 = (inp[10]) ? 3'b110 : node3824;
											assign node3824 = (inp[6]) ? 3'b110 : 3'b010;
										assign node3828 = (inp[1]) ? 3'b011 : node3829;
											assign node3829 = (inp[10]) ? node3833 : node3830;
												assign node3830 = (inp[6]) ? 3'b111 : 3'b011;
												assign node3833 = (inp[6]) ? 3'b011 : 3'b111;
									assign node3837 = (inp[1]) ? node3845 : node3838;
										assign node3838 = (inp[6]) ? node3842 : node3839;
											assign node3839 = (inp[10]) ? 3'b111 : 3'b011;
											assign node3842 = (inp[10]) ? 3'b011 : 3'b111;
										assign node3845 = (inp[10]) ? node3849 : node3846;
											assign node3846 = (inp[6]) ? 3'b111 : 3'b011;
											assign node3849 = (inp[6]) ? 3'b011 : 3'b111;
								assign node3852 = (inp[0]) ? node3874 : node3853;
									assign node3853 = (inp[2]) ? node3861 : node3854;
										assign node3854 = (inp[10]) ? node3858 : node3855;
											assign node3855 = (inp[6]) ? 3'b111 : 3'b011;
											assign node3858 = (inp[6]) ? 3'b011 : 3'b111;
										assign node3861 = (inp[1]) ? node3869 : node3862;
											assign node3862 = (inp[6]) ? node3866 : node3863;
												assign node3863 = (inp[10]) ? 3'b110 : 3'b010;
												assign node3866 = (inp[10]) ? 3'b010 : 3'b110;
											assign node3869 = (inp[6]) ? node3871 : 3'b110;
												assign node3871 = (inp[10]) ? 3'b010 : 3'b110;
									assign node3874 = (inp[2]) ? node3882 : node3875;
										assign node3875 = (inp[10]) ? node3879 : node3876;
											assign node3876 = (inp[6]) ? 3'b110 : 3'b010;
											assign node3879 = (inp[6]) ? 3'b010 : 3'b110;
										assign node3882 = (inp[1]) ? node3886 : node3883;
											assign node3883 = (inp[10]) ? 3'b110 : 3'b010;
											assign node3886 = (inp[10]) ? node3888 : 3'b110;
												assign node3888 = (inp[6]) ? 3'b010 : 3'b110;
						assign node3891 = (inp[10]) ? node3977 : node3892;
							assign node3892 = (inp[6]) ? node3934 : node3893;
								assign node3893 = (inp[1]) ? node3913 : node3894;
									assign node3894 = (inp[2]) ? node3904 : node3895;
										assign node3895 = (inp[0]) ? node3897 : 3'b010;
											assign node3897 = (inp[9]) ? node3901 : node3898;
												assign node3898 = (inp[7]) ? 3'b011 : 3'b010;
												assign node3901 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3904 = (inp[0]) ? 3'b010 : node3905;
											assign node3905 = (inp[7]) ? node3909 : node3906;
												assign node3906 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3909 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3913 = (inp[2]) ? node3927 : node3914;
										assign node3914 = (inp[9]) ? node3922 : node3915;
											assign node3915 = (inp[7]) ? node3919 : node3916;
												assign node3916 = (inp[0]) ? 3'b010 : 3'b011;
												assign node3919 = (inp[0]) ? 3'b011 : 3'b010;
											assign node3922 = (inp[7]) ? node3924 : 3'b010;
												assign node3924 = (inp[0]) ? 3'b010 : 3'b011;
										assign node3927 = (inp[9]) ? node3931 : node3928;
											assign node3928 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3931 = (inp[7]) ? 3'b010 : 3'b011;
								assign node3934 = (inp[1]) ? node3954 : node3935;
									assign node3935 = (inp[9]) ? node3943 : node3936;
										assign node3936 = (inp[7]) ? 3'b101 : node3937;
											assign node3937 = (inp[0]) ? 3'b100 : node3938;
												assign node3938 = (inp[2]) ? 3'b100 : 3'b101;
										assign node3943 = (inp[7]) ? node3949 : node3944;
											assign node3944 = (inp[0]) ? 3'b101 : node3945;
												assign node3945 = (inp[2]) ? 3'b101 : 3'b100;
											assign node3949 = (inp[0]) ? 3'b100 : node3950;
												assign node3950 = (inp[2]) ? 3'b100 : 3'b101;
									assign node3954 = (inp[0]) ? node3970 : node3955;
										assign node3955 = (inp[7]) ? node3963 : node3956;
											assign node3956 = (inp[2]) ? node3960 : node3957;
												assign node3957 = (inp[9]) ? 3'b100 : 3'b101;
												assign node3960 = (inp[9]) ? 3'b101 : 3'b100;
											assign node3963 = (inp[2]) ? node3967 : node3964;
												assign node3964 = (inp[9]) ? 3'b101 : 3'b100;
												assign node3967 = (inp[9]) ? 3'b100 : 3'b101;
										assign node3970 = (inp[9]) ? node3974 : node3971;
											assign node3971 = (inp[7]) ? 3'b101 : 3'b100;
											assign node3974 = (inp[7]) ? 3'b100 : 3'b101;
							assign node3977 = (inp[6]) ? node4001 : node3978;
								assign node3978 = (inp[9]) ? node3990 : node3979;
									assign node3979 = (inp[7]) ? node3985 : node3980;
										assign node3980 = (inp[0]) ? 3'b100 : node3981;
											assign node3981 = (inp[2]) ? 3'b100 : 3'b101;
										assign node3985 = (inp[0]) ? 3'b101 : node3986;
											assign node3986 = (inp[2]) ? 3'b101 : 3'b100;
									assign node3990 = (inp[7]) ? node3996 : node3991;
										assign node3991 = (inp[2]) ? 3'b101 : node3992;
											assign node3992 = (inp[0]) ? 3'b101 : 3'b100;
										assign node3996 = (inp[2]) ? 3'b100 : node3997;
											assign node3997 = (inp[0]) ? 3'b100 : 3'b101;
								assign node4001 = (inp[7]) ? node4013 : node4002;
									assign node4002 = (inp[9]) ? node4008 : node4003;
										assign node4003 = (inp[0]) ? 3'b000 : node4004;
											assign node4004 = (inp[2]) ? 3'b000 : 3'b001;
										assign node4008 = (inp[0]) ? 3'b001 : node4009;
											assign node4009 = (inp[2]) ? 3'b001 : 3'b000;
									assign node4013 = (inp[9]) ? node4019 : node4014;
										assign node4014 = (inp[0]) ? 3'b001 : node4015;
											assign node4015 = (inp[2]) ? 3'b001 : 3'b000;
										assign node4019 = (inp[2]) ? 3'b000 : node4020;
											assign node4020 = (inp[0]) ? 3'b000 : 3'b001;
			assign node4024 = (inp[6]) ? node4490 : node4025;
				assign node4025 = (inp[10]) ? node4299 : node4026;
					assign node4026 = (inp[8]) ? node4152 : node4027;
						assign node4027 = (inp[2]) ? node4071 : node4028;
							assign node4028 = (inp[7]) ? node4052 : node4029;
								assign node4029 = (inp[9]) ? node4039 : node4030;
									assign node4030 = (inp[4]) ? node4034 : node4031;
										assign node4031 = (inp[5]) ? 3'b001 : 3'b011;
										assign node4034 = (inp[5]) ? node4036 : 3'b001;
											assign node4036 = (inp[0]) ? 3'b010 : 3'b011;
									assign node4039 = (inp[0]) ? node4047 : node4040;
										assign node4040 = (inp[4]) ? node4044 : node4041;
											assign node4041 = (inp[5]) ? 3'b000 : 3'b010;
											assign node4044 = (inp[5]) ? 3'b010 : 3'b000;
										assign node4047 = (inp[4]) ? node4049 : 3'b000;
											assign node4049 = (inp[5]) ? 3'b011 : 3'b000;
								assign node4052 = (inp[9]) ? node4062 : node4053;
									assign node4053 = (inp[5]) ? node4057 : node4054;
										assign node4054 = (inp[4]) ? 3'b000 : 3'b010;
										assign node4057 = (inp[4]) ? node4059 : 3'b000;
											assign node4059 = (inp[0]) ? 3'b011 : 3'b010;
									assign node4062 = (inp[5]) ? node4066 : node4063;
										assign node4063 = (inp[4]) ? 3'b001 : 3'b011;
										assign node4066 = (inp[0]) ? 3'b010 : node4067;
											assign node4067 = (inp[4]) ? 3'b011 : 3'b001;
							assign node4071 = (inp[7]) ? node4109 : node4072;
								assign node4072 = (inp[9]) ? node4088 : node4073;
									assign node4073 = (inp[0]) ? node4081 : node4074;
										assign node4074 = (inp[5]) ? node4078 : node4075;
											assign node4075 = (inp[4]) ? 3'b001 : 3'b011;
											assign node4078 = (inp[4]) ? 3'b010 : 3'b001;
										assign node4081 = (inp[4]) ? node4085 : node4082;
											assign node4082 = (inp[5]) ? 3'b000 : 3'b010;
											assign node4085 = (inp[5]) ? 3'b010 : 3'b000;
									assign node4088 = (inp[0]) ? node4096 : node4089;
										assign node4089 = (inp[5]) ? node4093 : node4090;
											assign node4090 = (inp[4]) ? 3'b000 : 3'b010;
											assign node4093 = (inp[4]) ? 3'b011 : 3'b000;
										assign node4096 = (inp[1]) ? node4102 : node4097;
											assign node4097 = (inp[5]) ? node4099 : 3'b011;
												assign node4099 = (inp[4]) ? 3'b011 : 3'b001;
											assign node4102 = (inp[4]) ? node4106 : node4103;
												assign node4103 = (inp[5]) ? 3'b001 : 3'b011;
												assign node4106 = (inp[5]) ? 3'b011 : 3'b001;
								assign node4109 = (inp[9]) ? node4133 : node4110;
									assign node4110 = (inp[0]) ? node4118 : node4111;
										assign node4111 = (inp[5]) ? node4115 : node4112;
											assign node4112 = (inp[4]) ? 3'b000 : 3'b010;
											assign node4115 = (inp[4]) ? 3'b011 : 3'b000;
										assign node4118 = (inp[1]) ? node4126 : node4119;
											assign node4119 = (inp[5]) ? node4123 : node4120;
												assign node4120 = (inp[4]) ? 3'b001 : 3'b011;
												assign node4123 = (inp[4]) ? 3'b011 : 3'b001;
											assign node4126 = (inp[5]) ? node4130 : node4127;
												assign node4127 = (inp[4]) ? 3'b001 : 3'b011;
												assign node4130 = (inp[4]) ? 3'b011 : 3'b001;
									assign node4133 = (inp[0]) ? node4141 : node4134;
										assign node4134 = (inp[4]) ? node4138 : node4135;
											assign node4135 = (inp[5]) ? 3'b001 : 3'b011;
											assign node4138 = (inp[5]) ? 3'b010 : 3'b001;
										assign node4141 = (inp[1]) ? node4147 : node4142;
											assign node4142 = (inp[4]) ? node4144 : 3'b000;
												assign node4144 = (inp[5]) ? 3'b010 : 3'b000;
											assign node4147 = (inp[5]) ? node4149 : 3'b010;
												assign node4149 = (inp[4]) ? 3'b010 : 3'b000;
						assign node4152 = (inp[5]) ? node4214 : node4153;
							assign node4153 = (inp[4]) ? node4177 : node4154;
								assign node4154 = (inp[7]) ? node4166 : node4155;
									assign node4155 = (inp[9]) ? node4161 : node4156;
										assign node4156 = (inp[0]) ? node4158 : 3'b001;
											assign node4158 = (inp[2]) ? 3'b000 : 3'b001;
										assign node4161 = (inp[0]) ? node4163 : 3'b000;
											assign node4163 = (inp[2]) ? 3'b001 : 3'b000;
									assign node4166 = (inp[9]) ? node4172 : node4167;
										assign node4167 = (inp[2]) ? node4169 : 3'b000;
											assign node4169 = (inp[0]) ? 3'b001 : 3'b000;
										assign node4172 = (inp[0]) ? node4174 : 3'b001;
											assign node4174 = (inp[2]) ? 3'b000 : 3'b001;
								assign node4177 = (inp[0]) ? node4193 : node4178;
									assign node4178 = (inp[2]) ? node4186 : node4179;
										assign node4179 = (inp[7]) ? node4183 : node4180;
											assign node4180 = (inp[9]) ? 3'b010 : 3'b011;
											assign node4183 = (inp[9]) ? 3'b011 : 3'b010;
										assign node4186 = (inp[7]) ? node4190 : node4187;
											assign node4187 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4190 = (inp[9]) ? 3'b010 : 3'b011;
									assign node4193 = (inp[2]) ? node4207 : node4194;
										assign node4194 = (inp[1]) ? node4202 : node4195;
											assign node4195 = (inp[9]) ? node4199 : node4196;
												assign node4196 = (inp[7]) ? 3'b011 : 3'b010;
												assign node4199 = (inp[7]) ? 3'b010 : 3'b011;
											assign node4202 = (inp[9]) ? 3'b010 : node4203;
												assign node4203 = (inp[7]) ? 3'b011 : 3'b010;
										assign node4207 = (inp[9]) ? node4211 : node4208;
											assign node4208 = (inp[7]) ? 3'b011 : 3'b010;
											assign node4211 = (inp[7]) ? 3'b010 : 3'b011;
							assign node4214 = (inp[4]) ? node4268 : node4215;
								assign node4215 = (inp[2]) ? node4247 : node4216;
									assign node4216 = (inp[1]) ? node4232 : node4217;
										assign node4217 = (inp[9]) ? node4225 : node4218;
											assign node4218 = (inp[7]) ? node4222 : node4219;
												assign node4219 = (inp[0]) ? 3'b010 : 3'b011;
												assign node4222 = (inp[0]) ? 3'b011 : 3'b010;
											assign node4225 = (inp[7]) ? node4229 : node4226;
												assign node4226 = (inp[0]) ? 3'b011 : 3'b010;
												assign node4229 = (inp[0]) ? 3'b010 : 3'b011;
										assign node4232 = (inp[7]) ? node4240 : node4233;
											assign node4233 = (inp[9]) ? node4237 : node4234;
												assign node4234 = (inp[0]) ? 3'b010 : 3'b011;
												assign node4237 = (inp[0]) ? 3'b011 : 3'b010;
											assign node4240 = (inp[0]) ? node4244 : node4241;
												assign node4241 = (inp[9]) ? 3'b011 : 3'b010;
												assign node4244 = (inp[9]) ? 3'b010 : 3'b011;
									assign node4247 = (inp[1]) ? node4255 : node4248;
										assign node4248 = (inp[7]) ? node4252 : node4249;
											assign node4249 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4252 = (inp[9]) ? 3'b010 : 3'b011;
										assign node4255 = (inp[0]) ? node4263 : node4256;
											assign node4256 = (inp[7]) ? node4260 : node4257;
												assign node4257 = (inp[9]) ? 3'b011 : 3'b010;
												assign node4260 = (inp[9]) ? 3'b010 : 3'b011;
											assign node4263 = (inp[9]) ? 3'b010 : node4264;
												assign node4264 = (inp[7]) ? 3'b011 : 3'b010;
								assign node4268 = (inp[0]) ? node4284 : node4269;
									assign node4269 = (inp[9]) ? node4277 : node4270;
										assign node4270 = (inp[2]) ? node4274 : node4271;
											assign node4271 = (inp[7]) ? 3'b000 : 3'b001;
											assign node4274 = (inp[7]) ? 3'b001 : 3'b000;
										assign node4277 = (inp[7]) ? node4281 : node4278;
											assign node4278 = (inp[2]) ? 3'b001 : 3'b000;
											assign node4281 = (inp[2]) ? 3'b000 : 3'b001;
									assign node4284 = (inp[2]) ? node4292 : node4285;
										assign node4285 = (inp[9]) ? node4289 : node4286;
											assign node4286 = (inp[7]) ? 3'b001 : 3'b000;
											assign node4289 = (inp[7]) ? 3'b000 : 3'b001;
										assign node4292 = (inp[7]) ? node4296 : node4293;
											assign node4293 = (inp[9]) ? 3'b001 : 3'b000;
											assign node4296 = (inp[9]) ? 3'b000 : 3'b001;
					assign node4299 = (inp[0]) ? node4381 : node4300;
						assign node4300 = (inp[9]) ? node4350 : node4301;
							assign node4301 = (inp[7]) ? node4329 : node4302;
								assign node4302 = (inp[2]) ? node4322 : node4303;
									assign node4303 = (inp[1]) ? node4311 : node4304;
										assign node4304 = (inp[8]) ? node4308 : node4305;
											assign node4305 = (inp[4]) ? 3'b111 : 3'b101;
											assign node4308 = (inp[4]) ? 3'b101 : 3'b111;
										assign node4311 = (inp[5]) ? node4317 : node4312;
											assign node4312 = (inp[4]) ? node4314 : 3'b101;
												assign node4314 = (inp[8]) ? 3'b101 : 3'b111;
											assign node4317 = (inp[8]) ? node4319 : 3'b101;
												assign node4319 = (inp[4]) ? 3'b101 : 3'b111;
									assign node4322 = (inp[8]) ? node4326 : node4323;
										assign node4323 = (inp[4]) ? 3'b110 : 3'b101;
										assign node4326 = (inp[4]) ? 3'b100 : 3'b110;
								assign node4329 = (inp[2]) ? node4343 : node4330;
									assign node4330 = (inp[5]) ? node4338 : node4331;
										assign node4331 = (inp[4]) ? node4335 : node4332;
											assign node4332 = (inp[8]) ? 3'b110 : 3'b100;
											assign node4335 = (inp[8]) ? 3'b100 : 3'b110;
										assign node4338 = (inp[4]) ? node4340 : 3'b110;
											assign node4340 = (inp[8]) ? 3'b100 : 3'b110;
									assign node4343 = (inp[4]) ? node4347 : node4344;
										assign node4344 = (inp[8]) ? 3'b111 : 3'b100;
										assign node4347 = (inp[8]) ? 3'b101 : 3'b111;
							assign node4350 = (inp[7]) ? node4366 : node4351;
								assign node4351 = (inp[2]) ? node4359 : node4352;
									assign node4352 = (inp[8]) ? node4356 : node4353;
										assign node4353 = (inp[4]) ? 3'b110 : 3'b100;
										assign node4356 = (inp[4]) ? 3'b100 : 3'b110;
									assign node4359 = (inp[8]) ? node4363 : node4360;
										assign node4360 = (inp[4]) ? 3'b111 : 3'b100;
										assign node4363 = (inp[4]) ? 3'b101 : 3'b111;
								assign node4366 = (inp[2]) ? node4374 : node4367;
									assign node4367 = (inp[4]) ? node4371 : node4368;
										assign node4368 = (inp[8]) ? 3'b111 : 3'b101;
										assign node4371 = (inp[8]) ? 3'b101 : 3'b111;
									assign node4374 = (inp[4]) ? node4378 : node4375;
										assign node4375 = (inp[8]) ? 3'b110 : 3'b101;
										assign node4378 = (inp[8]) ? 3'b100 : 3'b110;
						assign node4381 = (inp[4]) ? node4437 : node4382;
							assign node4382 = (inp[8]) ? node4422 : node4383;
								assign node4383 = (inp[1]) ? node4401 : node4384;
									assign node4384 = (inp[7]) ? node4396 : node4385;
										assign node4385 = (inp[5]) ? node4391 : node4386;
											assign node4386 = (inp[2]) ? 3'b100 : node4387;
												assign node4387 = (inp[9]) ? 3'b100 : 3'b101;
											assign node4391 = (inp[9]) ? node4393 : 3'b100;
												assign node4393 = (inp[2]) ? 3'b101 : 3'b100;
										assign node4396 = (inp[2]) ? node4398 : 3'b101;
											assign node4398 = (inp[9]) ? 3'b100 : 3'b101;
									assign node4401 = (inp[7]) ? node4415 : node4402;
										assign node4402 = (inp[5]) ? node4410 : node4403;
											assign node4403 = (inp[9]) ? node4407 : node4404;
												assign node4404 = (inp[2]) ? 3'b100 : 3'b101;
												assign node4407 = (inp[2]) ? 3'b101 : 3'b100;
											assign node4410 = (inp[9]) ? node4412 : 3'b101;
												assign node4412 = (inp[2]) ? 3'b101 : 3'b100;
										assign node4415 = (inp[2]) ? node4419 : node4416;
											assign node4416 = (inp[9]) ? 3'b101 : 3'b100;
											assign node4419 = (inp[9]) ? 3'b100 : 3'b101;
								assign node4422 = (inp[1]) ? node4430 : node4423;
									assign node4423 = (inp[7]) ? node4427 : node4424;
										assign node4424 = (inp[9]) ? 3'b111 : 3'b110;
										assign node4427 = (inp[9]) ? 3'b110 : 3'b111;
									assign node4430 = (inp[7]) ? node4434 : node4431;
										assign node4431 = (inp[9]) ? 3'b111 : 3'b110;
										assign node4434 = (inp[9]) ? 3'b110 : 3'b111;
							assign node4437 = (inp[8]) ? node4461 : node4438;
								assign node4438 = (inp[5]) ? node4454 : node4439;
									assign node4439 = (inp[1]) ? node4447 : node4440;
										assign node4440 = (inp[9]) ? node4444 : node4441;
											assign node4441 = (inp[7]) ? 3'b111 : 3'b110;
											assign node4444 = (inp[7]) ? 3'b110 : 3'b111;
										assign node4447 = (inp[9]) ? node4451 : node4448;
											assign node4448 = (inp[7]) ? 3'b111 : 3'b110;
											assign node4451 = (inp[7]) ? 3'b110 : 3'b111;
									assign node4454 = (inp[7]) ? node4458 : node4455;
										assign node4455 = (inp[9]) ? 3'b111 : 3'b110;
										assign node4458 = (inp[9]) ? 3'b110 : 3'b111;
								assign node4461 = (inp[5]) ? node4483 : node4462;
									assign node4462 = (inp[2]) ? node4476 : node4463;
										assign node4463 = (inp[1]) ? node4471 : node4464;
											assign node4464 = (inp[9]) ? node4468 : node4465;
												assign node4465 = (inp[7]) ? 3'b101 : 3'b100;
												assign node4468 = (inp[7]) ? 3'b100 : 3'b101;
											assign node4471 = (inp[9]) ? node4473 : 3'b100;
												assign node4473 = (inp[7]) ? 3'b100 : 3'b101;
										assign node4476 = (inp[9]) ? node4480 : node4477;
											assign node4477 = (inp[7]) ? 3'b101 : 3'b100;
											assign node4480 = (inp[7]) ? 3'b100 : 3'b101;
									assign node4483 = (inp[7]) ? node4487 : node4484;
										assign node4484 = (inp[9]) ? 3'b101 : 3'b100;
										assign node4487 = (inp[9]) ? 3'b100 : 3'b101;
				assign node4490 = (inp[10]) ? node4642 : node4491;
					assign node4491 = (inp[9]) ? node4565 : node4492;
						assign node4492 = (inp[7]) ? node4524 : node4493;
							assign node4493 = (inp[2]) ? node4509 : node4494;
								assign node4494 = (inp[0]) ? node4502 : node4495;
									assign node4495 = (inp[8]) ? node4499 : node4496;
										assign node4496 = (inp[4]) ? 3'b111 : 3'b101;
										assign node4499 = (inp[4]) ? 3'b101 : 3'b111;
									assign node4502 = (inp[4]) ? node4506 : node4503;
										assign node4503 = (inp[8]) ? 3'b110 : 3'b101;
										assign node4506 = (inp[8]) ? 3'b100 : 3'b110;
								assign node4509 = (inp[0]) ? node4517 : node4510;
									assign node4510 = (inp[8]) ? node4514 : node4511;
										assign node4511 = (inp[4]) ? 3'b110 : 3'b101;
										assign node4514 = (inp[4]) ? 3'b100 : 3'b110;
									assign node4517 = (inp[4]) ? node4521 : node4518;
										assign node4518 = (inp[8]) ? 3'b110 : 3'b100;
										assign node4521 = (inp[8]) ? 3'b100 : 3'b110;
							assign node4524 = (inp[2]) ? node4556 : node4525;
								assign node4525 = (inp[0]) ? node4549 : node4526;
									assign node4526 = (inp[1]) ? node4534 : node4527;
										assign node4527 = (inp[8]) ? node4531 : node4528;
											assign node4528 = (inp[4]) ? 3'b110 : 3'b100;
											assign node4531 = (inp[4]) ? 3'b100 : 3'b110;
										assign node4534 = (inp[5]) ? node4542 : node4535;
											assign node4535 = (inp[4]) ? node4539 : node4536;
												assign node4536 = (inp[8]) ? 3'b110 : 3'b100;
												assign node4539 = (inp[8]) ? 3'b100 : 3'b110;
											assign node4542 = (inp[4]) ? node4546 : node4543;
												assign node4543 = (inp[8]) ? 3'b110 : 3'b100;
												assign node4546 = (inp[8]) ? 3'b100 : 3'b110;
									assign node4549 = (inp[8]) ? node4553 : node4550;
										assign node4550 = (inp[4]) ? 3'b111 : 3'b100;
										assign node4553 = (inp[4]) ? 3'b101 : 3'b111;
								assign node4556 = (inp[8]) ? node4562 : node4557;
									assign node4557 = (inp[4]) ? 3'b111 : node4558;
										assign node4558 = (inp[0]) ? 3'b101 : 3'b100;
									assign node4562 = (inp[4]) ? 3'b101 : 3'b111;
						assign node4565 = (inp[7]) ? node4603 : node4566;
							assign node4566 = (inp[2]) ? node4588 : node4567;
								assign node4567 = (inp[0]) ? node4581 : node4568;
									assign node4568 = (inp[1]) ? node4574 : node4569;
										assign node4569 = (inp[8]) ? 3'b100 : node4570;
											assign node4570 = (inp[4]) ? 3'b110 : 3'b100;
										assign node4574 = (inp[8]) ? node4578 : node4575;
											assign node4575 = (inp[4]) ? 3'b110 : 3'b100;
											assign node4578 = (inp[4]) ? 3'b100 : 3'b110;
									assign node4581 = (inp[8]) ? node4585 : node4582;
										assign node4582 = (inp[4]) ? 3'b111 : 3'b100;
										assign node4585 = (inp[4]) ? 3'b101 : 3'b111;
								assign node4588 = (inp[0]) ? node4596 : node4589;
									assign node4589 = (inp[8]) ? node4593 : node4590;
										assign node4590 = (inp[4]) ? 3'b111 : 3'b100;
										assign node4593 = (inp[4]) ? 3'b101 : 3'b111;
									assign node4596 = (inp[8]) ? node4600 : node4597;
										assign node4597 = (inp[4]) ? 3'b111 : 3'b101;
										assign node4600 = (inp[4]) ? 3'b101 : 3'b111;
							assign node4603 = (inp[0]) ? node4633 : node4604;
								assign node4604 = (inp[2]) ? node4626 : node4605;
									assign node4605 = (inp[1]) ? node4619 : node4606;
										assign node4606 = (inp[5]) ? node4614 : node4607;
											assign node4607 = (inp[8]) ? node4611 : node4608;
												assign node4608 = (inp[4]) ? 3'b111 : 3'b101;
												assign node4611 = (inp[4]) ? 3'b101 : 3'b111;
											assign node4614 = (inp[8]) ? node4616 : 3'b111;
												assign node4616 = (inp[4]) ? 3'b101 : 3'b111;
										assign node4619 = (inp[8]) ? node4623 : node4620;
											assign node4620 = (inp[4]) ? 3'b111 : 3'b101;
											assign node4623 = (inp[4]) ? 3'b101 : 3'b111;
									assign node4626 = (inp[8]) ? node4630 : node4627;
										assign node4627 = (inp[4]) ? 3'b110 : 3'b101;
										assign node4630 = (inp[4]) ? 3'b100 : 3'b110;
								assign node4633 = (inp[4]) ? node4639 : node4634;
									assign node4634 = (inp[8]) ? 3'b110 : node4635;
										assign node4635 = (inp[2]) ? 3'b100 : 3'b101;
									assign node4639 = (inp[8]) ? 3'b100 : 3'b110;
					assign node4642 = (inp[2]) ? node4722 : node4643;
						assign node4643 = (inp[9]) ? node4683 : node4644;
							assign node4644 = (inp[7]) ? node4660 : node4645;
								assign node4645 = (inp[0]) ? node4653 : node4646;
									assign node4646 = (inp[4]) ? node4650 : node4647;
										assign node4647 = (inp[8]) ? 3'b011 : 3'b001;
										assign node4650 = (inp[8]) ? 3'b001 : 3'b011;
									assign node4653 = (inp[8]) ? node4657 : node4654;
										assign node4654 = (inp[4]) ? 3'b010 : 3'b001;
										assign node4657 = (inp[4]) ? 3'b000 : 3'b010;
								assign node4660 = (inp[0]) ? node4676 : node4661;
									assign node4661 = (inp[1]) ? node4669 : node4662;
										assign node4662 = (inp[4]) ? node4666 : node4663;
											assign node4663 = (inp[8]) ? 3'b010 : 3'b000;
											assign node4666 = (inp[8]) ? 3'b000 : 3'b010;
										assign node4669 = (inp[8]) ? node4673 : node4670;
											assign node4670 = (inp[4]) ? 3'b010 : 3'b000;
											assign node4673 = (inp[4]) ? 3'b000 : 3'b010;
									assign node4676 = (inp[4]) ? node4680 : node4677;
										assign node4677 = (inp[8]) ? 3'b011 : 3'b000;
										assign node4680 = (inp[8]) ? 3'b001 : 3'b011;
							assign node4683 = (inp[7]) ? node4699 : node4684;
								assign node4684 = (inp[0]) ? node4692 : node4685;
									assign node4685 = (inp[8]) ? node4689 : node4686;
										assign node4686 = (inp[4]) ? 3'b010 : 3'b000;
										assign node4689 = (inp[4]) ? 3'b000 : 3'b010;
									assign node4692 = (inp[4]) ? node4696 : node4693;
										assign node4693 = (inp[8]) ? 3'b011 : 3'b000;
										assign node4696 = (inp[8]) ? 3'b001 : 3'b011;
								assign node4699 = (inp[0]) ? node4715 : node4700;
									assign node4700 = (inp[1]) ? node4708 : node4701;
										assign node4701 = (inp[8]) ? node4705 : node4702;
											assign node4702 = (inp[4]) ? 3'b011 : 3'b001;
											assign node4705 = (inp[4]) ? 3'b001 : 3'b011;
										assign node4708 = (inp[8]) ? node4712 : node4709;
											assign node4709 = (inp[4]) ? 3'b011 : 3'b001;
											assign node4712 = (inp[4]) ? 3'b001 : 3'b011;
									assign node4715 = (inp[4]) ? node4719 : node4716;
										assign node4716 = (inp[8]) ? 3'b010 : 3'b001;
										assign node4719 = (inp[8]) ? 3'b000 : 3'b010;
						assign node4722 = (inp[1]) ? node4770 : node4723;
							assign node4723 = (inp[4]) ? node4747 : node4724;
								assign node4724 = (inp[8]) ? node4740 : node4725;
									assign node4725 = (inp[0]) ? node4733 : node4726;
										assign node4726 = (inp[9]) ? node4730 : node4727;
											assign node4727 = (inp[7]) ? 3'b000 : 3'b001;
											assign node4730 = (inp[7]) ? 3'b001 : 3'b000;
										assign node4733 = (inp[9]) ? node4737 : node4734;
											assign node4734 = (inp[7]) ? 3'b001 : 3'b000;
											assign node4737 = (inp[7]) ? 3'b000 : 3'b001;
									assign node4740 = (inp[9]) ? node4744 : node4741;
										assign node4741 = (inp[7]) ? 3'b011 : 3'b010;
										assign node4744 = (inp[7]) ? 3'b010 : 3'b011;
								assign node4747 = (inp[8]) ? node4763 : node4748;
									assign node4748 = (inp[5]) ? node4756 : node4749;
										assign node4749 = (inp[7]) ? node4753 : node4750;
											assign node4750 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4753 = (inp[9]) ? 3'b010 : 3'b011;
										assign node4756 = (inp[7]) ? node4760 : node4757;
											assign node4757 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4760 = (inp[9]) ? 3'b010 : 3'b011;
									assign node4763 = (inp[9]) ? node4767 : node4764;
										assign node4764 = (inp[7]) ? 3'b001 : 3'b000;
										assign node4767 = (inp[7]) ? 3'b000 : 3'b001;
							assign node4770 = (inp[0]) ? node4804 : node4771;
								assign node4771 = (inp[4]) ? node4791 : node4772;
									assign node4772 = (inp[8]) ? node4784 : node4773;
										assign node4773 = (inp[5]) ? node4779 : node4774;
											assign node4774 = (inp[9]) ? node4776 : 3'b001;
												assign node4776 = (inp[7]) ? 3'b001 : 3'b000;
											assign node4779 = (inp[9]) ? 3'b000 : node4780;
												assign node4780 = (inp[7]) ? 3'b000 : 3'b001;
										assign node4784 = (inp[7]) ? node4788 : node4785;
											assign node4785 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4788 = (inp[9]) ? 3'b010 : 3'b011;
									assign node4791 = (inp[8]) ? node4797 : node4792;
										assign node4792 = (inp[9]) ? node4794 : 3'b010;
											assign node4794 = (inp[7]) ? 3'b010 : 3'b011;
										assign node4797 = (inp[9]) ? node4801 : node4798;
											assign node4798 = (inp[7]) ? 3'b001 : 3'b000;
											assign node4801 = (inp[7]) ? 3'b000 : 3'b001;
								assign node4804 = (inp[8]) ? node4820 : node4805;
									assign node4805 = (inp[4]) ? node4813 : node4806;
										assign node4806 = (inp[7]) ? node4810 : node4807;
											assign node4807 = (inp[9]) ? 3'b001 : 3'b000;
											assign node4810 = (inp[9]) ? 3'b000 : 3'b001;
										assign node4813 = (inp[7]) ? node4817 : node4814;
											assign node4814 = (inp[9]) ? 3'b011 : 3'b010;
											assign node4817 = (inp[9]) ? 3'b010 : 3'b011;
									assign node4820 = (inp[4]) ? node4828 : node4821;
										assign node4821 = (inp[9]) ? node4825 : node4822;
											assign node4822 = (inp[7]) ? 3'b011 : 3'b010;
											assign node4825 = (inp[7]) ? 3'b010 : 3'b011;
										assign node4828 = (inp[9]) ? node4832 : node4829;
											assign node4829 = (inp[7]) ? 3'b001 : 3'b000;
											assign node4832 = (inp[7]) ? 3'b000 : 3'b001;

endmodule