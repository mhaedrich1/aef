module dtc_split25_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node11;
	wire [9-1:0] node13;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node32;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node39;
	wire [9-1:0] node41;
	wire [9-1:0] node42;
	wire [9-1:0] node45;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node67;
	wire [9-1:0] node68;
	wire [9-1:0] node69;
	wire [9-1:0] node70;
	wire [9-1:0] node75;
	wire [9-1:0] node76;
	wire [9-1:0] node77;
	wire [9-1:0] node78;
	wire [9-1:0] node79;
	wire [9-1:0] node82;
	wire [9-1:0] node85;
	wire [9-1:0] node89;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node95;
	wire [9-1:0] node98;
	wire [9-1:0] node102;
	wire [9-1:0] node103;
	wire [9-1:0] node104;
	wire [9-1:0] node105;
	wire [9-1:0] node106;
	wire [9-1:0] node107;
	wire [9-1:0] node112;
	wire [9-1:0] node113;
	wire [9-1:0] node114;
	wire [9-1:0] node119;
	wire [9-1:0] node120;
	wire [9-1:0] node121;
	wire [9-1:0] node122;
	wire [9-1:0] node127;
	wire [9-1:0] node128;
	wire [9-1:0] node129;
	wire [9-1:0] node130;
	wire [9-1:0] node131;
	wire [9-1:0] node136;
	wire [9-1:0] node137;
	wire [9-1:0] node138;
	wire [9-1:0] node143;
	wire [9-1:0] node144;
	wire [9-1:0] node145;
	wire [9-1:0] node146;
	wire [9-1:0] node151;
	wire [9-1:0] node152;
	wire [9-1:0] node153;
	wire [9-1:0] node158;
	wire [9-1:0] node159;
	wire [9-1:0] node160;
	wire [9-1:0] node163;
	wire [9-1:0] node165;
	wire [9-1:0] node166;
	wire [9-1:0] node169;
	wire [9-1:0] node172;
	wire [9-1:0] node173;
	wire [9-1:0] node176;
	wire [9-1:0] node178;
	wire [9-1:0] node181;
	wire [9-1:0] node182;
	wire [9-1:0] node183;
	wire [9-1:0] node184;
	wire [9-1:0] node185;
	wire [9-1:0] node186;
	wire [9-1:0] node191;
	wire [9-1:0] node192;
	wire [9-1:0] node193;
	wire [9-1:0] node194;
	wire [9-1:0] node199;
	wire [9-1:0] node202;
	wire [9-1:0] node203;
	wire [9-1:0] node204;
	wire [9-1:0] node205;
	wire [9-1:0] node210;
	wire [9-1:0] node211;
	wire [9-1:0] node212;
	wire [9-1:0] node213;
	wire [9-1:0] node218;
	wire [9-1:0] node221;
	wire [9-1:0] node222;
	wire [9-1:0] node223;
	wire [9-1:0] node224;
	wire [9-1:0] node225;
	wire [9-1:0] node230;
	wire [9-1:0] node231;
	wire [9-1:0] node232;
	wire [9-1:0] node233;
	wire [9-1:0] node238;
	wire [9-1:0] node241;
	wire [9-1:0] node242;
	wire [9-1:0] node243;
	wire [9-1:0] node244;
	wire [9-1:0] node245;
	wire [9-1:0] node246;
	wire [9-1:0] node248;
	wire [9-1:0] node251;
	wire [9-1:0] node255;
	wire [9-1:0] node256;
	wire [9-1:0] node257;
	wire [9-1:0] node258;
	wire [9-1:0] node259;
	wire [9-1:0] node263;
	wire [9-1:0] node264;
	wire [9-1:0] node269;
	wire [9-1:0] node270;
	wire [9-1:0] node274;
	wire [9-1:0] node275;
	wire [9-1:0] node276;
	wire [9-1:0] node278;
	wire [9-1:0] node279;
	wire [9-1:0] node282;
	wire [9-1:0] node285;
	wire [9-1:0] node286;
	wire [9-1:0] node288;
	wire [9-1:0] node290;
	wire [9-1:0] node293;
	wire [9-1:0] node296;
	wire [9-1:0] node297;
	wire [9-1:0] node300;
	wire [9-1:0] node303;
	wire [9-1:0] node304;
	wire [9-1:0] node305;
	wire [9-1:0] node306;
	wire [9-1:0] node307;
	wire [9-1:0] node309;
	wire [9-1:0] node312;
	wire [9-1:0] node313;
	wire [9-1:0] node316;
	wire [9-1:0] node319;
	wire [9-1:0] node320;
	wire [9-1:0] node322;
	wire [9-1:0] node324;
	wire [9-1:0] node327;
	wire [9-1:0] node329;
	wire [9-1:0] node332;
	wire [9-1:0] node333;
	wire [9-1:0] node336;
	wire [9-1:0] node339;
	wire [9-1:0] node340;
	wire [9-1:0] node341;
	wire [9-1:0] node342;
	wire [9-1:0] node344;
	wire [9-1:0] node346;
	wire [9-1:0] node349;
	wire [9-1:0] node352;
	wire [9-1:0] node353;
	wire [9-1:0] node354;
	wire [9-1:0] node358;
	wire [9-1:0] node359;
	wire [9-1:0] node360;
	wire [9-1:0] node365;
	wire [9-1:0] node366;
	wire [9-1:0] node369;
	wire [9-1:0] node372;
	wire [9-1:0] node373;
	wire [9-1:0] node374;
	wire [9-1:0] node375;
	wire [9-1:0] node377;
	wire [9-1:0] node380;
	wire [9-1:0] node381;
	wire [9-1:0] node384;
	wire [9-1:0] node385;
	wire [9-1:0] node388;
	wire [9-1:0] node389;
	wire [9-1:0] node392;
	wire [9-1:0] node395;
	wire [9-1:0] node396;
	wire [9-1:0] node398;
	wire [9-1:0] node401;
	wire [9-1:0] node402;
	wire [9-1:0] node405;
	wire [9-1:0] node406;
	wire [9-1:0] node409;
	wire [9-1:0] node410;
	wire [9-1:0] node413;
	wire [9-1:0] node416;
	wire [9-1:0] node417;
	wire [9-1:0] node418;
	wire [9-1:0] node419;
	wire [9-1:0] node422;
	wire [9-1:0] node424;
	wire [9-1:0] node427;
	wire [9-1:0] node428;
	wire [9-1:0] node431;
	wire [9-1:0] node433;
	wire [9-1:0] node434;
	wire [9-1:0] node437;
	wire [9-1:0] node440;
	wire [9-1:0] node441;
	wire [9-1:0] node442;
	wire [9-1:0] node445;
	wire [9-1:0] node448;
	wire [9-1:0] node449;
	wire [9-1:0] node452;
	wire [9-1:0] node453;
	wire [9-1:0] node454;
	wire [9-1:0] node457;
	wire [9-1:0] node458;
	wire [9-1:0] node461;
	wire [9-1:0] node464;
	wire [9-1:0] node465;
	wire [9-1:0] node468;
	wire [9-1:0] node469;
	wire [9-1:0] node472;

	assign outp = (inp[12]) ? node48 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[9]) ? node11 : 9'b100010001;
							assign node11 = (inp[8]) ? node13 : 9'b100010001;
								assign node13 = (inp[4]) ? 9'b100010001 : node14;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[9]) ? node26 : 9'b101010101;
							assign node26 = (inp[4]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node39 : node30;
						assign node30 = (inp[8]) ? node32 : 9'b111010111;
							assign node32 = (inp[9]) ? node34 : 9'b101010111;
								assign node34 = (inp[4]) ? 9'b111010111 : node35;
									assign node35 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node39 = (inp[8]) ? node41 : 9'b011010111;
							assign node41 = (inp[4]) ? node45 : node42;
								assign node42 = (inp[9]) ? 9'b000010111 : 9'b001010111;
								assign node45 = (inp[9]) ? 9'b001010101 : 9'b001010111;
		assign node48 = (inp[8]) ? node372 : node49;
			assign node49 = (inp[6]) ? node181 : node50;
				assign node50 = (inp[7]) ? node102 : node51;
					assign node51 = (inp[13]) ? node67 : node52;
						assign node52 = (inp[11]) ? node60 : node53;
							assign node53 = (inp[9]) ? 9'b111011000 : node54;
								assign node54 = (inp[1]) ? 9'b111011000 : node55;
									assign node55 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node60 = (inp[9]) ? 9'b111011100 : node61;
								assign node61 = (inp[1]) ? 9'b111011100 : node62;
									assign node62 = (inp[2]) ? 9'b111111100 : 9'b111110100;
						assign node67 = (inp[3]) ? node75 : node68;
							assign node68 = (inp[9]) ? 9'b111011100 : node69;
								assign node69 = (inp[1]) ? 9'b111011100 : node70;
									assign node70 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node75 = (inp[14]) ? node89 : node76;
								assign node76 = (inp[9]) ? 9'b110011110 : node77;
									assign node77 = (inp[1]) ? node85 : node78;
										assign node78 = (inp[2]) ? node82 : node79;
											assign node79 = (inp[10]) ? 9'b110110110 : 9'b110110100;
											assign node82 = (inp[10]) ? 9'b110111110 : 9'b110111100;
										assign node85 = (inp[10]) ? 9'b110011110 : 9'b110011100;
								assign node89 = (inp[9]) ? 9'b111011110 : node90;
									assign node90 = (inp[1]) ? node98 : node91;
										assign node91 = (inp[10]) ? node95 : node92;
											assign node92 = (inp[2]) ? 9'b111111100 : 9'b111110100;
											assign node95 = (inp[2]) ? 9'b111111110 : 9'b111110110;
										assign node98 = (inp[10]) ? 9'b111011110 : 9'b111011100;
					assign node102 = (inp[4]) ? node158 : node103;
						assign node103 = (inp[13]) ? node119 : node104;
							assign node104 = (inp[11]) ? node112 : node105;
								assign node105 = (inp[2]) ? 9'b111111000 : node106;
									assign node106 = (inp[9]) ? 9'b111111000 : node107;
										assign node107 = (inp[1]) ? 9'b111111000 : 9'b111110000;
								assign node112 = (inp[2]) ? 9'b111111100 : node113;
									assign node113 = (inp[9]) ? 9'b111111100 : node114;
										assign node114 = (inp[1]) ? 9'b111111100 : 9'b111110100;
							assign node119 = (inp[3]) ? node127 : node120;
								assign node120 = (inp[1]) ? 9'b111111100 : node121;
									assign node121 = (inp[2]) ? 9'b111111100 : node122;
										assign node122 = (inp[9]) ? 9'b111111100 : 9'b111110100;
								assign node127 = (inp[14]) ? node143 : node128;
									assign node128 = (inp[10]) ? node136 : node129;
										assign node129 = (inp[9]) ? 9'b110111110 : node130;
											assign node130 = (inp[1]) ? 9'b110111100 : node131;
												assign node131 = (inp[2]) ? 9'b110111100 : 9'b110110100;
										assign node136 = (inp[11]) ? 9'b110111110 : node137;
											assign node137 = (inp[2]) ? 9'b110111110 : node138;
												assign node138 = (inp[1]) ? 9'b110111110 : 9'b110110110;
									assign node143 = (inp[10]) ? node151 : node144;
										assign node144 = (inp[9]) ? 9'b111111110 : node145;
											assign node145 = (inp[1]) ? 9'b111111100 : node146;
												assign node146 = (inp[2]) ? 9'b111111100 : 9'b111110100;
										assign node151 = (inp[1]) ? 9'b111111110 : node152;
											assign node152 = (inp[2]) ? 9'b111111110 : node153;
												assign node153 = (inp[5]) ? 9'b111110110 : 9'b111111110;
						assign node158 = (inp[9]) ? node172 : node159;
							assign node159 = (inp[13]) ? node163 : node160;
								assign node160 = (inp[11]) ? 9'b111110100 : 9'b111110000;
								assign node163 = (inp[3]) ? node165 : 9'b111110100;
									assign node165 = (inp[10]) ? node169 : node166;
										assign node166 = (inp[14]) ? 9'b111110100 : 9'b110110100;
										assign node169 = (inp[14]) ? 9'b111110110 : 9'b110110110;
							assign node172 = (inp[13]) ? node176 : node173;
								assign node173 = (inp[11]) ? 9'b111010100 : 9'b111010000;
								assign node176 = (inp[3]) ? node178 : 9'b111010100;
									assign node178 = (inp[14]) ? 9'b111010110 : 9'b110010110;
				assign node181 = (inp[13]) ? node221 : node182;
					assign node182 = (inp[11]) ? node202 : node183;
						assign node183 = (inp[7]) ? node191 : node184;
							assign node184 = (inp[9]) ? 9'b111011000 : node185;
								assign node185 = (inp[1]) ? 9'b111011000 : node186;
									assign node186 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node191 = (inp[4]) ? node199 : node192;
								assign node192 = (inp[1]) ? 9'b111111000 : node193;
									assign node193 = (inp[9]) ? 9'b111111000 : node194;
										assign node194 = (inp[2]) ? 9'b111111000 : 9'b111110000;
								assign node199 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node202 = (inp[7]) ? node210 : node203;
							assign node203 = (inp[1]) ? 9'b111011101 : node204;
								assign node204 = (inp[9]) ? 9'b111011101 : node205;
									assign node205 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node210 = (inp[4]) ? node218 : node211;
								assign node211 = (inp[1]) ? 9'b111111101 : node212;
									assign node212 = (inp[9]) ? 9'b111111101 : node213;
										assign node213 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node218 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node221 = (inp[3]) ? node241 : node222;
						assign node222 = (inp[7]) ? node230 : node223;
							assign node223 = (inp[1]) ? 9'b111011101 : node224;
								assign node224 = (inp[9]) ? 9'b111011101 : node225;
									assign node225 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node230 = (inp[4]) ? node238 : node231;
								assign node231 = (inp[2]) ? 9'b111111101 : node232;
									assign node232 = (inp[9]) ? 9'b111111101 : node233;
										assign node233 = (inp[1]) ? 9'b111111101 : 9'b111110101;
								assign node238 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node241 = (inp[14]) ? node303 : node242;
							assign node242 = (inp[5]) ? node274 : node243;
								assign node243 = (inp[7]) ? node255 : node244;
									assign node244 = (inp[9]) ? 9'b110001111 : node245;
										assign node245 = (inp[1]) ? node251 : node246;
											assign node246 = (inp[2]) ? node248 : 9'b110100101;
												assign node248 = (inp[10]) ? 9'b110101111 : 9'b110101101;
											assign node251 = (inp[10]) ? 9'b110001111 : 9'b110001101;
									assign node255 = (inp[4]) ? node269 : node256;
										assign node256 = (inp[9]) ? 9'b110101111 : node257;
											assign node257 = (inp[10]) ? node263 : node258;
												assign node258 = (inp[1]) ? 9'b110101101 : node259;
													assign node259 = (inp[0]) ? 9'b110100101 : 9'b110101101;
												assign node263 = (inp[1]) ? 9'b110101111 : node264;
													assign node264 = (inp[2]) ? 9'b110101111 : 9'b110100111;
										assign node269 = (inp[9]) ? 9'b110000111 : node270;
											assign node270 = (inp[10]) ? 9'b110100111 : 9'b110100101;
								assign node274 = (inp[9]) ? node296 : node275;
									assign node275 = (inp[10]) ? node285 : node276;
										assign node276 = (inp[11]) ? node278 : 9'b110110101;
											assign node278 = (inp[7]) ? node282 : node279;
												assign node279 = (inp[0]) ? 9'b110011101 : 9'b110111101;
												assign node282 = (inp[4]) ? 9'b110110101 : 9'b110111101;
										assign node285 = (inp[1]) ? node293 : node286;
											assign node286 = (inp[2]) ? node288 : 9'b110110111;
												assign node288 = (inp[7]) ? node290 : 9'b110111111;
													assign node290 = (inp[4]) ? 9'b110110111 : 9'b110111111;
											assign node293 = (inp[7]) ? 9'b110110111 : 9'b110011111;
									assign node296 = (inp[4]) ? node300 : node297;
										assign node297 = (inp[7]) ? 9'b110111111 : 9'b110011111;
										assign node300 = (inp[7]) ? 9'b110010111 : 9'b110011111;
							assign node303 = (inp[5]) ? node339 : node304;
								assign node304 = (inp[9]) ? node332 : node305;
									assign node305 = (inp[10]) ? node319 : node306;
										assign node306 = (inp[2]) ? node312 : node307;
											assign node307 = (inp[1]) ? node309 : 9'b111100101;
												assign node309 = (inp[7]) ? 9'b111100101 : 9'b111001101;
											assign node312 = (inp[7]) ? node316 : node313;
												assign node313 = (inp[1]) ? 9'b111001101 : 9'b111101101;
												assign node316 = (inp[11]) ? 9'b111100101 : 9'b111101101;
										assign node319 = (inp[1]) ? node327 : node320;
											assign node320 = (inp[2]) ? node322 : 9'b111100111;
												assign node322 = (inp[7]) ? node324 : 9'b111101111;
													assign node324 = (inp[4]) ? 9'b111100111 : 9'b111101111;
											assign node327 = (inp[7]) ? node329 : 9'b111001111;
												assign node329 = (inp[4]) ? 9'b111100111 : 9'b111101111;
									assign node332 = (inp[4]) ? node336 : node333;
										assign node333 = (inp[7]) ? 9'b111101111 : 9'b111001111;
										assign node336 = (inp[7]) ? 9'b111000111 : 9'b111001111;
								assign node339 = (inp[9]) ? node365 : node340;
									assign node340 = (inp[10]) ? node352 : node341;
										assign node341 = (inp[1]) ? node349 : node342;
											assign node342 = (inp[2]) ? node344 : 9'b111110101;
												assign node344 = (inp[11]) ? node346 : 9'b111111101;
													assign node346 = (inp[0]) ? 9'b111110101 : 9'b111111101;
											assign node349 = (inp[7]) ? 9'b111111101 : 9'b111011101;
										assign node352 = (inp[7]) ? node358 : node353;
											assign node353 = (inp[1]) ? 9'b111011111 : node354;
												assign node354 = (inp[2]) ? 9'b111111111 : 9'b111110111;
											assign node358 = (inp[4]) ? 9'b111110111 : node359;
												assign node359 = (inp[2]) ? 9'b111111111 : node360;
													assign node360 = (inp[1]) ? 9'b111111111 : 9'b111110111;
									assign node365 = (inp[4]) ? node369 : node366;
										assign node366 = (inp[7]) ? 9'b111111111 : 9'b111011111;
										assign node369 = (inp[7]) ? 9'b111010111 : 9'b111011111;
			assign node372 = (inp[9]) ? node416 : node373;
				assign node373 = (inp[4]) ? node395 : node374;
					assign node374 = (inp[13]) ? node380 : node375;
						assign node375 = (inp[11]) ? node377 : 9'b101111000;
							assign node377 = (inp[6]) ? 9'b101111101 : 9'b101111100;
						assign node380 = (inp[3]) ? node384 : node381;
							assign node381 = (inp[6]) ? 9'b101111101 : 9'b101111100;
							assign node384 = (inp[6]) ? node388 : node385;
								assign node385 = (inp[14]) ? 9'b101111110 : 9'b100111110;
								assign node388 = (inp[14]) ? node392 : node389;
									assign node389 = (inp[5]) ? 9'b100111111 : 9'b100101111;
									assign node392 = (inp[5]) ? 9'b101111111 : 9'b101101111;
					assign node395 = (inp[13]) ? node401 : node396;
						assign node396 = (inp[11]) ? node398 : 9'b101010000;
							assign node398 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node401 = (inp[3]) ? node405 : node402;
							assign node402 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node405 = (inp[6]) ? node409 : node406;
								assign node406 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node409 = (inp[14]) ? node413 : node410;
									assign node410 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node413 = (inp[5]) ? 9'b101010111 : 9'b101000111;
				assign node416 = (inp[6]) ? node440 : node417;
					assign node417 = (inp[4]) ? node427 : node418;
						assign node418 = (inp[13]) ? node422 : node419;
							assign node419 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node422 = (inp[3]) ? node424 : 9'b101010100;
								assign node424 = (inp[0]) ? 9'b100010110 : 9'b111010100;
						assign node427 = (inp[13]) ? node431 : node428;
							assign node428 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node431 = (inp[3]) ? node433 : 9'b111010100;
								assign node433 = (inp[0]) ? node437 : node434;
									assign node434 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node437 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node440 = (inp[13]) ? node448 : node441;
						assign node441 = (inp[11]) ? node445 : node442;
							assign node442 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node445 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node448 = (inp[3]) ? node452 : node449;
							assign node449 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node452 = (inp[0]) ? node464 : node453;
								assign node453 = (inp[4]) ? node457 : node454;
									assign node454 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node457 = (inp[5]) ? node461 : node458;
										assign node458 = (inp[14]) ? 9'b111000111 : 9'b110000111;
										assign node461 = (inp[14]) ? 9'b111010111 : 9'b110010111;
								assign node464 = (inp[4]) ? node468 : node465;
									assign node465 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node468 = (inp[14]) ? node472 : node469;
										assign node469 = (inp[5]) ? 9'b100010101 : 9'b100000101;
										assign node472 = (inp[5]) ? 9'b101010101 : 9'b101000101;

endmodule