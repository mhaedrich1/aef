module dtc_split66_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node505;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node705;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node745;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node764;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node786;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node974;

	assign outp = (inp[3]) ? node718 : node1;
		assign node1 = (inp[9]) ? node303 : node2;
			assign node2 = (inp[1]) ? node94 : node3;
				assign node3 = (inp[4]) ? node41 : node4;
					assign node4 = (inp[6]) ? node20 : node5;
						assign node5 = (inp[5]) ? node15 : node6;
							assign node6 = (inp[0]) ? node8 : 3'b001;
								assign node8 = (inp[8]) ? 3'b000 : node9;
									assign node9 = (inp[7]) ? 3'b000 : node10;
										assign node10 = (inp[2]) ? 3'b000 : 3'b001;
							assign node15 = (inp[0]) ? 3'b001 : node16;
								assign node16 = (inp[7]) ? 3'b001 : 3'b000;
						assign node20 = (inp[5]) ? node28 : node21;
							assign node21 = (inp[0]) ? node23 : 3'b000;
								assign node23 = (inp[10]) ? node25 : 3'b000;
									assign node25 = (inp[7]) ? 3'b001 : 3'b000;
							assign node28 = (inp[0]) ? node34 : node29;
								assign node29 = (inp[7]) ? node31 : 3'b001;
									assign node31 = (inp[8]) ? 3'b000 : 3'b001;
								assign node34 = (inp[10]) ? node36 : 3'b000;
									assign node36 = (inp[2]) ? node38 : 3'b000;
										assign node38 = (inp[7]) ? 3'b001 : 3'b000;
					assign node41 = (inp[6]) ? node61 : node42;
						assign node42 = (inp[0]) ? node44 : 3'b000;
							assign node44 = (inp[5]) ? node52 : node45;
								assign node45 = (inp[2]) ? 3'b001 : node46;
									assign node46 = (inp[7]) ? 3'b001 : node47;
										assign node47 = (inp[8]) ? 3'b001 : 3'b000;
								assign node52 = (inp[7]) ? 3'b000 : node53;
									assign node53 = (inp[11]) ? 3'b000 : node54;
										assign node54 = (inp[2]) ? 3'b000 : node55;
											assign node55 = (inp[8]) ? 3'b001 : 3'b000;
						assign node61 = (inp[5]) ? node75 : node62;
							assign node62 = (inp[0]) ? 3'b000 : node63;
								assign node63 = (inp[8]) ? node69 : node64;
									assign node64 = (inp[7]) ? node66 : 3'b000;
										assign node66 = (inp[10]) ? 3'b001 : 3'b000;
									assign node69 = (inp[10]) ? 3'b001 : node70;
										assign node70 = (inp[7]) ? 3'b000 : 3'b001;
							assign node75 = (inp[0]) ? 3'b001 : node76;
								assign node76 = (inp[10]) ? node82 : node77;
									assign node77 = (inp[8]) ? node79 : 3'b000;
										assign node79 = (inp[11]) ? 3'b000 : 3'b001;
									assign node82 = (inp[8]) ? node88 : node83;
										assign node83 = (inp[2]) ? node85 : 3'b000;
											assign node85 = (inp[7]) ? 3'b001 : 3'b000;
										assign node88 = (inp[7]) ? 3'b001 : node89;
											assign node89 = (inp[11]) ? 3'b000 : 3'b001;
				assign node94 = (inp[6]) ? node208 : node95;
					assign node95 = (inp[5]) ? node149 : node96;
						assign node96 = (inp[7]) ? node118 : node97;
							assign node97 = (inp[0]) ? node113 : node98;
								assign node98 = (inp[4]) ? node106 : node99;
									assign node99 = (inp[10]) ? 3'b001 : node100;
										assign node100 = (inp[2]) ? node102 : 3'b000;
											assign node102 = (inp[8]) ? 3'b000 : 3'b001;
									assign node106 = (inp[2]) ? node108 : 3'b001;
										assign node108 = (inp[8]) ? node110 : 3'b000;
											assign node110 = (inp[10]) ? 3'b000 : 3'b001;
								assign node113 = (inp[4]) ? node115 : 3'b000;
									assign node115 = (inp[8]) ? 3'b000 : 3'b001;
							assign node118 = (inp[8]) ? node138 : node119;
								assign node119 = (inp[2]) ? node129 : node120;
									assign node120 = (inp[4]) ? node124 : node121;
										assign node121 = (inp[10]) ? 3'b001 : 3'b000;
										assign node124 = (inp[10]) ? node126 : 3'b001;
											assign node126 = (inp[0]) ? 3'b001 : 3'b000;
									assign node129 = (inp[11]) ? 3'b000 : node130;
										assign node130 = (inp[10]) ? 3'b001 : node131;
											assign node131 = (inp[0]) ? 3'b000 : node132;
												assign node132 = (inp[4]) ? 3'b000 : 3'b001;
								assign node138 = (inp[0]) ? 3'b001 : node139;
									assign node139 = (inp[4]) ? node145 : node140;
										assign node140 = (inp[10]) ? 3'b000 : node141;
											assign node141 = (inp[2]) ? 3'b000 : 3'b001;
										assign node145 = (inp[2]) ? 3'b001 : 3'b000;
						assign node149 = (inp[0]) ? node193 : node150;
							assign node150 = (inp[4]) ? node174 : node151;
								assign node151 = (inp[11]) ? node167 : node152;
									assign node152 = (inp[7]) ? node158 : node153;
										assign node153 = (inp[2]) ? node155 : 3'b001;
											assign node155 = (inp[10]) ? 3'b001 : 3'b000;
										assign node158 = (inp[8]) ? 3'b000 : node159;
											assign node159 = (inp[2]) ? node163 : node160;
												assign node160 = (inp[10]) ? 3'b001 : 3'b000;
												assign node163 = (inp[10]) ? 3'b000 : 3'b001;
									assign node167 = (inp[10]) ? 3'b001 : node168;
										assign node168 = (inp[8]) ? 3'b001 : node169;
											assign node169 = (inp[7]) ? 3'b000 : 3'b001;
								assign node174 = (inp[7]) ? node184 : node175;
									assign node175 = (inp[11]) ? 3'b000 : node176;
										assign node176 = (inp[8]) ? node178 : 3'b000;
											assign node178 = (inp[2]) ? node180 : 3'b000;
												assign node180 = (inp[10]) ? 3'b000 : 3'b001;
									assign node184 = (inp[10]) ? node188 : node185;
										assign node185 = (inp[11]) ? 3'b001 : 3'b000;
										assign node188 = (inp[11]) ? 3'b000 : node189;
											assign node189 = (inp[2]) ? 3'b001 : 3'b000;
							assign node193 = (inp[7]) ? node201 : node194;
								assign node194 = (inp[11]) ? node196 : 3'b001;
									assign node196 = (inp[4]) ? node198 : 3'b001;
										assign node198 = (inp[8]) ? 3'b001 : 3'b000;
								assign node201 = (inp[4]) ? 3'b001 : node202;
									assign node202 = (inp[8]) ? node204 : 3'b000;
										assign node204 = (inp[11]) ? 3'b000 : 3'b001;
					assign node208 = (inp[5]) ? node236 : node209;
						assign node209 = (inp[4]) ? node227 : node210;
							assign node210 = (inp[0]) ? 3'b001 : node211;
								assign node211 = (inp[7]) ? node217 : node212;
									assign node212 = (inp[10]) ? 3'b000 : node213;
										assign node213 = (inp[8]) ? 3'b001 : 3'b000;
									assign node217 = (inp[10]) ? node221 : node218;
										assign node218 = (inp[8]) ? 3'b000 : 3'b001;
										assign node221 = (inp[8]) ? 3'b001 : node222;
											assign node222 = (inp[2]) ? 3'b000 : 3'b001;
							assign node227 = (inp[0]) ? 3'b000 : node228;
								assign node228 = (inp[8]) ? node230 : 3'b001;
									assign node230 = (inp[2]) ? node232 : 3'b001;
										assign node232 = (inp[7]) ? 3'b000 : 3'b001;
						assign node236 = (inp[4]) ? node256 : node237;
							assign node237 = (inp[8]) ? node245 : node238;
								assign node238 = (inp[0]) ? 3'b000 : node239;
									assign node239 = (inp[7]) ? node241 : 3'b000;
										assign node241 = (inp[11]) ? 3'b000 : 3'b001;
								assign node245 = (inp[0]) ? 3'b001 : node246;
									assign node246 = (inp[10]) ? 3'b000 : node247;
										assign node247 = (inp[7]) ? node249 : 3'b000;
											assign node249 = (inp[2]) ? node251 : 3'b001;
												assign node251 = (inp[11]) ? 3'b001 : 3'b000;
							assign node256 = (inp[11]) ? node264 : node257;
								assign node257 = (inp[7]) ? node261 : node258;
									assign node258 = (inp[0]) ? 3'b001 : 3'b000;
									assign node261 = (inp[0]) ? 3'b000 : 3'b001;
								assign node264 = (inp[8]) ? node280 : node265;
									assign node265 = (inp[10]) ? node273 : node266;
										assign node266 = (inp[7]) ? node270 : node267;
											assign node267 = (inp[0]) ? 3'b001 : 3'b000;
											assign node270 = (inp[0]) ? 3'b000 : 3'b001;
										assign node273 = (inp[0]) ? node277 : node274;
											assign node274 = (inp[7]) ? 3'b001 : 3'b000;
											assign node277 = (inp[7]) ? 3'b000 : 3'b001;
									assign node280 = (inp[10]) ? node290 : node281;
										assign node281 = (inp[2]) ? node283 : 3'b000;
											assign node283 = (inp[7]) ? node287 : node284;
												assign node284 = (inp[0]) ? 3'b001 : 3'b000;
												assign node287 = (inp[0]) ? 3'b000 : 3'b001;
										assign node290 = (inp[2]) ? node298 : node291;
											assign node291 = (inp[0]) ? node295 : node292;
												assign node292 = (inp[7]) ? 3'b001 : 3'b000;
												assign node295 = (inp[7]) ? 3'b000 : 3'b001;
											assign node298 = (inp[0]) ? 3'b000 : node299;
												assign node299 = (inp[7]) ? 3'b001 : 3'b000;
			assign node303 = (inp[4]) ? node533 : node304;
				assign node304 = (inp[6]) ? node414 : node305;
					assign node305 = (inp[0]) ? node359 : node306;
						assign node306 = (inp[1]) ? node314 : node307;
							assign node307 = (inp[5]) ? node311 : node308;
								assign node308 = (inp[7]) ? 3'b110 : 3'b010;
								assign node311 = (inp[7]) ? 3'b010 : 3'b100;
							assign node314 = (inp[5]) ? node336 : node315;
								assign node315 = (inp[7]) ? node323 : node316;
									assign node316 = (inp[10]) ? 3'b110 : node317;
										assign node317 = (inp[8]) ? 3'b101 : node318;
											assign node318 = (inp[2]) ? 3'b110 : 3'b101;
									assign node323 = (inp[2]) ? node331 : node324;
										assign node324 = (inp[11]) ? node326 : 3'b001;
											assign node326 = (inp[8]) ? 3'b010 : node327;
												assign node327 = (inp[10]) ? 3'b110 : 3'b101;
										assign node331 = (inp[8]) ? 3'b001 : node332;
											assign node332 = (inp[10]) ? 3'b001 : 3'b010;
								assign node336 = (inp[7]) ? node346 : node337;
									assign node337 = (inp[8]) ? node339 : 3'b010;
										assign node339 = (inp[11]) ? 3'b010 : node340;
											assign node340 = (inp[10]) ? 3'b010 : node341;
												assign node341 = (inp[2]) ? 3'b001 : 3'b010;
									assign node346 = (inp[8]) ? node352 : node347;
										assign node347 = (inp[2]) ? 3'b110 : node348;
											assign node348 = (inp[10]) ? 3'b010 : 3'b001;
										assign node352 = (inp[11]) ? node354 : 3'b101;
											assign node354 = (inp[10]) ? 3'b110 : node355;
												assign node355 = (inp[2]) ? 3'b110 : 3'b101;
						assign node359 = (inp[5]) ? node385 : node360;
							assign node360 = (inp[7]) ? node376 : node361;
								assign node361 = (inp[1]) ? node369 : node362;
									assign node362 = (inp[2]) ? 3'b001 : node363;
										assign node363 = (inp[8]) ? 3'b001 : node364;
											assign node364 = (inp[11]) ? 3'b110 : 3'b010;
									assign node369 = (inp[8]) ? node373 : node370;
										assign node370 = (inp[11]) ? 3'b001 : 3'b101;
										assign node373 = (inp[11]) ? 3'b000 : 3'b100;
								assign node376 = (inp[8]) ? node382 : node377;
									assign node377 = (inp[2]) ? 3'b101 : node378;
										assign node378 = (inp[1]) ? 3'b101 : 3'b001;
									assign node382 = (inp[1]) ? 3'b011 : 3'b001;
							assign node385 = (inp[1]) ? node401 : node386;
								assign node386 = (inp[8]) ? node392 : node387;
									assign node387 = (inp[7]) ? 3'b110 : node388;
										assign node388 = (inp[2]) ? 3'b110 : 3'b010;
									assign node392 = (inp[2]) ? node398 : node393;
										assign node393 = (inp[7]) ? 3'b110 : node394;
											assign node394 = (inp[11]) ? 3'b110 : 3'b101;
										assign node398 = (inp[7]) ? 3'b010 : 3'b110;
								assign node401 = (inp[7]) ? node407 : node402;
									assign node402 = (inp[11]) ? node404 : 3'b111;
										assign node404 = (inp[8]) ? 3'b111 : 3'b110;
									assign node407 = (inp[11]) ? node411 : node408;
										assign node408 = (inp[8]) ? 3'b111 : 3'b101;
										assign node411 = (inp[8]) ? 3'b101 : 3'b001;
					assign node414 = (inp[1]) ? node464 : node415;
						assign node415 = (inp[7]) ? node433 : node416;
							assign node416 = (inp[5]) ? node422 : node417;
								assign node417 = (inp[10]) ? node419 : 3'b101;
									assign node419 = (inp[0]) ? 3'b101 : 3'b001;
								assign node422 = (inp[0]) ? 3'b101 : node423;
									assign node423 = (inp[11]) ? node425 : 3'b110;
										assign node425 = (inp[8]) ? 3'b110 : node426;
											assign node426 = (inp[2]) ? 3'b110 : node427;
												assign node427 = (inp[10]) ? 3'b010 : 3'b110;
							assign node433 = (inp[10]) ? node447 : node434;
								assign node434 = (inp[0]) ? node440 : node435;
									assign node435 = (inp[8]) ? 3'b001 : node436;
										assign node436 = (inp[5]) ? 3'b010 : 3'b001;
									assign node440 = (inp[8]) ? 3'b101 : node441;
										assign node441 = (inp[2]) ? 3'b001 : node442;
											assign node442 = (inp[11]) ? 3'b101 : 3'b001;
								assign node447 = (inp[0]) ? node455 : node448;
									assign node448 = (inp[5]) ? node450 : 3'b101;
										assign node450 = (inp[8]) ? 3'b001 : node451;
											assign node451 = (inp[2]) ? 3'b010 : 3'b110;
									assign node455 = (inp[2]) ? node459 : node456;
										assign node456 = (inp[5]) ? 3'b101 : 3'b011;
										assign node459 = (inp[8]) ? node461 : 3'b011;
											assign node461 = (inp[5]) ? 3'b011 : 3'b111;
						assign node464 = (inp[5]) ? node496 : node465;
							assign node465 = (inp[0]) ? node487 : node466;
								assign node466 = (inp[10]) ? node476 : node467;
									assign node467 = (inp[7]) ? node473 : node468;
										assign node468 = (inp[2]) ? node470 : 3'b011;
											assign node470 = (inp[8]) ? 3'b011 : 3'b001;
										assign node473 = (inp[8]) ? 3'b001 : 3'b011;
									assign node476 = (inp[7]) ? node482 : node477;
										assign node477 = (inp[2]) ? 3'b101 : node478;
											assign node478 = (inp[8]) ? 3'b101 : 3'b001;
										assign node482 = (inp[8]) ? 3'b011 : node483;
											assign node483 = (inp[2]) ? 3'b001 : 3'b011;
								assign node487 = (inp[7]) ? 3'b111 : node488;
									assign node488 = (inp[10]) ? node490 : 3'b011;
										assign node490 = (inp[8]) ? node492 : 3'b011;
											assign node492 = (inp[2]) ? 3'b111 : 3'b011;
							assign node496 = (inp[8]) ? node516 : node497;
								assign node497 = (inp[10]) ? node505 : node498;
									assign node498 = (inp[7]) ? node500 : 3'b001;
										assign node500 = (inp[0]) ? 3'b001 : node501;
											assign node501 = (inp[11]) ? 3'b001 : 3'b011;
									assign node505 = (inp[2]) ? node507 : 3'b001;
										assign node507 = (inp[11]) ? node511 : node508;
											assign node508 = (inp[7]) ? 3'b101 : 3'b001;
											assign node511 = (inp[7]) ? node513 : 3'b101;
												assign node513 = (inp[0]) ? 3'b001 : 3'b101;
								assign node516 = (inp[0]) ? 3'b011 : node517;
									assign node517 = (inp[10]) ? node529 : node518;
										assign node518 = (inp[7]) ? node524 : node519;
											assign node519 = (inp[11]) ? 3'b001 : node520;
												assign node520 = (inp[2]) ? 3'b011 : 3'b001;
											assign node524 = (inp[2]) ? node526 : 3'b011;
												assign node526 = (inp[11]) ? 3'b011 : 3'b001;
										assign node529 = (inp[7]) ? 3'b101 : 3'b001;
				assign node533 = (inp[6]) ? node631 : node534;
					assign node534 = (inp[0]) ? node598 : node535;
						assign node535 = (inp[5]) ? node569 : node536;
							assign node536 = (inp[1]) ? node544 : node537;
								assign node537 = (inp[7]) ? 3'b100 : node538;
									assign node538 = (inp[10]) ? node540 : 3'b100;
										assign node540 = (inp[11]) ? 3'b000 : 3'b100;
								assign node544 = (inp[7]) ? node556 : node545;
									assign node545 = (inp[2]) ? node551 : node546;
										assign node546 = (inp[8]) ? 3'b110 : node547;
											assign node547 = (inp[10]) ? 3'b000 : 3'b010;
										assign node551 = (inp[8]) ? node553 : 3'b100;
											assign node553 = (inp[10]) ? 3'b100 : 3'b110;
									assign node556 = (inp[11]) ? 3'b010 : node557;
										assign node557 = (inp[10]) ? node563 : node558;
											assign node558 = (inp[2]) ? 3'b000 : node559;
												assign node559 = (inp[8]) ? 3'b000 : 3'b010;
											assign node563 = (inp[2]) ? 3'b010 : node564;
												assign node564 = (inp[8]) ? 3'b010 : 3'b000;
							assign node569 = (inp[1]) ? node571 : 3'b000;
								assign node571 = (inp[7]) ? node583 : node572;
									assign node572 = (inp[8]) ? node574 : 3'b000;
										assign node574 = (inp[2]) ? node578 : node575;
											assign node575 = (inp[11]) ? 3'b000 : 3'b100;
											assign node578 = (inp[10]) ? 3'b000 : node579;
												assign node579 = (inp[11]) ? 3'b000 : 3'b010;
									assign node583 = (inp[8]) ? node591 : node584;
										assign node584 = (inp[2]) ? node588 : node585;
											assign node585 = (inp[10]) ? 3'b000 : 3'b010;
											assign node588 = (inp[11]) ? 3'b110 : 3'b100;
										assign node591 = (inp[10]) ? node595 : node592;
											assign node592 = (inp[2]) ? 3'b100 : 3'b110;
											assign node595 = (inp[11]) ? 3'b100 : 3'b110;
						assign node598 = (inp[5]) ? node614 : node599;
							assign node599 = (inp[1]) ? node609 : node600;
								assign node600 = (inp[7]) ? 3'b010 : node601;
									assign node601 = (inp[2]) ? 3'b010 : node602;
										assign node602 = (inp[8]) ? 3'b010 : node603;
											assign node603 = (inp[11]) ? 3'b100 : 3'b000;
								assign node609 = (inp[7]) ? 3'b110 : node610;
									assign node610 = (inp[8]) ? 3'b100 : 3'b010;
							assign node614 = (inp[1]) ? node624 : node615;
								assign node615 = (inp[7]) ? 3'b100 : node616;
									assign node616 = (inp[8]) ? node620 : node617;
										assign node617 = (inp[2]) ? 3'b100 : 3'b000;
										assign node620 = (inp[2]) ? 3'b100 : 3'b110;
								assign node624 = (inp[11]) ? node626 : 3'b010;
									assign node626 = (inp[7]) ? 3'b010 : node627;
										assign node627 = (inp[8]) ? 3'b010 : 3'b100;
					assign node631 = (inp[0]) ? node699 : node632;
						assign node632 = (inp[8]) ? node656 : node633;
							assign node633 = (inp[7]) ? node639 : node634;
								assign node634 = (inp[1]) ? node636 : 3'b100;
									assign node636 = (inp[5]) ? 3'b100 : 3'b110;
								assign node639 = (inp[1]) ? node649 : node640;
									assign node640 = (inp[10]) ? node644 : node641;
										assign node641 = (inp[5]) ? 3'b100 : 3'b000;
										assign node644 = (inp[5]) ? node646 : 3'b010;
											assign node646 = (inp[2]) ? 3'b010 : 3'b000;
									assign node649 = (inp[5]) ? node651 : 3'b110;
										assign node651 = (inp[2]) ? node653 : 3'b010;
											assign node653 = (inp[11]) ? 3'b101 : 3'b110;
							assign node656 = (inp[10]) ? node674 : node657;
								assign node657 = (inp[7]) ? node665 : node658;
									assign node658 = (inp[5]) ? node660 : 3'b010;
										assign node660 = (inp[11]) ? 3'b100 : node661;
											assign node661 = (inp[1]) ? 3'b100 : 3'b010;
									assign node665 = (inp[5]) ? node671 : node666;
										assign node666 = (inp[1]) ? node668 : 3'b100;
											assign node668 = (inp[2]) ? 3'b001 : 3'b110;
										assign node671 = (inp[1]) ? 3'b010 : 3'b000;
								assign node674 = (inp[1]) ? node686 : node675;
									assign node675 = (inp[11]) ? node677 : 3'b010;
										assign node677 = (inp[2]) ? node681 : node678;
											assign node678 = (inp[5]) ? 3'b100 : 3'b010;
											assign node681 = (inp[5]) ? 3'b010 : node682;
												assign node682 = (inp[7]) ? 3'b110 : 3'b010;
									assign node686 = (inp[7]) ? node690 : node687;
										assign node687 = (inp[5]) ? 3'b100 : 3'b110;
										assign node690 = (inp[5]) ? node694 : node691;
											assign node691 = (inp[2]) ? 3'b001 : 3'b110;
											assign node694 = (inp[2]) ? node696 : 3'b010;
												assign node696 = (inp[11]) ? 3'b110 : 3'b010;
						assign node699 = (inp[5]) ? node709 : node700;
							assign node700 = (inp[7]) ? node702 : 3'b001;
								assign node702 = (inp[1]) ? 3'b101 : node703;
									assign node703 = (inp[10]) ? node705 : 3'b001;
										assign node705 = (inp[2]) ? 3'b101 : 3'b001;
							assign node709 = (inp[7]) ? node713 : node710;
								assign node710 = (inp[1]) ? 3'b110 : 3'b010;
								assign node713 = (inp[1]) ? 3'b001 : node714;
									assign node714 = (inp[10]) ? 3'b110 : 3'b010;
		assign node718 = (inp[6]) ? node740 : node719;
			assign node719 = (inp[0]) ? node721 : 3'b000;
				assign node721 = (inp[9]) ? node723 : 3'b000;
					assign node723 = (inp[1]) ? node725 : 3'b000;
						assign node725 = (inp[4]) ? 3'b000 : node726;
							assign node726 = (inp[5]) ? node732 : node727;
								assign node727 = (inp[8]) ? 3'b100 : node728;
									assign node728 = (inp[7]) ? 3'b100 : 3'b000;
								assign node732 = (inp[11]) ? 3'b000 : node733;
									assign node733 = (inp[7]) ? 3'b000 : node734;
										assign node734 = (inp[8]) ? 3'b100 : 3'b000;
			assign node740 = (inp[9]) ? node892 : node741;
				assign node741 = (inp[4]) ? node771 : node742;
					assign node742 = (inp[0]) ? node764 : node743;
						assign node743 = (inp[2]) ? node745 : 3'b010;
							assign node745 = (inp[7]) ? node747 : 3'b010;
								assign node747 = (inp[1]) ? node749 : 3'b010;
									assign node749 = (inp[11]) ? node755 : node750;
										assign node750 = (inp[8]) ? node752 : 3'b010;
											assign node752 = (inp[5]) ? 3'b010 : 3'b011;
										assign node755 = (inp[10]) ? 3'b011 : node756;
											assign node756 = (inp[5]) ? node760 : node757;
												assign node757 = (inp[8]) ? 3'b011 : 3'b010;
												assign node760 = (inp[8]) ? 3'b010 : 3'b011;
						assign node764 = (inp[5]) ? node766 : 3'b011;
							assign node766 = (inp[1]) ? node768 : 3'b010;
								assign node768 = (inp[7]) ? 3'b011 : 3'b010;
					assign node771 = (inp[0]) ? node823 : node772;
						assign node772 = (inp[10]) ? node806 : node773;
							assign node773 = (inp[5]) ? node791 : node774;
								assign node774 = (inp[7]) ? node778 : node775;
									assign node775 = (inp[1]) ? 3'b000 : 3'b010;
									assign node778 = (inp[11]) ? node780 : 3'b010;
										assign node780 = (inp[2]) ? node786 : node781;
											assign node781 = (inp[1]) ? 3'b010 : node782;
												assign node782 = (inp[8]) ? 3'b010 : 3'b110;
											assign node786 = (inp[1]) ? node788 : 3'b010;
												assign node788 = (inp[8]) ? 3'b100 : 3'b010;
								assign node791 = (inp[7]) ? node797 : node792;
									assign node792 = (inp[1]) ? node794 : 3'b000;
										assign node794 = (inp[11]) ? 3'b100 : 3'b000;
									assign node797 = (inp[11]) ? 3'b100 : node798;
										assign node798 = (inp[1]) ? 3'b010 : node799;
											assign node799 = (inp[8]) ? node801 : 3'b100;
												assign node801 = (inp[2]) ? 3'b010 : 3'b000;
							assign node806 = (inp[1]) ? node808 : 3'b000;
								assign node808 = (inp[5]) ? node816 : node809;
									assign node809 = (inp[8]) ? 3'b000 : node810;
										assign node810 = (inp[11]) ? node812 : 3'b000;
											assign node812 = (inp[2]) ? 3'b000 : 3'b100;
									assign node816 = (inp[8]) ? 3'b100 : node817;
										assign node817 = (inp[11]) ? node819 : 3'b000;
											assign node819 = (inp[7]) ? 3'b000 : 3'b100;
						assign node823 = (inp[7]) ? node855 : node824;
							assign node824 = (inp[10]) ? node846 : node825;
								assign node825 = (inp[1]) ? node837 : node826;
									assign node826 = (inp[11]) ? node832 : node827;
										assign node827 = (inp[8]) ? 3'b010 : node828;
											assign node828 = (inp[2]) ? 3'b100 : 3'b010;
										assign node832 = (inp[5]) ? 3'b100 : node833;
											assign node833 = (inp[8]) ? 3'b010 : 3'b100;
									assign node837 = (inp[11]) ? node843 : node838;
										assign node838 = (inp[8]) ? 3'b110 : node839;
											assign node839 = (inp[2]) ? 3'b110 : 3'b010;
										assign node843 = (inp[5]) ? 3'b010 : 3'b110;
								assign node846 = (inp[8]) ? node848 : 3'b100;
									assign node848 = (inp[1]) ? node850 : 3'b100;
										assign node850 = (inp[2]) ? 3'b010 : node851;
											assign node851 = (inp[5]) ? 3'b100 : 3'b010;
							assign node855 = (inp[10]) ? node881 : node856;
								assign node856 = (inp[1]) ? node866 : node857;
									assign node857 = (inp[2]) ? node861 : node858;
										assign node858 = (inp[8]) ? 3'b110 : 3'b010;
										assign node861 = (inp[8]) ? node863 : 3'b110;
											assign node863 = (inp[5]) ? 3'b110 : 3'b010;
									assign node866 = (inp[5]) ? node874 : node867;
										assign node867 = (inp[11]) ? node869 : 3'b101;
											assign node869 = (inp[2]) ? 3'b101 : node870;
												assign node870 = (inp[8]) ? 3'b001 : 3'b101;
										assign node874 = (inp[11]) ? 3'b110 : node875;
											assign node875 = (inp[2]) ? node877 : 3'b110;
												assign node877 = (inp[8]) ? 3'b001 : 3'b110;
								assign node881 = (inp[2]) ? node887 : node882;
									assign node882 = (inp[1]) ? node884 : 3'b100;
										assign node884 = (inp[5]) ? 3'b010 : 3'b110;
									assign node887 = (inp[8]) ? node889 : 3'b010;
										assign node889 = (inp[1]) ? 3'b110 : 3'b010;
				assign node892 = (inp[0]) ? node924 : node893;
					assign node893 = (inp[4]) ? 3'b000 : node894;
						assign node894 = (inp[10]) ? node904 : node895;
							assign node895 = (inp[7]) ? node897 : 3'b000;
								assign node897 = (inp[8]) ? 3'b000 : node898;
									assign node898 = (inp[5]) ? node900 : 3'b000;
										assign node900 = (inp[2]) ? 3'b010 : 3'b000;
							assign node904 = (inp[1]) ? node912 : node905;
								assign node905 = (inp[7]) ? node907 : 3'b000;
									assign node907 = (inp[5]) ? 3'b000 : node908;
										assign node908 = (inp[8]) ? 3'b100 : 3'b000;
								assign node912 = (inp[2]) ? node918 : node913;
									assign node913 = (inp[5]) ? 3'b000 : node914;
										assign node914 = (inp[7]) ? 3'b100 : 3'b000;
									assign node918 = (inp[8]) ? node920 : 3'b100;
										assign node920 = (inp[11]) ? 3'b100 : 3'b000;
					assign node924 = (inp[4]) ? node936 : node925;
						assign node925 = (inp[5]) ? node931 : node926;
							assign node926 = (inp[1]) ? node928 : 3'b010;
								assign node928 = (inp[7]) ? 3'b110 : 3'b010;
							assign node931 = (inp[7]) ? node933 : 3'b100;
								assign node933 = (inp[1]) ? 3'b010 : 3'b100;
						assign node936 = (inp[1]) ? node946 : node937;
							assign node937 = (inp[7]) ? node939 : 3'b000;
								assign node939 = (inp[10]) ? 3'b000 : node940;
									assign node940 = (inp[8]) ? node942 : 3'b000;
										assign node942 = (inp[11]) ? 3'b000 : 3'b100;
							assign node946 = (inp[10]) ? node962 : node947;
								assign node947 = (inp[7]) ? node955 : node948;
									assign node948 = (inp[5]) ? node950 : 3'b100;
										assign node950 = (inp[8]) ? node952 : 3'b000;
											assign node952 = (inp[11]) ? 3'b000 : 3'b100;
									assign node955 = (inp[5]) ? 3'b100 : node956;
										assign node956 = (inp[11]) ? node958 : 3'b010;
											assign node958 = (inp[2]) ? 3'b100 : 3'b110;
								assign node962 = (inp[7]) ? node964 : 3'b000;
									assign node964 = (inp[5]) ? node970 : node965;
										assign node965 = (inp[11]) ? 3'b100 : node966;
											assign node966 = (inp[2]) ? 3'b000 : 3'b100;
										assign node970 = (inp[8]) ? node972 : 3'b000;
											assign node972 = (inp[2]) ? node974 : 3'b000;
												assign node974 = (inp[11]) ? 3'b000 : 3'b100;

endmodule