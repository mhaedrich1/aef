module dtc_split25_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node10;
	wire [15-1:0] node11;
	wire [15-1:0] node12;
	wire [15-1:0] node16;
	wire [15-1:0] node17;
	wire [15-1:0] node20;
	wire [15-1:0] node23;
	wire [15-1:0] node24;
	wire [15-1:0] node26;
	wire [15-1:0] node29;
	wire [15-1:0] node30;
	wire [15-1:0] node34;
	wire [15-1:0] node35;
	wire [15-1:0] node36;
	wire [15-1:0] node38;
	wire [15-1:0] node41;
	wire [15-1:0] node44;
	wire [15-1:0] node45;
	wire [15-1:0] node47;
	wire [15-1:0] node50;
	wire [15-1:0] node53;
	wire [15-1:0] node54;
	wire [15-1:0] node55;
	wire [15-1:0] node56;
	wire [15-1:0] node57;
	wire [15-1:0] node61;
	wire [15-1:0] node62;
	wire [15-1:0] node66;
	wire [15-1:0] node67;
	wire [15-1:0] node69;
	wire [15-1:0] node72;
	wire [15-1:0] node73;
	wire [15-1:0] node77;
	wire [15-1:0] node78;
	wire [15-1:0] node79;
	wire [15-1:0] node82;
	wire [15-1:0] node83;
	wire [15-1:0] node87;
	wire [15-1:0] node89;
	wire [15-1:0] node90;
	wire [15-1:0] node94;
	wire [15-1:0] node95;
	wire [15-1:0] node96;
	wire [15-1:0] node97;
	wire [15-1:0] node98;
	wire [15-1:0] node101;
	wire [15-1:0] node103;
	wire [15-1:0] node106;
	wire [15-1:0] node107;
	wire [15-1:0] node108;
	wire [15-1:0] node111;
	wire [15-1:0] node114;
	wire [15-1:0] node115;
	wire [15-1:0] node119;
	wire [15-1:0] node120;
	wire [15-1:0] node121;
	wire [15-1:0] node122;
	wire [15-1:0] node126;
	wire [15-1:0] node127;
	wire [15-1:0] node130;
	wire [15-1:0] node133;
	wire [15-1:0] node134;
	wire [15-1:0] node136;
	wire [15-1:0] node139;
	wire [15-1:0] node140;
	wire [15-1:0] node143;
	wire [15-1:0] node146;
	wire [15-1:0] node147;
	wire [15-1:0] node148;
	wire [15-1:0] node149;
	wire [15-1:0] node151;
	wire [15-1:0] node154;
	wire [15-1:0] node156;
	wire [15-1:0] node159;
	wire [15-1:0] node160;
	wire [15-1:0] node161;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node169;
	wire [15-1:0] node172;
	wire [15-1:0] node173;
	wire [15-1:0] node174;
	wire [15-1:0] node178;
	wire [15-1:0] node179;
	wire [15-1:0] node180;
	wire [15-1:0] node184;
	wire [15-1:0] node187;
	wire [15-1:0] node188;
	wire [15-1:0] node189;
	wire [15-1:0] node190;
	wire [15-1:0] node191;
	wire [15-1:0] node192;
	wire [15-1:0] node193;
	wire [15-1:0] node198;
	wire [15-1:0] node199;
	wire [15-1:0] node200;
	wire [15-1:0] node203;
	wire [15-1:0] node206;
	wire [15-1:0] node207;
	wire [15-1:0] node211;
	wire [15-1:0] node212;
	wire [15-1:0] node214;
	wire [15-1:0] node215;
	wire [15-1:0] node219;
	wire [15-1:0] node220;
	wire [15-1:0] node222;
	wire [15-1:0] node225;
	wire [15-1:0] node226;
	wire [15-1:0] node229;
	wire [15-1:0] node232;
	wire [15-1:0] node233;
	wire [15-1:0] node234;
	wire [15-1:0] node236;
	wire [15-1:0] node237;
	wire [15-1:0] node240;
	wire [15-1:0] node243;
	wire [15-1:0] node244;
	wire [15-1:0] node246;
	wire [15-1:0] node249;
	wire [15-1:0] node252;
	wire [15-1:0] node253;
	wire [15-1:0] node254;
	wire [15-1:0] node257;
	wire [15-1:0] node260;
	wire [15-1:0] node263;
	wire [15-1:0] node264;
	wire [15-1:0] node265;
	wire [15-1:0] node266;
	wire [15-1:0] node267;
	wire [15-1:0] node268;
	wire [15-1:0] node271;
	wire [15-1:0] node275;
	wire [15-1:0] node276;
	wire [15-1:0] node277;
	wire [15-1:0] node281;
	wire [15-1:0] node283;
	wire [15-1:0] node286;
	wire [15-1:0] node287;
	wire [15-1:0] node288;
	wire [15-1:0] node290;
	wire [15-1:0] node293;
	wire [15-1:0] node296;
	wire [15-1:0] node297;
	wire [15-1:0] node299;
	wire [15-1:0] node303;
	wire [15-1:0] node304;
	wire [15-1:0] node305;
	wire [15-1:0] node306;
	wire [15-1:0] node307;
	wire [15-1:0] node310;
	wire [15-1:0] node313;
	wire [15-1:0] node315;
	wire [15-1:0] node318;
	wire [15-1:0] node319;
	wire [15-1:0] node320;
	wire [15-1:0] node323;
	wire [15-1:0] node326;
	wire [15-1:0] node328;
	wire [15-1:0] node331;
	wire [15-1:0] node332;
	wire [15-1:0] node333;
	wire [15-1:0] node336;
	wire [15-1:0] node339;
	wire [15-1:0] node341;
	wire [15-1:0] node343;
	wire [15-1:0] node346;
	wire [15-1:0] node347;
	wire [15-1:0] node348;
	wire [15-1:0] node349;
	wire [15-1:0] node350;
	wire [15-1:0] node351;
	wire [15-1:0] node352;
	wire [15-1:0] node353;
	wire [15-1:0] node357;
	wire [15-1:0] node358;
	wire [15-1:0] node362;
	wire [15-1:0] node364;
	wire [15-1:0] node365;
	wire [15-1:0] node369;
	wire [15-1:0] node370;
	wire [15-1:0] node371;
	wire [15-1:0] node373;
	wire [15-1:0] node376;
	wire [15-1:0] node377;
	wire [15-1:0] node380;
	wire [15-1:0] node383;
	wire [15-1:0] node385;
	wire [15-1:0] node386;
	wire [15-1:0] node390;
	wire [15-1:0] node391;
	wire [15-1:0] node392;
	wire [15-1:0] node393;
	wire [15-1:0] node396;
	wire [15-1:0] node397;
	wire [15-1:0] node401;
	wire [15-1:0] node403;
	wire [15-1:0] node404;
	wire [15-1:0] node407;
	wire [15-1:0] node410;
	wire [15-1:0] node411;
	wire [15-1:0] node412;
	wire [15-1:0] node414;
	wire [15-1:0] node417;
	wire [15-1:0] node418;
	wire [15-1:0] node422;
	wire [15-1:0] node423;
	wire [15-1:0] node424;
	wire [15-1:0] node427;
	wire [15-1:0] node430;
	wire [15-1:0] node432;
	wire [15-1:0] node435;
	wire [15-1:0] node436;
	wire [15-1:0] node437;
	wire [15-1:0] node438;
	wire [15-1:0] node439;
	wire [15-1:0] node440;
	wire [15-1:0] node443;
	wire [15-1:0] node447;
	wire [15-1:0] node448;
	wire [15-1:0] node449;
	wire [15-1:0] node452;
	wire [15-1:0] node456;
	wire [15-1:0] node457;
	wire [15-1:0] node458;
	wire [15-1:0] node459;
	wire [15-1:0] node462;
	wire [15-1:0] node466;
	wire [15-1:0] node468;
	wire [15-1:0] node470;
	wire [15-1:0] node473;
	wire [15-1:0] node474;
	wire [15-1:0] node475;
	wire [15-1:0] node477;
	wire [15-1:0] node480;
	wire [15-1:0] node481;
	wire [15-1:0] node482;
	wire [15-1:0] node487;
	wire [15-1:0] node488;
	wire [15-1:0] node489;
	wire [15-1:0] node493;
	wire [15-1:0] node494;
	wire [15-1:0] node495;
	wire [15-1:0] node499;
	wire [15-1:0] node501;
	wire [15-1:0] node504;
	wire [15-1:0] node505;
	wire [15-1:0] node506;
	wire [15-1:0] node507;
	wire [15-1:0] node508;
	wire [15-1:0] node509;
	wire [15-1:0] node512;
	wire [15-1:0] node514;
	wire [15-1:0] node517;
	wire [15-1:0] node519;
	wire [15-1:0] node522;
	wire [15-1:0] node523;
	wire [15-1:0] node524;
	wire [15-1:0] node526;
	wire [15-1:0] node529;
	wire [15-1:0] node533;
	wire [15-1:0] node534;
	wire [15-1:0] node535;
	wire [15-1:0] node538;
	wire [15-1:0] node539;
	wire [15-1:0] node540;
	wire [15-1:0] node544;
	wire [15-1:0] node547;
	wire [15-1:0] node548;
	wire [15-1:0] node549;
	wire [15-1:0] node550;
	wire [15-1:0] node553;
	wire [15-1:0] node556;
	wire [15-1:0] node558;
	wire [15-1:0] node561;
	wire [15-1:0] node562;
	wire [15-1:0] node564;
	wire [15-1:0] node567;
	wire [15-1:0] node569;
	wire [15-1:0] node572;
	wire [15-1:0] node573;
	wire [15-1:0] node574;
	wire [15-1:0] node575;
	wire [15-1:0] node577;
	wire [15-1:0] node578;
	wire [15-1:0] node583;
	wire [15-1:0] node584;
	wire [15-1:0] node585;
	wire [15-1:0] node589;
	wire [15-1:0] node592;
	wire [15-1:0] node593;
	wire [15-1:0] node594;
	wire [15-1:0] node595;
	wire [15-1:0] node597;
	wire [15-1:0] node600;
	wire [15-1:0] node601;
	wire [15-1:0] node604;
	wire [15-1:0] node607;
	wire [15-1:0] node608;
	wire [15-1:0] node610;
	wire [15-1:0] node613;
	wire [15-1:0] node615;
	wire [15-1:0] node618;
	wire [15-1:0] node619;
	wire [15-1:0] node622;
	wire [15-1:0] node623;
	wire [15-1:0] node625;
	wire [15-1:0] node628;
	wire [15-1:0] node629;
	wire [15-1:0] node633;
	wire [15-1:0] node634;
	wire [15-1:0] node635;
	wire [15-1:0] node636;
	wire [15-1:0] node637;
	wire [15-1:0] node638;
	wire [15-1:0] node639;
	wire [15-1:0] node640;
	wire [15-1:0] node641;
	wire [15-1:0] node644;
	wire [15-1:0] node647;
	wire [15-1:0] node648;
	wire [15-1:0] node652;
	wire [15-1:0] node653;
	wire [15-1:0] node654;
	wire [15-1:0] node658;
	wire [15-1:0] node659;
	wire [15-1:0] node663;
	wire [15-1:0] node664;
	wire [15-1:0] node665;
	wire [15-1:0] node667;
	wire [15-1:0] node671;
	wire [15-1:0] node672;
	wire [15-1:0] node674;
	wire [15-1:0] node678;
	wire [15-1:0] node679;
	wire [15-1:0] node680;
	wire [15-1:0] node681;
	wire [15-1:0] node682;
	wire [15-1:0] node686;
	wire [15-1:0] node687;
	wire [15-1:0] node690;
	wire [15-1:0] node693;
	wire [15-1:0] node694;
	wire [15-1:0] node696;
	wire [15-1:0] node700;
	wire [15-1:0] node701;
	wire [15-1:0] node703;
	wire [15-1:0] node705;
	wire [15-1:0] node708;
	wire [15-1:0] node709;
	wire [15-1:0] node710;
	wire [15-1:0] node713;
	wire [15-1:0] node716;
	wire [15-1:0] node717;
	wire [15-1:0] node720;
	wire [15-1:0] node723;
	wire [15-1:0] node724;
	wire [15-1:0] node725;
	wire [15-1:0] node726;
	wire [15-1:0] node727;
	wire [15-1:0] node729;
	wire [15-1:0] node733;
	wire [15-1:0] node734;
	wire [15-1:0] node735;
	wire [15-1:0] node738;
	wire [15-1:0] node741;
	wire [15-1:0] node743;
	wire [15-1:0] node746;
	wire [15-1:0] node747;
	wire [15-1:0] node748;
	wire [15-1:0] node749;
	wire [15-1:0] node752;
	wire [15-1:0] node755;
	wire [15-1:0] node756;
	wire [15-1:0] node759;
	wire [15-1:0] node762;
	wire [15-1:0] node763;
	wire [15-1:0] node767;
	wire [15-1:0] node768;
	wire [15-1:0] node769;
	wire [15-1:0] node770;
	wire [15-1:0] node771;
	wire [15-1:0] node776;
	wire [15-1:0] node778;
	wire [15-1:0] node781;
	wire [15-1:0] node782;
	wire [15-1:0] node783;
	wire [15-1:0] node784;
	wire [15-1:0] node788;
	wire [15-1:0] node791;
	wire [15-1:0] node794;
	wire [15-1:0] node795;
	wire [15-1:0] node796;
	wire [15-1:0] node797;
	wire [15-1:0] node798;
	wire [15-1:0] node800;
	wire [15-1:0] node801;
	wire [15-1:0] node804;
	wire [15-1:0] node807;
	wire [15-1:0] node808;
	wire [15-1:0] node809;
	wire [15-1:0] node812;
	wire [15-1:0] node815;
	wire [15-1:0] node817;
	wire [15-1:0] node820;
	wire [15-1:0] node821;
	wire [15-1:0] node822;
	wire [15-1:0] node824;
	wire [15-1:0] node828;
	wire [15-1:0] node829;
	wire [15-1:0] node831;
	wire [15-1:0] node834;
	wire [15-1:0] node837;
	wire [15-1:0] node838;
	wire [15-1:0] node839;
	wire [15-1:0] node841;
	wire [15-1:0] node842;
	wire [15-1:0] node846;
	wire [15-1:0] node847;
	wire [15-1:0] node849;
	wire [15-1:0] node852;
	wire [15-1:0] node853;
	wire [15-1:0] node856;
	wire [15-1:0] node859;
	wire [15-1:0] node860;
	wire [15-1:0] node861;
	wire [15-1:0] node863;
	wire [15-1:0] node866;
	wire [15-1:0] node869;
	wire [15-1:0] node870;
	wire [15-1:0] node871;
	wire [15-1:0] node874;
	wire [15-1:0] node877;
	wire [15-1:0] node879;
	wire [15-1:0] node882;
	wire [15-1:0] node883;
	wire [15-1:0] node884;
	wire [15-1:0] node885;
	wire [15-1:0] node887;
	wire [15-1:0] node888;
	wire [15-1:0] node891;
	wire [15-1:0] node894;
	wire [15-1:0] node896;
	wire [15-1:0] node897;
	wire [15-1:0] node901;
	wire [15-1:0] node902;
	wire [15-1:0] node903;
	wire [15-1:0] node906;
	wire [15-1:0] node908;
	wire [15-1:0] node911;
	wire [15-1:0] node912;
	wire [15-1:0] node914;
	wire [15-1:0] node917;
	wire [15-1:0] node920;
	wire [15-1:0] node921;
	wire [15-1:0] node922;
	wire [15-1:0] node924;
	wire [15-1:0] node927;
	wire [15-1:0] node928;
	wire [15-1:0] node930;
	wire [15-1:0] node934;
	wire [15-1:0] node935;
	wire [15-1:0] node936;
	wire [15-1:0] node939;
	wire [15-1:0] node941;
	wire [15-1:0] node944;
	wire [15-1:0] node947;
	wire [15-1:0] node948;
	wire [15-1:0] node949;
	wire [15-1:0] node950;
	wire [15-1:0] node951;
	wire [15-1:0] node952;
	wire [15-1:0] node953;
	wire [15-1:0] node954;
	wire [15-1:0] node958;
	wire [15-1:0] node961;
	wire [15-1:0] node962;
	wire [15-1:0] node963;
	wire [15-1:0] node966;
	wire [15-1:0] node970;
	wire [15-1:0] node971;
	wire [15-1:0] node972;
	wire [15-1:0] node974;
	wire [15-1:0] node977;
	wire [15-1:0] node978;
	wire [15-1:0] node982;
	wire [15-1:0] node983;
	wire [15-1:0] node985;
	wire [15-1:0] node988;
	wire [15-1:0] node989;
	wire [15-1:0] node993;
	wire [15-1:0] node994;
	wire [15-1:0] node995;
	wire [15-1:0] node996;
	wire [15-1:0] node997;
	wire [15-1:0] node1000;
	wire [15-1:0] node1003;
	wire [15-1:0] node1004;
	wire [15-1:0] node1007;
	wire [15-1:0] node1010;
	wire [15-1:0] node1011;
	wire [15-1:0] node1012;
	wire [15-1:0] node1015;
	wire [15-1:0] node1018;
	wire [15-1:0] node1019;
	wire [15-1:0] node1023;
	wire [15-1:0] node1024;
	wire [15-1:0] node1025;
	wire [15-1:0] node1026;
	wire [15-1:0] node1030;
	wire [15-1:0] node1031;
	wire [15-1:0] node1034;
	wire [15-1:0] node1037;
	wire [15-1:0] node1038;
	wire [15-1:0] node1040;
	wire [15-1:0] node1043;
	wire [15-1:0] node1044;
	wire [15-1:0] node1048;
	wire [15-1:0] node1049;
	wire [15-1:0] node1050;
	wire [15-1:0] node1051;
	wire [15-1:0] node1053;
	wire [15-1:0] node1054;
	wire [15-1:0] node1057;
	wire [15-1:0] node1060;
	wire [15-1:0] node1062;
	wire [15-1:0] node1065;
	wire [15-1:0] node1066;
	wire [15-1:0] node1067;
	wire [15-1:0] node1068;
	wire [15-1:0] node1072;
	wire [15-1:0] node1074;
	wire [15-1:0] node1077;
	wire [15-1:0] node1078;
	wire [15-1:0] node1079;
	wire [15-1:0] node1082;
	wire [15-1:0] node1086;
	wire [15-1:0] node1087;
	wire [15-1:0] node1088;
	wire [15-1:0] node1089;
	wire [15-1:0] node1091;
	wire [15-1:0] node1094;
	wire [15-1:0] node1095;
	wire [15-1:0] node1099;
	wire [15-1:0] node1100;
	wire [15-1:0] node1101;
	wire [15-1:0] node1104;
	wire [15-1:0] node1107;
	wire [15-1:0] node1108;
	wire [15-1:0] node1111;
	wire [15-1:0] node1114;
	wire [15-1:0] node1115;
	wire [15-1:0] node1116;
	wire [15-1:0] node1117;
	wire [15-1:0] node1121;
	wire [15-1:0] node1122;
	wire [15-1:0] node1125;
	wire [15-1:0] node1128;
	wire [15-1:0] node1129;
	wire [15-1:0] node1133;
	wire [15-1:0] node1134;
	wire [15-1:0] node1135;
	wire [15-1:0] node1136;
	wire [15-1:0] node1137;
	wire [15-1:0] node1138;
	wire [15-1:0] node1139;
	wire [15-1:0] node1144;
	wire [15-1:0] node1146;
	wire [15-1:0] node1148;
	wire [15-1:0] node1151;
	wire [15-1:0] node1152;
	wire [15-1:0] node1153;
	wire [15-1:0] node1155;
	wire [15-1:0] node1159;
	wire [15-1:0] node1161;
	wire [15-1:0] node1164;
	wire [15-1:0] node1165;
	wire [15-1:0] node1166;
	wire [15-1:0] node1167;
	wire [15-1:0] node1168;
	wire [15-1:0] node1172;
	wire [15-1:0] node1173;
	wire [15-1:0] node1176;
	wire [15-1:0] node1179;
	wire [15-1:0] node1180;
	wire [15-1:0] node1182;
	wire [15-1:0] node1185;
	wire [15-1:0] node1187;
	wire [15-1:0] node1190;
	wire [15-1:0] node1191;
	wire [15-1:0] node1193;
	wire [15-1:0] node1195;
	wire [15-1:0] node1198;
	wire [15-1:0] node1200;
	wire [15-1:0] node1203;
	wire [15-1:0] node1204;
	wire [15-1:0] node1205;
	wire [15-1:0] node1206;
	wire [15-1:0] node1209;
	wire [15-1:0] node1210;
	wire [15-1:0] node1211;
	wire [15-1:0] node1214;
	wire [15-1:0] node1217;
	wire [15-1:0] node1218;
	wire [15-1:0] node1221;
	wire [15-1:0] node1224;
	wire [15-1:0] node1225;
	wire [15-1:0] node1226;
	wire [15-1:0] node1228;
	wire [15-1:0] node1231;
	wire [15-1:0] node1232;
	wire [15-1:0] node1235;
	wire [15-1:0] node1238;
	wire [15-1:0] node1239;
	wire [15-1:0] node1240;
	wire [15-1:0] node1244;
	wire [15-1:0] node1246;
	wire [15-1:0] node1249;
	wire [15-1:0] node1250;
	wire [15-1:0] node1251;
	wire [15-1:0] node1252;
	wire [15-1:0] node1253;
	wire [15-1:0] node1256;
	wire [15-1:0] node1259;
	wire [15-1:0] node1261;
	wire [15-1:0] node1264;
	wire [15-1:0] node1265;
	wire [15-1:0] node1268;
	wire [15-1:0] node1270;
	wire [15-1:0] node1273;
	wire [15-1:0] node1274;
	wire [15-1:0] node1275;
	wire [15-1:0] node1277;
	wire [15-1:0] node1280;
	wire [15-1:0] node1282;
	wire [15-1:0] node1285;
	wire [15-1:0] node1286;
	wire [15-1:0] node1288;
	wire [15-1:0] node1291;
	wire [15-1:0] node1292;
	wire [15-1:0] node1295;
	wire [15-1:0] node1298;
	wire [15-1:0] node1299;
	wire [15-1:0] node1300;
	wire [15-1:0] node1301;
	wire [15-1:0] node1302;
	wire [15-1:0] node1303;
	wire [15-1:0] node1304;
	wire [15-1:0] node1305;
	wire [15-1:0] node1308;
	wire [15-1:0] node1309;
	wire [15-1:0] node1310;
	wire [15-1:0] node1313;
	wire [15-1:0] node1316;
	wire [15-1:0] node1317;
	wire [15-1:0] node1320;
	wire [15-1:0] node1323;
	wire [15-1:0] node1324;
	wire [15-1:0] node1325;
	wire [15-1:0] node1326;
	wire [15-1:0] node1329;
	wire [15-1:0] node1332;
	wire [15-1:0] node1334;
	wire [15-1:0] node1337;
	wire [15-1:0] node1338;
	wire [15-1:0] node1339;
	wire [15-1:0] node1342;
	wire [15-1:0] node1345;
	wire [15-1:0] node1346;
	wire [15-1:0] node1350;
	wire [15-1:0] node1351;
	wire [15-1:0] node1352;
	wire [15-1:0] node1353;
	wire [15-1:0] node1356;
	wire [15-1:0] node1359;
	wire [15-1:0] node1360;
	wire [15-1:0] node1361;
	wire [15-1:0] node1364;
	wire [15-1:0] node1368;
	wire [15-1:0] node1369;
	wire [15-1:0] node1370;
	wire [15-1:0] node1371;
	wire [15-1:0] node1374;
	wire [15-1:0] node1377;
	wire [15-1:0] node1378;
	wire [15-1:0] node1381;
	wire [15-1:0] node1384;
	wire [15-1:0] node1385;
	wire [15-1:0] node1387;
	wire [15-1:0] node1391;
	wire [15-1:0] node1392;
	wire [15-1:0] node1393;
	wire [15-1:0] node1394;
	wire [15-1:0] node1396;
	wire [15-1:0] node1399;
	wire [15-1:0] node1400;
	wire [15-1:0] node1401;
	wire [15-1:0] node1405;
	wire [15-1:0] node1408;
	wire [15-1:0] node1409;
	wire [15-1:0] node1410;
	wire [15-1:0] node1414;
	wire [15-1:0] node1416;
	wire [15-1:0] node1417;
	wire [15-1:0] node1421;
	wire [15-1:0] node1422;
	wire [15-1:0] node1423;
	wire [15-1:0] node1424;
	wire [15-1:0] node1425;
	wire [15-1:0] node1428;
	wire [15-1:0] node1431;
	wire [15-1:0] node1432;
	wire [15-1:0] node1435;
	wire [15-1:0] node1438;
	wire [15-1:0] node1439;
	wire [15-1:0] node1442;
	wire [15-1:0] node1443;
	wire [15-1:0] node1447;
	wire [15-1:0] node1448;
	wire [15-1:0] node1449;
	wire [15-1:0] node1452;
	wire [15-1:0] node1454;
	wire [15-1:0] node1457;
	wire [15-1:0] node1458;
	wire [15-1:0] node1462;
	wire [15-1:0] node1463;
	wire [15-1:0] node1464;
	wire [15-1:0] node1465;
	wire [15-1:0] node1466;
	wire [15-1:0] node1467;
	wire [15-1:0] node1469;
	wire [15-1:0] node1472;
	wire [15-1:0] node1474;
	wire [15-1:0] node1477;
	wire [15-1:0] node1478;
	wire [15-1:0] node1479;
	wire [15-1:0] node1483;
	wire [15-1:0] node1484;
	wire [15-1:0] node1487;
	wire [15-1:0] node1490;
	wire [15-1:0] node1491;
	wire [15-1:0] node1492;
	wire [15-1:0] node1493;
	wire [15-1:0] node1496;
	wire [15-1:0] node1499;
	wire [15-1:0] node1501;
	wire [15-1:0] node1504;
	wire [15-1:0] node1505;
	wire [15-1:0] node1506;
	wire [15-1:0] node1509;
	wire [15-1:0] node1513;
	wire [15-1:0] node1514;
	wire [15-1:0] node1515;
	wire [15-1:0] node1516;
	wire [15-1:0] node1518;
	wire [15-1:0] node1522;
	wire [15-1:0] node1523;
	wire [15-1:0] node1524;
	wire [15-1:0] node1527;
	wire [15-1:0] node1530;
	wire [15-1:0] node1531;
	wire [15-1:0] node1535;
	wire [15-1:0] node1536;
	wire [15-1:0] node1537;
	wire [15-1:0] node1540;
	wire [15-1:0] node1541;
	wire [15-1:0] node1545;
	wire [15-1:0] node1546;
	wire [15-1:0] node1547;
	wire [15-1:0] node1550;
	wire [15-1:0] node1553;
	wire [15-1:0] node1556;
	wire [15-1:0] node1557;
	wire [15-1:0] node1558;
	wire [15-1:0] node1559;
	wire [15-1:0] node1560;
	wire [15-1:0] node1561;
	wire [15-1:0] node1566;
	wire [15-1:0] node1567;
	wire [15-1:0] node1568;
	wire [15-1:0] node1572;
	wire [15-1:0] node1574;
	wire [15-1:0] node1577;
	wire [15-1:0] node1578;
	wire [15-1:0] node1579;
	wire [15-1:0] node1581;
	wire [15-1:0] node1585;
	wire [15-1:0] node1588;
	wire [15-1:0] node1589;
	wire [15-1:0] node1590;
	wire [15-1:0] node1591;
	wire [15-1:0] node1592;
	wire [15-1:0] node1595;
	wire [15-1:0] node1598;
	wire [15-1:0] node1600;
	wire [15-1:0] node1603;
	wire [15-1:0] node1605;
	wire [15-1:0] node1606;
	wire [15-1:0] node1610;
	wire [15-1:0] node1611;
	wire [15-1:0] node1613;
	wire [15-1:0] node1614;
	wire [15-1:0] node1618;
	wire [15-1:0] node1619;
	wire [15-1:0] node1621;
	wire [15-1:0] node1624;
	wire [15-1:0] node1625;
	wire [15-1:0] node1629;
	wire [15-1:0] node1630;
	wire [15-1:0] node1631;
	wire [15-1:0] node1632;
	wire [15-1:0] node1633;
	wire [15-1:0] node1634;
	wire [15-1:0] node1635;
	wire [15-1:0] node1637;
	wire [15-1:0] node1640;
	wire [15-1:0] node1641;
	wire [15-1:0] node1645;
	wire [15-1:0] node1646;
	wire [15-1:0] node1647;
	wire [15-1:0] node1650;
	wire [15-1:0] node1653;
	wire [15-1:0] node1656;
	wire [15-1:0] node1657;
	wire [15-1:0] node1658;
	wire [15-1:0] node1660;
	wire [15-1:0] node1663;
	wire [15-1:0] node1664;
	wire [15-1:0] node1667;
	wire [15-1:0] node1670;
	wire [15-1:0] node1671;
	wire [15-1:0] node1672;
	wire [15-1:0] node1675;
	wire [15-1:0] node1678;
	wire [15-1:0] node1679;
	wire [15-1:0] node1683;
	wire [15-1:0] node1684;
	wire [15-1:0] node1685;
	wire [15-1:0] node1686;
	wire [15-1:0] node1687;
	wire [15-1:0] node1690;
	wire [15-1:0] node1693;
	wire [15-1:0] node1694;
	wire [15-1:0] node1697;
	wire [15-1:0] node1700;
	wire [15-1:0] node1702;
	wire [15-1:0] node1705;
	wire [15-1:0] node1706;
	wire [15-1:0] node1708;
	wire [15-1:0] node1709;
	wire [15-1:0] node1713;
	wire [15-1:0] node1715;
	wire [15-1:0] node1716;
	wire [15-1:0] node1720;
	wire [15-1:0] node1721;
	wire [15-1:0] node1722;
	wire [15-1:0] node1723;
	wire [15-1:0] node1724;
	wire [15-1:0] node1725;
	wire [15-1:0] node1729;
	wire [15-1:0] node1732;
	wire [15-1:0] node1733;
	wire [15-1:0] node1734;
	wire [15-1:0] node1738;
	wire [15-1:0] node1739;
	wire [15-1:0] node1743;
	wire [15-1:0] node1744;
	wire [15-1:0] node1746;
	wire [15-1:0] node1747;
	wire [15-1:0] node1751;
	wire [15-1:0] node1752;
	wire [15-1:0] node1753;
	wire [15-1:0] node1756;
	wire [15-1:0] node1759;
	wire [15-1:0] node1760;
	wire [15-1:0] node1764;
	wire [15-1:0] node1765;
	wire [15-1:0] node1766;
	wire [15-1:0] node1768;
	wire [15-1:0] node1769;
	wire [15-1:0] node1773;
	wire [15-1:0] node1774;
	wire [15-1:0] node1775;
	wire [15-1:0] node1778;
	wire [15-1:0] node1781;
	wire [15-1:0] node1783;
	wire [15-1:0] node1786;
	wire [15-1:0] node1787;
	wire [15-1:0] node1789;
	wire [15-1:0] node1790;
	wire [15-1:0] node1794;
	wire [15-1:0] node1795;
	wire [15-1:0] node1798;
	wire [15-1:0] node1800;
	wire [15-1:0] node1803;
	wire [15-1:0] node1804;
	wire [15-1:0] node1805;
	wire [15-1:0] node1806;
	wire [15-1:0] node1807;
	wire [15-1:0] node1808;
	wire [15-1:0] node1810;
	wire [15-1:0] node1814;
	wire [15-1:0] node1815;
	wire [15-1:0] node1816;
	wire [15-1:0] node1819;
	wire [15-1:0] node1822;
	wire [15-1:0] node1823;
	wire [15-1:0] node1827;
	wire [15-1:0] node1828;
	wire [15-1:0] node1829;
	wire [15-1:0] node1831;
	wire [15-1:0] node1835;
	wire [15-1:0] node1836;
	wire [15-1:0] node1838;
	wire [15-1:0] node1842;
	wire [15-1:0] node1843;
	wire [15-1:0] node1844;
	wire [15-1:0] node1845;
	wire [15-1:0] node1846;
	wire [15-1:0] node1849;
	wire [15-1:0] node1852;
	wire [15-1:0] node1853;
	wire [15-1:0] node1856;
	wire [15-1:0] node1859;
	wire [15-1:0] node1861;
	wire [15-1:0] node1862;
	wire [15-1:0] node1865;
	wire [15-1:0] node1868;
	wire [15-1:0] node1869;
	wire [15-1:0] node1871;
	wire [15-1:0] node1874;
	wire [15-1:0] node1875;
	wire [15-1:0] node1878;
	wire [15-1:0] node1880;
	wire [15-1:0] node1883;
	wire [15-1:0] node1884;
	wire [15-1:0] node1885;
	wire [15-1:0] node1886;
	wire [15-1:0] node1887;
	wire [15-1:0] node1889;
	wire [15-1:0] node1892;
	wire [15-1:0] node1895;
	wire [15-1:0] node1896;
	wire [15-1:0] node1898;
	wire [15-1:0] node1901;
	wire [15-1:0] node1902;
	wire [15-1:0] node1906;
	wire [15-1:0] node1907;
	wire [15-1:0] node1908;
	wire [15-1:0] node1911;
	wire [15-1:0] node1912;
	wire [15-1:0] node1916;
	wire [15-1:0] node1917;
	wire [15-1:0] node1919;
	wire [15-1:0] node1923;
	wire [15-1:0] node1924;
	wire [15-1:0] node1925;
	wire [15-1:0] node1926;
	wire [15-1:0] node1927;
	wire [15-1:0] node1931;
	wire [15-1:0] node1934;
	wire [15-1:0] node1935;
	wire [15-1:0] node1937;
	wire [15-1:0] node1940;
	wire [15-1:0] node1941;
	wire [15-1:0] node1944;
	wire [15-1:0] node1947;
	wire [15-1:0] node1948;
	wire [15-1:0] node1949;
	wire [15-1:0] node1951;
	wire [15-1:0] node1954;
	wire [15-1:0] node1955;
	wire [15-1:0] node1958;
	wire [15-1:0] node1961;
	wire [15-1:0] node1963;
	wire [15-1:0] node1966;
	wire [15-1:0] node1967;
	wire [15-1:0] node1968;
	wire [15-1:0] node1969;
	wire [15-1:0] node1970;
	wire [15-1:0] node1971;
	wire [15-1:0] node1972;
	wire [15-1:0] node1973;
	wire [15-1:0] node1975;
	wire [15-1:0] node1978;
	wire [15-1:0] node1981;
	wire [15-1:0] node1982;
	wire [15-1:0] node1983;
	wire [15-1:0] node1986;
	wire [15-1:0] node1989;
	wire [15-1:0] node1992;
	wire [15-1:0] node1993;
	wire [15-1:0] node1995;
	wire [15-1:0] node1999;
	wire [15-1:0] node2000;
	wire [15-1:0] node2001;
	wire [15-1:0] node2002;
	wire [15-1:0] node2004;
	wire [15-1:0] node2007;
	wire [15-1:0] node2008;
	wire [15-1:0] node2012;
	wire [15-1:0] node2013;
	wire [15-1:0] node2016;
	wire [15-1:0] node2017;
	wire [15-1:0] node2021;
	wire [15-1:0] node2022;
	wire [15-1:0] node2023;
	wire [15-1:0] node2024;
	wire [15-1:0] node2027;
	wire [15-1:0] node2030;
	wire [15-1:0] node2033;
	wire [15-1:0] node2034;
	wire [15-1:0] node2038;
	wire [15-1:0] node2039;
	wire [15-1:0] node2040;
	wire [15-1:0] node2041;
	wire [15-1:0] node2042;
	wire [15-1:0] node2045;
	wire [15-1:0] node2046;
	wire [15-1:0] node2049;
	wire [15-1:0] node2052;
	wire [15-1:0] node2053;
	wire [15-1:0] node2055;
	wire [15-1:0] node2058;
	wire [15-1:0] node2059;
	wire [15-1:0] node2063;
	wire [15-1:0] node2064;
	wire [15-1:0] node2065;
	wire [15-1:0] node2067;
	wire [15-1:0] node2070;
	wire [15-1:0] node2073;
	wire [15-1:0] node2074;
	wire [15-1:0] node2075;
	wire [15-1:0] node2080;
	wire [15-1:0] node2081;
	wire [15-1:0] node2082;
	wire [15-1:0] node2083;
	wire [15-1:0] node2086;
	wire [15-1:0] node2087;
	wire [15-1:0] node2090;
	wire [15-1:0] node2093;
	wire [15-1:0] node2094;
	wire [15-1:0] node2096;
	wire [15-1:0] node2099;
	wire [15-1:0] node2100;
	wire [15-1:0] node2104;
	wire [15-1:0] node2105;
	wire [15-1:0] node2108;
	wire [15-1:0] node2110;
	wire [15-1:0] node2111;
	wire [15-1:0] node2115;
	wire [15-1:0] node2116;
	wire [15-1:0] node2117;
	wire [15-1:0] node2118;
	wire [15-1:0] node2119;
	wire [15-1:0] node2121;
	wire [15-1:0] node2122;
	wire [15-1:0] node2125;
	wire [15-1:0] node2128;
	wire [15-1:0] node2130;
	wire [15-1:0] node2131;
	wire [15-1:0] node2135;
	wire [15-1:0] node2136;
	wire [15-1:0] node2137;
	wire [15-1:0] node2139;
	wire [15-1:0] node2142;
	wire [15-1:0] node2143;
	wire [15-1:0] node2147;
	wire [15-1:0] node2148;
	wire [15-1:0] node2152;
	wire [15-1:0] node2153;
	wire [15-1:0] node2154;
	wire [15-1:0] node2155;
	wire [15-1:0] node2157;
	wire [15-1:0] node2161;
	wire [15-1:0] node2163;
	wire [15-1:0] node2166;
	wire [15-1:0] node2167;
	wire [15-1:0] node2168;
	wire [15-1:0] node2169;
	wire [15-1:0] node2173;
	wire [15-1:0] node2175;
	wire [15-1:0] node2178;
	wire [15-1:0] node2179;
	wire [15-1:0] node2181;
	wire [15-1:0] node2184;
	wire [15-1:0] node2187;
	wire [15-1:0] node2188;
	wire [15-1:0] node2189;
	wire [15-1:0] node2190;
	wire [15-1:0] node2191;
	wire [15-1:0] node2192;
	wire [15-1:0] node2195;
	wire [15-1:0] node2198;
	wire [15-1:0] node2199;
	wire [15-1:0] node2203;
	wire [15-1:0] node2205;
	wire [15-1:0] node2206;
	wire [15-1:0] node2209;
	wire [15-1:0] node2212;
	wire [15-1:0] node2213;
	wire [15-1:0] node2214;
	wire [15-1:0] node2215;
	wire [15-1:0] node2218;
	wire [15-1:0] node2221;
	wire [15-1:0] node2223;
	wire [15-1:0] node2226;
	wire [15-1:0] node2227;
	wire [15-1:0] node2229;
	wire [15-1:0] node2232;
	wire [15-1:0] node2234;
	wire [15-1:0] node2237;
	wire [15-1:0] node2238;
	wire [15-1:0] node2239;
	wire [15-1:0] node2241;
	wire [15-1:0] node2244;
	wire [15-1:0] node2245;
	wire [15-1:0] node2246;
	wire [15-1:0] node2250;
	wire [15-1:0] node2253;
	wire [15-1:0] node2254;
	wire [15-1:0] node2255;
	wire [15-1:0] node2256;
	wire [15-1:0] node2260;
	wire [15-1:0] node2261;
	wire [15-1:0] node2265;
	wire [15-1:0] node2266;
	wire [15-1:0] node2269;
	wire [15-1:0] node2270;
	wire [15-1:0] node2274;
	wire [15-1:0] node2275;
	wire [15-1:0] node2276;
	wire [15-1:0] node2277;
	wire [15-1:0] node2278;
	wire [15-1:0] node2279;
	wire [15-1:0] node2280;
	wire [15-1:0] node2283;
	wire [15-1:0] node2284;
	wire [15-1:0] node2288;
	wire [15-1:0] node2289;
	wire [15-1:0] node2291;
	wire [15-1:0] node2295;
	wire [15-1:0] node2296;
	wire [15-1:0] node2297;
	wire [15-1:0] node2300;
	wire [15-1:0] node2302;
	wire [15-1:0] node2305;
	wire [15-1:0] node2307;
	wire [15-1:0] node2308;
	wire [15-1:0] node2312;
	wire [15-1:0] node2313;
	wire [15-1:0] node2314;
	wire [15-1:0] node2315;
	wire [15-1:0] node2317;
	wire [15-1:0] node2320;
	wire [15-1:0] node2321;
	wire [15-1:0] node2324;
	wire [15-1:0] node2327;
	wire [15-1:0] node2329;
	wire [15-1:0] node2330;
	wire [15-1:0] node2334;
	wire [15-1:0] node2335;
	wire [15-1:0] node2337;
	wire [15-1:0] node2338;
	wire [15-1:0] node2342;
	wire [15-1:0] node2343;
	wire [15-1:0] node2346;
	wire [15-1:0] node2348;
	wire [15-1:0] node2351;
	wire [15-1:0] node2352;
	wire [15-1:0] node2353;
	wire [15-1:0] node2354;
	wire [15-1:0] node2355;
	wire [15-1:0] node2357;
	wire [15-1:0] node2360;
	wire [15-1:0] node2363;
	wire [15-1:0] node2364;
	wire [15-1:0] node2366;
	wire [15-1:0] node2369;
	wire [15-1:0] node2371;
	wire [15-1:0] node2374;
	wire [15-1:0] node2375;
	wire [15-1:0] node2377;
	wire [15-1:0] node2378;
	wire [15-1:0] node2382;
	wire [15-1:0] node2383;
	wire [15-1:0] node2385;
	wire [15-1:0] node2388;
	wire [15-1:0] node2391;
	wire [15-1:0] node2392;
	wire [15-1:0] node2393;
	wire [15-1:0] node2395;
	wire [15-1:0] node2396;
	wire [15-1:0] node2399;
	wire [15-1:0] node2402;
	wire [15-1:0] node2403;
	wire [15-1:0] node2405;
	wire [15-1:0] node2408;
	wire [15-1:0] node2411;
	wire [15-1:0] node2412;
	wire [15-1:0] node2413;
	wire [15-1:0] node2416;
	wire [15-1:0] node2418;
	wire [15-1:0] node2421;
	wire [15-1:0] node2422;
	wire [15-1:0] node2424;
	wire [15-1:0] node2427;
	wire [15-1:0] node2429;
	wire [15-1:0] node2432;
	wire [15-1:0] node2433;
	wire [15-1:0] node2434;
	wire [15-1:0] node2435;
	wire [15-1:0] node2436;
	wire [15-1:0] node2439;
	wire [15-1:0] node2440;
	wire [15-1:0] node2442;
	wire [15-1:0] node2445;
	wire [15-1:0] node2448;
	wire [15-1:0] node2449;
	wire [15-1:0] node2451;
	wire [15-1:0] node2452;
	wire [15-1:0] node2456;
	wire [15-1:0] node2457;
	wire [15-1:0] node2458;
	wire [15-1:0] node2461;
	wire [15-1:0] node2464;
	wire [15-1:0] node2466;
	wire [15-1:0] node2469;
	wire [15-1:0] node2470;
	wire [15-1:0] node2471;
	wire [15-1:0] node2472;
	wire [15-1:0] node2474;
	wire [15-1:0] node2477;
	wire [15-1:0] node2478;
	wire [15-1:0] node2481;
	wire [15-1:0] node2484;
	wire [15-1:0] node2485;
	wire [15-1:0] node2486;
	wire [15-1:0] node2489;
	wire [15-1:0] node2492;
	wire [15-1:0] node2494;
	wire [15-1:0] node2497;
	wire [15-1:0] node2498;
	wire [15-1:0] node2499;
	wire [15-1:0] node2501;
	wire [15-1:0] node2505;
	wire [15-1:0] node2506;
	wire [15-1:0] node2509;
	wire [15-1:0] node2510;
	wire [15-1:0] node2514;
	wire [15-1:0] node2515;
	wire [15-1:0] node2516;
	wire [15-1:0] node2517;
	wire [15-1:0] node2518;
	wire [15-1:0] node2521;
	wire [15-1:0] node2523;
	wire [15-1:0] node2526;
	wire [15-1:0] node2527;
	wire [15-1:0] node2530;
	wire [15-1:0] node2532;
	wire [15-1:0] node2535;
	wire [15-1:0] node2536;
	wire [15-1:0] node2538;
	wire [15-1:0] node2540;
	wire [15-1:0] node2543;
	wire [15-1:0] node2545;
	wire [15-1:0] node2546;
	wire [15-1:0] node2550;
	wire [15-1:0] node2551;
	wire [15-1:0] node2552;
	wire [15-1:0] node2553;
	wire [15-1:0] node2556;
	wire [15-1:0] node2559;
	wire [15-1:0] node2560;
	wire [15-1:0] node2562;
	wire [15-1:0] node2566;
	wire [15-1:0] node2567;
	wire [15-1:0] node2568;
	wire [15-1:0] node2571;
	wire [15-1:0] node2574;
	wire [15-1:0] node2575;
	wire [15-1:0] node2576;
	wire [15-1:0] node2580;
	wire [15-1:0] node2583;
	wire [15-1:0] node2584;
	wire [15-1:0] node2585;
	wire [15-1:0] node2586;
	wire [15-1:0] node2587;
	wire [15-1:0] node2588;
	wire [15-1:0] node2589;
	wire [15-1:0] node2590;
	wire [15-1:0] node2591;
	wire [15-1:0] node2592;
	wire [15-1:0] node2593;
	wire [15-1:0] node2597;
	wire [15-1:0] node2598;
	wire [15-1:0] node2602;
	wire [15-1:0] node2603;
	wire [15-1:0] node2605;
	wire [15-1:0] node2608;
	wire [15-1:0] node2609;
	wire [15-1:0] node2612;
	wire [15-1:0] node2615;
	wire [15-1:0] node2616;
	wire [15-1:0] node2617;
	wire [15-1:0] node2620;
	wire [15-1:0] node2622;
	wire [15-1:0] node2625;
	wire [15-1:0] node2626;
	wire [15-1:0] node2627;
	wire [15-1:0] node2630;
	wire [15-1:0] node2633;
	wire [15-1:0] node2634;
	wire [15-1:0] node2638;
	wire [15-1:0] node2639;
	wire [15-1:0] node2640;
	wire [15-1:0] node2641;
	wire [15-1:0] node2643;
	wire [15-1:0] node2646;
	wire [15-1:0] node2648;
	wire [15-1:0] node2651;
	wire [15-1:0] node2652;
	wire [15-1:0] node2653;
	wire [15-1:0] node2656;
	wire [15-1:0] node2659;
	wire [15-1:0] node2660;
	wire [15-1:0] node2663;
	wire [15-1:0] node2666;
	wire [15-1:0] node2667;
	wire [15-1:0] node2668;
	wire [15-1:0] node2669;
	wire [15-1:0] node2672;
	wire [15-1:0] node2675;
	wire [15-1:0] node2678;
	wire [15-1:0] node2679;
	wire [15-1:0] node2683;
	wire [15-1:0] node2684;
	wire [15-1:0] node2685;
	wire [15-1:0] node2686;
	wire [15-1:0] node2688;
	wire [15-1:0] node2689;
	wire [15-1:0] node2693;
	wire [15-1:0] node2694;
	wire [15-1:0] node2695;
	wire [15-1:0] node2699;
	wire [15-1:0] node2700;
	wire [15-1:0] node2704;
	wire [15-1:0] node2705;
	wire [15-1:0] node2706;
	wire [15-1:0] node2707;
	wire [15-1:0] node2710;
	wire [15-1:0] node2713;
	wire [15-1:0] node2714;
	wire [15-1:0] node2718;
	wire [15-1:0] node2719;
	wire [15-1:0] node2721;
	wire [15-1:0] node2724;
	wire [15-1:0] node2725;
	wire [15-1:0] node2728;
	wire [15-1:0] node2731;
	wire [15-1:0] node2732;
	wire [15-1:0] node2733;
	wire [15-1:0] node2734;
	wire [15-1:0] node2735;
	wire [15-1:0] node2740;
	wire [15-1:0] node2742;
	wire [15-1:0] node2743;
	wire [15-1:0] node2746;
	wire [15-1:0] node2749;
	wire [15-1:0] node2750;
	wire [15-1:0] node2751;
	wire [15-1:0] node2753;
	wire [15-1:0] node2756;
	wire [15-1:0] node2757;
	wire [15-1:0] node2761;
	wire [15-1:0] node2764;
	wire [15-1:0] node2765;
	wire [15-1:0] node2766;
	wire [15-1:0] node2767;
	wire [15-1:0] node2768;
	wire [15-1:0] node2769;
	wire [15-1:0] node2770;
	wire [15-1:0] node2774;
	wire [15-1:0] node2777;
	wire [15-1:0] node2778;
	wire [15-1:0] node2779;
	wire [15-1:0] node2783;
	wire [15-1:0] node2785;
	wire [15-1:0] node2788;
	wire [15-1:0] node2789;
	wire [15-1:0] node2790;
	wire [15-1:0] node2791;
	wire [15-1:0] node2795;
	wire [15-1:0] node2796;
	wire [15-1:0] node2800;
	wire [15-1:0] node2801;
	wire [15-1:0] node2802;
	wire [15-1:0] node2806;
	wire [15-1:0] node2809;
	wire [15-1:0] node2810;
	wire [15-1:0] node2811;
	wire [15-1:0] node2812;
	wire [15-1:0] node2813;
	wire [15-1:0] node2816;
	wire [15-1:0] node2819;
	wire [15-1:0] node2822;
	wire [15-1:0] node2823;
	wire [15-1:0] node2824;
	wire [15-1:0] node2827;
	wire [15-1:0] node2830;
	wire [15-1:0] node2831;
	wire [15-1:0] node2835;
	wire [15-1:0] node2836;
	wire [15-1:0] node2837;
	wire [15-1:0] node2839;
	wire [15-1:0] node2843;
	wire [15-1:0] node2845;
	wire [15-1:0] node2846;
	wire [15-1:0] node2850;
	wire [15-1:0] node2851;
	wire [15-1:0] node2852;
	wire [15-1:0] node2853;
	wire [15-1:0] node2854;
	wire [15-1:0] node2856;
	wire [15-1:0] node2859;
	wire [15-1:0] node2860;
	wire [15-1:0] node2864;
	wire [15-1:0] node2867;
	wire [15-1:0] node2868;
	wire [15-1:0] node2869;
	wire [15-1:0] node2871;
	wire [15-1:0] node2874;
	wire [15-1:0] node2875;
	wire [15-1:0] node2879;
	wire [15-1:0] node2880;
	wire [15-1:0] node2883;
	wire [15-1:0] node2884;
	wire [15-1:0] node2888;
	wire [15-1:0] node2889;
	wire [15-1:0] node2890;
	wire [15-1:0] node2891;
	wire [15-1:0] node2893;
	wire [15-1:0] node2896;
	wire [15-1:0] node2898;
	wire [15-1:0] node2901;
	wire [15-1:0] node2903;
	wire [15-1:0] node2904;
	wire [15-1:0] node2907;
	wire [15-1:0] node2910;
	wire [15-1:0] node2911;
	wire [15-1:0] node2912;
	wire [15-1:0] node2914;
	wire [15-1:0] node2918;
	wire [15-1:0] node2919;
	wire [15-1:0] node2920;
	wire [15-1:0] node2923;
	wire [15-1:0] node2926;
	wire [15-1:0] node2927;
	wire [15-1:0] node2930;
	wire [15-1:0] node2933;
	wire [15-1:0] node2934;
	wire [15-1:0] node2935;
	wire [15-1:0] node2936;
	wire [15-1:0] node2937;
	wire [15-1:0] node2938;
	wire [15-1:0] node2939;
	wire [15-1:0] node2942;
	wire [15-1:0] node2944;
	wire [15-1:0] node2947;
	wire [15-1:0] node2948;
	wire [15-1:0] node2950;
	wire [15-1:0] node2953;
	wire [15-1:0] node2954;
	wire [15-1:0] node2958;
	wire [15-1:0] node2959;
	wire [15-1:0] node2961;
	wire [15-1:0] node2963;
	wire [15-1:0] node2966;
	wire [15-1:0] node2967;
	wire [15-1:0] node2968;
	wire [15-1:0] node2971;
	wire [15-1:0] node2975;
	wire [15-1:0] node2976;
	wire [15-1:0] node2977;
	wire [15-1:0] node2978;
	wire [15-1:0] node2979;
	wire [15-1:0] node2984;
	wire [15-1:0] node2985;
	wire [15-1:0] node2987;
	wire [15-1:0] node2991;
	wire [15-1:0] node2992;
	wire [15-1:0] node2993;
	wire [15-1:0] node2995;
	wire [15-1:0] node2999;
	wire [15-1:0] node3002;
	wire [15-1:0] node3003;
	wire [15-1:0] node3004;
	wire [15-1:0] node3005;
	wire [15-1:0] node3006;
	wire [15-1:0] node3007;
	wire [15-1:0] node3010;
	wire [15-1:0] node3013;
	wire [15-1:0] node3014;
	wire [15-1:0] node3017;
	wire [15-1:0] node3020;
	wire [15-1:0] node3021;
	wire [15-1:0] node3022;
	wire [15-1:0] node3025;
	wire [15-1:0] node3028;
	wire [15-1:0] node3029;
	wire [15-1:0] node3032;
	wire [15-1:0] node3035;
	wire [15-1:0] node3036;
	wire [15-1:0] node3037;
	wire [15-1:0] node3039;
	wire [15-1:0] node3042;
	wire [15-1:0] node3043;
	wire [15-1:0] node3047;
	wire [15-1:0] node3048;
	wire [15-1:0] node3050;
	wire [15-1:0] node3054;
	wire [15-1:0] node3055;
	wire [15-1:0] node3056;
	wire [15-1:0] node3057;
	wire [15-1:0] node3059;
	wire [15-1:0] node3062;
	wire [15-1:0] node3065;
	wire [15-1:0] node3066;
	wire [15-1:0] node3067;
	wire [15-1:0] node3070;
	wire [15-1:0] node3073;
	wire [15-1:0] node3074;
	wire [15-1:0] node3078;
	wire [15-1:0] node3079;
	wire [15-1:0] node3080;
	wire [15-1:0] node3081;
	wire [15-1:0] node3084;
	wire [15-1:0] node3087;
	wire [15-1:0] node3090;
	wire [15-1:0] node3092;
	wire [15-1:0] node3095;
	wire [15-1:0] node3096;
	wire [15-1:0] node3097;
	wire [15-1:0] node3098;
	wire [15-1:0] node3099;
	wire [15-1:0] node3100;
	wire [15-1:0] node3103;
	wire [15-1:0] node3104;
	wire [15-1:0] node3108;
	wire [15-1:0] node3109;
	wire [15-1:0] node3112;
	wire [15-1:0] node3115;
	wire [15-1:0] node3116;
	wire [15-1:0] node3117;
	wire [15-1:0] node3121;
	wire [15-1:0] node3122;
	wire [15-1:0] node3123;
	wire [15-1:0] node3126;
	wire [15-1:0] node3130;
	wire [15-1:0] node3131;
	wire [15-1:0] node3132;
	wire [15-1:0] node3133;
	wire [15-1:0] node3136;
	wire [15-1:0] node3139;
	wire [15-1:0] node3140;
	wire [15-1:0] node3143;
	wire [15-1:0] node3144;
	wire [15-1:0] node3148;
	wire [15-1:0] node3149;
	wire [15-1:0] node3150;
	wire [15-1:0] node3151;
	wire [15-1:0] node3154;
	wire [15-1:0] node3158;
	wire [15-1:0] node3159;
	wire [15-1:0] node3161;
	wire [15-1:0] node3164;
	wire [15-1:0] node3165;
	wire [15-1:0] node3169;
	wire [15-1:0] node3170;
	wire [15-1:0] node3171;
	wire [15-1:0] node3172;
	wire [15-1:0] node3173;
	wire [15-1:0] node3175;
	wire [15-1:0] node3179;
	wire [15-1:0] node3180;
	wire [15-1:0] node3184;
	wire [15-1:0] node3185;
	wire [15-1:0] node3186;
	wire [15-1:0] node3188;
	wire [15-1:0] node3191;
	wire [15-1:0] node3192;
	wire [15-1:0] node3196;
	wire [15-1:0] node3197;
	wire [15-1:0] node3200;
	wire [15-1:0] node3201;
	wire [15-1:0] node3205;
	wire [15-1:0] node3206;
	wire [15-1:0] node3207;
	wire [15-1:0] node3208;
	wire [15-1:0] node3209;
	wire [15-1:0] node3213;
	wire [15-1:0] node3214;
	wire [15-1:0] node3217;
	wire [15-1:0] node3220;
	wire [15-1:0] node3221;
	wire [15-1:0] node3223;
	wire [15-1:0] node3226;
	wire [15-1:0] node3227;
	wire [15-1:0] node3231;
	wire [15-1:0] node3232;
	wire [15-1:0] node3234;
	wire [15-1:0] node3237;
	wire [15-1:0] node3238;
	wire [15-1:0] node3240;
	wire [15-1:0] node3244;
	wire [15-1:0] node3245;
	wire [15-1:0] node3246;
	wire [15-1:0] node3247;
	wire [15-1:0] node3248;
	wire [15-1:0] node3249;
	wire [15-1:0] node3250;
	wire [15-1:0] node3251;
	wire [15-1:0] node3252;
	wire [15-1:0] node3256;
	wire [15-1:0] node3257;
	wire [15-1:0] node3261;
	wire [15-1:0] node3262;
	wire [15-1:0] node3263;
	wire [15-1:0] node3267;
	wire [15-1:0] node3268;
	wire [15-1:0] node3272;
	wire [15-1:0] node3273;
	wire [15-1:0] node3274;
	wire [15-1:0] node3276;
	wire [15-1:0] node3279;
	wire [15-1:0] node3280;
	wire [15-1:0] node3284;
	wire [15-1:0] node3285;
	wire [15-1:0] node3287;
	wire [15-1:0] node3290;
	wire [15-1:0] node3291;
	wire [15-1:0] node3295;
	wire [15-1:0] node3296;
	wire [15-1:0] node3297;
	wire [15-1:0] node3298;
	wire [15-1:0] node3299;
	wire [15-1:0] node3303;
	wire [15-1:0] node3306;
	wire [15-1:0] node3307;
	wire [15-1:0] node3309;
	wire [15-1:0] node3313;
	wire [15-1:0] node3314;
	wire [15-1:0] node3315;
	wire [15-1:0] node3318;
	wire [15-1:0] node3319;
	wire [15-1:0] node3322;
	wire [15-1:0] node3325;
	wire [15-1:0] node3326;
	wire [15-1:0] node3328;
	wire [15-1:0] node3331;
	wire [15-1:0] node3332;
	wire [15-1:0] node3336;
	wire [15-1:0] node3337;
	wire [15-1:0] node3338;
	wire [15-1:0] node3339;
	wire [15-1:0] node3340;
	wire [15-1:0] node3341;
	wire [15-1:0] node3344;
	wire [15-1:0] node3347;
	wire [15-1:0] node3348;
	wire [15-1:0] node3352;
	wire [15-1:0] node3353;
	wire [15-1:0] node3354;
	wire [15-1:0] node3357;
	wire [15-1:0] node3360;
	wire [15-1:0] node3363;
	wire [15-1:0] node3364;
	wire [15-1:0] node3365;
	wire [15-1:0] node3366;
	wire [15-1:0] node3369;
	wire [15-1:0] node3372;
	wire [15-1:0] node3373;
	wire [15-1:0] node3376;
	wire [15-1:0] node3379;
	wire [15-1:0] node3380;
	wire [15-1:0] node3382;
	wire [15-1:0] node3386;
	wire [15-1:0] node3387;
	wire [15-1:0] node3388;
	wire [15-1:0] node3390;
	wire [15-1:0] node3391;
	wire [15-1:0] node3395;
	wire [15-1:0] node3396;
	wire [15-1:0] node3398;
	wire [15-1:0] node3401;
	wire [15-1:0] node3402;
	wire [15-1:0] node3405;
	wire [15-1:0] node3408;
	wire [15-1:0] node3409;
	wire [15-1:0] node3411;
	wire [15-1:0] node3414;
	wire [15-1:0] node3415;
	wire [15-1:0] node3419;
	wire [15-1:0] node3420;
	wire [15-1:0] node3421;
	wire [15-1:0] node3422;
	wire [15-1:0] node3423;
	wire [15-1:0] node3424;
	wire [15-1:0] node3425;
	wire [15-1:0] node3429;
	wire [15-1:0] node3432;
	wire [15-1:0] node3433;
	wire [15-1:0] node3434;
	wire [15-1:0] node3438;
	wire [15-1:0] node3441;
	wire [15-1:0] node3442;
	wire [15-1:0] node3445;
	wire [15-1:0] node3446;
	wire [15-1:0] node3447;
	wire [15-1:0] node3452;
	wire [15-1:0] node3453;
	wire [15-1:0] node3454;
	wire [15-1:0] node3456;
	wire [15-1:0] node3459;
	wire [15-1:0] node3460;
	wire [15-1:0] node3461;
	wire [15-1:0] node3464;
	wire [15-1:0] node3467;
	wire [15-1:0] node3469;
	wire [15-1:0] node3472;
	wire [15-1:0] node3473;
	wire [15-1:0] node3474;
	wire [15-1:0] node3476;
	wire [15-1:0] node3479;
	wire [15-1:0] node3481;
	wire [15-1:0] node3484;
	wire [15-1:0] node3485;
	wire [15-1:0] node3486;
	wire [15-1:0] node3491;
	wire [15-1:0] node3492;
	wire [15-1:0] node3493;
	wire [15-1:0] node3494;
	wire [15-1:0] node3496;
	wire [15-1:0] node3498;
	wire [15-1:0] node3501;
	wire [15-1:0] node3502;
	wire [15-1:0] node3504;
	wire [15-1:0] node3507;
	wire [15-1:0] node3508;
	wire [15-1:0] node3511;
	wire [15-1:0] node3514;
	wire [15-1:0] node3515;
	wire [15-1:0] node3516;
	wire [15-1:0] node3518;
	wire [15-1:0] node3521;
	wire [15-1:0] node3524;
	wire [15-1:0] node3525;
	wire [15-1:0] node3526;
	wire [15-1:0] node3529;
	wire [15-1:0] node3532;
	wire [15-1:0] node3533;
	wire [15-1:0] node3536;
	wire [15-1:0] node3539;
	wire [15-1:0] node3540;
	wire [15-1:0] node3541;
	wire [15-1:0] node3543;
	wire [15-1:0] node3544;
	wire [15-1:0] node3547;
	wire [15-1:0] node3550;
	wire [15-1:0] node3551;
	wire [15-1:0] node3554;
	wire [15-1:0] node3555;
	wire [15-1:0] node3559;
	wire [15-1:0] node3560;
	wire [15-1:0] node3563;
	wire [15-1:0] node3564;
	wire [15-1:0] node3566;
	wire [15-1:0] node3569;
	wire [15-1:0] node3570;
	wire [15-1:0] node3573;
	wire [15-1:0] node3576;
	wire [15-1:0] node3577;
	wire [15-1:0] node3578;
	wire [15-1:0] node3579;
	wire [15-1:0] node3580;
	wire [15-1:0] node3581;
	wire [15-1:0] node3582;
	wire [15-1:0] node3583;
	wire [15-1:0] node3586;
	wire [15-1:0] node3589;
	wire [15-1:0] node3590;
	wire [15-1:0] node3594;
	wire [15-1:0] node3595;
	wire [15-1:0] node3596;
	wire [15-1:0] node3600;
	wire [15-1:0] node3601;
	wire [15-1:0] node3605;
	wire [15-1:0] node3606;
	wire [15-1:0] node3607;
	wire [15-1:0] node3609;
	wire [15-1:0] node3612;
	wire [15-1:0] node3613;
	wire [15-1:0] node3617;
	wire [15-1:0] node3618;
	wire [15-1:0] node3619;
	wire [15-1:0] node3622;
	wire [15-1:0] node3625;
	wire [15-1:0] node3626;
	wire [15-1:0] node3629;
	wire [15-1:0] node3632;
	wire [15-1:0] node3633;
	wire [15-1:0] node3634;
	wire [15-1:0] node3635;
	wire [15-1:0] node3639;
	wire [15-1:0] node3641;
	wire [15-1:0] node3644;
	wire [15-1:0] node3645;
	wire [15-1:0] node3647;
	wire [15-1:0] node3648;
	wire [15-1:0] node3652;
	wire [15-1:0] node3653;
	wire [15-1:0] node3656;
	wire [15-1:0] node3657;
	wire [15-1:0] node3660;
	wire [15-1:0] node3663;
	wire [15-1:0] node3664;
	wire [15-1:0] node3665;
	wire [15-1:0] node3666;
	wire [15-1:0] node3667;
	wire [15-1:0] node3669;
	wire [15-1:0] node3672;
	wire [15-1:0] node3674;
	wire [15-1:0] node3677;
	wire [15-1:0] node3678;
	wire [15-1:0] node3681;
	wire [15-1:0] node3683;
	wire [15-1:0] node3686;
	wire [15-1:0] node3687;
	wire [15-1:0] node3688;
	wire [15-1:0] node3689;
	wire [15-1:0] node3694;
	wire [15-1:0] node3695;
	wire [15-1:0] node3697;
	wire [15-1:0] node3701;
	wire [15-1:0] node3702;
	wire [15-1:0] node3703;
	wire [15-1:0] node3705;
	wire [15-1:0] node3707;
	wire [15-1:0] node3710;
	wire [15-1:0] node3711;
	wire [15-1:0] node3713;
	wire [15-1:0] node3717;
	wire [15-1:0] node3718;
	wire [15-1:0] node3719;
	wire [15-1:0] node3722;
	wire [15-1:0] node3724;
	wire [15-1:0] node3727;
	wire [15-1:0] node3728;
	wire [15-1:0] node3730;
	wire [15-1:0] node3733;
	wire [15-1:0] node3736;
	wire [15-1:0] node3737;
	wire [15-1:0] node3738;
	wire [15-1:0] node3739;
	wire [15-1:0] node3740;
	wire [15-1:0] node3742;
	wire [15-1:0] node3743;
	wire [15-1:0] node3747;
	wire [15-1:0] node3748;
	wire [15-1:0] node3749;
	wire [15-1:0] node3752;
	wire [15-1:0] node3755;
	wire [15-1:0] node3757;
	wire [15-1:0] node3760;
	wire [15-1:0] node3761;
	wire [15-1:0] node3762;
	wire [15-1:0] node3764;
	wire [15-1:0] node3768;
	wire [15-1:0] node3769;
	wire [15-1:0] node3770;
	wire [15-1:0] node3774;
	wire [15-1:0] node3775;
	wire [15-1:0] node3779;
	wire [15-1:0] node3780;
	wire [15-1:0] node3781;
	wire [15-1:0] node3782;
	wire [15-1:0] node3783;
	wire [15-1:0] node3787;
	wire [15-1:0] node3788;
	wire [15-1:0] node3792;
	wire [15-1:0] node3795;
	wire [15-1:0] node3796;
	wire [15-1:0] node3797;
	wire [15-1:0] node3800;
	wire [15-1:0] node3801;
	wire [15-1:0] node3804;
	wire [15-1:0] node3807;
	wire [15-1:0] node3808;
	wire [15-1:0] node3810;
	wire [15-1:0] node3813;
	wire [15-1:0] node3815;
	wire [15-1:0] node3818;
	wire [15-1:0] node3819;
	wire [15-1:0] node3820;
	wire [15-1:0] node3821;
	wire [15-1:0] node3822;
	wire [15-1:0] node3824;
	wire [15-1:0] node3828;
	wire [15-1:0] node3830;
	wire [15-1:0] node3833;
	wire [15-1:0] node3834;
	wire [15-1:0] node3835;
	wire [15-1:0] node3836;
	wire [15-1:0] node3841;
	wire [15-1:0] node3842;
	wire [15-1:0] node3843;
	wire [15-1:0] node3846;
	wire [15-1:0] node3849;
	wire [15-1:0] node3851;
	wire [15-1:0] node3854;
	wire [15-1:0] node3855;
	wire [15-1:0] node3856;
	wire [15-1:0] node3857;
	wire [15-1:0] node3858;
	wire [15-1:0] node3862;
	wire [15-1:0] node3863;
	wire [15-1:0] node3866;
	wire [15-1:0] node3869;
	wire [15-1:0] node3870;
	wire [15-1:0] node3872;
	wire [15-1:0] node3875;
	wire [15-1:0] node3877;
	wire [15-1:0] node3880;
	wire [15-1:0] node3881;
	wire [15-1:0] node3882;
	wire [15-1:0] node3885;
	wire [15-1:0] node3886;
	wire [15-1:0] node3889;
	wire [15-1:0] node3892;
	wire [15-1:0] node3893;
	wire [15-1:0] node3896;
	wire [15-1:0] node3897;
	wire [15-1:0] node3900;
	wire [15-1:0] node3903;
	wire [15-1:0] node3904;
	wire [15-1:0] node3905;
	wire [15-1:0] node3906;
	wire [15-1:0] node3907;
	wire [15-1:0] node3908;
	wire [15-1:0] node3909;
	wire [15-1:0] node3910;
	wire [15-1:0] node3911;
	wire [15-1:0] node3912;
	wire [15-1:0] node3915;
	wire [15-1:0] node3918;
	wire [15-1:0] node3919;
	wire [15-1:0] node3922;
	wire [15-1:0] node3925;
	wire [15-1:0] node3926;
	wire [15-1:0] node3929;
	wire [15-1:0] node3932;
	wire [15-1:0] node3933;
	wire [15-1:0] node3934;
	wire [15-1:0] node3936;
	wire [15-1:0] node3939;
	wire [15-1:0] node3940;
	wire [15-1:0] node3944;
	wire [15-1:0] node3945;
	wire [15-1:0] node3946;
	wire [15-1:0] node3949;
	wire [15-1:0] node3953;
	wire [15-1:0] node3954;
	wire [15-1:0] node3955;
	wire [15-1:0] node3956;
	wire [15-1:0] node3957;
	wire [15-1:0] node3961;
	wire [15-1:0] node3962;
	wire [15-1:0] node3966;
	wire [15-1:0] node3967;
	wire [15-1:0] node3970;
	wire [15-1:0] node3971;
	wire [15-1:0] node3974;
	wire [15-1:0] node3977;
	wire [15-1:0] node3978;
	wire [15-1:0] node3979;
	wire [15-1:0] node3981;
	wire [15-1:0] node3985;
	wire [15-1:0] node3986;
	wire [15-1:0] node3989;
	wire [15-1:0] node3990;
	wire [15-1:0] node3993;
	wire [15-1:0] node3996;
	wire [15-1:0] node3997;
	wire [15-1:0] node3998;
	wire [15-1:0] node3999;
	wire [15-1:0] node4000;
	wire [15-1:0] node4001;
	wire [15-1:0] node4004;
	wire [15-1:0] node4007;
	wire [15-1:0] node4008;
	wire [15-1:0] node4011;
	wire [15-1:0] node4014;
	wire [15-1:0] node4015;
	wire [15-1:0] node4016;
	wire [15-1:0] node4019;
	wire [15-1:0] node4022;
	wire [15-1:0] node4023;
	wire [15-1:0] node4027;
	wire [15-1:0] node4028;
	wire [15-1:0] node4030;
	wire [15-1:0] node4032;
	wire [15-1:0] node4035;
	wire [15-1:0] node4037;
	wire [15-1:0] node4038;
	wire [15-1:0] node4042;
	wire [15-1:0] node4043;
	wire [15-1:0] node4044;
	wire [15-1:0] node4045;
	wire [15-1:0] node4047;
	wire [15-1:0] node4051;
	wire [15-1:0] node4052;
	wire [15-1:0] node4054;
	wire [15-1:0] node4057;
	wire [15-1:0] node4058;
	wire [15-1:0] node4061;
	wire [15-1:0] node4064;
	wire [15-1:0] node4065;
	wire [15-1:0] node4066;
	wire [15-1:0] node4068;
	wire [15-1:0] node4071;
	wire [15-1:0] node4073;
	wire [15-1:0] node4076;
	wire [15-1:0] node4078;
	wire [15-1:0] node4079;
	wire [15-1:0] node4082;
	wire [15-1:0] node4085;
	wire [15-1:0] node4086;
	wire [15-1:0] node4087;
	wire [15-1:0] node4088;
	wire [15-1:0] node4089;
	wire [15-1:0] node4090;
	wire [15-1:0] node4091;
	wire [15-1:0] node4094;
	wire [15-1:0] node4097;
	wire [15-1:0] node4098;
	wire [15-1:0] node4102;
	wire [15-1:0] node4103;
	wire [15-1:0] node4104;
	wire [15-1:0] node4107;
	wire [15-1:0] node4110;
	wire [15-1:0] node4112;
	wire [15-1:0] node4115;
	wire [15-1:0] node4116;
	wire [15-1:0] node4117;
	wire [15-1:0] node4119;
	wire [15-1:0] node4123;
	wire [15-1:0] node4124;
	wire [15-1:0] node4126;
	wire [15-1:0] node4129;
	wire [15-1:0] node4131;
	wire [15-1:0] node4134;
	wire [15-1:0] node4135;
	wire [15-1:0] node4136;
	wire [15-1:0] node4138;
	wire [15-1:0] node4139;
	wire [15-1:0] node4142;
	wire [15-1:0] node4145;
	wire [15-1:0] node4146;
	wire [15-1:0] node4148;
	wire [15-1:0] node4151;
	wire [15-1:0] node4153;
	wire [15-1:0] node4156;
	wire [15-1:0] node4157;
	wire [15-1:0] node4158;
	wire [15-1:0] node4159;
	wire [15-1:0] node4163;
	wire [15-1:0] node4164;
	wire [15-1:0] node4167;
	wire [15-1:0] node4170;
	wire [15-1:0] node4171;
	wire [15-1:0] node4175;
	wire [15-1:0] node4176;
	wire [15-1:0] node4177;
	wire [15-1:0] node4178;
	wire [15-1:0] node4180;
	wire [15-1:0] node4181;
	wire [15-1:0] node4184;
	wire [15-1:0] node4187;
	wire [15-1:0] node4188;
	wire [15-1:0] node4191;
	wire [15-1:0] node4194;
	wire [15-1:0] node4195;
	wire [15-1:0] node4197;
	wire [15-1:0] node4198;
	wire [15-1:0] node4202;
	wire [15-1:0] node4204;
	wire [15-1:0] node4205;
	wire [15-1:0] node4209;
	wire [15-1:0] node4210;
	wire [15-1:0] node4211;
	wire [15-1:0] node4212;
	wire [15-1:0] node4215;
	wire [15-1:0] node4216;
	wire [15-1:0] node4219;
	wire [15-1:0] node4222;
	wire [15-1:0] node4223;
	wire [15-1:0] node4224;
	wire [15-1:0] node4227;
	wire [15-1:0] node4230;
	wire [15-1:0] node4231;
	wire [15-1:0] node4234;
	wire [15-1:0] node4237;
	wire [15-1:0] node4238;
	wire [15-1:0] node4239;
	wire [15-1:0] node4242;
	wire [15-1:0] node4243;
	wire [15-1:0] node4247;
	wire [15-1:0] node4248;
	wire [15-1:0] node4250;
	wire [15-1:0] node4253;
	wire [15-1:0] node4254;
	wire [15-1:0] node4258;
	wire [15-1:0] node4259;
	wire [15-1:0] node4260;
	wire [15-1:0] node4261;
	wire [15-1:0] node4262;
	wire [15-1:0] node4263;
	wire [15-1:0] node4264;
	wire [15-1:0] node4265;
	wire [15-1:0] node4269;
	wire [15-1:0] node4270;
	wire [15-1:0] node4274;
	wire [15-1:0] node4275;
	wire [15-1:0] node4279;
	wire [15-1:0] node4280;
	wire [15-1:0] node4281;
	wire [15-1:0] node4283;
	wire [15-1:0] node4287;
	wire [15-1:0] node4289;
	wire [15-1:0] node4290;
	wire [15-1:0] node4294;
	wire [15-1:0] node4295;
	wire [15-1:0] node4296;
	wire [15-1:0] node4297;
	wire [15-1:0] node4298;
	wire [15-1:0] node4302;
	wire [15-1:0] node4303;
	wire [15-1:0] node4307;
	wire [15-1:0] node4309;
	wire [15-1:0] node4312;
	wire [15-1:0] node4313;
	wire [15-1:0] node4315;
	wire [15-1:0] node4317;
	wire [15-1:0] node4320;
	wire [15-1:0] node4321;
	wire [15-1:0] node4322;
	wire [15-1:0] node4326;
	wire [15-1:0] node4327;
	wire [15-1:0] node4331;
	wire [15-1:0] node4332;
	wire [15-1:0] node4333;
	wire [15-1:0] node4334;
	wire [15-1:0] node4335;
	wire [15-1:0] node4336;
	wire [15-1:0] node4339;
	wire [15-1:0] node4342;
	wire [15-1:0] node4344;
	wire [15-1:0] node4347;
	wire [15-1:0] node4348;
	wire [15-1:0] node4350;
	wire [15-1:0] node4353;
	wire [15-1:0] node4354;
	wire [15-1:0] node4358;
	wire [15-1:0] node4359;
	wire [15-1:0] node4360;
	wire [15-1:0] node4361;
	wire [15-1:0] node4365;
	wire [15-1:0] node4366;
	wire [15-1:0] node4369;
	wire [15-1:0] node4372;
	wire [15-1:0] node4373;
	wire [15-1:0] node4375;
	wire [15-1:0] node4379;
	wire [15-1:0] node4380;
	wire [15-1:0] node4381;
	wire [15-1:0] node4382;
	wire [15-1:0] node4383;
	wire [15-1:0] node4386;
	wire [15-1:0] node4389;
	wire [15-1:0] node4392;
	wire [15-1:0] node4393;
	wire [15-1:0] node4394;
	wire [15-1:0] node4399;
	wire [15-1:0] node4400;
	wire [15-1:0] node4401;
	wire [15-1:0] node4405;
	wire [15-1:0] node4406;
	wire [15-1:0] node4408;
	wire [15-1:0] node4411;
	wire [15-1:0] node4414;
	wire [15-1:0] node4415;
	wire [15-1:0] node4416;
	wire [15-1:0] node4417;
	wire [15-1:0] node4418;
	wire [15-1:0] node4419;
	wire [15-1:0] node4420;
	wire [15-1:0] node4423;
	wire [15-1:0] node4426;
	wire [15-1:0] node4427;
	wire [15-1:0] node4431;
	wire [15-1:0] node4432;
	wire [15-1:0] node4434;
	wire [15-1:0] node4438;
	wire [15-1:0] node4439;
	wire [15-1:0] node4440;
	wire [15-1:0] node4443;
	wire [15-1:0] node4446;
	wire [15-1:0] node4449;
	wire [15-1:0] node4450;
	wire [15-1:0] node4451;
	wire [15-1:0] node4452;
	wire [15-1:0] node4456;
	wire [15-1:0] node4458;
	wire [15-1:0] node4459;
	wire [15-1:0] node4463;
	wire [15-1:0] node4464;
	wire [15-1:0] node4465;
	wire [15-1:0] node4466;
	wire [15-1:0] node4469;
	wire [15-1:0] node4472;
	wire [15-1:0] node4473;
	wire [15-1:0] node4476;
	wire [15-1:0] node4479;
	wire [15-1:0] node4480;
	wire [15-1:0] node4481;
	wire [15-1:0] node4484;
	wire [15-1:0] node4487;
	wire [15-1:0] node4489;
	wire [15-1:0] node4492;
	wire [15-1:0] node4493;
	wire [15-1:0] node4494;
	wire [15-1:0] node4495;
	wire [15-1:0] node4496;
	wire [15-1:0] node4500;
	wire [15-1:0] node4501;
	wire [15-1:0] node4502;
	wire [15-1:0] node4505;
	wire [15-1:0] node4508;
	wire [15-1:0] node4510;
	wire [15-1:0] node4513;
	wire [15-1:0] node4514;
	wire [15-1:0] node4516;
	wire [15-1:0] node4517;
	wire [15-1:0] node4521;
	wire [15-1:0] node4522;
	wire [15-1:0] node4523;
	wire [15-1:0] node4526;
	wire [15-1:0] node4529;
	wire [15-1:0] node4530;
	wire [15-1:0] node4533;
	wire [15-1:0] node4536;
	wire [15-1:0] node4537;
	wire [15-1:0] node4538;
	wire [15-1:0] node4539;
	wire [15-1:0] node4540;
	wire [15-1:0] node4543;
	wire [15-1:0] node4546;
	wire [15-1:0] node4549;
	wire [15-1:0] node4550;
	wire [15-1:0] node4551;
	wire [15-1:0] node4554;
	wire [15-1:0] node4558;
	wire [15-1:0] node4559;
	wire [15-1:0] node4560;
	wire [15-1:0] node4562;
	wire [15-1:0] node4565;
	wire [15-1:0] node4566;
	wire [15-1:0] node4569;
	wire [15-1:0] node4572;
	wire [15-1:0] node4573;
	wire [15-1:0] node4575;
	wire [15-1:0] node4578;
	wire [15-1:0] node4580;
	wire [15-1:0] node4583;
	wire [15-1:0] node4584;
	wire [15-1:0] node4585;
	wire [15-1:0] node4586;
	wire [15-1:0] node4587;
	wire [15-1:0] node4588;
	wire [15-1:0] node4589;
	wire [15-1:0] node4590;
	wire [15-1:0] node4591;
	wire [15-1:0] node4595;
	wire [15-1:0] node4598;
	wire [15-1:0] node4600;
	wire [15-1:0] node4601;
	wire [15-1:0] node4605;
	wire [15-1:0] node4606;
	wire [15-1:0] node4609;
	wire [15-1:0] node4612;
	wire [15-1:0] node4613;
	wire [15-1:0] node4614;
	wire [15-1:0] node4615;
	wire [15-1:0] node4616;
	wire [15-1:0] node4620;
	wire [15-1:0] node4621;
	wire [15-1:0] node4625;
	wire [15-1:0] node4627;
	wire [15-1:0] node4628;
	wire [15-1:0] node4632;
	wire [15-1:0] node4633;
	wire [15-1:0] node4634;
	wire [15-1:0] node4636;
	wire [15-1:0] node4640;
	wire [15-1:0] node4641;
	wire [15-1:0] node4643;
	wire [15-1:0] node4646;
	wire [15-1:0] node4649;
	wire [15-1:0] node4650;
	wire [15-1:0] node4651;
	wire [15-1:0] node4652;
	wire [15-1:0] node4653;
	wire [15-1:0] node4654;
	wire [15-1:0] node4658;
	wire [15-1:0] node4661;
	wire [15-1:0] node4662;
	wire [15-1:0] node4664;
	wire [15-1:0] node4668;
	wire [15-1:0] node4669;
	wire [15-1:0] node4670;
	wire [15-1:0] node4671;
	wire [15-1:0] node4675;
	wire [15-1:0] node4676;
	wire [15-1:0] node4679;
	wire [15-1:0] node4682;
	wire [15-1:0] node4684;
	wire [15-1:0] node4685;
	wire [15-1:0] node4689;
	wire [15-1:0] node4690;
	wire [15-1:0] node4691;
	wire [15-1:0] node4694;
	wire [15-1:0] node4695;
	wire [15-1:0] node4697;
	wire [15-1:0] node4701;
	wire [15-1:0] node4702;
	wire [15-1:0] node4705;
	wire [15-1:0] node4706;
	wire [15-1:0] node4707;
	wire [15-1:0] node4711;
	wire [15-1:0] node4713;
	wire [15-1:0] node4716;
	wire [15-1:0] node4717;
	wire [15-1:0] node4718;
	wire [15-1:0] node4719;
	wire [15-1:0] node4720;
	wire [15-1:0] node4721;
	wire [15-1:0] node4723;
	wire [15-1:0] node4726;
	wire [15-1:0] node4727;
	wire [15-1:0] node4730;
	wire [15-1:0] node4733;
	wire [15-1:0] node4734;
	wire [15-1:0] node4736;
	wire [15-1:0] node4739;
	wire [15-1:0] node4742;
	wire [15-1:0] node4743;
	wire [15-1:0] node4744;
	wire [15-1:0] node4748;
	wire [15-1:0] node4750;
	wire [15-1:0] node4752;
	wire [15-1:0] node4755;
	wire [15-1:0] node4756;
	wire [15-1:0] node4757;
	wire [15-1:0] node4759;
	wire [15-1:0] node4762;
	wire [15-1:0] node4763;
	wire [15-1:0] node4765;
	wire [15-1:0] node4768;
	wire [15-1:0] node4769;
	wire [15-1:0] node4773;
	wire [15-1:0] node4774;
	wire [15-1:0] node4775;
	wire [15-1:0] node4778;
	wire [15-1:0] node4780;
	wire [15-1:0] node4783;
	wire [15-1:0] node4784;
	wire [15-1:0] node4785;
	wire [15-1:0] node4788;
	wire [15-1:0] node4791;
	wire [15-1:0] node4793;
	wire [15-1:0] node4796;
	wire [15-1:0] node4797;
	wire [15-1:0] node4798;
	wire [15-1:0] node4799;
	wire [15-1:0] node4800;
	wire [15-1:0] node4801;
	wire [15-1:0] node4805;
	wire [15-1:0] node4808;
	wire [15-1:0] node4810;
	wire [15-1:0] node4811;
	wire [15-1:0] node4815;
	wire [15-1:0] node4816;
	wire [15-1:0] node4817;
	wire [15-1:0] node4818;
	wire [15-1:0] node4822;
	wire [15-1:0] node4823;
	wire [15-1:0] node4827;
	wire [15-1:0] node4828;
	wire [15-1:0] node4830;
	wire [15-1:0] node4833;
	wire [15-1:0] node4835;
	wire [15-1:0] node4838;
	wire [15-1:0] node4839;
	wire [15-1:0] node4840;
	wire [15-1:0] node4841;
	wire [15-1:0] node4843;
	wire [15-1:0] node4846;
	wire [15-1:0] node4847;
	wire [15-1:0] node4851;
	wire [15-1:0] node4852;
	wire [15-1:0] node4855;
	wire [15-1:0] node4858;
	wire [15-1:0] node4859;
	wire [15-1:0] node4861;
	wire [15-1:0] node4862;
	wire [15-1:0] node4865;
	wire [15-1:0] node4868;
	wire [15-1:0] node4869;
	wire [15-1:0] node4870;
	wire [15-1:0] node4874;
	wire [15-1:0] node4876;
	wire [15-1:0] node4879;
	wire [15-1:0] node4880;
	wire [15-1:0] node4881;
	wire [15-1:0] node4882;
	wire [15-1:0] node4883;
	wire [15-1:0] node4884;
	wire [15-1:0] node4885;
	wire [15-1:0] node4886;
	wire [15-1:0] node4891;
	wire [15-1:0] node4893;
	wire [15-1:0] node4895;
	wire [15-1:0] node4898;
	wire [15-1:0] node4899;
	wire [15-1:0] node4901;
	wire [15-1:0] node4902;
	wire [15-1:0] node4905;
	wire [15-1:0] node4908;
	wire [15-1:0] node4910;
	wire [15-1:0] node4911;
	wire [15-1:0] node4914;
	wire [15-1:0] node4917;
	wire [15-1:0] node4918;
	wire [15-1:0] node4919;
	wire [15-1:0] node4920;
	wire [15-1:0] node4923;
	wire [15-1:0] node4926;
	wire [15-1:0] node4928;
	wire [15-1:0] node4929;
	wire [15-1:0] node4932;
	wire [15-1:0] node4935;
	wire [15-1:0] node4936;
	wire [15-1:0] node4937;
	wire [15-1:0] node4939;
	wire [15-1:0] node4943;
	wire [15-1:0] node4945;
	wire [15-1:0] node4946;
	wire [15-1:0] node4949;
	wire [15-1:0] node4952;
	wire [15-1:0] node4953;
	wire [15-1:0] node4954;
	wire [15-1:0] node4955;
	wire [15-1:0] node4957;
	wire [15-1:0] node4960;
	wire [15-1:0] node4961;
	wire [15-1:0] node4962;
	wire [15-1:0] node4965;
	wire [15-1:0] node4968;
	wire [15-1:0] node4969;
	wire [15-1:0] node4973;
	wire [15-1:0] node4974;
	wire [15-1:0] node4975;
	wire [15-1:0] node4977;
	wire [15-1:0] node4980;
	wire [15-1:0] node4981;
	wire [15-1:0] node4984;
	wire [15-1:0] node4987;
	wire [15-1:0] node4988;
	wire [15-1:0] node4990;
	wire [15-1:0] node4993;
	wire [15-1:0] node4995;
	wire [15-1:0] node4998;
	wire [15-1:0] node4999;
	wire [15-1:0] node5000;
	wire [15-1:0] node5001;
	wire [15-1:0] node5003;
	wire [15-1:0] node5006;
	wire [15-1:0] node5007;
	wire [15-1:0] node5011;
	wire [15-1:0] node5012;
	wire [15-1:0] node5016;
	wire [15-1:0] node5017;
	wire [15-1:0] node5018;
	wire [15-1:0] node5019;
	wire [15-1:0] node5022;
	wire [15-1:0] node5025;
	wire [15-1:0] node5026;
	wire [15-1:0] node5029;
	wire [15-1:0] node5032;
	wire [15-1:0] node5033;
	wire [15-1:0] node5036;
	wire [15-1:0] node5038;
	wire [15-1:0] node5041;
	wire [15-1:0] node5042;
	wire [15-1:0] node5043;
	wire [15-1:0] node5044;
	wire [15-1:0] node5045;
	wire [15-1:0] node5046;
	wire [15-1:0] node5047;
	wire [15-1:0] node5051;
	wire [15-1:0] node5054;
	wire [15-1:0] node5055;
	wire [15-1:0] node5057;
	wire [15-1:0] node5060;
	wire [15-1:0] node5061;
	wire [15-1:0] node5065;
	wire [15-1:0] node5066;
	wire [15-1:0] node5067;
	wire [15-1:0] node5068;
	wire [15-1:0] node5073;
	wire [15-1:0] node5074;
	wire [15-1:0] node5076;
	wire [15-1:0] node5079;
	wire [15-1:0] node5080;
	wire [15-1:0] node5084;
	wire [15-1:0] node5085;
	wire [15-1:0] node5086;
	wire [15-1:0] node5087;
	wire [15-1:0] node5090;
	wire [15-1:0] node5091;
	wire [15-1:0] node5094;
	wire [15-1:0] node5097;
	wire [15-1:0] node5098;
	wire [15-1:0] node5100;
	wire [15-1:0] node5103;
	wire [15-1:0] node5104;
	wire [15-1:0] node5107;
	wire [15-1:0] node5110;
	wire [15-1:0] node5111;
	wire [15-1:0] node5112;
	wire [15-1:0] node5114;
	wire [15-1:0] node5117;
	wire [15-1:0] node5119;
	wire [15-1:0] node5122;
	wire [15-1:0] node5123;
	wire [15-1:0] node5127;
	wire [15-1:0] node5128;
	wire [15-1:0] node5129;
	wire [15-1:0] node5130;
	wire [15-1:0] node5131;
	wire [15-1:0] node5132;
	wire [15-1:0] node5137;
	wire [15-1:0] node5138;
	wire [15-1:0] node5139;
	wire [15-1:0] node5142;
	wire [15-1:0] node5145;
	wire [15-1:0] node5147;
	wire [15-1:0] node5150;
	wire [15-1:0] node5151;
	wire [15-1:0] node5152;
	wire [15-1:0] node5153;
	wire [15-1:0] node5157;
	wire [15-1:0] node5158;
	wire [15-1:0] node5161;
	wire [15-1:0] node5164;
	wire [15-1:0] node5165;
	wire [15-1:0] node5167;
	wire [15-1:0] node5170;
	wire [15-1:0] node5171;
	wire [15-1:0] node5174;
	wire [15-1:0] node5177;
	wire [15-1:0] node5178;
	wire [15-1:0] node5179;
	wire [15-1:0] node5180;
	wire [15-1:0] node5182;
	wire [15-1:0] node5185;
	wire [15-1:0] node5188;
	wire [15-1:0] node5190;
	wire [15-1:0] node5191;
	wire [15-1:0] node5194;
	wire [15-1:0] node5197;
	wire [15-1:0] node5198;
	wire [15-1:0] node5199;
	wire [15-1:0] node5203;
	wire [15-1:0] node5204;
	wire [15-1:0] node5205;
	wire [15-1:0] node5209;
	wire [15-1:0] node5210;
	wire [15-1:0] node5214;
	wire [15-1:0] node5215;
	wire [15-1:0] node5216;
	wire [15-1:0] node5217;
	wire [15-1:0] node5218;
	wire [15-1:0] node5219;
	wire [15-1:0] node5220;
	wire [15-1:0] node5221;
	wire [15-1:0] node5222;
	wire [15-1:0] node5223;
	wire [15-1:0] node5224;
	wire [15-1:0] node5225;
	wire [15-1:0] node5228;
	wire [15-1:0] node5232;
	wire [15-1:0] node5233;
	wire [15-1:0] node5234;
	wire [15-1:0] node5238;
	wire [15-1:0] node5239;
	wire [15-1:0] node5242;
	wire [15-1:0] node5245;
	wire [15-1:0] node5246;
	wire [15-1:0] node5248;
	wire [15-1:0] node5249;
	wire [15-1:0] node5252;
	wire [15-1:0] node5255;
	wire [15-1:0] node5257;
	wire [15-1:0] node5259;
	wire [15-1:0] node5262;
	wire [15-1:0] node5263;
	wire [15-1:0] node5264;
	wire [15-1:0] node5265;
	wire [15-1:0] node5268;
	wire [15-1:0] node5269;
	wire [15-1:0] node5273;
	wire [15-1:0] node5274;
	wire [15-1:0] node5276;
	wire [15-1:0] node5279;
	wire [15-1:0] node5280;
	wire [15-1:0] node5283;
	wire [15-1:0] node5286;
	wire [15-1:0] node5287;
	wire [15-1:0] node5288;
	wire [15-1:0] node5290;
	wire [15-1:0] node5294;
	wire [15-1:0] node5295;
	wire [15-1:0] node5296;
	wire [15-1:0] node5299;
	wire [15-1:0] node5303;
	wire [15-1:0] node5304;
	wire [15-1:0] node5305;
	wire [15-1:0] node5306;
	wire [15-1:0] node5308;
	wire [15-1:0] node5309;
	wire [15-1:0] node5313;
	wire [15-1:0] node5314;
	wire [15-1:0] node5316;
	wire [15-1:0] node5320;
	wire [15-1:0] node5321;
	wire [15-1:0] node5322;
	wire [15-1:0] node5323;
	wire [15-1:0] node5327;
	wire [15-1:0] node5328;
	wire [15-1:0] node5331;
	wire [15-1:0] node5334;
	wire [15-1:0] node5335;
	wire [15-1:0] node5337;
	wire [15-1:0] node5340;
	wire [15-1:0] node5341;
	wire [15-1:0] node5345;
	wire [15-1:0] node5346;
	wire [15-1:0] node5347;
	wire [15-1:0] node5348;
	wire [15-1:0] node5350;
	wire [15-1:0] node5353;
	wire [15-1:0] node5356;
	wire [15-1:0] node5358;
	wire [15-1:0] node5361;
	wire [15-1:0] node5362;
	wire [15-1:0] node5363;
	wire [15-1:0] node5365;
	wire [15-1:0] node5368;
	wire [15-1:0] node5371;
	wire [15-1:0] node5373;
	wire [15-1:0] node5374;
	wire [15-1:0] node5378;
	wire [15-1:0] node5379;
	wire [15-1:0] node5380;
	wire [15-1:0] node5381;
	wire [15-1:0] node5382;
	wire [15-1:0] node5383;
	wire [15-1:0] node5385;
	wire [15-1:0] node5388;
	wire [15-1:0] node5389;
	wire [15-1:0] node5392;
	wire [15-1:0] node5395;
	wire [15-1:0] node5396;
	wire [15-1:0] node5397;
	wire [15-1:0] node5400;
	wire [15-1:0] node5404;
	wire [15-1:0] node5405;
	wire [15-1:0] node5406;
	wire [15-1:0] node5407;
	wire [15-1:0] node5411;
	wire [15-1:0] node5412;
	wire [15-1:0] node5415;
	wire [15-1:0] node5418;
	wire [15-1:0] node5419;
	wire [15-1:0] node5420;
	wire [15-1:0] node5423;
	wire [15-1:0] node5426;
	wire [15-1:0] node5427;
	wire [15-1:0] node5431;
	wire [15-1:0] node5432;
	wire [15-1:0] node5433;
	wire [15-1:0] node5435;
	wire [15-1:0] node5437;
	wire [15-1:0] node5440;
	wire [15-1:0] node5441;
	wire [15-1:0] node5442;
	wire [15-1:0] node5445;
	wire [15-1:0] node5448;
	wire [15-1:0] node5450;
	wire [15-1:0] node5453;
	wire [15-1:0] node5454;
	wire [15-1:0] node5455;
	wire [15-1:0] node5458;
	wire [15-1:0] node5459;
	wire [15-1:0] node5462;
	wire [15-1:0] node5465;
	wire [15-1:0] node5467;
	wire [15-1:0] node5470;
	wire [15-1:0] node5471;
	wire [15-1:0] node5472;
	wire [15-1:0] node5473;
	wire [15-1:0] node5474;
	wire [15-1:0] node5476;
	wire [15-1:0] node5480;
	wire [15-1:0] node5481;
	wire [15-1:0] node5482;
	wire [15-1:0] node5487;
	wire [15-1:0] node5488;
	wire [15-1:0] node5489;
	wire [15-1:0] node5492;
	wire [15-1:0] node5493;
	wire [15-1:0] node5497;
	wire [15-1:0] node5498;
	wire [15-1:0] node5499;
	wire [15-1:0] node5503;
	wire [15-1:0] node5504;
	wire [15-1:0] node5508;
	wire [15-1:0] node5509;
	wire [15-1:0] node5510;
	wire [15-1:0] node5512;
	wire [15-1:0] node5513;
	wire [15-1:0] node5517;
	wire [15-1:0] node5518;
	wire [15-1:0] node5519;
	wire [15-1:0] node5522;
	wire [15-1:0] node5526;
	wire [15-1:0] node5527;
	wire [15-1:0] node5530;
	wire [15-1:0] node5531;
	wire [15-1:0] node5533;
	wire [15-1:0] node5536;
	wire [15-1:0] node5538;
	wire [15-1:0] node5541;
	wire [15-1:0] node5542;
	wire [15-1:0] node5543;
	wire [15-1:0] node5544;
	wire [15-1:0] node5545;
	wire [15-1:0] node5546;
	wire [15-1:0] node5547;
	wire [15-1:0] node5548;
	wire [15-1:0] node5551;
	wire [15-1:0] node5554;
	wire [15-1:0] node5555;
	wire [15-1:0] node5559;
	wire [15-1:0] node5560;
	wire [15-1:0] node5563;
	wire [15-1:0] node5564;
	wire [15-1:0] node5567;
	wire [15-1:0] node5570;
	wire [15-1:0] node5571;
	wire [15-1:0] node5572;
	wire [15-1:0] node5573;
	wire [15-1:0] node5576;
	wire [15-1:0] node5579;
	wire [15-1:0] node5580;
	wire [15-1:0] node5583;
	wire [15-1:0] node5586;
	wire [15-1:0] node5588;
	wire [15-1:0] node5591;
	wire [15-1:0] node5592;
	wire [15-1:0] node5593;
	wire [15-1:0] node5594;
	wire [15-1:0] node5595;
	wire [15-1:0] node5598;
	wire [15-1:0] node5601;
	wire [15-1:0] node5602;
	wire [15-1:0] node5606;
	wire [15-1:0] node5607;
	wire [15-1:0] node5608;
	wire [15-1:0] node5611;
	wire [15-1:0] node5614;
	wire [15-1:0] node5615;
	wire [15-1:0] node5619;
	wire [15-1:0] node5620;
	wire [15-1:0] node5621;
	wire [15-1:0] node5622;
	wire [15-1:0] node5625;
	wire [15-1:0] node5628;
	wire [15-1:0] node5630;
	wire [15-1:0] node5633;
	wire [15-1:0] node5635;
	wire [15-1:0] node5636;
	wire [15-1:0] node5639;
	wire [15-1:0] node5642;
	wire [15-1:0] node5643;
	wire [15-1:0] node5644;
	wire [15-1:0] node5645;
	wire [15-1:0] node5646;
	wire [15-1:0] node5647;
	wire [15-1:0] node5650;
	wire [15-1:0] node5653;
	wire [15-1:0] node5654;
	wire [15-1:0] node5658;
	wire [15-1:0] node5660;
	wire [15-1:0] node5661;
	wire [15-1:0] node5665;
	wire [15-1:0] node5666;
	wire [15-1:0] node5667;
	wire [15-1:0] node5669;
	wire [15-1:0] node5672;
	wire [15-1:0] node5673;
	wire [15-1:0] node5676;
	wire [15-1:0] node5679;
	wire [15-1:0] node5680;
	wire [15-1:0] node5682;
	wire [15-1:0] node5685;
	wire [15-1:0] node5686;
	wire [15-1:0] node5690;
	wire [15-1:0] node5691;
	wire [15-1:0] node5692;
	wire [15-1:0] node5693;
	wire [15-1:0] node5695;
	wire [15-1:0] node5699;
	wire [15-1:0] node5700;
	wire [15-1:0] node5704;
	wire [15-1:0] node5705;
	wire [15-1:0] node5706;
	wire [15-1:0] node5708;
	wire [15-1:0] node5711;
	wire [15-1:0] node5712;
	wire [15-1:0] node5715;
	wire [15-1:0] node5718;
	wire [15-1:0] node5720;
	wire [15-1:0] node5723;
	wire [15-1:0] node5724;
	wire [15-1:0] node5725;
	wire [15-1:0] node5726;
	wire [15-1:0] node5727;
	wire [15-1:0] node5728;
	wire [15-1:0] node5730;
	wire [15-1:0] node5733;
	wire [15-1:0] node5734;
	wire [15-1:0] node5738;
	wire [15-1:0] node5739;
	wire [15-1:0] node5740;
	wire [15-1:0] node5743;
	wire [15-1:0] node5746;
	wire [15-1:0] node5748;
	wire [15-1:0] node5751;
	wire [15-1:0] node5752;
	wire [15-1:0] node5753;
	wire [15-1:0] node5755;
	wire [15-1:0] node5758;
	wire [15-1:0] node5759;
	wire [15-1:0] node5763;
	wire [15-1:0] node5764;
	wire [15-1:0] node5766;
	wire [15-1:0] node5769;
	wire [15-1:0] node5772;
	wire [15-1:0] node5773;
	wire [15-1:0] node5774;
	wire [15-1:0] node5775;
	wire [15-1:0] node5777;
	wire [15-1:0] node5781;
	wire [15-1:0] node5782;
	wire [15-1:0] node5784;
	wire [15-1:0] node5787;
	wire [15-1:0] node5790;
	wire [15-1:0] node5791;
	wire [15-1:0] node5792;
	wire [15-1:0] node5795;
	wire [15-1:0] node5796;
	wire [15-1:0] node5799;
	wire [15-1:0] node5802;
	wire [15-1:0] node5803;
	wire [15-1:0] node5804;
	wire [15-1:0] node5807;
	wire [15-1:0] node5810;
	wire [15-1:0] node5813;
	wire [15-1:0] node5814;
	wire [15-1:0] node5815;
	wire [15-1:0] node5816;
	wire [15-1:0] node5817;
	wire [15-1:0] node5820;
	wire [15-1:0] node5821;
	wire [15-1:0] node5825;
	wire [15-1:0] node5826;
	wire [15-1:0] node5828;
	wire [15-1:0] node5831;
	wire [15-1:0] node5833;
	wire [15-1:0] node5836;
	wire [15-1:0] node5837;
	wire [15-1:0] node5839;
	wire [15-1:0] node5840;
	wire [15-1:0] node5844;
	wire [15-1:0] node5845;
	wire [15-1:0] node5846;
	wire [15-1:0] node5850;
	wire [15-1:0] node5851;
	wire [15-1:0] node5855;
	wire [15-1:0] node5856;
	wire [15-1:0] node5857;
	wire [15-1:0] node5858;
	wire [15-1:0] node5859;
	wire [15-1:0] node5863;
	wire [15-1:0] node5865;
	wire [15-1:0] node5868;
	wire [15-1:0] node5869;
	wire [15-1:0] node5871;
	wire [15-1:0] node5874;
	wire [15-1:0] node5875;
	wire [15-1:0] node5878;
	wire [15-1:0] node5881;
	wire [15-1:0] node5882;
	wire [15-1:0] node5883;
	wire [15-1:0] node5885;
	wire [15-1:0] node5888;
	wire [15-1:0] node5890;
	wire [15-1:0] node5893;
	wire [15-1:0] node5894;
	wire [15-1:0] node5895;
	wire [15-1:0] node5898;
	wire [15-1:0] node5901;
	wire [15-1:0] node5902;
	wire [15-1:0] node5906;
	wire [15-1:0] node5907;
	wire [15-1:0] node5908;
	wire [15-1:0] node5909;
	wire [15-1:0] node5910;
	wire [15-1:0] node5911;
	wire [15-1:0] node5912;
	wire [15-1:0] node5913;
	wire [15-1:0] node5914;
	wire [15-1:0] node5917;
	wire [15-1:0] node5921;
	wire [15-1:0] node5922;
	wire [15-1:0] node5923;
	wire [15-1:0] node5927;
	wire [15-1:0] node5930;
	wire [15-1:0] node5931;
	wire [15-1:0] node5932;
	wire [15-1:0] node5935;
	wire [15-1:0] node5937;
	wire [15-1:0] node5940;
	wire [15-1:0] node5941;
	wire [15-1:0] node5943;
	wire [15-1:0] node5947;
	wire [15-1:0] node5948;
	wire [15-1:0] node5949;
	wire [15-1:0] node5950;
	wire [15-1:0] node5954;
	wire [15-1:0] node5955;
	wire [15-1:0] node5956;
	wire [15-1:0] node5959;
	wire [15-1:0] node5962;
	wire [15-1:0] node5963;
	wire [15-1:0] node5967;
	wire [15-1:0] node5968;
	wire [15-1:0] node5969;
	wire [15-1:0] node5970;
	wire [15-1:0] node5973;
	wire [15-1:0] node5976;
	wire [15-1:0] node5978;
	wire [15-1:0] node5981;
	wire [15-1:0] node5982;
	wire [15-1:0] node5984;
	wire [15-1:0] node5987;
	wire [15-1:0] node5988;
	wire [15-1:0] node5991;
	wire [15-1:0] node5994;
	wire [15-1:0] node5995;
	wire [15-1:0] node5996;
	wire [15-1:0] node5997;
	wire [15-1:0] node5998;
	wire [15-1:0] node6001;
	wire [15-1:0] node6002;
	wire [15-1:0] node6006;
	wire [15-1:0] node6007;
	wire [15-1:0] node6008;
	wire [15-1:0] node6011;
	wire [15-1:0] node6014;
	wire [15-1:0] node6017;
	wire [15-1:0] node6018;
	wire [15-1:0] node6019;
	wire [15-1:0] node6021;
	wire [15-1:0] node6024;
	wire [15-1:0] node6026;
	wire [15-1:0] node6029;
	wire [15-1:0] node6030;
	wire [15-1:0] node6034;
	wire [15-1:0] node6035;
	wire [15-1:0] node6036;
	wire [15-1:0] node6037;
	wire [15-1:0] node6039;
	wire [15-1:0] node6043;
	wire [15-1:0] node6044;
	wire [15-1:0] node6045;
	wire [15-1:0] node6048;
	wire [15-1:0] node6051;
	wire [15-1:0] node6054;
	wire [15-1:0] node6055;
	wire [15-1:0] node6057;
	wire [15-1:0] node6058;
	wire [15-1:0] node6061;
	wire [15-1:0] node6064;
	wire [15-1:0] node6066;
	wire [15-1:0] node6069;
	wire [15-1:0] node6070;
	wire [15-1:0] node6071;
	wire [15-1:0] node6072;
	wire [15-1:0] node6073;
	wire [15-1:0] node6074;
	wire [15-1:0] node6075;
	wire [15-1:0] node6078;
	wire [15-1:0] node6081;
	wire [15-1:0] node6082;
	wire [15-1:0] node6086;
	wire [15-1:0] node6087;
	wire [15-1:0] node6091;
	wire [15-1:0] node6092;
	wire [15-1:0] node6094;
	wire [15-1:0] node6097;
	wire [15-1:0] node6098;
	wire [15-1:0] node6099;
	wire [15-1:0] node6103;
	wire [15-1:0] node6104;
	wire [15-1:0] node6108;
	wire [15-1:0] node6109;
	wire [15-1:0] node6110;
	wire [15-1:0] node6111;
	wire [15-1:0] node6115;
	wire [15-1:0] node6116;
	wire [15-1:0] node6119;
	wire [15-1:0] node6120;
	wire [15-1:0] node6124;
	wire [15-1:0] node6125;
	wire [15-1:0] node6126;
	wire [15-1:0] node6128;
	wire [15-1:0] node6132;
	wire [15-1:0] node6133;
	wire [15-1:0] node6135;
	wire [15-1:0] node6139;
	wire [15-1:0] node6140;
	wire [15-1:0] node6141;
	wire [15-1:0] node6142;
	wire [15-1:0] node6143;
	wire [15-1:0] node6146;
	wire [15-1:0] node6148;
	wire [15-1:0] node6151;
	wire [15-1:0] node6152;
	wire [15-1:0] node6153;
	wire [15-1:0] node6156;
	wire [15-1:0] node6160;
	wire [15-1:0] node6161;
	wire [15-1:0] node6162;
	wire [15-1:0] node6164;
	wire [15-1:0] node6167;
	wire [15-1:0] node6168;
	wire [15-1:0] node6171;
	wire [15-1:0] node6174;
	wire [15-1:0] node6175;
	wire [15-1:0] node6176;
	wire [15-1:0] node6180;
	wire [15-1:0] node6182;
	wire [15-1:0] node6185;
	wire [15-1:0] node6186;
	wire [15-1:0] node6187;
	wire [15-1:0] node6189;
	wire [15-1:0] node6190;
	wire [15-1:0] node6194;
	wire [15-1:0] node6195;
	wire [15-1:0] node6196;
	wire [15-1:0] node6199;
	wire [15-1:0] node6202;
	wire [15-1:0] node6203;
	wire [15-1:0] node6207;
	wire [15-1:0] node6208;
	wire [15-1:0] node6209;
	wire [15-1:0] node6211;
	wire [15-1:0] node6215;
	wire [15-1:0] node6216;
	wire [15-1:0] node6218;
	wire [15-1:0] node6222;
	wire [15-1:0] node6223;
	wire [15-1:0] node6224;
	wire [15-1:0] node6225;
	wire [15-1:0] node6226;
	wire [15-1:0] node6227;
	wire [15-1:0] node6228;
	wire [15-1:0] node6229;
	wire [15-1:0] node6233;
	wire [15-1:0] node6234;
	wire [15-1:0] node6238;
	wire [15-1:0] node6239;
	wire [15-1:0] node6240;
	wire [15-1:0] node6244;
	wire [15-1:0] node6245;
	wire [15-1:0] node6249;
	wire [15-1:0] node6250;
	wire [15-1:0] node6251;
	wire [15-1:0] node6252;
	wire [15-1:0] node6256;
	wire [15-1:0] node6258;
	wire [15-1:0] node6261;
	wire [15-1:0] node6262;
	wire [15-1:0] node6263;
	wire [15-1:0] node6267;
	wire [15-1:0] node6268;
	wire [15-1:0] node6272;
	wire [15-1:0] node6273;
	wire [15-1:0] node6274;
	wire [15-1:0] node6276;
	wire [15-1:0] node6277;
	wire [15-1:0] node6281;
	wire [15-1:0] node6282;
	wire [15-1:0] node6283;
	wire [15-1:0] node6286;
	wire [15-1:0] node6289;
	wire [15-1:0] node6290;
	wire [15-1:0] node6293;
	wire [15-1:0] node6296;
	wire [15-1:0] node6297;
	wire [15-1:0] node6298;
	wire [15-1:0] node6300;
	wire [15-1:0] node6303;
	wire [15-1:0] node6305;
	wire [15-1:0] node6308;
	wire [15-1:0] node6309;
	wire [15-1:0] node6310;
	wire [15-1:0] node6313;
	wire [15-1:0] node6317;
	wire [15-1:0] node6318;
	wire [15-1:0] node6319;
	wire [15-1:0] node6320;
	wire [15-1:0] node6321;
	wire [15-1:0] node6322;
	wire [15-1:0] node6325;
	wire [15-1:0] node6328;
	wire [15-1:0] node6329;
	wire [15-1:0] node6333;
	wire [15-1:0] node6334;
	wire [15-1:0] node6337;
	wire [15-1:0] node6338;
	wire [15-1:0] node6342;
	wire [15-1:0] node6343;
	wire [15-1:0] node6344;
	wire [15-1:0] node6346;
	wire [15-1:0] node6349;
	wire [15-1:0] node6350;
	wire [15-1:0] node6354;
	wire [15-1:0] node6356;
	wire [15-1:0] node6357;
	wire [15-1:0] node6361;
	wire [15-1:0] node6362;
	wire [15-1:0] node6363;
	wire [15-1:0] node6364;
	wire [15-1:0] node6366;
	wire [15-1:0] node6370;
	wire [15-1:0] node6371;
	wire [15-1:0] node6374;
	wire [15-1:0] node6375;
	wire [15-1:0] node6378;
	wire [15-1:0] node6381;
	wire [15-1:0] node6382;
	wire [15-1:0] node6383;
	wire [15-1:0] node6384;
	wire [15-1:0] node6389;
	wire [15-1:0] node6390;
	wire [15-1:0] node6391;
	wire [15-1:0] node6394;
	wire [15-1:0] node6398;
	wire [15-1:0] node6399;
	wire [15-1:0] node6400;
	wire [15-1:0] node6401;
	wire [15-1:0] node6402;
	wire [15-1:0] node6404;
	wire [15-1:0] node6407;
	wire [15-1:0] node6408;
	wire [15-1:0] node6409;
	wire [15-1:0] node6413;
	wire [15-1:0] node6416;
	wire [15-1:0] node6417;
	wire [15-1:0] node6418;
	wire [15-1:0] node6420;
	wire [15-1:0] node6423;
	wire [15-1:0] node6424;
	wire [15-1:0] node6428;
	wire [15-1:0] node6429;
	wire [15-1:0] node6430;
	wire [15-1:0] node6434;
	wire [15-1:0] node6435;
	wire [15-1:0] node6439;
	wire [15-1:0] node6440;
	wire [15-1:0] node6441;
	wire [15-1:0] node6442;
	wire [15-1:0] node6443;
	wire [15-1:0] node6446;
	wire [15-1:0] node6449;
	wire [15-1:0] node6451;
	wire [15-1:0] node6454;
	wire [15-1:0] node6455;
	wire [15-1:0] node6457;
	wire [15-1:0] node6460;
	wire [15-1:0] node6462;
	wire [15-1:0] node6465;
	wire [15-1:0] node6466;
	wire [15-1:0] node6467;
	wire [15-1:0] node6471;
	wire [15-1:0] node6472;
	wire [15-1:0] node6475;
	wire [15-1:0] node6476;
	wire [15-1:0] node6480;
	wire [15-1:0] node6481;
	wire [15-1:0] node6482;
	wire [15-1:0] node6483;
	wire [15-1:0] node6484;
	wire [15-1:0] node6485;
	wire [15-1:0] node6490;
	wire [15-1:0] node6491;
	wire [15-1:0] node6492;
	wire [15-1:0] node6496;
	wire [15-1:0] node6498;
	wire [15-1:0] node6501;
	wire [15-1:0] node6502;
	wire [15-1:0] node6503;
	wire [15-1:0] node6506;
	wire [15-1:0] node6507;
	wire [15-1:0] node6511;
	wire [15-1:0] node6512;
	wire [15-1:0] node6514;
	wire [15-1:0] node6517;
	wire [15-1:0] node6518;
	wire [15-1:0] node6521;
	wire [15-1:0] node6524;
	wire [15-1:0] node6525;
	wire [15-1:0] node6526;
	wire [15-1:0] node6528;
	wire [15-1:0] node6529;
	wire [15-1:0] node6533;
	wire [15-1:0] node6535;
	wire [15-1:0] node6537;
	wire [15-1:0] node6540;
	wire [15-1:0] node6541;
	wire [15-1:0] node6542;
	wire [15-1:0] node6543;
	wire [15-1:0] node6546;
	wire [15-1:0] node6549;
	wire [15-1:0] node6550;
	wire [15-1:0] node6553;
	wire [15-1:0] node6556;
	wire [15-1:0] node6557;
	wire [15-1:0] node6559;
	wire [15-1:0] node6562;
	wire [15-1:0] node6563;
	wire [15-1:0] node6567;
	wire [15-1:0] node6568;
	wire [15-1:0] node6569;
	wire [15-1:0] node6570;
	wire [15-1:0] node6571;
	wire [15-1:0] node6572;
	wire [15-1:0] node6573;
	wire [15-1:0] node6574;
	wire [15-1:0] node6575;
	wire [15-1:0] node6576;
	wire [15-1:0] node6579;
	wire [15-1:0] node6582;
	wire [15-1:0] node6583;
	wire [15-1:0] node6587;
	wire [15-1:0] node6588;
	wire [15-1:0] node6589;
	wire [15-1:0] node6592;
	wire [15-1:0] node6595;
	wire [15-1:0] node6598;
	wire [15-1:0] node6599;
	wire [15-1:0] node6600;
	wire [15-1:0] node6602;
	wire [15-1:0] node6605;
	wire [15-1:0] node6607;
	wire [15-1:0] node6610;
	wire [15-1:0] node6612;
	wire [15-1:0] node6613;
	wire [15-1:0] node6616;
	wire [15-1:0] node6619;
	wire [15-1:0] node6620;
	wire [15-1:0] node6621;
	wire [15-1:0] node6622;
	wire [15-1:0] node6624;
	wire [15-1:0] node6627;
	wire [15-1:0] node6628;
	wire [15-1:0] node6632;
	wire [15-1:0] node6634;
	wire [15-1:0] node6635;
	wire [15-1:0] node6639;
	wire [15-1:0] node6640;
	wire [15-1:0] node6641;
	wire [15-1:0] node6642;
	wire [15-1:0] node6645;
	wire [15-1:0] node6648;
	wire [15-1:0] node6649;
	wire [15-1:0] node6653;
	wire [15-1:0] node6655;
	wire [15-1:0] node6656;
	wire [15-1:0] node6659;
	wire [15-1:0] node6662;
	wire [15-1:0] node6663;
	wire [15-1:0] node6664;
	wire [15-1:0] node6665;
	wire [15-1:0] node6666;
	wire [15-1:0] node6669;
	wire [15-1:0] node6670;
	wire [15-1:0] node6673;
	wire [15-1:0] node6676;
	wire [15-1:0] node6677;
	wire [15-1:0] node6679;
	wire [15-1:0] node6682;
	wire [15-1:0] node6683;
	wire [15-1:0] node6686;
	wire [15-1:0] node6689;
	wire [15-1:0] node6690;
	wire [15-1:0] node6692;
	wire [15-1:0] node6693;
	wire [15-1:0] node6697;
	wire [15-1:0] node6698;
	wire [15-1:0] node6699;
	wire [15-1:0] node6702;
	wire [15-1:0] node6705;
	wire [15-1:0] node6708;
	wire [15-1:0] node6709;
	wire [15-1:0] node6710;
	wire [15-1:0] node6711;
	wire [15-1:0] node6713;
	wire [15-1:0] node6716;
	wire [15-1:0] node6717;
	wire [15-1:0] node6721;
	wire [15-1:0] node6722;
	wire [15-1:0] node6723;
	wire [15-1:0] node6726;
	wire [15-1:0] node6729;
	wire [15-1:0] node6730;
	wire [15-1:0] node6734;
	wire [15-1:0] node6735;
	wire [15-1:0] node6736;
	wire [15-1:0] node6739;
	wire [15-1:0] node6741;
	wire [15-1:0] node6744;
	wire [15-1:0] node6745;
	wire [15-1:0] node6748;
	wire [15-1:0] node6749;
	wire [15-1:0] node6752;
	wire [15-1:0] node6755;
	wire [15-1:0] node6756;
	wire [15-1:0] node6757;
	wire [15-1:0] node6758;
	wire [15-1:0] node6759;
	wire [15-1:0] node6761;
	wire [15-1:0] node6762;
	wire [15-1:0] node6765;
	wire [15-1:0] node6768;
	wire [15-1:0] node6770;
	wire [15-1:0] node6772;
	wire [15-1:0] node6775;
	wire [15-1:0] node6776;
	wire [15-1:0] node6778;
	wire [15-1:0] node6779;
	wire [15-1:0] node6783;
	wire [15-1:0] node6784;
	wire [15-1:0] node6786;
	wire [15-1:0] node6789;
	wire [15-1:0] node6792;
	wire [15-1:0] node6793;
	wire [15-1:0] node6794;
	wire [15-1:0] node6795;
	wire [15-1:0] node6796;
	wire [15-1:0] node6800;
	wire [15-1:0] node6802;
	wire [15-1:0] node6805;
	wire [15-1:0] node6806;
	wire [15-1:0] node6808;
	wire [15-1:0] node6812;
	wire [15-1:0] node6813;
	wire [15-1:0] node6814;
	wire [15-1:0] node6815;
	wire [15-1:0] node6818;
	wire [15-1:0] node6822;
	wire [15-1:0] node6823;
	wire [15-1:0] node6825;
	wire [15-1:0] node6828;
	wire [15-1:0] node6831;
	wire [15-1:0] node6832;
	wire [15-1:0] node6833;
	wire [15-1:0] node6834;
	wire [15-1:0] node6835;
	wire [15-1:0] node6836;
	wire [15-1:0] node6841;
	wire [15-1:0] node6842;
	wire [15-1:0] node6843;
	wire [15-1:0] node6847;
	wire [15-1:0] node6849;
	wire [15-1:0] node6852;
	wire [15-1:0] node6853;
	wire [15-1:0] node6854;
	wire [15-1:0] node6855;
	wire [15-1:0] node6858;
	wire [15-1:0] node6861;
	wire [15-1:0] node6863;
	wire [15-1:0] node6866;
	wire [15-1:0] node6868;
	wire [15-1:0] node6870;
	wire [15-1:0] node6873;
	wire [15-1:0] node6874;
	wire [15-1:0] node6876;
	wire [15-1:0] node6877;
	wire [15-1:0] node6879;
	wire [15-1:0] node6882;
	wire [15-1:0] node6883;
	wire [15-1:0] node6887;
	wire [15-1:0] node6888;
	wire [15-1:0] node6889;
	wire [15-1:0] node6891;
	wire [15-1:0] node6895;
	wire [15-1:0] node6896;
	wire [15-1:0] node6897;
	wire [15-1:0] node6900;
	wire [15-1:0] node6904;
	wire [15-1:0] node6905;
	wire [15-1:0] node6906;
	wire [15-1:0] node6907;
	wire [15-1:0] node6908;
	wire [15-1:0] node6909;
	wire [15-1:0] node6910;
	wire [15-1:0] node6911;
	wire [15-1:0] node6914;
	wire [15-1:0] node6917;
	wire [15-1:0] node6918;
	wire [15-1:0] node6921;
	wire [15-1:0] node6924;
	wire [15-1:0] node6925;
	wire [15-1:0] node6926;
	wire [15-1:0] node6930;
	wire [15-1:0] node6933;
	wire [15-1:0] node6934;
	wire [15-1:0] node6935;
	wire [15-1:0] node6938;
	wire [15-1:0] node6939;
	wire [15-1:0] node6942;
	wire [15-1:0] node6945;
	wire [15-1:0] node6946;
	wire [15-1:0] node6948;
	wire [15-1:0] node6952;
	wire [15-1:0] node6953;
	wire [15-1:0] node6954;
	wire [15-1:0] node6955;
	wire [15-1:0] node6956;
	wire [15-1:0] node6960;
	wire [15-1:0] node6963;
	wire [15-1:0] node6964;
	wire [15-1:0] node6966;
	wire [15-1:0] node6970;
	wire [15-1:0] node6971;
	wire [15-1:0] node6972;
	wire [15-1:0] node6973;
	wire [15-1:0] node6977;
	wire [15-1:0] node6978;
	wire [15-1:0] node6982;
	wire [15-1:0] node6983;
	wire [15-1:0] node6984;
	wire [15-1:0] node6988;
	wire [15-1:0] node6991;
	wire [15-1:0] node6992;
	wire [15-1:0] node6993;
	wire [15-1:0] node6994;
	wire [15-1:0] node6996;
	wire [15-1:0] node6998;
	wire [15-1:0] node7001;
	wire [15-1:0] node7002;
	wire [15-1:0] node7003;
	wire [15-1:0] node7006;
	wire [15-1:0] node7009;
	wire [15-1:0] node7011;
	wire [15-1:0] node7014;
	wire [15-1:0] node7015;
	wire [15-1:0] node7016;
	wire [15-1:0] node7018;
	wire [15-1:0] node7021;
	wire [15-1:0] node7022;
	wire [15-1:0] node7025;
	wire [15-1:0] node7028;
	wire [15-1:0] node7029;
	wire [15-1:0] node7030;
	wire [15-1:0] node7034;
	wire [15-1:0] node7036;
	wire [15-1:0] node7039;
	wire [15-1:0] node7040;
	wire [15-1:0] node7041;
	wire [15-1:0] node7043;
	wire [15-1:0] node7046;
	wire [15-1:0] node7048;
	wire [15-1:0] node7049;
	wire [15-1:0] node7053;
	wire [15-1:0] node7054;
	wire [15-1:0] node7055;
	wire [15-1:0] node7057;
	wire [15-1:0] node7060;
	wire [15-1:0] node7061;
	wire [15-1:0] node7064;
	wire [15-1:0] node7067;
	wire [15-1:0] node7069;
	wire [15-1:0] node7071;
	wire [15-1:0] node7074;
	wire [15-1:0] node7075;
	wire [15-1:0] node7076;
	wire [15-1:0] node7077;
	wire [15-1:0] node7078;
	wire [15-1:0] node7079;
	wire [15-1:0] node7080;
	wire [15-1:0] node7084;
	wire [15-1:0] node7085;
	wire [15-1:0] node7089;
	wire [15-1:0] node7091;
	wire [15-1:0] node7093;
	wire [15-1:0] node7096;
	wire [15-1:0] node7097;
	wire [15-1:0] node7098;
	wire [15-1:0] node7099;
	wire [15-1:0] node7102;
	wire [15-1:0] node7105;
	wire [15-1:0] node7106;
	wire [15-1:0] node7110;
	wire [15-1:0] node7111;
	wire [15-1:0] node7113;
	wire [15-1:0] node7116;
	wire [15-1:0] node7117;
	wire [15-1:0] node7120;
	wire [15-1:0] node7123;
	wire [15-1:0] node7124;
	wire [15-1:0] node7125;
	wire [15-1:0] node7126;
	wire [15-1:0] node7128;
	wire [15-1:0] node7131;
	wire [15-1:0] node7132;
	wire [15-1:0] node7135;
	wire [15-1:0] node7138;
	wire [15-1:0] node7139;
	wire [15-1:0] node7141;
	wire [15-1:0] node7144;
	wire [15-1:0] node7145;
	wire [15-1:0] node7149;
	wire [15-1:0] node7150;
	wire [15-1:0] node7151;
	wire [15-1:0] node7155;
	wire [15-1:0] node7157;
	wire [15-1:0] node7158;
	wire [15-1:0] node7162;
	wire [15-1:0] node7163;
	wire [15-1:0] node7164;
	wire [15-1:0] node7165;
	wire [15-1:0] node7166;
	wire [15-1:0] node7167;
	wire [15-1:0] node7171;
	wire [15-1:0] node7172;
	wire [15-1:0] node7176;
	wire [15-1:0] node7177;
	wire [15-1:0] node7180;
	wire [15-1:0] node7182;
	wire [15-1:0] node7185;
	wire [15-1:0] node7186;
	wire [15-1:0] node7187;
	wire [15-1:0] node7189;
	wire [15-1:0] node7193;
	wire [15-1:0] node7194;
	wire [15-1:0] node7195;
	wire [15-1:0] node7198;
	wire [15-1:0] node7202;
	wire [15-1:0] node7203;
	wire [15-1:0] node7204;
	wire [15-1:0] node7205;
	wire [15-1:0] node7207;
	wire [15-1:0] node7211;
	wire [15-1:0] node7212;
	wire [15-1:0] node7213;
	wire [15-1:0] node7216;
	wire [15-1:0] node7219;
	wire [15-1:0] node7220;
	wire [15-1:0] node7223;
	wire [15-1:0] node7226;
	wire [15-1:0] node7227;
	wire [15-1:0] node7228;
	wire [15-1:0] node7229;
	wire [15-1:0] node7232;
	wire [15-1:0] node7236;
	wire [15-1:0] node7237;
	wire [15-1:0] node7240;
	wire [15-1:0] node7241;
	wire [15-1:0] node7245;
	wire [15-1:0] node7246;
	wire [15-1:0] node7247;
	wire [15-1:0] node7248;
	wire [15-1:0] node7249;
	wire [15-1:0] node7250;
	wire [15-1:0] node7251;
	wire [15-1:0] node7252;
	wire [15-1:0] node7253;
	wire [15-1:0] node7256;
	wire [15-1:0] node7259;
	wire [15-1:0] node7262;
	wire [15-1:0] node7263;
	wire [15-1:0] node7264;
	wire [15-1:0] node7268;
	wire [15-1:0] node7269;
	wire [15-1:0] node7272;
	wire [15-1:0] node7275;
	wire [15-1:0] node7276;
	wire [15-1:0] node7278;
	wire [15-1:0] node7279;
	wire [15-1:0] node7283;
	wire [15-1:0] node7284;
	wire [15-1:0] node7285;
	wire [15-1:0] node7289;
	wire [15-1:0] node7291;
	wire [15-1:0] node7294;
	wire [15-1:0] node7295;
	wire [15-1:0] node7296;
	wire [15-1:0] node7297;
	wire [15-1:0] node7298;
	wire [15-1:0] node7303;
	wire [15-1:0] node7305;
	wire [15-1:0] node7306;
	wire [15-1:0] node7310;
	wire [15-1:0] node7311;
	wire [15-1:0] node7314;
	wire [15-1:0] node7315;
	wire [15-1:0] node7317;
	wire [15-1:0] node7320;
	wire [15-1:0] node7323;
	wire [15-1:0] node7324;
	wire [15-1:0] node7325;
	wire [15-1:0] node7326;
	wire [15-1:0] node7327;
	wire [15-1:0] node7331;
	wire [15-1:0] node7333;
	wire [15-1:0] node7336;
	wire [15-1:0] node7337;
	wire [15-1:0] node7339;
	wire [15-1:0] node7340;
	wire [15-1:0] node7343;
	wire [15-1:0] node7346;
	wire [15-1:0] node7347;
	wire [15-1:0] node7348;
	wire [15-1:0] node7352;
	wire [15-1:0] node7355;
	wire [15-1:0] node7356;
	wire [15-1:0] node7357;
	wire [15-1:0] node7358;
	wire [15-1:0] node7360;
	wire [15-1:0] node7363;
	wire [15-1:0] node7364;
	wire [15-1:0] node7368;
	wire [15-1:0] node7369;
	wire [15-1:0] node7371;
	wire [15-1:0] node7374;
	wire [15-1:0] node7375;
	wire [15-1:0] node7379;
	wire [15-1:0] node7380;
	wire [15-1:0] node7382;
	wire [15-1:0] node7383;
	wire [15-1:0] node7387;
	wire [15-1:0] node7388;
	wire [15-1:0] node7391;
	wire [15-1:0] node7392;
	wire [15-1:0] node7395;
	wire [15-1:0] node7398;
	wire [15-1:0] node7399;
	wire [15-1:0] node7400;
	wire [15-1:0] node7401;
	wire [15-1:0] node7402;
	wire [15-1:0] node7403;
	wire [15-1:0] node7404;
	wire [15-1:0] node7407;
	wire [15-1:0] node7410;
	wire [15-1:0] node7412;
	wire [15-1:0] node7415;
	wire [15-1:0] node7417;
	wire [15-1:0] node7420;
	wire [15-1:0] node7421;
	wire [15-1:0] node7422;
	wire [15-1:0] node7423;
	wire [15-1:0] node7428;
	wire [15-1:0] node7430;
	wire [15-1:0] node7433;
	wire [15-1:0] node7434;
	wire [15-1:0] node7435;
	wire [15-1:0] node7436;
	wire [15-1:0] node7437;
	wire [15-1:0] node7441;
	wire [15-1:0] node7442;
	wire [15-1:0] node7446;
	wire [15-1:0] node7447;
	wire [15-1:0] node7449;
	wire [15-1:0] node7452;
	wire [15-1:0] node7455;
	wire [15-1:0] node7456;
	wire [15-1:0] node7457;
	wire [15-1:0] node7459;
	wire [15-1:0] node7462;
	wire [15-1:0] node7463;
	wire [15-1:0] node7466;
	wire [15-1:0] node7469;
	wire [15-1:0] node7470;
	wire [15-1:0] node7473;
	wire [15-1:0] node7475;
	wire [15-1:0] node7478;
	wire [15-1:0] node7479;
	wire [15-1:0] node7480;
	wire [15-1:0] node7481;
	wire [15-1:0] node7482;
	wire [15-1:0] node7483;
	wire [15-1:0] node7486;
	wire [15-1:0] node7489;
	wire [15-1:0] node7491;
	wire [15-1:0] node7494;
	wire [15-1:0] node7495;
	wire [15-1:0] node7498;
	wire [15-1:0] node7500;
	wire [15-1:0] node7503;
	wire [15-1:0] node7504;
	wire [15-1:0] node7505;
	wire [15-1:0] node7507;
	wire [15-1:0] node7510;
	wire [15-1:0] node7511;
	wire [15-1:0] node7514;
	wire [15-1:0] node7517;
	wire [15-1:0] node7519;
	wire [15-1:0] node7520;
	wire [15-1:0] node7523;
	wire [15-1:0] node7526;
	wire [15-1:0] node7527;
	wire [15-1:0] node7528;
	wire [15-1:0] node7529;
	wire [15-1:0] node7530;
	wire [15-1:0] node7534;
	wire [15-1:0] node7536;
	wire [15-1:0] node7539;
	wire [15-1:0] node7541;
	wire [15-1:0] node7544;
	wire [15-1:0] node7545;
	wire [15-1:0] node7546;
	wire [15-1:0] node7548;
	wire [15-1:0] node7551;
	wire [15-1:0] node7553;
	wire [15-1:0] node7556;
	wire [15-1:0] node7557;
	wire [15-1:0] node7558;
	wire [15-1:0] node7561;
	wire [15-1:0] node7564;
	wire [15-1:0] node7566;
	wire [15-1:0] node7569;
	wire [15-1:0] node7570;
	wire [15-1:0] node7571;
	wire [15-1:0] node7572;
	wire [15-1:0] node7573;
	wire [15-1:0] node7574;
	wire [15-1:0] node7575;
	wire [15-1:0] node7577;
	wire [15-1:0] node7580;
	wire [15-1:0] node7582;
	wire [15-1:0] node7585;
	wire [15-1:0] node7586;
	wire [15-1:0] node7587;
	wire [15-1:0] node7592;
	wire [15-1:0] node7594;
	wire [15-1:0] node7597;
	wire [15-1:0] node7598;
	wire [15-1:0] node7599;
	wire [15-1:0] node7600;
	wire [15-1:0] node7602;
	wire [15-1:0] node7605;
	wire [15-1:0] node7608;
	wire [15-1:0] node7609;
	wire [15-1:0] node7611;
	wire [15-1:0] node7614;
	wire [15-1:0] node7617;
	wire [15-1:0] node7618;
	wire [15-1:0] node7620;
	wire [15-1:0] node7621;
	wire [15-1:0] node7624;
	wire [15-1:0] node7627;
	wire [15-1:0] node7629;
	wire [15-1:0] node7630;
	wire [15-1:0] node7634;
	wire [15-1:0] node7635;
	wire [15-1:0] node7636;
	wire [15-1:0] node7637;
	wire [15-1:0] node7638;
	wire [15-1:0] node7642;
	wire [15-1:0] node7645;
	wire [15-1:0] node7646;
	wire [15-1:0] node7648;
	wire [15-1:0] node7649;
	wire [15-1:0] node7653;
	wire [15-1:0] node7655;
	wire [15-1:0] node7656;
	wire [15-1:0] node7660;
	wire [15-1:0] node7661;
	wire [15-1:0] node7662;
	wire [15-1:0] node7663;
	wire [15-1:0] node7666;
	wire [15-1:0] node7669;
	wire [15-1:0] node7671;
	wire [15-1:0] node7672;
	wire [15-1:0] node7675;
	wire [15-1:0] node7678;
	wire [15-1:0] node7679;
	wire [15-1:0] node7680;
	wire [15-1:0] node7684;
	wire [15-1:0] node7685;
	wire [15-1:0] node7686;
	wire [15-1:0] node7689;
	wire [15-1:0] node7692;
	wire [15-1:0] node7693;
	wire [15-1:0] node7696;
	wire [15-1:0] node7699;
	wire [15-1:0] node7700;
	wire [15-1:0] node7701;
	wire [15-1:0] node7702;
	wire [15-1:0] node7703;
	wire [15-1:0] node7704;
	wire [15-1:0] node7705;
	wire [15-1:0] node7708;
	wire [15-1:0] node7711;
	wire [15-1:0] node7714;
	wire [15-1:0] node7715;
	wire [15-1:0] node7718;
	wire [15-1:0] node7719;
	wire [15-1:0] node7723;
	wire [15-1:0] node7724;
	wire [15-1:0] node7725;
	wire [15-1:0] node7726;
	wire [15-1:0] node7729;
	wire [15-1:0] node7732;
	wire [15-1:0] node7735;
	wire [15-1:0] node7736;
	wire [15-1:0] node7737;
	wire [15-1:0] node7741;
	wire [15-1:0] node7743;
	wire [15-1:0] node7746;
	wire [15-1:0] node7747;
	wire [15-1:0] node7748;
	wire [15-1:0] node7749;
	wire [15-1:0] node7750;
	wire [15-1:0] node7755;
	wire [15-1:0] node7756;
	wire [15-1:0] node7759;
	wire [15-1:0] node7760;
	wire [15-1:0] node7763;
	wire [15-1:0] node7766;
	wire [15-1:0] node7767;
	wire [15-1:0] node7768;
	wire [15-1:0] node7770;
	wire [15-1:0] node7773;
	wire [15-1:0] node7775;
	wire [15-1:0] node7778;
	wire [15-1:0] node7779;
	wire [15-1:0] node7780;
	wire [15-1:0] node7783;
	wire [15-1:0] node7786;
	wire [15-1:0] node7787;
	wire [15-1:0] node7790;
	wire [15-1:0] node7793;
	wire [15-1:0] node7794;
	wire [15-1:0] node7795;
	wire [15-1:0] node7796;
	wire [15-1:0] node7797;
	wire [15-1:0] node7798;
	wire [15-1:0] node7801;
	wire [15-1:0] node7804;
	wire [15-1:0] node7805;
	wire [15-1:0] node7809;
	wire [15-1:0] node7810;
	wire [15-1:0] node7811;
	wire [15-1:0] node7815;
	wire [15-1:0] node7817;
	wire [15-1:0] node7820;
	wire [15-1:0] node7821;
	wire [15-1:0] node7822;
	wire [15-1:0] node7824;
	wire [15-1:0] node7827;
	wire [15-1:0] node7829;
	wire [15-1:0] node7832;
	wire [15-1:0] node7833;
	wire [15-1:0] node7834;
	wire [15-1:0] node7838;
	wire [15-1:0] node7841;
	wire [15-1:0] node7842;
	wire [15-1:0] node7843;
	wire [15-1:0] node7844;
	wire [15-1:0] node7845;
	wire [15-1:0] node7848;
	wire [15-1:0] node7851;
	wire [15-1:0] node7852;
	wire [15-1:0] node7855;
	wire [15-1:0] node7858;
	wire [15-1:0] node7859;
	wire [15-1:0] node7861;
	wire [15-1:0] node7864;
	wire [15-1:0] node7865;
	wire [15-1:0] node7868;
	wire [15-1:0] node7871;
	wire [15-1:0] node7872;
	wire [15-1:0] node7873;
	wire [15-1:0] node7875;
	wire [15-1:0] node7878;
	wire [15-1:0] node7879;
	wire [15-1:0] node7883;
	wire [15-1:0] node7884;
	wire [15-1:0] node7887;
	wire [15-1:0] node7889;
	wire [15-1:0] node7892;
	wire [15-1:0] node7893;
	wire [15-1:0] node7894;
	wire [15-1:0] node7895;
	wire [15-1:0] node7896;
	wire [15-1:0] node7897;
	wire [15-1:0] node7898;
	wire [15-1:0] node7899;
	wire [15-1:0] node7900;
	wire [15-1:0] node7901;
	wire [15-1:0] node7902;
	wire [15-1:0] node7906;
	wire [15-1:0] node7907;
	wire [15-1:0] node7911;
	wire [15-1:0] node7912;
	wire [15-1:0] node7913;
	wire [15-1:0] node7917;
	wire [15-1:0] node7918;
	wire [15-1:0] node7922;
	wire [15-1:0] node7923;
	wire [15-1:0] node7924;
	wire [15-1:0] node7925;
	wire [15-1:0] node7928;
	wire [15-1:0] node7931;
	wire [15-1:0] node7932;
	wire [15-1:0] node7935;
	wire [15-1:0] node7938;
	wire [15-1:0] node7939;
	wire [15-1:0] node7943;
	wire [15-1:0] node7944;
	wire [15-1:0] node7945;
	wire [15-1:0] node7946;
	wire [15-1:0] node7947;
	wire [15-1:0] node7951;
	wire [15-1:0] node7953;
	wire [15-1:0] node7956;
	wire [15-1:0] node7957;
	wire [15-1:0] node7960;
	wire [15-1:0] node7961;
	wire [15-1:0] node7964;
	wire [15-1:0] node7967;
	wire [15-1:0] node7968;
	wire [15-1:0] node7969;
	wire [15-1:0] node7970;
	wire [15-1:0] node7974;
	wire [15-1:0] node7977;
	wire [15-1:0] node7979;
	wire [15-1:0] node7980;
	wire [15-1:0] node7984;
	wire [15-1:0] node7985;
	wire [15-1:0] node7986;
	wire [15-1:0] node7987;
	wire [15-1:0] node7988;
	wire [15-1:0] node7989;
	wire [15-1:0] node7993;
	wire [15-1:0] node7994;
	wire [15-1:0] node7997;
	wire [15-1:0] node8000;
	wire [15-1:0] node8002;
	wire [15-1:0] node8003;
	wire [15-1:0] node8006;
	wire [15-1:0] node8009;
	wire [15-1:0] node8010;
	wire [15-1:0] node8012;
	wire [15-1:0] node8014;
	wire [15-1:0] node8017;
	wire [15-1:0] node8018;
	wire [15-1:0] node8021;
	wire [15-1:0] node8024;
	wire [15-1:0] node8025;
	wire [15-1:0] node8026;
	wire [15-1:0] node8027;
	wire [15-1:0] node8031;
	wire [15-1:0] node8032;
	wire [15-1:0] node8033;
	wire [15-1:0] node8038;
	wire [15-1:0] node8039;
	wire [15-1:0] node8040;
	wire [15-1:0] node8044;
	wire [15-1:0] node8046;
	wire [15-1:0] node8049;
	wire [15-1:0] node8050;
	wire [15-1:0] node8051;
	wire [15-1:0] node8052;
	wire [15-1:0] node8053;
	wire [15-1:0] node8054;
	wire [15-1:0] node8058;
	wire [15-1:0] node8059;
	wire [15-1:0] node8060;
	wire [15-1:0] node8063;
	wire [15-1:0] node8066;
	wire [15-1:0] node8067;
	wire [15-1:0] node8071;
	wire [15-1:0] node8072;
	wire [15-1:0] node8074;
	wire [15-1:0] node8075;
	wire [15-1:0] node8079;
	wire [15-1:0] node8080;
	wire [15-1:0] node8081;
	wire [15-1:0] node8085;
	wire [15-1:0] node8086;
	wire [15-1:0] node8089;
	wire [15-1:0] node8092;
	wire [15-1:0] node8093;
	wire [15-1:0] node8094;
	wire [15-1:0] node8095;
	wire [15-1:0] node8099;
	wire [15-1:0] node8100;
	wire [15-1:0] node8101;
	wire [15-1:0] node8105;
	wire [15-1:0] node8107;
	wire [15-1:0] node8110;
	wire [15-1:0] node8111;
	wire [15-1:0] node8113;
	wire [15-1:0] node8114;
	wire [15-1:0] node8118;
	wire [15-1:0] node8119;
	wire [15-1:0] node8121;
	wire [15-1:0] node8125;
	wire [15-1:0] node8126;
	wire [15-1:0] node8127;
	wire [15-1:0] node8128;
	wire [15-1:0] node8131;
	wire [15-1:0] node8132;
	wire [15-1:0] node8135;
	wire [15-1:0] node8138;
	wire [15-1:0] node8139;
	wire [15-1:0] node8140;
	wire [15-1:0] node8143;
	wire [15-1:0] node8144;
	wire [15-1:0] node8147;
	wire [15-1:0] node8150;
	wire [15-1:0] node8151;
	wire [15-1:0] node8154;
	wire [15-1:0] node8157;
	wire [15-1:0] node8158;
	wire [15-1:0] node8159;
	wire [15-1:0] node8160;
	wire [15-1:0] node8161;
	wire [15-1:0] node8164;
	wire [15-1:0] node8167;
	wire [15-1:0] node8169;
	wire [15-1:0] node8172;
	wire [15-1:0] node8173;
	wire [15-1:0] node8177;
	wire [15-1:0] node8178;
	wire [15-1:0] node8179;
	wire [15-1:0] node8183;
	wire [15-1:0] node8184;
	wire [15-1:0] node8186;
	wire [15-1:0] node8189;
	wire [15-1:0] node8190;
	wire [15-1:0] node8193;
	wire [15-1:0] node8196;
	wire [15-1:0] node8197;
	wire [15-1:0] node8198;
	wire [15-1:0] node8199;
	wire [15-1:0] node8200;
	wire [15-1:0] node8201;
	wire [15-1:0] node8202;
	wire [15-1:0] node8205;
	wire [15-1:0] node8206;
	wire [15-1:0] node8210;
	wire [15-1:0] node8211;
	wire [15-1:0] node8213;
	wire [15-1:0] node8217;
	wire [15-1:0] node8218;
	wire [15-1:0] node8220;
	wire [15-1:0] node8221;
	wire [15-1:0] node8224;
	wire [15-1:0] node8227;
	wire [15-1:0] node8228;
	wire [15-1:0] node8229;
	wire [15-1:0] node8233;
	wire [15-1:0] node8236;
	wire [15-1:0] node8237;
	wire [15-1:0] node8238;
	wire [15-1:0] node8240;
	wire [15-1:0] node8243;
	wire [15-1:0] node8245;
	wire [15-1:0] node8246;
	wire [15-1:0] node8250;
	wire [15-1:0] node8251;
	wire [15-1:0] node8252;
	wire [15-1:0] node8253;
	wire [15-1:0] node8256;
	wire [15-1:0] node8260;
	wire [15-1:0] node8261;
	wire [15-1:0] node8262;
	wire [15-1:0] node8267;
	wire [15-1:0] node8268;
	wire [15-1:0] node8269;
	wire [15-1:0] node8270;
	wire [15-1:0] node8271;
	wire [15-1:0] node8273;
	wire [15-1:0] node8276;
	wire [15-1:0] node8277;
	wire [15-1:0] node8280;
	wire [15-1:0] node8283;
	wire [15-1:0] node8284;
	wire [15-1:0] node8287;
	wire [15-1:0] node8288;
	wire [15-1:0] node8292;
	wire [15-1:0] node8293;
	wire [15-1:0] node8294;
	wire [15-1:0] node8295;
	wire [15-1:0] node8299;
	wire [15-1:0] node8300;
	wire [15-1:0] node8304;
	wire [15-1:0] node8306;
	wire [15-1:0] node8307;
	wire [15-1:0] node8311;
	wire [15-1:0] node8312;
	wire [15-1:0] node8313;
	wire [15-1:0] node8315;
	wire [15-1:0] node8316;
	wire [15-1:0] node8320;
	wire [15-1:0] node8321;
	wire [15-1:0] node8323;
	wire [15-1:0] node8326;
	wire [15-1:0] node8328;
	wire [15-1:0] node8331;
	wire [15-1:0] node8332;
	wire [15-1:0] node8333;
	wire [15-1:0] node8335;
	wire [15-1:0] node8338;
	wire [15-1:0] node8339;
	wire [15-1:0] node8343;
	wire [15-1:0] node8344;
	wire [15-1:0] node8346;
	wire [15-1:0] node8350;
	wire [15-1:0] node8351;
	wire [15-1:0] node8352;
	wire [15-1:0] node8353;
	wire [15-1:0] node8354;
	wire [15-1:0] node8355;
	wire [15-1:0] node8356;
	wire [15-1:0] node8361;
	wire [15-1:0] node8362;
	wire [15-1:0] node8363;
	wire [15-1:0] node8366;
	wire [15-1:0] node8369;
	wire [15-1:0] node8370;
	wire [15-1:0] node8374;
	wire [15-1:0] node8375;
	wire [15-1:0] node8376;
	wire [15-1:0] node8377;
	wire [15-1:0] node8380;
	wire [15-1:0] node8383;
	wire [15-1:0] node8386;
	wire [15-1:0] node8389;
	wire [15-1:0] node8390;
	wire [15-1:0] node8391;
	wire [15-1:0] node8392;
	wire [15-1:0] node8395;
	wire [15-1:0] node8398;
	wire [15-1:0] node8399;
	wire [15-1:0] node8400;
	wire [15-1:0] node8403;
	wire [15-1:0] node8406;
	wire [15-1:0] node8408;
	wire [15-1:0] node8411;
	wire [15-1:0] node8412;
	wire [15-1:0] node8413;
	wire [15-1:0] node8415;
	wire [15-1:0] node8418;
	wire [15-1:0] node8421;
	wire [15-1:0] node8422;
	wire [15-1:0] node8424;
	wire [15-1:0] node8428;
	wire [15-1:0] node8429;
	wire [15-1:0] node8430;
	wire [15-1:0] node8431;
	wire [15-1:0] node8432;
	wire [15-1:0] node8435;
	wire [15-1:0] node8437;
	wire [15-1:0] node8440;
	wire [15-1:0] node8442;
	wire [15-1:0] node8444;
	wire [15-1:0] node8447;
	wire [15-1:0] node8448;
	wire [15-1:0] node8449;
	wire [15-1:0] node8453;
	wire [15-1:0] node8455;
	wire [15-1:0] node8456;
	wire [15-1:0] node8460;
	wire [15-1:0] node8461;
	wire [15-1:0] node8462;
	wire [15-1:0] node8463;
	wire [15-1:0] node8464;
	wire [15-1:0] node8468;
	wire [15-1:0] node8470;
	wire [15-1:0] node8473;
	wire [15-1:0] node8474;
	wire [15-1:0] node8476;
	wire [15-1:0] node8479;
	wire [15-1:0] node8480;
	wire [15-1:0] node8484;
	wire [15-1:0] node8485;
	wire [15-1:0] node8486;
	wire [15-1:0] node8489;
	wire [15-1:0] node8491;
	wire [15-1:0] node8494;
	wire [15-1:0] node8495;
	wire [15-1:0] node8497;
	wire [15-1:0] node8500;
	wire [15-1:0] node8501;
	wire [15-1:0] node8504;
	wire [15-1:0] node8507;
	wire [15-1:0] node8508;
	wire [15-1:0] node8509;
	wire [15-1:0] node8510;
	wire [15-1:0] node8511;
	wire [15-1:0] node8512;
	wire [15-1:0] node8513;
	wire [15-1:0] node8514;
	wire [15-1:0] node8517;
	wire [15-1:0] node8519;
	wire [15-1:0] node8522;
	wire [15-1:0] node8523;
	wire [15-1:0] node8524;
	wire [15-1:0] node8529;
	wire [15-1:0] node8530;
	wire [15-1:0] node8531;
	wire [15-1:0] node8532;
	wire [15-1:0] node8535;
	wire [15-1:0] node8538;
	wire [15-1:0] node8541;
	wire [15-1:0] node8542;
	wire [15-1:0] node8543;
	wire [15-1:0] node8546;
	wire [15-1:0] node8549;
	wire [15-1:0] node8550;
	wire [15-1:0] node8553;
	wire [15-1:0] node8556;
	wire [15-1:0] node8557;
	wire [15-1:0] node8558;
	wire [15-1:0] node8559;
	wire [15-1:0] node8560;
	wire [15-1:0] node8564;
	wire [15-1:0] node8567;
	wire [15-1:0] node8569;
	wire [15-1:0] node8570;
	wire [15-1:0] node8573;
	wire [15-1:0] node8576;
	wire [15-1:0] node8577;
	wire [15-1:0] node8578;
	wire [15-1:0] node8580;
	wire [15-1:0] node8584;
	wire [15-1:0] node8585;
	wire [15-1:0] node8587;
	wire [15-1:0] node8590;
	wire [15-1:0] node8593;
	wire [15-1:0] node8594;
	wire [15-1:0] node8595;
	wire [15-1:0] node8596;
	wire [15-1:0] node8597;
	wire [15-1:0] node8599;
	wire [15-1:0] node8602;
	wire [15-1:0] node8603;
	wire [15-1:0] node8606;
	wire [15-1:0] node8609;
	wire [15-1:0] node8610;
	wire [15-1:0] node8612;
	wire [15-1:0] node8615;
	wire [15-1:0] node8616;
	wire [15-1:0] node8620;
	wire [15-1:0] node8621;
	wire [15-1:0] node8622;
	wire [15-1:0] node8623;
	wire [15-1:0] node8627;
	wire [15-1:0] node8629;
	wire [15-1:0] node8632;
	wire [15-1:0] node8634;
	wire [15-1:0] node8635;
	wire [15-1:0] node8639;
	wire [15-1:0] node8640;
	wire [15-1:0] node8641;
	wire [15-1:0] node8643;
	wire [15-1:0] node8646;
	wire [15-1:0] node8647;
	wire [15-1:0] node8649;
	wire [15-1:0] node8652;
	wire [15-1:0] node8653;
	wire [15-1:0] node8656;
	wire [15-1:0] node8659;
	wire [15-1:0] node8660;
	wire [15-1:0] node8661;
	wire [15-1:0] node8662;
	wire [15-1:0] node8666;
	wire [15-1:0] node8668;
	wire [15-1:0] node8671;
	wire [15-1:0] node8673;
	wire [15-1:0] node8675;
	wire [15-1:0] node8678;
	wire [15-1:0] node8679;
	wire [15-1:0] node8680;
	wire [15-1:0] node8681;
	wire [15-1:0] node8682;
	wire [15-1:0] node8683;
	wire [15-1:0] node8684;
	wire [15-1:0] node8688;
	wire [15-1:0] node8689;
	wire [15-1:0] node8693;
	wire [15-1:0] node8696;
	wire [15-1:0] node8697;
	wire [15-1:0] node8700;
	wire [15-1:0] node8702;
	wire [15-1:0] node8705;
	wire [15-1:0] node8706;
	wire [15-1:0] node8707;
	wire [15-1:0] node8708;
	wire [15-1:0] node8710;
	wire [15-1:0] node8713;
	wire [15-1:0] node8714;
	wire [15-1:0] node8718;
	wire [15-1:0] node8719;
	wire [15-1:0] node8720;
	wire [15-1:0] node8723;
	wire [15-1:0] node8727;
	wire [15-1:0] node8728;
	wire [15-1:0] node8729;
	wire [15-1:0] node8733;
	wire [15-1:0] node8734;
	wire [15-1:0] node8735;
	wire [15-1:0] node8739;
	wire [15-1:0] node8741;
	wire [15-1:0] node8744;
	wire [15-1:0] node8745;
	wire [15-1:0] node8746;
	wire [15-1:0] node8747;
	wire [15-1:0] node8749;
	wire [15-1:0] node8750;
	wire [15-1:0] node8754;
	wire [15-1:0] node8755;
	wire [15-1:0] node8757;
	wire [15-1:0] node8761;
	wire [15-1:0] node8762;
	wire [15-1:0] node8764;
	wire [15-1:0] node8766;
	wire [15-1:0] node8769;
	wire [15-1:0] node8770;
	wire [15-1:0] node8771;
	wire [15-1:0] node8775;
	wire [15-1:0] node8777;
	wire [15-1:0] node8780;
	wire [15-1:0] node8781;
	wire [15-1:0] node8782;
	wire [15-1:0] node8783;
	wire [15-1:0] node8785;
	wire [15-1:0] node8788;
	wire [15-1:0] node8789;
	wire [15-1:0] node8793;
	wire [15-1:0] node8794;
	wire [15-1:0] node8795;
	wire [15-1:0] node8798;
	wire [15-1:0] node8801;
	wire [15-1:0] node8802;
	wire [15-1:0] node8805;
	wire [15-1:0] node8808;
	wire [15-1:0] node8809;
	wire [15-1:0] node8810;
	wire [15-1:0] node8812;
	wire [15-1:0] node8815;
	wire [15-1:0] node8816;
	wire [15-1:0] node8820;
	wire [15-1:0] node8821;
	wire [15-1:0] node8822;
	wire [15-1:0] node8825;
	wire [15-1:0] node8828;
	wire [15-1:0] node8829;
	wire [15-1:0] node8833;
	wire [15-1:0] node8834;
	wire [15-1:0] node8835;
	wire [15-1:0] node8836;
	wire [15-1:0] node8837;
	wire [15-1:0] node8838;
	wire [15-1:0] node8839;
	wire [15-1:0] node8840;
	wire [15-1:0] node8843;
	wire [15-1:0] node8847;
	wire [15-1:0] node8850;
	wire [15-1:0] node8851;
	wire [15-1:0] node8852;
	wire [15-1:0] node8853;
	wire [15-1:0] node8858;
	wire [15-1:0] node8859;
	wire [15-1:0] node8860;
	wire [15-1:0] node8863;
	wire [15-1:0] node8866;
	wire [15-1:0] node8868;
	wire [15-1:0] node8871;
	wire [15-1:0] node8872;
	wire [15-1:0] node8873;
	wire [15-1:0] node8874;
	wire [15-1:0] node8877;
	wire [15-1:0] node8878;
	wire [15-1:0] node8881;
	wire [15-1:0] node8884;
	wire [15-1:0] node8886;
	wire [15-1:0] node8887;
	wire [15-1:0] node8891;
	wire [15-1:0] node8892;
	wire [15-1:0] node8893;
	wire [15-1:0] node8894;
	wire [15-1:0] node8898;
	wire [15-1:0] node8899;
	wire [15-1:0] node8902;
	wire [15-1:0] node8905;
	wire [15-1:0] node8906;
	wire [15-1:0] node8907;
	wire [15-1:0] node8910;
	wire [15-1:0] node8913;
	wire [15-1:0] node8914;
	wire [15-1:0] node8917;
	wire [15-1:0] node8920;
	wire [15-1:0] node8921;
	wire [15-1:0] node8922;
	wire [15-1:0] node8923;
	wire [15-1:0] node8924;
	wire [15-1:0] node8925;
	wire [15-1:0] node8928;
	wire [15-1:0] node8932;
	wire [15-1:0] node8933;
	wire [15-1:0] node8935;
	wire [15-1:0] node8939;
	wire [15-1:0] node8940;
	wire [15-1:0] node8941;
	wire [15-1:0] node8943;
	wire [15-1:0] node8946;
	wire [15-1:0] node8947;
	wire [15-1:0] node8951;
	wire [15-1:0] node8952;
	wire [15-1:0] node8954;
	wire [15-1:0] node8957;
	wire [15-1:0] node8958;
	wire [15-1:0] node8962;
	wire [15-1:0] node8963;
	wire [15-1:0] node8964;
	wire [15-1:0] node8965;
	wire [15-1:0] node8969;
	wire [15-1:0] node8970;
	wire [15-1:0] node8973;
	wire [15-1:0] node8974;
	wire [15-1:0] node8978;
	wire [15-1:0] node8979;
	wire [15-1:0] node8980;
	wire [15-1:0] node8982;
	wire [15-1:0] node8986;
	wire [15-1:0] node8988;
	wire [15-1:0] node8989;
	wire [15-1:0] node8992;
	wire [15-1:0] node8995;
	wire [15-1:0] node8996;
	wire [15-1:0] node8997;
	wire [15-1:0] node8998;
	wire [15-1:0] node8999;
	wire [15-1:0] node9000;
	wire [15-1:0] node9003;
	wire [15-1:0] node9005;
	wire [15-1:0] node9008;
	wire [15-1:0] node9009;
	wire [15-1:0] node9010;
	wire [15-1:0] node9013;
	wire [15-1:0] node9016;
	wire [15-1:0] node9017;
	wire [15-1:0] node9021;
	wire [15-1:0] node9022;
	wire [15-1:0] node9023;
	wire [15-1:0] node9026;
	wire [15-1:0] node9028;
	wire [15-1:0] node9031;
	wire [15-1:0] node9032;
	wire [15-1:0] node9033;
	wire [15-1:0] node9036;
	wire [15-1:0] node9039;
	wire [15-1:0] node9040;
	wire [15-1:0] node9044;
	wire [15-1:0] node9045;
	wire [15-1:0] node9046;
	wire [15-1:0] node9047;
	wire [15-1:0] node9048;
	wire [15-1:0] node9052;
	wire [15-1:0] node9055;
	wire [15-1:0] node9056;
	wire [15-1:0] node9057;
	wire [15-1:0] node9060;
	wire [15-1:0] node9063;
	wire [15-1:0] node9064;
	wire [15-1:0] node9067;
	wire [15-1:0] node9070;
	wire [15-1:0] node9071;
	wire [15-1:0] node9072;
	wire [15-1:0] node9073;
	wire [15-1:0] node9076;
	wire [15-1:0] node9079;
	wire [15-1:0] node9081;
	wire [15-1:0] node9084;
	wire [15-1:0] node9085;
	wire [15-1:0] node9086;
	wire [15-1:0] node9089;
	wire [15-1:0] node9092;
	wire [15-1:0] node9093;
	wire [15-1:0] node9097;
	wire [15-1:0] node9098;
	wire [15-1:0] node9099;
	wire [15-1:0] node9100;
	wire [15-1:0] node9101;
	wire [15-1:0] node9103;
	wire [15-1:0] node9106;
	wire [15-1:0] node9109;
	wire [15-1:0] node9110;
	wire [15-1:0] node9112;
	wire [15-1:0] node9115;
	wire [15-1:0] node9117;
	wire [15-1:0] node9120;
	wire [15-1:0] node9121;
	wire [15-1:0] node9122;
	wire [15-1:0] node9125;
	wire [15-1:0] node9126;
	wire [15-1:0] node9129;
	wire [15-1:0] node9132;
	wire [15-1:0] node9133;
	wire [15-1:0] node9134;
	wire [15-1:0] node9137;
	wire [15-1:0] node9140;
	wire [15-1:0] node9141;
	wire [15-1:0] node9144;
	wire [15-1:0] node9147;
	wire [15-1:0] node9148;
	wire [15-1:0] node9149;
	wire [15-1:0] node9150;
	wire [15-1:0] node9153;
	wire [15-1:0] node9155;
	wire [15-1:0] node9158;
	wire [15-1:0] node9159;
	wire [15-1:0] node9161;
	wire [15-1:0] node9164;
	wire [15-1:0] node9165;
	wire [15-1:0] node9169;
	wire [15-1:0] node9170;
	wire [15-1:0] node9171;
	wire [15-1:0] node9172;
	wire [15-1:0] node9175;
	wire [15-1:0] node9178;
	wire [15-1:0] node9179;
	wire [15-1:0] node9182;
	wire [15-1:0] node9185;
	wire [15-1:0] node9186;
	wire [15-1:0] node9187;
	wire [15-1:0] node9191;
	wire [15-1:0] node9193;
	wire [15-1:0] node9196;
	wire [15-1:0] node9197;
	wire [15-1:0] node9198;
	wire [15-1:0] node9199;
	wire [15-1:0] node9200;
	wire [15-1:0] node9201;
	wire [15-1:0] node9202;
	wire [15-1:0] node9203;
	wire [15-1:0] node9204;
	wire [15-1:0] node9205;
	wire [15-1:0] node9209;
	wire [15-1:0] node9210;
	wire [15-1:0] node9214;
	wire [15-1:0] node9215;
	wire [15-1:0] node9216;
	wire [15-1:0] node9219;
	wire [15-1:0] node9222;
	wire [15-1:0] node9224;
	wire [15-1:0] node9227;
	wire [15-1:0] node9228;
	wire [15-1:0] node9230;
	wire [15-1:0] node9233;
	wire [15-1:0] node9234;
	wire [15-1:0] node9236;
	wire [15-1:0] node9239;
	wire [15-1:0] node9240;
	wire [15-1:0] node9244;
	wire [15-1:0] node9245;
	wire [15-1:0] node9246;
	wire [15-1:0] node9247;
	wire [15-1:0] node9248;
	wire [15-1:0] node9251;
	wire [15-1:0] node9254;
	wire [15-1:0] node9255;
	wire [15-1:0] node9258;
	wire [15-1:0] node9261;
	wire [15-1:0] node9262;
	wire [15-1:0] node9263;
	wire [15-1:0] node9266;
	wire [15-1:0] node9270;
	wire [15-1:0] node9271;
	wire [15-1:0] node9272;
	wire [15-1:0] node9274;
	wire [15-1:0] node9277;
	wire [15-1:0] node9279;
	wire [15-1:0] node9282;
	wire [15-1:0] node9283;
	wire [15-1:0] node9284;
	wire [15-1:0] node9287;
	wire [15-1:0] node9290;
	wire [15-1:0] node9293;
	wire [15-1:0] node9294;
	wire [15-1:0] node9295;
	wire [15-1:0] node9296;
	wire [15-1:0] node9297;
	wire [15-1:0] node9299;
	wire [15-1:0] node9303;
	wire [15-1:0] node9304;
	wire [15-1:0] node9306;
	wire [15-1:0] node9309;
	wire [15-1:0] node9310;
	wire [15-1:0] node9314;
	wire [15-1:0] node9315;
	wire [15-1:0] node9317;
	wire [15-1:0] node9318;
	wire [15-1:0] node9322;
	wire [15-1:0] node9323;
	wire [15-1:0] node9324;
	wire [15-1:0] node9328;
	wire [15-1:0] node9330;
	wire [15-1:0] node9333;
	wire [15-1:0] node9334;
	wire [15-1:0] node9335;
	wire [15-1:0] node9336;
	wire [15-1:0] node9339;
	wire [15-1:0] node9340;
	wire [15-1:0] node9343;
	wire [15-1:0] node9346;
	wire [15-1:0] node9347;
	wire [15-1:0] node9348;
	wire [15-1:0] node9351;
	wire [15-1:0] node9354;
	wire [15-1:0] node9355;
	wire [15-1:0] node9358;
	wire [15-1:0] node9361;
	wire [15-1:0] node9362;
	wire [15-1:0] node9363;
	wire [15-1:0] node9366;
	wire [15-1:0] node9367;
	wire [15-1:0] node9371;
	wire [15-1:0] node9372;
	wire [15-1:0] node9374;
	wire [15-1:0] node9377;
	wire [15-1:0] node9378;
	wire [15-1:0] node9381;
	wire [15-1:0] node9384;
	wire [15-1:0] node9385;
	wire [15-1:0] node9386;
	wire [15-1:0] node9387;
	wire [15-1:0] node9388;
	wire [15-1:0] node9390;
	wire [15-1:0] node9391;
	wire [15-1:0] node9395;
	wire [15-1:0] node9397;
	wire [15-1:0] node9398;
	wire [15-1:0] node9402;
	wire [15-1:0] node9403;
	wire [15-1:0] node9404;
	wire [15-1:0] node9405;
	wire [15-1:0] node9410;
	wire [15-1:0] node9411;
	wire [15-1:0] node9415;
	wire [15-1:0] node9416;
	wire [15-1:0] node9417;
	wire [15-1:0] node9418;
	wire [15-1:0] node9420;
	wire [15-1:0] node9424;
	wire [15-1:0] node9426;
	wire [15-1:0] node9429;
	wire [15-1:0] node9430;
	wire [15-1:0] node9431;
	wire [15-1:0] node9433;
	wire [15-1:0] node9436;
	wire [15-1:0] node9437;
	wire [15-1:0] node9440;
	wire [15-1:0] node9443;
	wire [15-1:0] node9445;
	wire [15-1:0] node9446;
	wire [15-1:0] node9450;
	wire [15-1:0] node9451;
	wire [15-1:0] node9452;
	wire [15-1:0] node9453;
	wire [15-1:0] node9454;
	wire [15-1:0] node9455;
	wire [15-1:0] node9459;
	wire [15-1:0] node9462;
	wire [15-1:0] node9463;
	wire [15-1:0] node9464;
	wire [15-1:0] node9468;
	wire [15-1:0] node9469;
	wire [15-1:0] node9472;
	wire [15-1:0] node9475;
	wire [15-1:0] node9476;
	wire [15-1:0] node9477;
	wire [15-1:0] node9480;
	wire [15-1:0] node9482;
	wire [15-1:0] node9485;
	wire [15-1:0] node9486;
	wire [15-1:0] node9488;
	wire [15-1:0] node9491;
	wire [15-1:0] node9493;
	wire [15-1:0] node9496;
	wire [15-1:0] node9497;
	wire [15-1:0] node9498;
	wire [15-1:0] node9501;
	wire [15-1:0] node9502;
	wire [15-1:0] node9506;
	wire [15-1:0] node9507;
	wire [15-1:0] node9508;
	wire [15-1:0] node9510;
	wire [15-1:0] node9514;
	wire [15-1:0] node9515;
	wire [15-1:0] node9516;
	wire [15-1:0] node9520;
	wire [15-1:0] node9521;
	wire [15-1:0] node9524;
	wire [15-1:0] node9527;
	wire [15-1:0] node9528;
	wire [15-1:0] node9529;
	wire [15-1:0] node9530;
	wire [15-1:0] node9531;
	wire [15-1:0] node9532;
	wire [15-1:0] node9533;
	wire [15-1:0] node9534;
	wire [15-1:0] node9538;
	wire [15-1:0] node9541;
	wire [15-1:0] node9542;
	wire [15-1:0] node9544;
	wire [15-1:0] node9547;
	wire [15-1:0] node9548;
	wire [15-1:0] node9552;
	wire [15-1:0] node9553;
	wire [15-1:0] node9555;
	wire [15-1:0] node9556;
	wire [15-1:0] node9560;
	wire [15-1:0] node9561;
	wire [15-1:0] node9564;
	wire [15-1:0] node9567;
	wire [15-1:0] node9568;
	wire [15-1:0] node9569;
	wire [15-1:0] node9571;
	wire [15-1:0] node9572;
	wire [15-1:0] node9576;
	wire [15-1:0] node9577;
	wire [15-1:0] node9581;
	wire [15-1:0] node9582;
	wire [15-1:0] node9584;
	wire [15-1:0] node9586;
	wire [15-1:0] node9589;
	wire [15-1:0] node9590;
	wire [15-1:0] node9592;
	wire [15-1:0] node9595;
	wire [15-1:0] node9598;
	wire [15-1:0] node9599;
	wire [15-1:0] node9600;
	wire [15-1:0] node9601;
	wire [15-1:0] node9602;
	wire [15-1:0] node9604;
	wire [15-1:0] node9607;
	wire [15-1:0] node9610;
	wire [15-1:0] node9611;
	wire [15-1:0] node9614;
	wire [15-1:0] node9616;
	wire [15-1:0] node9619;
	wire [15-1:0] node9620;
	wire [15-1:0] node9621;
	wire [15-1:0] node9623;
	wire [15-1:0] node9626;
	wire [15-1:0] node9628;
	wire [15-1:0] node9631;
	wire [15-1:0] node9632;
	wire [15-1:0] node9634;
	wire [15-1:0] node9637;
	wire [15-1:0] node9639;
	wire [15-1:0] node9642;
	wire [15-1:0] node9643;
	wire [15-1:0] node9644;
	wire [15-1:0] node9647;
	wire [15-1:0] node9648;
	wire [15-1:0] node9650;
	wire [15-1:0] node9653;
	wire [15-1:0] node9654;
	wire [15-1:0] node9658;
	wire [15-1:0] node9659;
	wire [15-1:0] node9660;
	wire [15-1:0] node9663;
	wire [15-1:0] node9665;
	wire [15-1:0] node9668;
	wire [15-1:0] node9669;
	wire [15-1:0] node9670;
	wire [15-1:0] node9673;
	wire [15-1:0] node9676;
	wire [15-1:0] node9677;
	wire [15-1:0] node9681;
	wire [15-1:0] node9682;
	wire [15-1:0] node9683;
	wire [15-1:0] node9684;
	wire [15-1:0] node9685;
	wire [15-1:0] node9687;
	wire [15-1:0] node9690;
	wire [15-1:0] node9691;
	wire [15-1:0] node9692;
	wire [15-1:0] node9696;
	wire [15-1:0] node9697;
	wire [15-1:0] node9700;
	wire [15-1:0] node9703;
	wire [15-1:0] node9704;
	wire [15-1:0] node9706;
	wire [15-1:0] node9707;
	wire [15-1:0] node9710;
	wire [15-1:0] node9713;
	wire [15-1:0] node9714;
	wire [15-1:0] node9716;
	wire [15-1:0] node9719;
	wire [15-1:0] node9721;
	wire [15-1:0] node9724;
	wire [15-1:0] node9725;
	wire [15-1:0] node9726;
	wire [15-1:0] node9727;
	wire [15-1:0] node9728;
	wire [15-1:0] node9731;
	wire [15-1:0] node9734;
	wire [15-1:0] node9736;
	wire [15-1:0] node9739;
	wire [15-1:0] node9740;
	wire [15-1:0] node9741;
	wire [15-1:0] node9744;
	wire [15-1:0] node9747;
	wire [15-1:0] node9748;
	wire [15-1:0] node9751;
	wire [15-1:0] node9754;
	wire [15-1:0] node9755;
	wire [15-1:0] node9756;
	wire [15-1:0] node9760;
	wire [15-1:0] node9761;
	wire [15-1:0] node9762;
	wire [15-1:0] node9766;
	wire [15-1:0] node9767;
	wire [15-1:0] node9770;
	wire [15-1:0] node9773;
	wire [15-1:0] node9774;
	wire [15-1:0] node9775;
	wire [15-1:0] node9776;
	wire [15-1:0] node9777;
	wire [15-1:0] node9780;
	wire [15-1:0] node9781;
	wire [15-1:0] node9785;
	wire [15-1:0] node9787;
	wire [15-1:0] node9788;
	wire [15-1:0] node9791;
	wire [15-1:0] node9794;
	wire [15-1:0] node9795;
	wire [15-1:0] node9796;
	wire [15-1:0] node9798;
	wire [15-1:0] node9802;
	wire [15-1:0] node9803;
	wire [15-1:0] node9804;
	wire [15-1:0] node9808;
	wire [15-1:0] node9809;
	wire [15-1:0] node9812;
	wire [15-1:0] node9815;
	wire [15-1:0] node9816;
	wire [15-1:0] node9817;
	wire [15-1:0] node9818;
	wire [15-1:0] node9819;
	wire [15-1:0] node9822;
	wire [15-1:0] node9825;
	wire [15-1:0] node9826;
	wire [15-1:0] node9830;
	wire [15-1:0] node9831;
	wire [15-1:0] node9833;
	wire [15-1:0] node9836;
	wire [15-1:0] node9837;
	wire [15-1:0] node9840;
	wire [15-1:0] node9843;
	wire [15-1:0] node9844;
	wire [15-1:0] node9845;
	wire [15-1:0] node9847;
	wire [15-1:0] node9850;
	wire [15-1:0] node9851;
	wire [15-1:0] node9854;
	wire [15-1:0] node9857;
	wire [15-1:0] node9859;
	wire [15-1:0] node9860;
	wire [15-1:0] node9863;
	wire [15-1:0] node9866;
	wire [15-1:0] node9867;
	wire [15-1:0] node9868;
	wire [15-1:0] node9869;
	wire [15-1:0] node9870;
	wire [15-1:0] node9871;
	wire [15-1:0] node9872;
	wire [15-1:0] node9873;
	wire [15-1:0] node9876;
	wire [15-1:0] node9879;
	wire [15-1:0] node9880;
	wire [15-1:0] node9881;
	wire [15-1:0] node9885;
	wire [15-1:0] node9887;
	wire [15-1:0] node9890;
	wire [15-1:0] node9891;
	wire [15-1:0] node9892;
	wire [15-1:0] node9894;
	wire [15-1:0] node9897;
	wire [15-1:0] node9898;
	wire [15-1:0] node9901;
	wire [15-1:0] node9904;
	wire [15-1:0] node9906;
	wire [15-1:0] node9907;
	wire [15-1:0] node9911;
	wire [15-1:0] node9912;
	wire [15-1:0] node9913;
	wire [15-1:0] node9916;
	wire [15-1:0] node9917;
	wire [15-1:0] node9921;
	wire [15-1:0] node9922;
	wire [15-1:0] node9923;
	wire [15-1:0] node9925;
	wire [15-1:0] node9928;
	wire [15-1:0] node9931;
	wire [15-1:0] node9932;
	wire [15-1:0] node9935;
	wire [15-1:0] node9937;
	wire [15-1:0] node9940;
	wire [15-1:0] node9941;
	wire [15-1:0] node9942;
	wire [15-1:0] node9943;
	wire [15-1:0] node9944;
	wire [15-1:0] node9947;
	wire [15-1:0] node9948;
	wire [15-1:0] node9951;
	wire [15-1:0] node9954;
	wire [15-1:0] node9955;
	wire [15-1:0] node9958;
	wire [15-1:0] node9959;
	wire [15-1:0] node9962;
	wire [15-1:0] node9965;
	wire [15-1:0] node9966;
	wire [15-1:0] node9967;
	wire [15-1:0] node9969;
	wire [15-1:0] node9972;
	wire [15-1:0] node9973;
	wire [15-1:0] node9977;
	wire [15-1:0] node9978;
	wire [15-1:0] node9979;
	wire [15-1:0] node9984;
	wire [15-1:0] node9985;
	wire [15-1:0] node9986;
	wire [15-1:0] node9987;
	wire [15-1:0] node9989;
	wire [15-1:0] node9992;
	wire [15-1:0] node9993;
	wire [15-1:0] node9997;
	wire [15-1:0] node9998;
	wire [15-1:0] node10000;
	wire [15-1:0] node10003;
	wire [15-1:0] node10004;
	wire [15-1:0] node10008;
	wire [15-1:0] node10009;
	wire [15-1:0] node10010;
	wire [15-1:0] node10011;
	wire [15-1:0] node10015;
	wire [15-1:0] node10017;
	wire [15-1:0] node10020;
	wire [15-1:0] node10021;
	wire [15-1:0] node10023;
	wire [15-1:0] node10026;
	wire [15-1:0] node10028;
	wire [15-1:0] node10031;
	wire [15-1:0] node10032;
	wire [15-1:0] node10033;
	wire [15-1:0] node10034;
	wire [15-1:0] node10035;
	wire [15-1:0] node10036;
	wire [15-1:0] node10037;
	wire [15-1:0] node10041;
	wire [15-1:0] node10043;
	wire [15-1:0] node10046;
	wire [15-1:0] node10047;
	wire [15-1:0] node10048;
	wire [15-1:0] node10051;
	wire [15-1:0] node10055;
	wire [15-1:0] node10056;
	wire [15-1:0] node10058;
	wire [15-1:0] node10059;
	wire [15-1:0] node10063;
	wire [15-1:0] node10064;
	wire [15-1:0] node10065;
	wire [15-1:0] node10069;
	wire [15-1:0] node10071;
	wire [15-1:0] node10074;
	wire [15-1:0] node10075;
	wire [15-1:0] node10076;
	wire [15-1:0] node10077;
	wire [15-1:0] node10079;
	wire [15-1:0] node10082;
	wire [15-1:0] node10084;
	wire [15-1:0] node10087;
	wire [15-1:0] node10088;
	wire [15-1:0] node10089;
	wire [15-1:0] node10092;
	wire [15-1:0] node10095;
	wire [15-1:0] node10096;
	wire [15-1:0] node10099;
	wire [15-1:0] node10102;
	wire [15-1:0] node10103;
	wire [15-1:0] node10104;
	wire [15-1:0] node10106;
	wire [15-1:0] node10109;
	wire [15-1:0] node10110;
	wire [15-1:0] node10114;
	wire [15-1:0] node10115;
	wire [15-1:0] node10116;
	wire [15-1:0] node10119;
	wire [15-1:0] node10122;
	wire [15-1:0] node10123;
	wire [15-1:0] node10126;
	wire [15-1:0] node10129;
	wire [15-1:0] node10130;
	wire [15-1:0] node10131;
	wire [15-1:0] node10132;
	wire [15-1:0] node10133;
	wire [15-1:0] node10136;
	wire [15-1:0] node10138;
	wire [15-1:0] node10141;
	wire [15-1:0] node10142;
	wire [15-1:0] node10144;
	wire [15-1:0] node10147;
	wire [15-1:0] node10148;
	wire [15-1:0] node10152;
	wire [15-1:0] node10153;
	wire [15-1:0] node10154;
	wire [15-1:0] node10155;
	wire [15-1:0] node10159;
	wire [15-1:0] node10160;
	wire [15-1:0] node10164;
	wire [15-1:0] node10165;
	wire [15-1:0] node10168;
	wire [15-1:0] node10170;
	wire [15-1:0] node10173;
	wire [15-1:0] node10174;
	wire [15-1:0] node10175;
	wire [15-1:0] node10176;
	wire [15-1:0] node10177;
	wire [15-1:0] node10180;
	wire [15-1:0] node10184;
	wire [15-1:0] node10185;
	wire [15-1:0] node10187;
	wire [15-1:0] node10190;
	wire [15-1:0] node10193;
	wire [15-1:0] node10194;
	wire [15-1:0] node10195;
	wire [15-1:0] node10197;
	wire [15-1:0] node10200;
	wire [15-1:0] node10202;
	wire [15-1:0] node10205;
	wire [15-1:0] node10207;
	wire [15-1:0] node10209;
	wire [15-1:0] node10212;
	wire [15-1:0] node10213;
	wire [15-1:0] node10214;
	wire [15-1:0] node10215;
	wire [15-1:0] node10216;
	wire [15-1:0] node10217;
	wire [15-1:0] node10218;
	wire [15-1:0] node10221;
	wire [15-1:0] node10222;
	wire [15-1:0] node10226;
	wire [15-1:0] node10228;
	wire [15-1:0] node10229;
	wire [15-1:0] node10232;
	wire [15-1:0] node10235;
	wire [15-1:0] node10236;
	wire [15-1:0] node10237;
	wire [15-1:0] node10240;
	wire [15-1:0] node10243;
	wire [15-1:0] node10245;
	wire [15-1:0] node10246;
	wire [15-1:0] node10250;
	wire [15-1:0] node10251;
	wire [15-1:0] node10252;
	wire [15-1:0] node10253;
	wire [15-1:0] node10255;
	wire [15-1:0] node10258;
	wire [15-1:0] node10259;
	wire [15-1:0] node10263;
	wire [15-1:0] node10264;
	wire [15-1:0] node10267;
	wire [15-1:0] node10268;
	wire [15-1:0] node10271;
	wire [15-1:0] node10274;
	wire [15-1:0] node10275;
	wire [15-1:0] node10277;
	wire [15-1:0] node10278;
	wire [15-1:0] node10282;
	wire [15-1:0] node10283;
	wire [15-1:0] node10284;
	wire [15-1:0] node10288;
	wire [15-1:0] node10291;
	wire [15-1:0] node10292;
	wire [15-1:0] node10293;
	wire [15-1:0] node10294;
	wire [15-1:0] node10295;
	wire [15-1:0] node10296;
	wire [15-1:0] node10300;
	wire [15-1:0] node10301;
	wire [15-1:0] node10305;
	wire [15-1:0] node10306;
	wire [15-1:0] node10307;
	wire [15-1:0] node10310;
	wire [15-1:0] node10313;
	wire [15-1:0] node10314;
	wire [15-1:0] node10317;
	wire [15-1:0] node10320;
	wire [15-1:0] node10321;
	wire [15-1:0] node10322;
	wire [15-1:0] node10323;
	wire [15-1:0] node10327;
	wire [15-1:0] node10329;
	wire [15-1:0] node10332;
	wire [15-1:0] node10333;
	wire [15-1:0] node10337;
	wire [15-1:0] node10338;
	wire [15-1:0] node10339;
	wire [15-1:0] node10340;
	wire [15-1:0] node10341;
	wire [15-1:0] node10345;
	wire [15-1:0] node10346;
	wire [15-1:0] node10350;
	wire [15-1:0] node10351;
	wire [15-1:0] node10353;
	wire [15-1:0] node10356;
	wire [15-1:0] node10359;
	wire [15-1:0] node10360;
	wire [15-1:0] node10361;
	wire [15-1:0] node10365;
	wire [15-1:0] node10366;
	wire [15-1:0] node10368;
	wire [15-1:0] node10371;
	wire [15-1:0] node10372;
	wire [15-1:0] node10375;
	wire [15-1:0] node10378;
	wire [15-1:0] node10379;
	wire [15-1:0] node10380;
	wire [15-1:0] node10381;
	wire [15-1:0] node10382;
	wire [15-1:0] node10384;
	wire [15-1:0] node10385;
	wire [15-1:0] node10389;
	wire [15-1:0] node10391;
	wire [15-1:0] node10394;
	wire [15-1:0] node10395;
	wire [15-1:0] node10396;
	wire [15-1:0] node10397;
	wire [15-1:0] node10400;
	wire [15-1:0] node10403;
	wire [15-1:0] node10404;
	wire [15-1:0] node10407;
	wire [15-1:0] node10410;
	wire [15-1:0] node10411;
	wire [15-1:0] node10414;
	wire [15-1:0] node10416;
	wire [15-1:0] node10419;
	wire [15-1:0] node10420;
	wire [15-1:0] node10421;
	wire [15-1:0] node10422;
	wire [15-1:0] node10425;
	wire [15-1:0] node10427;
	wire [15-1:0] node10430;
	wire [15-1:0] node10431;
	wire [15-1:0] node10432;
	wire [15-1:0] node10435;
	wire [15-1:0] node10438;
	wire [15-1:0] node10439;
	wire [15-1:0] node10442;
	wire [15-1:0] node10445;
	wire [15-1:0] node10446;
	wire [15-1:0] node10447;
	wire [15-1:0] node10448;
	wire [15-1:0] node10452;
	wire [15-1:0] node10453;
	wire [15-1:0] node10457;
	wire [15-1:0] node10458;
	wire [15-1:0] node10462;
	wire [15-1:0] node10463;
	wire [15-1:0] node10464;
	wire [15-1:0] node10465;
	wire [15-1:0] node10466;
	wire [15-1:0] node10467;
	wire [15-1:0] node10470;
	wire [15-1:0] node10474;
	wire [15-1:0] node10475;
	wire [15-1:0] node10477;
	wire [15-1:0] node10480;
	wire [15-1:0] node10482;
	wire [15-1:0] node10485;
	wire [15-1:0] node10486;
	wire [15-1:0] node10487;
	wire [15-1:0] node10489;
	wire [15-1:0] node10492;
	wire [15-1:0] node10493;
	wire [15-1:0] node10496;
	wire [15-1:0] node10499;
	wire [15-1:0] node10501;
	wire [15-1:0] node10502;
	wire [15-1:0] node10506;
	wire [15-1:0] node10507;
	wire [15-1:0] node10508;
	wire [15-1:0] node10509;
	wire [15-1:0] node10512;
	wire [15-1:0] node10513;
	wire [15-1:0] node10517;
	wire [15-1:0] node10518;
	wire [15-1:0] node10519;
	wire [15-1:0] node10522;
	wire [15-1:0] node10526;
	wire [15-1:0] node10527;
	wire [15-1:0] node10528;
	wire [15-1:0] node10529;
	wire [15-1:0] node10532;
	wire [15-1:0] node10535;
	wire [15-1:0] node10537;
	wire [15-1:0] node10540;
	wire [15-1:0] node10541;
	wire [15-1:0] node10542;
	wire [15-1:0] node10545;
	wire [15-1:0] node10548;
	wire [15-1:0] node10550;

	assign outp = (inp[11]) ? node5214 : node1;
		assign node1 = (inp[12]) ? node2583 : node2;
			assign node2 = (inp[5]) ? node1298 : node3;
				assign node3 = (inp[2]) ? node633 : node4;
					assign node4 = (inp[0]) ? node346 : node5;
						assign node5 = (inp[6]) ? node187 : node6;
							assign node6 = (inp[13]) ? node94 : node7;
								assign node7 = (inp[4]) ? node53 : node8;
									assign node8 = (inp[9]) ? node34 : node9;
										assign node9 = (inp[8]) ? node23 : node10;
											assign node10 = (inp[3]) ? node16 : node11;
												assign node11 = (inp[1]) ? 15'b001111111111111 : node12;
													assign node12 = (inp[10]) ? 15'b000111111111111 : 15'b011111111111111;
												assign node16 = (inp[1]) ? node20 : node17;
													assign node17 = (inp[10]) ? 15'b000111111111111 : 15'b011111111111111;
													assign node20 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node23 = (inp[10]) ? node29 : node24;
												assign node24 = (inp[7]) ? node26 : 15'b000111111111111;
													assign node26 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node29 = (inp[14]) ? 15'b000001111111111 : node30;
													assign node30 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node34 = (inp[3]) ? node44 : node35;
											assign node35 = (inp[14]) ? node41 : node36;
												assign node36 = (inp[7]) ? node38 : 15'b001111111111111;
													assign node38 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node41 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node44 = (inp[8]) ? node50 : node45;
												assign node45 = (inp[1]) ? node47 : 15'b000011111111111;
													assign node47 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node50 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node53 = (inp[10]) ? node77 : node54;
										assign node54 = (inp[14]) ? node66 : node55;
											assign node55 = (inp[1]) ? node61 : node56;
												assign node56 = (inp[3]) ? 15'b000011111111111 : node57;
													assign node57 = (inp[7]) ? 15'b001111111111111 : 15'b001111111111111;
												assign node61 = (inp[9]) ? 15'b000001111111111 : node62;
													assign node62 = (inp[8]) ? 15'b000111111111111 : 15'b000011111111111;
											assign node66 = (inp[8]) ? node72 : node67;
												assign node67 = (inp[7]) ? node69 : 15'b000011111111111;
													assign node69 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node72 = (inp[9]) ? 15'b000001111111111 : node73;
													assign node73 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node77 = (inp[14]) ? node87 : node78;
											assign node78 = (inp[3]) ? node82 : node79;
												assign node79 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node82 = (inp[1]) ? 15'b000001111111111 : node83;
													assign node83 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node87 = (inp[7]) ? node89 : 15'b000011111111111;
												assign node89 = (inp[9]) ? 15'b000000111111111 : node90;
													assign node90 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node94 = (inp[7]) ? node146 : node95;
									assign node95 = (inp[14]) ? node119 : node96;
										assign node96 = (inp[8]) ? node106 : node97;
											assign node97 = (inp[4]) ? node101 : node98;
												assign node98 = (inp[10]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node101 = (inp[3]) ? node103 : 15'b000111111111111;
													assign node103 = (inp[10]) ? 15'b000011111111111 : 15'b000011111111111;
											assign node106 = (inp[3]) ? node114 : node107;
												assign node107 = (inp[4]) ? node111 : node108;
													assign node108 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node111 = (inp[1]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node114 = (inp[9]) ? 15'b000001111111111 : node115;
													assign node115 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node119 = (inp[4]) ? node133 : node120;
											assign node120 = (inp[3]) ? node126 : node121;
												assign node121 = (inp[8]) ? 15'b000011111111111 : node122;
													assign node122 = (inp[10]) ? 15'b000011111111111 : 15'b001111111111111;
												assign node126 = (inp[10]) ? node130 : node127;
													assign node127 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node130 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node133 = (inp[10]) ? node139 : node134;
												assign node134 = (inp[1]) ? node136 : 15'b000001111111111;
													assign node136 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node139 = (inp[8]) ? node143 : node140;
													assign node140 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node143 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node146 = (inp[4]) ? node172 : node147;
										assign node147 = (inp[8]) ? node159 : node148;
											assign node148 = (inp[14]) ? node154 : node149;
												assign node149 = (inp[3]) ? node151 : 15'b000011111111111;
													assign node151 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node154 = (inp[1]) ? node156 : 15'b000011111111111;
													assign node156 = (inp[3]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node159 = (inp[1]) ? node165 : node160;
												assign node160 = (inp[9]) ? 15'b000011111111111 : node161;
													assign node161 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node165 = (inp[14]) ? node169 : node166;
													assign node166 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node169 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node172 = (inp[10]) ? node178 : node173;
											assign node173 = (inp[9]) ? 15'b000000111111111 : node174;
												assign node174 = (inp[14]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node178 = (inp[8]) ? node184 : node179;
												assign node179 = (inp[14]) ? 15'b000000011111111 : node180;
													assign node180 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node184 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
							assign node187 = (inp[3]) ? node263 : node188;
								assign node188 = (inp[10]) ? node232 : node189;
									assign node189 = (inp[14]) ? node211 : node190;
										assign node190 = (inp[9]) ? node198 : node191;
											assign node191 = (inp[1]) ? 15'b000011111111111 : node192;
												assign node192 = (inp[8]) ? 15'b000011111111111 : node193;
													assign node193 = (inp[7]) ? 15'b000111111111111 : 15'b000111111111111;
											assign node198 = (inp[13]) ? node206 : node199;
												assign node199 = (inp[4]) ? node203 : node200;
													assign node200 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node203 = (inp[1]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node206 = (inp[8]) ? 15'b000001111111111 : node207;
													assign node207 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node211 = (inp[13]) ? node219 : node212;
											assign node212 = (inp[8]) ? node214 : 15'b000011111111111;
												assign node214 = (inp[4]) ? 15'b000001111111111 : node215;
													assign node215 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node219 = (inp[1]) ? node225 : node220;
												assign node220 = (inp[8]) ? node222 : 15'b000011111111111;
													assign node222 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node225 = (inp[8]) ? node229 : node226;
													assign node226 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node229 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node232 = (inp[14]) ? node252 : node233;
										assign node233 = (inp[7]) ? node243 : node234;
											assign node234 = (inp[1]) ? node236 : 15'b000011111111111;
												assign node236 = (inp[8]) ? node240 : node237;
													assign node237 = (inp[4]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node240 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node243 = (inp[1]) ? node249 : node244;
												assign node244 = (inp[8]) ? node246 : 15'b000011111111111;
													assign node246 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node249 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node252 = (inp[7]) ? node260 : node253;
											assign node253 = (inp[8]) ? node257 : node254;
												assign node254 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node257 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node260 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node263 = (inp[13]) ? node303 : node264;
									assign node264 = (inp[10]) ? node286 : node265;
										assign node265 = (inp[7]) ? node275 : node266;
											assign node266 = (inp[8]) ? 15'b000001111111111 : node267;
												assign node267 = (inp[4]) ? node271 : node268;
													assign node268 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node271 = (inp[9]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node275 = (inp[1]) ? node281 : node276;
												assign node276 = (inp[8]) ? 15'b000001111111111 : node277;
													assign node277 = (inp[4]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node281 = (inp[14]) ? node283 : 15'b000001111111111;
													assign node283 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node286 = (inp[1]) ? node296 : node287;
											assign node287 = (inp[8]) ? node293 : node288;
												assign node288 = (inp[4]) ? node290 : 15'b000001111111111;
													assign node290 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node293 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node296 = (inp[7]) ? 15'b000000011111111 : node297;
												assign node297 = (inp[8]) ? node299 : 15'b000000111111111;
													assign node299 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
									assign node303 = (inp[10]) ? node331 : node304;
										assign node304 = (inp[9]) ? node318 : node305;
											assign node305 = (inp[1]) ? node313 : node306;
												assign node306 = (inp[8]) ? node310 : node307;
													assign node307 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node310 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node313 = (inp[4]) ? node315 : 15'b000000111111111;
													assign node315 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node318 = (inp[14]) ? node326 : node319;
												assign node319 = (inp[1]) ? node323 : node320;
													assign node320 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node323 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node326 = (inp[8]) ? node328 : 15'b000000011111111;
													assign node328 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node331 = (inp[14]) ? node339 : node332;
											assign node332 = (inp[1]) ? node336 : node333;
												assign node333 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node336 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node339 = (inp[8]) ? node341 : 15'b000000111111111;
												assign node341 = (inp[9]) ? node343 : 15'b000000001111111;
													assign node343 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
						assign node346 = (inp[1]) ? node504 : node347;
							assign node347 = (inp[13]) ? node435 : node348;
								assign node348 = (inp[14]) ? node390 : node349;
									assign node349 = (inp[9]) ? node369 : node350;
										assign node350 = (inp[8]) ? node362 : node351;
											assign node351 = (inp[3]) ? node357 : node352;
												assign node352 = (inp[6]) ? 15'b000011111111111 : node353;
													assign node353 = (inp[4]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node357 = (inp[4]) ? 15'b000011111111111 : node358;
													assign node358 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node362 = (inp[10]) ? node364 : 15'b000011111111111;
												assign node364 = (inp[7]) ? 15'b000000111111111 : node365;
													assign node365 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node369 = (inp[10]) ? node383 : node370;
											assign node370 = (inp[3]) ? node376 : node371;
												assign node371 = (inp[6]) ? node373 : 15'b000011111111111;
													assign node373 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node376 = (inp[4]) ? node380 : node377;
													assign node377 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node380 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node383 = (inp[6]) ? node385 : 15'b000001111111111;
												assign node385 = (inp[4]) ? 15'b000000001111111 : node386;
													assign node386 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node390 = (inp[3]) ? node410 : node391;
										assign node391 = (inp[7]) ? node401 : node392;
											assign node392 = (inp[6]) ? node396 : node393;
												assign node393 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node396 = (inp[9]) ? 15'b000001111111111 : node397;
													assign node397 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node401 = (inp[6]) ? node403 : 15'b000001111111111;
												assign node403 = (inp[10]) ? node407 : node404;
													assign node404 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node407 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node410 = (inp[6]) ? node422 : node411;
											assign node411 = (inp[8]) ? node417 : node412;
												assign node412 = (inp[9]) ? node414 : 15'b000001111111111;
													assign node414 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node417 = (inp[10]) ? 15'b000000111111111 : node418;
													assign node418 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node422 = (inp[4]) ? node430 : node423;
												assign node423 = (inp[10]) ? node427 : node424;
													assign node424 = (inp[8]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node427 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node430 = (inp[7]) ? node432 : 15'b000000111111111;
													assign node432 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node435 = (inp[4]) ? node473 : node436;
									assign node436 = (inp[6]) ? node456 : node437;
										assign node437 = (inp[10]) ? node447 : node438;
											assign node438 = (inp[8]) ? 15'b000001111111111 : node439;
												assign node439 = (inp[14]) ? node443 : node440;
													assign node440 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node443 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node447 = (inp[9]) ? 15'b000000111111111 : node448;
												assign node448 = (inp[8]) ? node452 : node449;
													assign node449 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node452 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node456 = (inp[3]) ? node466 : node457;
											assign node457 = (inp[7]) ? 15'b000000111111111 : node458;
												assign node458 = (inp[8]) ? node462 : node459;
													assign node459 = (inp[9]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node462 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node466 = (inp[14]) ? node468 : 15'b000000011111111;
												assign node468 = (inp[10]) ? node470 : 15'b000000111111111;
													assign node470 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node473 = (inp[10]) ? node487 : node474;
										assign node474 = (inp[6]) ? node480 : node475;
											assign node475 = (inp[9]) ? node477 : 15'b000000111111111;
												assign node477 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node480 = (inp[8]) ? 15'b000000111111111 : node481;
												assign node481 = (inp[14]) ? 15'b000000111111111 : node482;
													assign node482 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node487 = (inp[3]) ? node493 : node488;
											assign node488 = (inp[8]) ? 15'b000000011111111 : node489;
												assign node489 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node493 = (inp[8]) ? node499 : node494;
												assign node494 = (inp[6]) ? 15'b000000001111111 : node495;
													assign node495 = (inp[9]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node499 = (inp[9]) ? node501 : 15'b000000011111111;
													assign node501 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node504 = (inp[6]) ? node572 : node505;
								assign node505 = (inp[10]) ? node533 : node506;
									assign node506 = (inp[3]) ? node522 : node507;
										assign node507 = (inp[4]) ? node517 : node508;
											assign node508 = (inp[8]) ? node512 : node509;
												assign node509 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node512 = (inp[14]) ? node514 : 15'b000011111111111;
													assign node514 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node517 = (inp[13]) ? node519 : 15'b000001111111111;
												assign node519 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node522 = (inp[7]) ? 15'b000000011111111 : node523;
											assign node523 = (inp[4]) ? node529 : node524;
												assign node524 = (inp[8]) ? node526 : 15'b000011111111111;
													assign node526 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node529 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node533 = (inp[9]) ? node547 : node534;
										assign node534 = (inp[14]) ? node538 : node535;
											assign node535 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node538 = (inp[13]) ? node544 : node539;
												assign node539 = (inp[7]) ? 15'b000000111111111 : node540;
													assign node540 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node544 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node547 = (inp[3]) ? node561 : node548;
											assign node548 = (inp[8]) ? node556 : node549;
												assign node549 = (inp[14]) ? node553 : node550;
													assign node550 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node553 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node556 = (inp[13]) ? node558 : 15'b000000011111111;
													assign node558 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node561 = (inp[8]) ? node567 : node562;
												assign node562 = (inp[13]) ? node564 : 15'b000000111111111;
													assign node564 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node567 = (inp[13]) ? node569 : 15'b000000001111111;
													assign node569 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node572 = (inp[4]) ? node592 : node573;
									assign node573 = (inp[8]) ? node583 : node574;
										assign node574 = (inp[9]) ? 15'b000000001111111 : node575;
											assign node575 = (inp[7]) ? node577 : 15'b000001111111111;
												assign node577 = (inp[3]) ? 15'b000000111111111 : node578;
													assign node578 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node583 = (inp[10]) ? node589 : node584;
											assign node584 = (inp[7]) ? 15'b000000011111111 : node585;
												assign node585 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node589 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node592 = (inp[3]) ? node618 : node593;
										assign node593 = (inp[8]) ? node607 : node594;
											assign node594 = (inp[9]) ? node600 : node595;
												assign node595 = (inp[7]) ? node597 : 15'b000000111111111;
													assign node597 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node600 = (inp[10]) ? node604 : node601;
													assign node601 = (inp[13]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node604 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node607 = (inp[10]) ? node613 : node608;
												assign node608 = (inp[13]) ? node610 : 15'b000000111111111;
													assign node610 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node613 = (inp[7]) ? node615 : 15'b000000001111111;
													assign node615 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node618 = (inp[14]) ? node622 : node619;
											assign node619 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node622 = (inp[13]) ? node628 : node623;
												assign node623 = (inp[8]) ? node625 : 15'b000000011111111;
													assign node625 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node628 = (inp[8]) ? 15'b000000000011111 : node629;
													assign node629 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node633 = (inp[9]) ? node947 : node634;
						assign node634 = (inp[0]) ? node794 : node635;
							assign node635 = (inp[6]) ? node723 : node636;
								assign node636 = (inp[3]) ? node678 : node637;
									assign node637 = (inp[7]) ? node663 : node638;
										assign node638 = (inp[4]) ? node652 : node639;
											assign node639 = (inp[13]) ? node647 : node640;
												assign node640 = (inp[14]) ? node644 : node641;
													assign node641 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node644 = (inp[10]) ? 15'b000111111111111 : 15'b000111111111111;
												assign node647 = (inp[1]) ? 15'b000011111111111 : node648;
													assign node648 = (inp[14]) ? 15'b000011111111111 : 15'b001111111111111;
											assign node652 = (inp[13]) ? node658 : node653;
												assign node653 = (inp[8]) ? 15'b000001111111111 : node654;
													assign node654 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node658 = (inp[8]) ? 15'b000001111111111 : node659;
													assign node659 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node663 = (inp[1]) ? node671 : node664;
											assign node664 = (inp[13]) ? 15'b000001111111111 : node665;
												assign node665 = (inp[14]) ? node667 : 15'b000111111111111;
													assign node667 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node671 = (inp[10]) ? 15'b000000111111111 : node672;
												assign node672 = (inp[13]) ? node674 : 15'b000001111111111;
													assign node674 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node678 = (inp[8]) ? node700 : node679;
										assign node679 = (inp[10]) ? node693 : node680;
											assign node680 = (inp[13]) ? node686 : node681;
												assign node681 = (inp[1]) ? 15'b000011111111111 : node682;
													assign node682 = (inp[7]) ? 15'b000011111111111 : 15'b001111111111111;
												assign node686 = (inp[7]) ? node690 : node687;
													assign node687 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node690 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node693 = (inp[7]) ? 15'b000000111111111 : node694;
												assign node694 = (inp[1]) ? node696 : 15'b000001111111111;
													assign node696 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node700 = (inp[13]) ? node708 : node701;
											assign node701 = (inp[4]) ? node703 : 15'b000001111111111;
												assign node703 = (inp[14]) ? node705 : 15'b000001111111111;
													assign node705 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node708 = (inp[1]) ? node716 : node709;
												assign node709 = (inp[4]) ? node713 : node710;
													assign node710 = (inp[10]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node713 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node716 = (inp[14]) ? node720 : node717;
													assign node717 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node720 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node723 = (inp[13]) ? node767 : node724;
									assign node724 = (inp[4]) ? node746 : node725;
										assign node725 = (inp[8]) ? node733 : node726;
											assign node726 = (inp[10]) ? 15'b000001111111111 : node727;
												assign node727 = (inp[3]) ? node729 : 15'b000111111111111;
													assign node729 = (inp[14]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node733 = (inp[10]) ? node741 : node734;
												assign node734 = (inp[1]) ? node738 : node735;
													assign node735 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node738 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node741 = (inp[3]) ? node743 : 15'b000000111111111;
													assign node743 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node746 = (inp[10]) ? node762 : node747;
											assign node747 = (inp[8]) ? node755 : node748;
												assign node748 = (inp[14]) ? node752 : node749;
													assign node749 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node752 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node755 = (inp[1]) ? node759 : node756;
													assign node756 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node759 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node762 = (inp[14]) ? 15'b000000011111111 : node763;
												assign node763 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
									assign node767 = (inp[7]) ? node781 : node768;
										assign node768 = (inp[3]) ? node776 : node769;
											assign node769 = (inp[14]) ? 15'b000000111111111 : node770;
												assign node770 = (inp[10]) ? 15'b000000111111111 : node771;
													assign node771 = (inp[4]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node776 = (inp[4]) ? node778 : 15'b000001111111111;
												assign node778 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node781 = (inp[10]) ? node791 : node782;
											assign node782 = (inp[8]) ? node788 : node783;
												assign node783 = (inp[3]) ? 15'b000001111111111 : node784;
													assign node784 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node788 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node791 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node794 = (inp[8]) ? node882 : node795;
								assign node795 = (inp[13]) ? node837 : node796;
									assign node796 = (inp[1]) ? node820 : node797;
										assign node797 = (inp[4]) ? node807 : node798;
											assign node798 = (inp[14]) ? node800 : 15'b000011111111111;
												assign node800 = (inp[3]) ? node804 : node801;
													assign node801 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node804 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node807 = (inp[14]) ? node815 : node808;
												assign node808 = (inp[7]) ? node812 : node809;
													assign node809 = (inp[3]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node812 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node815 = (inp[7]) ? node817 : 15'b000000111111111;
													assign node817 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node820 = (inp[3]) ? node828 : node821;
											assign node821 = (inp[10]) ? 15'b000000111111111 : node822;
												assign node822 = (inp[6]) ? node824 : 15'b000001111111111;
													assign node824 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node828 = (inp[4]) ? node834 : node829;
												assign node829 = (inp[10]) ? node831 : 15'b000000111111111;
													assign node831 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node834 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node837 = (inp[14]) ? node859 : node838;
										assign node838 = (inp[3]) ? node846 : node839;
											assign node839 = (inp[10]) ? node841 : 15'b000001111111111;
												assign node841 = (inp[6]) ? 15'b000000011111111 : node842;
													assign node842 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node846 = (inp[7]) ? node852 : node847;
												assign node847 = (inp[6]) ? node849 : 15'b000000111111111;
													assign node849 = (inp[10]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node852 = (inp[1]) ? node856 : node853;
													assign node853 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node856 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node859 = (inp[6]) ? node869 : node860;
											assign node860 = (inp[4]) ? node866 : node861;
												assign node861 = (inp[1]) ? node863 : 15'b000000111111111;
													assign node863 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node866 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node869 = (inp[7]) ? node877 : node870;
												assign node870 = (inp[3]) ? node874 : node871;
													assign node871 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node874 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node877 = (inp[10]) ? node879 : 15'b000000011111111;
													assign node879 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node882 = (inp[7]) ? node920 : node883;
									assign node883 = (inp[1]) ? node901 : node884;
										assign node884 = (inp[10]) ? node894 : node885;
											assign node885 = (inp[3]) ? node887 : 15'b000001111111111;
												assign node887 = (inp[14]) ? node891 : node888;
													assign node888 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node891 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node894 = (inp[14]) ? node896 : 15'b000000111111111;
												assign node896 = (inp[4]) ? 15'b000000011111111 : node897;
													assign node897 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node901 = (inp[10]) ? node911 : node902;
											assign node902 = (inp[6]) ? node906 : node903;
												assign node903 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node906 = (inp[3]) ? node908 : 15'b000000111111111;
													assign node908 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node911 = (inp[4]) ? node917 : node912;
												assign node912 = (inp[14]) ? node914 : 15'b000000011111111;
													assign node914 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node917 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node920 = (inp[14]) ? node934 : node921;
										assign node921 = (inp[13]) ? node927 : node922;
											assign node922 = (inp[3]) ? node924 : 15'b000000111111111;
												assign node924 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node927 = (inp[6]) ? 15'b000000001111111 : node928;
												assign node928 = (inp[3]) ? node930 : 15'b000000011111111;
													assign node930 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node934 = (inp[4]) ? node944 : node935;
											assign node935 = (inp[6]) ? node939 : node936;
												assign node936 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node939 = (inp[3]) ? node941 : 15'b000000001111111;
													assign node941 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node944 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node947 = (inp[7]) ? node1133 : node948;
							assign node948 = (inp[14]) ? node1048 : node949;
								assign node949 = (inp[8]) ? node993 : node950;
									assign node950 = (inp[13]) ? node970 : node951;
										assign node951 = (inp[6]) ? node961 : node952;
											assign node952 = (inp[3]) ? node958 : node953;
												assign node953 = (inp[0]) ? 15'b000011111111111 : node954;
													assign node954 = (inp[4]) ? 15'b000111111111111 : 15'b000111111111111;
												assign node958 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node961 = (inp[4]) ? 15'b000000111111111 : node962;
												assign node962 = (inp[10]) ? node966 : node963;
													assign node963 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node966 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node970 = (inp[6]) ? node982 : node971;
											assign node971 = (inp[1]) ? node977 : node972;
												assign node972 = (inp[10]) ? node974 : 15'b000001111111111;
													assign node974 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node977 = (inp[10]) ? 15'b000000111111111 : node978;
													assign node978 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node982 = (inp[4]) ? node988 : node983;
												assign node983 = (inp[10]) ? node985 : 15'b000001111111111;
													assign node985 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node988 = (inp[1]) ? 15'b000000011111111 : node989;
													assign node989 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node993 = (inp[0]) ? node1023 : node994;
										assign node994 = (inp[3]) ? node1010 : node995;
											assign node995 = (inp[13]) ? node1003 : node996;
												assign node996 = (inp[6]) ? node1000 : node997;
													assign node997 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node1000 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1003 = (inp[10]) ? node1007 : node1004;
													assign node1004 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1007 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node1010 = (inp[10]) ? node1018 : node1011;
												assign node1011 = (inp[13]) ? node1015 : node1012;
													assign node1012 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1015 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1018 = (inp[1]) ? 15'b000000001111111 : node1019;
													assign node1019 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1023 = (inp[1]) ? node1037 : node1024;
											assign node1024 = (inp[4]) ? node1030 : node1025;
												assign node1025 = (inp[3]) ? 15'b000000111111111 : node1026;
													assign node1026 = (inp[10]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node1030 = (inp[10]) ? node1034 : node1031;
													assign node1031 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1034 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1037 = (inp[10]) ? node1043 : node1038;
												assign node1038 = (inp[13]) ? node1040 : 15'b000000011111111;
													assign node1040 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1043 = (inp[13]) ? 15'b000000000111111 : node1044;
													assign node1044 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1048 = (inp[8]) ? node1086 : node1049;
									assign node1049 = (inp[1]) ? node1065 : node1050;
										assign node1050 = (inp[13]) ? node1060 : node1051;
											assign node1051 = (inp[0]) ? node1053 : 15'b000001111111111;
												assign node1053 = (inp[4]) ? node1057 : node1054;
													assign node1054 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1057 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1060 = (inp[3]) ? node1062 : 15'b000000111111111;
												assign node1062 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1065 = (inp[10]) ? node1077 : node1066;
											assign node1066 = (inp[0]) ? node1072 : node1067;
												assign node1067 = (inp[6]) ? 15'b000000111111111 : node1068;
													assign node1068 = (inp[3]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node1072 = (inp[4]) ? node1074 : 15'b000000111111111;
													assign node1074 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1077 = (inp[4]) ? 15'b000000001111111 : node1078;
												assign node1078 = (inp[13]) ? node1082 : node1079;
													assign node1079 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1082 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1086 = (inp[1]) ? node1114 : node1087;
										assign node1087 = (inp[13]) ? node1099 : node1088;
											assign node1088 = (inp[10]) ? node1094 : node1089;
												assign node1089 = (inp[3]) ? node1091 : 15'b000011111111111;
													assign node1091 = (inp[6]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node1094 = (inp[6]) ? 15'b000000011111111 : node1095;
													assign node1095 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1099 = (inp[10]) ? node1107 : node1100;
												assign node1100 = (inp[0]) ? node1104 : node1101;
													assign node1101 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1104 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1107 = (inp[4]) ? node1111 : node1108;
													assign node1108 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1111 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1114 = (inp[3]) ? node1128 : node1115;
											assign node1115 = (inp[6]) ? node1121 : node1116;
												assign node1116 = (inp[4]) ? 15'b000000011111111 : node1117;
													assign node1117 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1121 = (inp[13]) ? node1125 : node1122;
													assign node1122 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1125 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1128 = (inp[10]) ? 15'b000000000111111 : node1129;
												assign node1129 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1133 = (inp[6]) ? node1203 : node1134;
								assign node1134 = (inp[13]) ? node1164 : node1135;
									assign node1135 = (inp[10]) ? node1151 : node1136;
										assign node1136 = (inp[3]) ? node1144 : node1137;
											assign node1137 = (inp[1]) ? 15'b000000011111111 : node1138;
												assign node1138 = (inp[4]) ? 15'b000001111111111 : node1139;
													assign node1139 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1144 = (inp[14]) ? node1146 : 15'b000000111111111;
												assign node1146 = (inp[1]) ? node1148 : 15'b000000111111111;
													assign node1148 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1151 = (inp[3]) ? node1159 : node1152;
											assign node1152 = (inp[0]) ? 15'b000000011111111 : node1153;
												assign node1153 = (inp[1]) ? node1155 : 15'b000001111111111;
													assign node1155 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node1159 = (inp[1]) ? node1161 : 15'b000000011111111;
												assign node1161 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1164 = (inp[10]) ? node1190 : node1165;
										assign node1165 = (inp[1]) ? node1179 : node1166;
											assign node1166 = (inp[0]) ? node1172 : node1167;
												assign node1167 = (inp[4]) ? 15'b000000111111111 : node1168;
													assign node1168 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1172 = (inp[14]) ? node1176 : node1173;
													assign node1173 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1176 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1179 = (inp[14]) ? node1185 : node1180;
												assign node1180 = (inp[8]) ? node1182 : 15'b000000011111111;
													assign node1182 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node1185 = (inp[3]) ? node1187 : 15'b000000001111111;
													assign node1187 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1190 = (inp[4]) ? node1198 : node1191;
											assign node1191 = (inp[14]) ? node1193 : 15'b000000011111111;
												assign node1193 = (inp[1]) ? node1195 : 15'b000000001111111;
													assign node1195 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node1198 = (inp[3]) ? node1200 : 15'b000000001111111;
												assign node1200 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1203 = (inp[13]) ? node1249 : node1204;
									assign node1204 = (inp[0]) ? node1224 : node1205;
										assign node1205 = (inp[1]) ? node1209 : node1206;
											assign node1206 = (inp[4]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node1209 = (inp[8]) ? node1217 : node1210;
												assign node1210 = (inp[10]) ? node1214 : node1211;
													assign node1211 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1214 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1217 = (inp[10]) ? node1221 : node1218;
													assign node1218 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1221 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1224 = (inp[1]) ? node1238 : node1225;
											assign node1225 = (inp[8]) ? node1231 : node1226;
												assign node1226 = (inp[10]) ? node1228 : 15'b000000011111111;
													assign node1228 = (inp[3]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node1231 = (inp[3]) ? node1235 : node1232;
													assign node1232 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1235 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1238 = (inp[14]) ? node1244 : node1239;
												assign node1239 = (inp[3]) ? 15'b000000001111111 : node1240;
													assign node1240 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1244 = (inp[8]) ? node1246 : 15'b000000000011111;
													assign node1246 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node1249 = (inp[10]) ? node1273 : node1250;
										assign node1250 = (inp[14]) ? node1264 : node1251;
											assign node1251 = (inp[8]) ? node1259 : node1252;
												assign node1252 = (inp[0]) ? node1256 : node1253;
													assign node1253 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1256 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1259 = (inp[3]) ? node1261 : 15'b000000011111111;
													assign node1261 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1264 = (inp[3]) ? node1268 : node1265;
												assign node1265 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1268 = (inp[8]) ? node1270 : 15'b000000001111111;
													assign node1270 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1273 = (inp[4]) ? node1285 : node1274;
											assign node1274 = (inp[1]) ? node1280 : node1275;
												assign node1275 = (inp[8]) ? node1277 : 15'b000000011111111;
													assign node1277 = (inp[14]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node1280 = (inp[14]) ? node1282 : 15'b000000000111111;
													assign node1282 = (inp[3]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node1285 = (inp[3]) ? node1291 : node1286;
												assign node1286 = (inp[14]) ? node1288 : 15'b000000000111111;
													assign node1288 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node1291 = (inp[14]) ? node1295 : node1292;
													assign node1292 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node1295 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node1298 = (inp[1]) ? node1966 : node1299;
					assign node1299 = (inp[2]) ? node1629 : node1300;
						assign node1300 = (inp[8]) ? node1462 : node1301;
							assign node1301 = (inp[9]) ? node1391 : node1302;
								assign node1302 = (inp[14]) ? node1350 : node1303;
									assign node1303 = (inp[4]) ? node1323 : node1304;
										assign node1304 = (inp[6]) ? node1308 : node1305;
											assign node1305 = (inp[13]) ? 15'b000111111111111 : 15'b001111111111111;
											assign node1308 = (inp[3]) ? node1316 : node1309;
												assign node1309 = (inp[7]) ? node1313 : node1310;
													assign node1310 = (inp[13]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node1313 = (inp[13]) ? 15'b000011111111111 : 15'b000011111111111;
												assign node1316 = (inp[13]) ? node1320 : node1317;
													assign node1317 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1320 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1323 = (inp[6]) ? node1337 : node1324;
											assign node1324 = (inp[10]) ? node1332 : node1325;
												assign node1325 = (inp[3]) ? node1329 : node1326;
													assign node1326 = (inp[7]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node1329 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1332 = (inp[13]) ? node1334 : 15'b000011111111111;
													assign node1334 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1337 = (inp[13]) ? node1345 : node1338;
												assign node1338 = (inp[0]) ? node1342 : node1339;
													assign node1339 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1342 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1345 = (inp[3]) ? 15'b000000111111111 : node1346;
													assign node1346 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1350 = (inp[3]) ? node1368 : node1351;
										assign node1351 = (inp[13]) ? node1359 : node1352;
											assign node1352 = (inp[0]) ? node1356 : node1353;
												assign node1353 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1356 = (inp[7]) ? 15'b000011111111111 : 15'b000001111111111;
											assign node1359 = (inp[4]) ? 15'b000000111111111 : node1360;
												assign node1360 = (inp[7]) ? node1364 : node1361;
													assign node1361 = (inp[0]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node1364 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1368 = (inp[0]) ? node1384 : node1369;
											assign node1369 = (inp[6]) ? node1377 : node1370;
												assign node1370 = (inp[13]) ? node1374 : node1371;
													assign node1371 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1374 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1377 = (inp[4]) ? node1381 : node1378;
													assign node1378 = (inp[7]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node1381 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1384 = (inp[10]) ? 15'b000000001111111 : node1385;
												assign node1385 = (inp[4]) ? node1387 : 15'b000000111111111;
													assign node1387 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1391 = (inp[10]) ? node1421 : node1392;
									assign node1392 = (inp[3]) ? node1408 : node1393;
										assign node1393 = (inp[6]) ? node1399 : node1394;
											assign node1394 = (inp[14]) ? node1396 : 15'b000111111111111;
												assign node1396 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1399 = (inp[4]) ? node1405 : node1400;
												assign node1400 = (inp[14]) ? 15'b000001111111111 : node1401;
													assign node1401 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1405 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1408 = (inp[7]) ? node1414 : node1409;
											assign node1409 = (inp[14]) ? 15'b000000111111111 : node1410;
												assign node1410 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
											assign node1414 = (inp[0]) ? node1416 : 15'b000001111111111;
												assign node1416 = (inp[13]) ? 15'b000000011111111 : node1417;
													assign node1417 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
									assign node1421 = (inp[4]) ? node1447 : node1422;
										assign node1422 = (inp[7]) ? node1438 : node1423;
											assign node1423 = (inp[6]) ? node1431 : node1424;
												assign node1424 = (inp[0]) ? node1428 : node1425;
													assign node1425 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1428 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1431 = (inp[0]) ? node1435 : node1432;
													assign node1432 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node1435 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1438 = (inp[14]) ? node1442 : node1439;
												assign node1439 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1442 = (inp[0]) ? 15'b000000011111111 : node1443;
													assign node1443 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1447 = (inp[7]) ? node1457 : node1448;
											assign node1448 = (inp[14]) ? node1452 : node1449;
												assign node1449 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1452 = (inp[3]) ? node1454 : 15'b000000011111111;
													assign node1454 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1457 = (inp[3]) ? 15'b000000001111111 : node1458;
												assign node1458 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1462 = (inp[3]) ? node1556 : node1463;
								assign node1463 = (inp[6]) ? node1513 : node1464;
									assign node1464 = (inp[0]) ? node1490 : node1465;
										assign node1465 = (inp[10]) ? node1477 : node1466;
											assign node1466 = (inp[7]) ? node1472 : node1467;
												assign node1467 = (inp[9]) ? node1469 : 15'b000011111111111;
													assign node1469 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1472 = (inp[9]) ? node1474 : 15'b000011111111111;
													assign node1474 = (inp[13]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node1477 = (inp[4]) ? node1483 : node1478;
												assign node1478 = (inp[7]) ? 15'b000001111111111 : node1479;
													assign node1479 = (inp[13]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node1483 = (inp[9]) ? node1487 : node1484;
													assign node1484 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1487 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1490 = (inp[9]) ? node1504 : node1491;
											assign node1491 = (inp[10]) ? node1499 : node1492;
												assign node1492 = (inp[4]) ? node1496 : node1493;
													assign node1493 = (inp[14]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node1496 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1499 = (inp[13]) ? node1501 : 15'b000001111111111;
													assign node1501 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1504 = (inp[13]) ? 15'b000000011111111 : node1505;
												assign node1505 = (inp[14]) ? node1509 : node1506;
													assign node1506 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1509 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1513 = (inp[14]) ? node1535 : node1514;
										assign node1514 = (inp[0]) ? node1522 : node1515;
											assign node1515 = (inp[10]) ? 15'b000000111111111 : node1516;
												assign node1516 = (inp[4]) ? node1518 : 15'b000001111111111;
													assign node1518 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1522 = (inp[10]) ? node1530 : node1523;
												assign node1523 = (inp[4]) ? node1527 : node1524;
													assign node1524 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node1527 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1530 = (inp[9]) ? 15'b000000011111111 : node1531;
													assign node1531 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1535 = (inp[0]) ? node1545 : node1536;
											assign node1536 = (inp[13]) ? node1540 : node1537;
												assign node1537 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1540 = (inp[9]) ? 15'b000000001111111 : node1541;
													assign node1541 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node1545 = (inp[7]) ? node1553 : node1546;
												assign node1546 = (inp[10]) ? node1550 : node1547;
													assign node1547 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1550 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1553 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1556 = (inp[4]) ? node1588 : node1557;
									assign node1557 = (inp[0]) ? node1577 : node1558;
										assign node1558 = (inp[10]) ? node1566 : node1559;
											assign node1559 = (inp[7]) ? 15'b000000111111111 : node1560;
												assign node1560 = (inp[13]) ? 15'b000001111111111 : node1561;
													assign node1561 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1566 = (inp[14]) ? node1572 : node1567;
												assign node1567 = (inp[13]) ? 15'b000000011111111 : node1568;
													assign node1568 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1572 = (inp[7]) ? node1574 : 15'b000000111111111;
													assign node1574 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1577 = (inp[9]) ? node1585 : node1578;
											assign node1578 = (inp[10]) ? 15'b000000011111111 : node1579;
												assign node1579 = (inp[6]) ? node1581 : 15'b000000111111111;
													assign node1581 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1585 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1588 = (inp[9]) ? node1610 : node1589;
										assign node1589 = (inp[13]) ? node1603 : node1590;
											assign node1590 = (inp[0]) ? node1598 : node1591;
												assign node1591 = (inp[10]) ? node1595 : node1592;
													assign node1592 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1595 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node1598 = (inp[14]) ? node1600 : 15'b000000011111111;
													assign node1600 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1603 = (inp[7]) ? node1605 : 15'b000000011111111;
												assign node1605 = (inp[10]) ? 15'b000000001111111 : node1606;
													assign node1606 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1610 = (inp[6]) ? node1618 : node1611;
											assign node1611 = (inp[7]) ? node1613 : 15'b000000011111111;
												assign node1613 = (inp[0]) ? 15'b000000001111111 : node1614;
													assign node1614 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1618 = (inp[10]) ? node1624 : node1619;
												assign node1619 = (inp[14]) ? node1621 : 15'b000000011111111;
													assign node1621 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1624 = (inp[14]) ? 15'b000000000011111 : node1625;
													assign node1625 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
						assign node1629 = (inp[13]) ? node1803 : node1630;
							assign node1630 = (inp[8]) ? node1720 : node1631;
								assign node1631 = (inp[14]) ? node1683 : node1632;
									assign node1632 = (inp[9]) ? node1656 : node1633;
										assign node1633 = (inp[0]) ? node1645 : node1634;
											assign node1634 = (inp[10]) ? node1640 : node1635;
												assign node1635 = (inp[3]) ? node1637 : 15'b000111111111111;
													assign node1637 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1640 = (inp[3]) ? 15'b000001111111111 : node1641;
													assign node1641 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1645 = (inp[10]) ? node1653 : node1646;
												assign node1646 = (inp[6]) ? node1650 : node1647;
													assign node1647 = (inp[7]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node1650 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1653 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node1656 = (inp[6]) ? node1670 : node1657;
											assign node1657 = (inp[4]) ? node1663 : node1658;
												assign node1658 = (inp[10]) ? node1660 : 15'b000011111111111;
													assign node1660 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1663 = (inp[10]) ? node1667 : node1664;
													assign node1664 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1667 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1670 = (inp[10]) ? node1678 : node1671;
												assign node1671 = (inp[7]) ? node1675 : node1672;
													assign node1672 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1675 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1678 = (inp[0]) ? 15'b000000011111111 : node1679;
													assign node1679 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1683 = (inp[3]) ? node1705 : node1684;
										assign node1684 = (inp[0]) ? node1700 : node1685;
											assign node1685 = (inp[4]) ? node1693 : node1686;
												assign node1686 = (inp[10]) ? node1690 : node1687;
													assign node1687 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1690 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1693 = (inp[9]) ? node1697 : node1694;
													assign node1694 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1697 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1700 = (inp[9]) ? node1702 : 15'b000000111111111;
												assign node1702 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1705 = (inp[4]) ? node1713 : node1706;
											assign node1706 = (inp[9]) ? node1708 : 15'b000000111111111;
												assign node1708 = (inp[7]) ? 15'b000000001111111 : node1709;
													assign node1709 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1713 = (inp[10]) ? node1715 : 15'b000000011111111;
												assign node1715 = (inp[9]) ? 15'b000000000011111 : node1716;
													assign node1716 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1720 = (inp[10]) ? node1764 : node1721;
									assign node1721 = (inp[3]) ? node1743 : node1722;
										assign node1722 = (inp[6]) ? node1732 : node1723;
											assign node1723 = (inp[4]) ? node1729 : node1724;
												assign node1724 = (inp[7]) ? 15'b000001111111111 : node1725;
													assign node1725 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1729 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1732 = (inp[9]) ? node1738 : node1733;
												assign node1733 = (inp[14]) ? 15'b000000111111111 : node1734;
													assign node1734 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1738 = (inp[4]) ? 15'b000000011111111 : node1739;
													assign node1739 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node1743 = (inp[4]) ? node1751 : node1744;
											assign node1744 = (inp[0]) ? node1746 : 15'b000000111111111;
												assign node1746 = (inp[9]) ? 15'b000000011111111 : node1747;
													assign node1747 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1751 = (inp[7]) ? node1759 : node1752;
												assign node1752 = (inp[9]) ? node1756 : node1753;
													assign node1753 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1756 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1759 = (inp[9]) ? 15'b000000000111111 : node1760;
													assign node1760 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1764 = (inp[9]) ? node1786 : node1765;
										assign node1765 = (inp[7]) ? node1773 : node1766;
											assign node1766 = (inp[4]) ? node1768 : 15'b000001111111111;
												assign node1768 = (inp[6]) ? 15'b000000011111111 : node1769;
													assign node1769 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1773 = (inp[6]) ? node1781 : node1774;
												assign node1774 = (inp[4]) ? node1778 : node1775;
													assign node1775 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1778 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1781 = (inp[14]) ? node1783 : 15'b000000001111111;
													assign node1783 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1786 = (inp[7]) ? node1794 : node1787;
											assign node1787 = (inp[14]) ? node1789 : 15'b000000011111111;
												assign node1789 = (inp[6]) ? 15'b000000001111111 : node1790;
													assign node1790 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1794 = (inp[3]) ? node1798 : node1795;
												assign node1795 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node1798 = (inp[0]) ? node1800 : 15'b000000001111111;
													assign node1800 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1803 = (inp[7]) ? node1883 : node1804;
								assign node1804 = (inp[6]) ? node1842 : node1805;
									assign node1805 = (inp[0]) ? node1827 : node1806;
										assign node1806 = (inp[14]) ? node1814 : node1807;
											assign node1807 = (inp[9]) ? 15'b000000111111111 : node1808;
												assign node1808 = (inp[10]) ? node1810 : 15'b000001111111111;
													assign node1810 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1814 = (inp[10]) ? node1822 : node1815;
												assign node1815 = (inp[3]) ? node1819 : node1816;
													assign node1816 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1819 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1822 = (inp[3]) ? 15'b000000001111111 : node1823;
													assign node1823 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1827 = (inp[9]) ? node1835 : node1828;
											assign node1828 = (inp[3]) ? 15'b000000011111111 : node1829;
												assign node1829 = (inp[14]) ? node1831 : 15'b000000111111111;
													assign node1831 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1835 = (inp[3]) ? 15'b000000001111111 : node1836;
												assign node1836 = (inp[8]) ? node1838 : 15'b000000011111111;
													assign node1838 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1842 = (inp[8]) ? node1868 : node1843;
										assign node1843 = (inp[3]) ? node1859 : node1844;
											assign node1844 = (inp[14]) ? node1852 : node1845;
												assign node1845 = (inp[10]) ? node1849 : node1846;
													assign node1846 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1849 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node1852 = (inp[9]) ? node1856 : node1853;
													assign node1853 = (inp[4]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node1856 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1859 = (inp[9]) ? node1861 : 15'b000000011111111;
												assign node1861 = (inp[14]) ? node1865 : node1862;
													assign node1862 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1865 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node1868 = (inp[9]) ? node1874 : node1869;
											assign node1869 = (inp[4]) ? node1871 : 15'b000000011111111;
												assign node1871 = (inp[3]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node1874 = (inp[3]) ? node1878 : node1875;
												assign node1875 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1878 = (inp[0]) ? node1880 : 15'b000000000111111;
													assign node1880 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1883 = (inp[3]) ? node1923 : node1884;
									assign node1884 = (inp[6]) ? node1906 : node1885;
										assign node1885 = (inp[0]) ? node1895 : node1886;
											assign node1886 = (inp[8]) ? node1892 : node1887;
												assign node1887 = (inp[14]) ? node1889 : 15'b000000111111111;
													assign node1889 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node1892 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1895 = (inp[10]) ? node1901 : node1896;
												assign node1896 = (inp[4]) ? node1898 : 15'b000000111111111;
													assign node1898 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1901 = (inp[9]) ? 15'b000000001111111 : node1902;
													assign node1902 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1906 = (inp[8]) ? node1916 : node1907;
											assign node1907 = (inp[4]) ? node1911 : node1908;
												assign node1908 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1911 = (inp[9]) ? 15'b000000001111111 : node1912;
													assign node1912 = (inp[0]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node1916 = (inp[10]) ? 15'b000000000001111 : node1917;
												assign node1917 = (inp[4]) ? node1919 : 15'b000000001111111;
													assign node1919 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1923 = (inp[10]) ? node1947 : node1924;
										assign node1924 = (inp[0]) ? node1934 : node1925;
											assign node1925 = (inp[9]) ? node1931 : node1926;
												assign node1926 = (inp[6]) ? 15'b000000011111111 : node1927;
													assign node1927 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1931 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1934 = (inp[4]) ? node1940 : node1935;
												assign node1935 = (inp[9]) ? node1937 : 15'b000000011111111;
													assign node1937 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1940 = (inp[6]) ? node1944 : node1941;
													assign node1941 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node1944 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node1947 = (inp[0]) ? node1961 : node1948;
											assign node1948 = (inp[9]) ? node1954 : node1949;
												assign node1949 = (inp[4]) ? node1951 : 15'b000000001111111;
													assign node1951 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1954 = (inp[8]) ? node1958 : node1955;
													assign node1955 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1958 = (inp[4]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node1961 = (inp[14]) ? node1963 : 15'b000000000111111;
												assign node1963 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node1966 = (inp[14]) ? node2274 : node1967;
						assign node1967 = (inp[3]) ? node2115 : node1968;
							assign node1968 = (inp[4]) ? node2038 : node1969;
								assign node1969 = (inp[9]) ? node1999 : node1970;
									assign node1970 = (inp[2]) ? node1992 : node1971;
										assign node1971 = (inp[6]) ? node1981 : node1972;
											assign node1972 = (inp[7]) ? node1978 : node1973;
												assign node1973 = (inp[10]) ? node1975 : 15'b000111111111111;
													assign node1975 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1978 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1981 = (inp[10]) ? node1989 : node1982;
												assign node1982 = (inp[8]) ? node1986 : node1983;
													assign node1983 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1986 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1989 = (inp[0]) ? 15'b000001111111111 : 15'b000000111111111;
										assign node1992 = (inp[6]) ? 15'b000000011111111 : node1993;
											assign node1993 = (inp[7]) ? node1995 : 15'b000001111111111;
												assign node1995 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1999 = (inp[8]) ? node2021 : node2000;
										assign node2000 = (inp[13]) ? node2012 : node2001;
											assign node2001 = (inp[7]) ? node2007 : node2002;
												assign node2002 = (inp[10]) ? node2004 : 15'b000001111111111;
													assign node2004 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2007 = (inp[6]) ? 15'b000000111111111 : node2008;
													assign node2008 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2012 = (inp[7]) ? node2016 : node2013;
												assign node2013 = (inp[0]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node2016 = (inp[2]) ? 15'b000000011111111 : node2017;
													assign node2017 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2021 = (inp[6]) ? node2033 : node2022;
											assign node2022 = (inp[7]) ? node2030 : node2023;
												assign node2023 = (inp[2]) ? node2027 : node2024;
													assign node2024 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2027 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2030 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2033 = (inp[2]) ? 15'b000000001111111 : node2034;
												assign node2034 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2038 = (inp[0]) ? node2080 : node2039;
									assign node2039 = (inp[13]) ? node2063 : node2040;
										assign node2040 = (inp[8]) ? node2052 : node2041;
											assign node2041 = (inp[7]) ? node2045 : node2042;
												assign node2042 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2045 = (inp[10]) ? node2049 : node2046;
													assign node2046 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2049 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2052 = (inp[9]) ? node2058 : node2053;
												assign node2053 = (inp[6]) ? node2055 : 15'b000001111111111;
													assign node2055 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2058 = (inp[6]) ? 15'b000000001111111 : node2059;
													assign node2059 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2063 = (inp[9]) ? node2073 : node2064;
											assign node2064 = (inp[2]) ? node2070 : node2065;
												assign node2065 = (inp[10]) ? node2067 : 15'b000000111111111;
													assign node2067 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2070 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2073 = (inp[6]) ? 15'b000000000111111 : node2074;
												assign node2074 = (inp[8]) ? 15'b000000011111111 : node2075;
													assign node2075 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2080 = (inp[9]) ? node2104 : node2081;
										assign node2081 = (inp[2]) ? node2093 : node2082;
											assign node2082 = (inp[8]) ? node2086 : node2083;
												assign node2083 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2086 = (inp[7]) ? node2090 : node2087;
													assign node2087 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2090 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2093 = (inp[10]) ? node2099 : node2094;
												assign node2094 = (inp[8]) ? node2096 : 15'b000000011111111;
													assign node2096 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2099 = (inp[8]) ? 15'b000000000111111 : node2100;
													assign node2100 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2104 = (inp[13]) ? node2108 : node2105;
											assign node2105 = (inp[2]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node2108 = (inp[2]) ? node2110 : 15'b000000001111111;
												assign node2110 = (inp[8]) ? 15'b000000000011111 : node2111;
													assign node2111 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2115 = (inp[2]) ? node2187 : node2116;
								assign node2116 = (inp[6]) ? node2152 : node2117;
									assign node2117 = (inp[13]) ? node2135 : node2118;
										assign node2118 = (inp[0]) ? node2128 : node2119;
											assign node2119 = (inp[7]) ? node2121 : 15'b000001111111111;
												assign node2121 = (inp[9]) ? node2125 : node2122;
													assign node2122 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2125 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2128 = (inp[7]) ? node2130 : 15'b000000111111111;
												assign node2130 = (inp[4]) ? 15'b000000011111111 : node2131;
													assign node2131 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2135 = (inp[8]) ? node2147 : node2136;
											assign node2136 = (inp[10]) ? node2142 : node2137;
												assign node2137 = (inp[4]) ? node2139 : 15'b000000111111111;
													assign node2139 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2142 = (inp[7]) ? 15'b000000011111111 : node2143;
													assign node2143 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2147 = (inp[9]) ? 15'b000000000111111 : node2148;
												assign node2148 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node2152 = (inp[7]) ? node2166 : node2153;
										assign node2153 = (inp[10]) ? node2161 : node2154;
											assign node2154 = (inp[4]) ? 15'b000000011111111 : node2155;
												assign node2155 = (inp[9]) ? node2157 : 15'b000000111111111;
													assign node2157 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2161 = (inp[9]) ? node2163 : 15'b000000011111111;
												assign node2163 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2166 = (inp[8]) ? node2178 : node2167;
											assign node2167 = (inp[10]) ? node2173 : node2168;
												assign node2168 = (inp[13]) ? 15'b000000011111111 : node2169;
													assign node2169 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2173 = (inp[0]) ? node2175 : 15'b000000011111111;
													assign node2175 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2178 = (inp[10]) ? node2184 : node2179;
												assign node2179 = (inp[0]) ? node2181 : 15'b000000001111111;
													assign node2181 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2184 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2187 = (inp[4]) ? node2237 : node2188;
									assign node2188 = (inp[13]) ? node2212 : node2189;
										assign node2189 = (inp[6]) ? node2203 : node2190;
											assign node2190 = (inp[0]) ? node2198 : node2191;
												assign node2191 = (inp[9]) ? node2195 : node2192;
													assign node2192 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2195 = (inp[7]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node2198 = (inp[7]) ? 15'b000000011111111 : node2199;
													assign node2199 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2203 = (inp[10]) ? node2205 : 15'b000000011111111;
												assign node2205 = (inp[7]) ? node2209 : node2206;
													assign node2206 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2209 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2212 = (inp[0]) ? node2226 : node2213;
											assign node2213 = (inp[6]) ? node2221 : node2214;
												assign node2214 = (inp[8]) ? node2218 : node2215;
													assign node2215 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2218 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2221 = (inp[7]) ? node2223 : 15'b000000011111111;
													assign node2223 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2226 = (inp[6]) ? node2232 : node2227;
												assign node2227 = (inp[7]) ? node2229 : 15'b000000011111111;
													assign node2229 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2232 = (inp[10]) ? node2234 : 15'b000000000111111;
													assign node2234 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2237 = (inp[7]) ? node2253 : node2238;
										assign node2238 = (inp[8]) ? node2244 : node2239;
											assign node2239 = (inp[13]) ? node2241 : 15'b000000011111111;
												assign node2241 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node2244 = (inp[6]) ? node2250 : node2245;
												assign node2245 = (inp[0]) ? 15'b000000000111111 : node2246;
													assign node2246 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node2250 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2253 = (inp[13]) ? node2265 : node2254;
											assign node2254 = (inp[9]) ? node2260 : node2255;
												assign node2255 = (inp[8]) ? 15'b000000000111111 : node2256;
													assign node2256 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2260 = (inp[0]) ? 15'b000000000011111 : node2261;
													assign node2261 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2265 = (inp[0]) ? node2269 : node2266;
												assign node2266 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node2269 = (inp[6]) ? 15'b000000000000111 : node2270;
													assign node2270 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node2274 = (inp[8]) ? node2432 : node2275;
							assign node2275 = (inp[7]) ? node2351 : node2276;
								assign node2276 = (inp[4]) ? node2312 : node2277;
									assign node2277 = (inp[13]) ? node2295 : node2278;
										assign node2278 = (inp[6]) ? node2288 : node2279;
											assign node2279 = (inp[10]) ? node2283 : node2280;
												assign node2280 = (inp[0]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node2283 = (inp[9]) ? 15'b000000111111111 : node2284;
													assign node2284 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2288 = (inp[2]) ? 15'b000000001111111 : node2289;
												assign node2289 = (inp[3]) ? node2291 : 15'b000001111111111;
													assign node2291 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2295 = (inp[2]) ? node2305 : node2296;
											assign node2296 = (inp[9]) ? node2300 : node2297;
												assign node2297 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2300 = (inp[10]) ? node2302 : 15'b000001111111111;
													assign node2302 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2305 = (inp[10]) ? node2307 : 15'b000000011111111;
												assign node2307 = (inp[0]) ? 15'b000000000111111 : node2308;
													assign node2308 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2312 = (inp[9]) ? node2334 : node2313;
										assign node2313 = (inp[10]) ? node2327 : node2314;
											assign node2314 = (inp[13]) ? node2320 : node2315;
												assign node2315 = (inp[6]) ? node2317 : 15'b000000111111111;
													assign node2317 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2320 = (inp[6]) ? node2324 : node2321;
													assign node2321 = (inp[3]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node2324 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2327 = (inp[0]) ? node2329 : 15'b000000011111111;
												assign node2329 = (inp[3]) ? 15'b000000001111111 : node2330;
													assign node2330 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2334 = (inp[3]) ? node2342 : node2335;
											assign node2335 = (inp[13]) ? node2337 : 15'b000000011111111;
												assign node2337 = (inp[2]) ? 15'b000000001111111 : node2338;
													assign node2338 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2342 = (inp[2]) ? node2346 : node2343;
												assign node2343 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node2346 = (inp[0]) ? node2348 : 15'b000000000111111;
													assign node2348 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2351 = (inp[6]) ? node2391 : node2352;
									assign node2352 = (inp[0]) ? node2374 : node2353;
										assign node2353 = (inp[10]) ? node2363 : node2354;
											assign node2354 = (inp[4]) ? node2360 : node2355;
												assign node2355 = (inp[9]) ? node2357 : 15'b000000111111111;
													assign node2357 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2360 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2363 = (inp[9]) ? node2369 : node2364;
												assign node2364 = (inp[2]) ? node2366 : 15'b000000011111111;
													assign node2366 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2369 = (inp[13]) ? node2371 : 15'b000000001111111;
													assign node2371 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2374 = (inp[9]) ? node2382 : node2375;
											assign node2375 = (inp[10]) ? node2377 : 15'b000000111111111;
												assign node2377 = (inp[2]) ? 15'b000000001111111 : node2378;
													assign node2378 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2382 = (inp[4]) ? node2388 : node2383;
												assign node2383 = (inp[3]) ? node2385 : 15'b000000001111111;
													assign node2385 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2388 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node2391 = (inp[4]) ? node2411 : node2392;
										assign node2392 = (inp[13]) ? node2402 : node2393;
											assign node2393 = (inp[2]) ? node2395 : 15'b000000011111111;
												assign node2395 = (inp[0]) ? node2399 : node2396;
													assign node2396 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node2399 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2402 = (inp[9]) ? node2408 : node2403;
												assign node2403 = (inp[10]) ? node2405 : 15'b000000001111111;
													assign node2405 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2408 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2411 = (inp[10]) ? node2421 : node2412;
											assign node2412 = (inp[2]) ? node2416 : node2413;
												assign node2413 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2416 = (inp[3]) ? node2418 : 15'b000000000111111;
													assign node2418 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2421 = (inp[9]) ? node2427 : node2422;
												assign node2422 = (inp[2]) ? node2424 : 15'b000000000111111;
													assign node2424 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node2427 = (inp[3]) ? node2429 : 15'b000000000011111;
													assign node2429 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node2432 = (inp[0]) ? node2514 : node2433;
								assign node2433 = (inp[10]) ? node2469 : node2434;
									assign node2434 = (inp[9]) ? node2448 : node2435;
										assign node2435 = (inp[7]) ? node2439 : node2436;
											assign node2436 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2439 = (inp[6]) ? node2445 : node2440;
												assign node2440 = (inp[3]) ? node2442 : 15'b000000011111111;
													assign node2442 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2445 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node2448 = (inp[2]) ? node2456 : node2449;
											assign node2449 = (inp[6]) ? node2451 : 15'b000000011111111;
												assign node2451 = (inp[13]) ? 15'b000000000111111 : node2452;
													assign node2452 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2456 = (inp[6]) ? node2464 : node2457;
												assign node2457 = (inp[7]) ? node2461 : node2458;
													assign node2458 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2461 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2464 = (inp[4]) ? node2466 : 15'b000000000111111;
													assign node2466 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2469 = (inp[2]) ? node2497 : node2470;
										assign node2470 = (inp[9]) ? node2484 : node2471;
											assign node2471 = (inp[3]) ? node2477 : node2472;
												assign node2472 = (inp[7]) ? node2474 : 15'b000000011111111;
													assign node2474 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2477 = (inp[4]) ? node2481 : node2478;
													assign node2478 = (inp[6]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node2481 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2484 = (inp[7]) ? node2492 : node2485;
												assign node2485 = (inp[4]) ? node2489 : node2486;
													assign node2486 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2489 = (inp[13]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node2492 = (inp[4]) ? node2494 : 15'b000000000111111;
													assign node2494 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2497 = (inp[13]) ? node2505 : node2498;
											assign node2498 = (inp[7]) ? 15'b000000000111111 : node2499;
												assign node2499 = (inp[3]) ? node2501 : 15'b000000111111111;
													assign node2501 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2505 = (inp[3]) ? node2509 : node2506;
												assign node2506 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2509 = (inp[9]) ? 15'b000000000001111 : node2510;
													assign node2510 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2514 = (inp[10]) ? node2550 : node2515;
									assign node2515 = (inp[2]) ? node2535 : node2516;
										assign node2516 = (inp[9]) ? node2526 : node2517;
											assign node2517 = (inp[13]) ? node2521 : node2518;
												assign node2518 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2521 = (inp[3]) ? node2523 : 15'b000000001111111;
													assign node2523 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2526 = (inp[3]) ? node2530 : node2527;
												assign node2527 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2530 = (inp[6]) ? node2532 : 15'b000000000111111;
													assign node2532 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2535 = (inp[3]) ? node2543 : node2536;
											assign node2536 = (inp[4]) ? node2538 : 15'b000000011111111;
												assign node2538 = (inp[9]) ? node2540 : 15'b000000001111111;
													assign node2540 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2543 = (inp[9]) ? node2545 : 15'b000000000011111;
												assign node2545 = (inp[7]) ? 15'b000000000011111 : node2546;
													assign node2546 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2550 = (inp[6]) ? node2566 : node2551;
										assign node2551 = (inp[7]) ? node2559 : node2552;
											assign node2552 = (inp[3]) ? node2556 : node2553;
												assign node2553 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2556 = (inp[4]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node2559 = (inp[4]) ? 15'b000000000011111 : node2560;
												assign node2560 = (inp[9]) ? node2562 : 15'b000000000111111;
													assign node2562 = (inp[13]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node2566 = (inp[13]) ? node2574 : node2567;
											assign node2567 = (inp[4]) ? node2571 : node2568;
												assign node2568 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2571 = (inp[7]) ? 15'b000000000011111 : 15'b000000000001111;
											assign node2574 = (inp[2]) ? node2580 : node2575;
												assign node2575 = (inp[3]) ? 15'b000000000001111 : node2576;
													assign node2576 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node2580 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
			assign node2583 = (inp[14]) ? node3903 : node2584;
				assign node2584 = (inp[5]) ? node3244 : node2585;
					assign node2585 = (inp[7]) ? node2933 : node2586;
						assign node2586 = (inp[9]) ? node2764 : node2587;
							assign node2587 = (inp[0]) ? node2683 : node2588;
								assign node2588 = (inp[13]) ? node2638 : node2589;
									assign node2589 = (inp[4]) ? node2615 : node2590;
										assign node2590 = (inp[3]) ? node2602 : node2591;
											assign node2591 = (inp[1]) ? node2597 : node2592;
												assign node2592 = (inp[8]) ? 15'b000111111111111 : node2593;
													assign node2593 = (inp[6]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node2597 = (inp[6]) ? 15'b000001111111111 : node2598;
													assign node2598 = (inp[2]) ? 15'b000001111111111 : 15'b000111111111111;
											assign node2602 = (inp[8]) ? node2608 : node2603;
												assign node2603 = (inp[10]) ? node2605 : 15'b000111111111111;
													assign node2605 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2608 = (inp[1]) ? node2612 : node2609;
													assign node2609 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2612 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2615 = (inp[10]) ? node2625 : node2616;
											assign node2616 = (inp[1]) ? node2620 : node2617;
												assign node2617 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2620 = (inp[6]) ? node2622 : 15'b000001111111111;
													assign node2622 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2625 = (inp[2]) ? node2633 : node2626;
												assign node2626 = (inp[8]) ? node2630 : node2627;
													assign node2627 = (inp[3]) ? 15'b000011111111111 : 15'b000001111111111;
													assign node2630 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2633 = (inp[1]) ? 15'b000000011111111 : node2634;
													assign node2634 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2638 = (inp[3]) ? node2666 : node2639;
										assign node2639 = (inp[2]) ? node2651 : node2640;
											assign node2640 = (inp[10]) ? node2646 : node2641;
												assign node2641 = (inp[4]) ? node2643 : 15'b000111111111111;
													assign node2643 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2646 = (inp[1]) ? node2648 : 15'b000001111111111;
													assign node2648 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2651 = (inp[1]) ? node2659 : node2652;
												assign node2652 = (inp[8]) ? node2656 : node2653;
													assign node2653 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2656 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2659 = (inp[10]) ? node2663 : node2660;
													assign node2660 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2663 = (inp[4]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node2666 = (inp[8]) ? node2678 : node2667;
											assign node2667 = (inp[4]) ? node2675 : node2668;
												assign node2668 = (inp[2]) ? node2672 : node2669;
													assign node2669 = (inp[10]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node2672 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2675 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2678 = (inp[10]) ? 15'b000000111111111 : node2679;
												assign node2679 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node2683 = (inp[13]) ? node2731 : node2684;
									assign node2684 = (inp[4]) ? node2704 : node2685;
										assign node2685 = (inp[10]) ? node2693 : node2686;
											assign node2686 = (inp[2]) ? node2688 : 15'b000011111111111;
												assign node2688 = (inp[8]) ? 15'b000000011111111 : node2689;
													assign node2689 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2693 = (inp[8]) ? node2699 : node2694;
												assign node2694 = (inp[1]) ? 15'b000001111111111 : node2695;
													assign node2695 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2699 = (inp[6]) ? 15'b000000111111111 : node2700;
													assign node2700 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2704 = (inp[1]) ? node2718 : node2705;
											assign node2705 = (inp[8]) ? node2713 : node2706;
												assign node2706 = (inp[10]) ? node2710 : node2707;
													assign node2707 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2710 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2713 = (inp[2]) ? 15'b000000011111111 : node2714;
													assign node2714 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2718 = (inp[2]) ? node2724 : node2719;
												assign node2719 = (inp[3]) ? node2721 : 15'b000000111111111;
													assign node2721 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2724 = (inp[6]) ? node2728 : node2725;
													assign node2725 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2728 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2731 = (inp[2]) ? node2749 : node2732;
										assign node2732 = (inp[10]) ? node2740 : node2733;
											assign node2733 = (inp[4]) ? 15'b000000111111111 : node2734;
												assign node2734 = (inp[6]) ? 15'b000001111111111 : node2735;
													assign node2735 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2740 = (inp[3]) ? node2742 : 15'b000000111111111;
												assign node2742 = (inp[6]) ? node2746 : node2743;
													assign node2743 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2746 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2749 = (inp[6]) ? node2761 : node2750;
											assign node2750 = (inp[10]) ? node2756 : node2751;
												assign node2751 = (inp[1]) ? node2753 : 15'b000000111111111;
													assign node2753 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2756 = (inp[4]) ? 15'b000000011111111 : node2757;
													assign node2757 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2761 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node2764 = (inp[10]) ? node2850 : node2765;
								assign node2765 = (inp[0]) ? node2809 : node2766;
									assign node2766 = (inp[13]) ? node2788 : node2767;
										assign node2767 = (inp[3]) ? node2777 : node2768;
											assign node2768 = (inp[1]) ? node2774 : node2769;
												assign node2769 = (inp[4]) ? 15'b000011111111111 : node2770;
													assign node2770 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2774 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2777 = (inp[6]) ? node2783 : node2778;
												assign node2778 = (inp[1]) ? 15'b000001111111111 : node2779;
													assign node2779 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2783 = (inp[2]) ? node2785 : 15'b000001111111111;
													assign node2785 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2788 = (inp[2]) ? node2800 : node2789;
											assign node2789 = (inp[8]) ? node2795 : node2790;
												assign node2790 = (inp[4]) ? 15'b000001111111111 : node2791;
													assign node2791 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2795 = (inp[4]) ? 15'b000000111111111 : node2796;
													assign node2796 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node2800 = (inp[8]) ? node2806 : node2801;
												assign node2801 = (inp[6]) ? 15'b000000111111111 : node2802;
													assign node2802 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2806 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2809 = (inp[13]) ? node2835 : node2810;
										assign node2810 = (inp[4]) ? node2822 : node2811;
											assign node2811 = (inp[8]) ? node2819 : node2812;
												assign node2812 = (inp[1]) ? node2816 : node2813;
													assign node2813 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2816 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2819 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node2822 = (inp[6]) ? node2830 : node2823;
												assign node2823 = (inp[3]) ? node2827 : node2824;
													assign node2824 = (inp[1]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node2827 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2830 = (inp[2]) ? 15'b000000001111111 : node2831;
													assign node2831 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2835 = (inp[2]) ? node2843 : node2836;
											assign node2836 = (inp[3]) ? 15'b000000011111111 : node2837;
												assign node2837 = (inp[8]) ? node2839 : 15'b000011111111111;
													assign node2839 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2843 = (inp[8]) ? node2845 : 15'b000000001111111;
												assign node2845 = (inp[1]) ? 15'b000000001111111 : node2846;
													assign node2846 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
								assign node2850 = (inp[6]) ? node2888 : node2851;
									assign node2851 = (inp[3]) ? node2867 : node2852;
										assign node2852 = (inp[13]) ? node2864 : node2853;
											assign node2853 = (inp[0]) ? node2859 : node2854;
												assign node2854 = (inp[2]) ? node2856 : 15'b000001111111111;
													assign node2856 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2859 = (inp[4]) ? 15'b000000001111111 : node2860;
													assign node2860 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2864 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node2867 = (inp[1]) ? node2879 : node2868;
											assign node2868 = (inp[2]) ? node2874 : node2869;
												assign node2869 = (inp[13]) ? node2871 : 15'b000001111111111;
													assign node2871 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2874 = (inp[13]) ? 15'b000000011111111 : node2875;
													assign node2875 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2879 = (inp[8]) ? node2883 : node2880;
												assign node2880 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2883 = (inp[4]) ? 15'b000000001111111 : node2884;
													assign node2884 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2888 = (inp[13]) ? node2910 : node2889;
										assign node2889 = (inp[1]) ? node2901 : node2890;
											assign node2890 = (inp[8]) ? node2896 : node2891;
												assign node2891 = (inp[3]) ? node2893 : 15'b000001111111111;
													assign node2893 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2896 = (inp[4]) ? node2898 : 15'b000000011111111;
													assign node2898 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2901 = (inp[8]) ? node2903 : 15'b000000011111111;
												assign node2903 = (inp[3]) ? node2907 : node2904;
													assign node2904 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2907 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node2910 = (inp[3]) ? node2918 : node2911;
											assign node2911 = (inp[1]) ? 15'b000000001111111 : node2912;
												assign node2912 = (inp[0]) ? node2914 : 15'b000000001111111;
													assign node2914 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2918 = (inp[0]) ? node2926 : node2919;
												assign node2919 = (inp[2]) ? node2923 : node2920;
													assign node2920 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2923 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2926 = (inp[8]) ? node2930 : node2927;
													assign node2927 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2930 = (inp[2]) ? 15'b000000000011111 : 15'b000000000011111;
						assign node2933 = (inp[4]) ? node3095 : node2934;
							assign node2934 = (inp[0]) ? node3002 : node2935;
								assign node2935 = (inp[1]) ? node2975 : node2936;
									assign node2936 = (inp[8]) ? node2958 : node2937;
										assign node2937 = (inp[6]) ? node2947 : node2938;
											assign node2938 = (inp[3]) ? node2942 : node2939;
												assign node2939 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2942 = (inp[9]) ? node2944 : 15'b000011111111111;
													assign node2944 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2947 = (inp[9]) ? node2953 : node2948;
												assign node2948 = (inp[13]) ? node2950 : 15'b000001111111111;
													assign node2950 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2953 = (inp[10]) ? 15'b000000111111111 : node2954;
													assign node2954 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2958 = (inp[13]) ? node2966 : node2959;
											assign node2959 = (inp[3]) ? node2961 : 15'b000001111111111;
												assign node2961 = (inp[2]) ? node2963 : 15'b000001111111111;
													assign node2963 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node2966 = (inp[6]) ? 15'b000000011111111 : node2967;
												assign node2967 = (inp[10]) ? node2971 : node2968;
													assign node2968 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2971 = (inp[9]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node2975 = (inp[3]) ? node2991 : node2976;
										assign node2976 = (inp[10]) ? node2984 : node2977;
											assign node2977 = (inp[8]) ? 15'b000000111111111 : node2978;
												assign node2978 = (inp[6]) ? 15'b000001111111111 : node2979;
													assign node2979 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node2984 = (inp[2]) ? 15'b000000011111111 : node2985;
												assign node2985 = (inp[13]) ? node2987 : 15'b000011111111111;
													assign node2987 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2991 = (inp[6]) ? node2999 : node2992;
											assign node2992 = (inp[10]) ? 15'b000000011111111 : node2993;
												assign node2993 = (inp[9]) ? node2995 : 15'b000000111111111;
													assign node2995 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2999 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node3002 = (inp[6]) ? node3054 : node3003;
									assign node3003 = (inp[3]) ? node3035 : node3004;
										assign node3004 = (inp[1]) ? node3020 : node3005;
											assign node3005 = (inp[8]) ? node3013 : node3006;
												assign node3006 = (inp[2]) ? node3010 : node3007;
													assign node3007 = (inp[10]) ? 15'b000011111111111 : 15'b000011111111111;
													assign node3010 = (inp[13]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node3013 = (inp[13]) ? node3017 : node3014;
													assign node3014 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3017 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3020 = (inp[9]) ? node3028 : node3021;
												assign node3021 = (inp[2]) ? node3025 : node3022;
													assign node3022 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3025 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3028 = (inp[13]) ? node3032 : node3029;
													assign node3029 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3032 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3035 = (inp[8]) ? node3047 : node3036;
											assign node3036 = (inp[10]) ? node3042 : node3037;
												assign node3037 = (inp[13]) ? node3039 : 15'b000000111111111;
													assign node3039 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3042 = (inp[1]) ? 15'b000000011111111 : node3043;
													assign node3043 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3047 = (inp[1]) ? 15'b000000000111111 : node3048;
												assign node3048 = (inp[2]) ? node3050 : 15'b000000011111111;
													assign node3050 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3054 = (inp[2]) ? node3078 : node3055;
										assign node3055 = (inp[9]) ? node3065 : node3056;
											assign node3056 = (inp[13]) ? node3062 : node3057;
												assign node3057 = (inp[1]) ? node3059 : 15'b000001111111111;
													assign node3059 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3062 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3065 = (inp[10]) ? node3073 : node3066;
												assign node3066 = (inp[13]) ? node3070 : node3067;
													assign node3067 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3070 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3073 = (inp[3]) ? 15'b000000001111111 : node3074;
													assign node3074 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3078 = (inp[1]) ? node3090 : node3079;
											assign node3079 = (inp[3]) ? node3087 : node3080;
												assign node3080 = (inp[10]) ? node3084 : node3081;
													assign node3081 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3084 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3087 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node3090 = (inp[9]) ? node3092 : 15'b000000001111111;
												assign node3092 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
							assign node3095 = (inp[1]) ? node3169 : node3096;
								assign node3096 = (inp[3]) ? node3130 : node3097;
									assign node3097 = (inp[6]) ? node3115 : node3098;
										assign node3098 = (inp[8]) ? node3108 : node3099;
											assign node3099 = (inp[9]) ? node3103 : node3100;
												assign node3100 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3103 = (inp[13]) ? 15'b000000111111111 : node3104;
													assign node3104 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3108 = (inp[13]) ? node3112 : node3109;
												assign node3109 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3112 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3115 = (inp[9]) ? node3121 : node3116;
											assign node3116 = (inp[13]) ? 15'b000000011111111 : node3117;
												assign node3117 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3121 = (inp[2]) ? 15'b000000001111111 : node3122;
												assign node3122 = (inp[0]) ? node3126 : node3123;
													assign node3123 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3126 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3130 = (inp[2]) ? node3148 : node3131;
										assign node3131 = (inp[13]) ? node3139 : node3132;
											assign node3132 = (inp[10]) ? node3136 : node3133;
												assign node3133 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3136 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3139 = (inp[10]) ? node3143 : node3140;
												assign node3140 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node3143 = (inp[0]) ? 15'b000000001111111 : node3144;
													assign node3144 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3148 = (inp[9]) ? node3158 : node3149;
											assign node3149 = (inp[6]) ? 15'b000000001111111 : node3150;
												assign node3150 = (inp[10]) ? node3154 : node3151;
													assign node3151 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3154 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3158 = (inp[8]) ? node3164 : node3159;
												assign node3159 = (inp[0]) ? node3161 : 15'b000000011111111;
													assign node3161 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node3164 = (inp[10]) ? 15'b000000000011111 : node3165;
													assign node3165 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3169 = (inp[6]) ? node3205 : node3170;
									assign node3170 = (inp[8]) ? node3184 : node3171;
										assign node3171 = (inp[0]) ? node3179 : node3172;
											assign node3172 = (inp[13]) ? 15'b000000111111111 : node3173;
												assign node3173 = (inp[2]) ? node3175 : 15'b000011111111111;
													assign node3175 = (inp[3]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node3179 = (inp[2]) ? 15'b000000001111111 : node3180;
												assign node3180 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3184 = (inp[10]) ? node3196 : node3185;
											assign node3185 = (inp[13]) ? node3191 : node3186;
												assign node3186 = (inp[0]) ? node3188 : 15'b000000111111111;
													assign node3188 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3191 = (inp[2]) ? 15'b000000001111111 : node3192;
													assign node3192 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3196 = (inp[3]) ? node3200 : node3197;
												assign node3197 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3200 = (inp[9]) ? 15'b000000000011111 : node3201;
													assign node3201 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3205 = (inp[8]) ? node3231 : node3206;
										assign node3206 = (inp[3]) ? node3220 : node3207;
											assign node3207 = (inp[13]) ? node3213 : node3208;
												assign node3208 = (inp[10]) ? 15'b000000011111111 : node3209;
													assign node3209 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3213 = (inp[9]) ? node3217 : node3214;
													assign node3214 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3217 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3220 = (inp[10]) ? node3226 : node3221;
												assign node3221 = (inp[0]) ? node3223 : 15'b000000001111111;
													assign node3223 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3226 = (inp[0]) ? 15'b000000000001111 : node3227;
													assign node3227 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3231 = (inp[2]) ? node3237 : node3232;
											assign node3232 = (inp[0]) ? node3234 : 15'b000000000111111;
												assign node3234 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3237 = (inp[10]) ? 15'b000000000011111 : node3238;
												assign node3238 = (inp[13]) ? node3240 : 15'b000000000111111;
													assign node3240 = (inp[3]) ? 15'b000000000011111 : 15'b000000000011111;
					assign node3244 = (inp[2]) ? node3576 : node3245;
						assign node3245 = (inp[9]) ? node3419 : node3246;
							assign node3246 = (inp[4]) ? node3336 : node3247;
								assign node3247 = (inp[7]) ? node3295 : node3248;
									assign node3248 = (inp[1]) ? node3272 : node3249;
										assign node3249 = (inp[13]) ? node3261 : node3250;
											assign node3250 = (inp[6]) ? node3256 : node3251;
												assign node3251 = (inp[10]) ? 15'b000011111111111 : node3252;
													assign node3252 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node3256 = (inp[3]) ? 15'b000001111111111 : node3257;
													assign node3257 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node3261 = (inp[10]) ? node3267 : node3262;
												assign node3262 = (inp[3]) ? 15'b000001111111111 : node3263;
													assign node3263 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3267 = (inp[0]) ? 15'b000000001111111 : node3268;
													assign node3268 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3272 = (inp[8]) ? node3284 : node3273;
											assign node3273 = (inp[0]) ? node3279 : node3274;
												assign node3274 = (inp[10]) ? node3276 : 15'b000111111111111;
													assign node3276 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3279 = (inp[13]) ? 15'b000000111111111 : node3280;
													assign node3280 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3284 = (inp[3]) ? node3290 : node3285;
												assign node3285 = (inp[13]) ? node3287 : 15'b000001111111111;
													assign node3287 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node3290 = (inp[10]) ? 15'b000000001111111 : node3291;
													assign node3291 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
									assign node3295 = (inp[0]) ? node3313 : node3296;
										assign node3296 = (inp[10]) ? node3306 : node3297;
											assign node3297 = (inp[3]) ? node3303 : node3298;
												assign node3298 = (inp[13]) ? 15'b000001111111111 : node3299;
													assign node3299 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3303 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3306 = (inp[13]) ? 15'b000000011111111 : node3307;
												assign node3307 = (inp[6]) ? node3309 : 15'b000001111111111;
													assign node3309 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3313 = (inp[1]) ? node3325 : node3314;
											assign node3314 = (inp[3]) ? node3318 : node3315;
												assign node3315 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3318 = (inp[10]) ? node3322 : node3319;
													assign node3319 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3322 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node3325 = (inp[3]) ? node3331 : node3326;
												assign node3326 = (inp[13]) ? node3328 : 15'b000000111111111;
													assign node3328 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3331 = (inp[6]) ? 15'b000000000111111 : node3332;
													assign node3332 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3336 = (inp[0]) ? node3386 : node3337;
									assign node3337 = (inp[1]) ? node3363 : node3338;
										assign node3338 = (inp[13]) ? node3352 : node3339;
											assign node3339 = (inp[10]) ? node3347 : node3340;
												assign node3340 = (inp[8]) ? node3344 : node3341;
													assign node3341 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3344 = (inp[7]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node3347 = (inp[7]) ? 15'b000000111111111 : node3348;
													assign node3348 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3352 = (inp[3]) ? node3360 : node3353;
												assign node3353 = (inp[8]) ? node3357 : node3354;
													assign node3354 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3357 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3360 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3363 = (inp[7]) ? node3379 : node3364;
											assign node3364 = (inp[6]) ? node3372 : node3365;
												assign node3365 = (inp[8]) ? node3369 : node3366;
													assign node3366 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3369 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3372 = (inp[3]) ? node3376 : node3373;
													assign node3373 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3376 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3379 = (inp[10]) ? 15'b000000001111111 : node3380;
												assign node3380 = (inp[3]) ? node3382 : 15'b000000011111111;
													assign node3382 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
									assign node3386 = (inp[6]) ? node3408 : node3387;
										assign node3387 = (inp[13]) ? node3395 : node3388;
											assign node3388 = (inp[3]) ? node3390 : 15'b000000011111111;
												assign node3390 = (inp[1]) ? 15'b000000011111111 : node3391;
													assign node3391 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3395 = (inp[8]) ? node3401 : node3396;
												assign node3396 = (inp[10]) ? node3398 : 15'b000000111111111;
													assign node3398 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3401 = (inp[3]) ? node3405 : node3402;
													assign node3402 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3405 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3408 = (inp[8]) ? node3414 : node3409;
											assign node3409 = (inp[3]) ? node3411 : 15'b000000011111111;
												assign node3411 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3414 = (inp[1]) ? 15'b000000000111111 : node3415;
												assign node3415 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node3419 = (inp[1]) ? node3491 : node3420;
								assign node3420 = (inp[4]) ? node3452 : node3421;
									assign node3421 = (inp[3]) ? node3441 : node3422;
										assign node3422 = (inp[8]) ? node3432 : node3423;
											assign node3423 = (inp[13]) ? node3429 : node3424;
												assign node3424 = (inp[0]) ? 15'b000001111111111 : node3425;
													assign node3425 = (inp[6]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node3429 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3432 = (inp[6]) ? node3438 : node3433;
												assign node3433 = (inp[7]) ? 15'b000000111111111 : node3434;
													assign node3434 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3438 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3441 = (inp[8]) ? node3445 : node3442;
											assign node3442 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3445 = (inp[7]) ? 15'b000000001111111 : node3446;
												assign node3446 = (inp[10]) ? 15'b000000001111111 : node3447;
													assign node3447 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
									assign node3452 = (inp[10]) ? node3472 : node3453;
										assign node3453 = (inp[8]) ? node3459 : node3454;
											assign node3454 = (inp[7]) ? node3456 : 15'b000000111111111;
												assign node3456 = (inp[3]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node3459 = (inp[6]) ? node3467 : node3460;
												assign node3460 = (inp[3]) ? node3464 : node3461;
													assign node3461 = (inp[13]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3464 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3467 = (inp[0]) ? node3469 : 15'b000000001111111;
													assign node3469 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3472 = (inp[0]) ? node3484 : node3473;
											assign node3473 = (inp[6]) ? node3479 : node3474;
												assign node3474 = (inp[13]) ? node3476 : 15'b000000011111111;
													assign node3476 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3479 = (inp[13]) ? node3481 : 15'b000000001111111;
													assign node3481 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3484 = (inp[13]) ? 15'b000000000011111 : node3485;
												assign node3485 = (inp[3]) ? 15'b000000000111111 : node3486;
													assign node3486 = (inp[8]) ? 15'b000000011111111 : 15'b000000001111111;
								assign node3491 = (inp[13]) ? node3539 : node3492;
									assign node3492 = (inp[8]) ? node3514 : node3493;
										assign node3493 = (inp[6]) ? node3501 : node3494;
											assign node3494 = (inp[7]) ? node3496 : 15'b000000111111111;
												assign node3496 = (inp[4]) ? node3498 : 15'b000000011111111;
													assign node3498 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3501 = (inp[3]) ? node3507 : node3502;
												assign node3502 = (inp[10]) ? node3504 : 15'b000000011111111;
													assign node3504 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node3507 = (inp[0]) ? node3511 : node3508;
													assign node3508 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3511 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3514 = (inp[10]) ? node3524 : node3515;
											assign node3515 = (inp[0]) ? node3521 : node3516;
												assign node3516 = (inp[7]) ? node3518 : 15'b000000011111111;
													assign node3518 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3521 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3524 = (inp[7]) ? node3532 : node3525;
												assign node3525 = (inp[3]) ? node3529 : node3526;
													assign node3526 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3529 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3532 = (inp[3]) ? node3536 : node3533;
													assign node3533 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3536 = (inp[0]) ? 15'b000000000111111 : 15'b000000000011111;
									assign node3539 = (inp[3]) ? node3559 : node3540;
										assign node3540 = (inp[0]) ? node3550 : node3541;
											assign node3541 = (inp[7]) ? node3543 : 15'b000000011111111;
												assign node3543 = (inp[10]) ? node3547 : node3544;
													assign node3544 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3547 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3550 = (inp[4]) ? node3554 : node3551;
												assign node3551 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3554 = (inp[7]) ? 15'b000000000011111 : node3555;
													assign node3555 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node3559 = (inp[7]) ? node3563 : node3560;
											assign node3560 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3563 = (inp[8]) ? node3569 : node3564;
												assign node3564 = (inp[0]) ? node3566 : 15'b000000000111111;
													assign node3566 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3569 = (inp[4]) ? node3573 : node3570;
													assign node3570 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node3573 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node3576 = (inp[3]) ? node3736 : node3577;
							assign node3577 = (inp[9]) ? node3663 : node3578;
								assign node3578 = (inp[8]) ? node3632 : node3579;
									assign node3579 = (inp[10]) ? node3605 : node3580;
										assign node3580 = (inp[6]) ? node3594 : node3581;
											assign node3581 = (inp[7]) ? node3589 : node3582;
												assign node3582 = (inp[0]) ? node3586 : node3583;
													assign node3583 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3586 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3589 = (inp[13]) ? 15'b000000011111111 : node3590;
													assign node3590 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3594 = (inp[1]) ? node3600 : node3595;
												assign node3595 = (inp[0]) ? 15'b000000111111111 : node3596;
													assign node3596 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3600 = (inp[4]) ? 15'b000000011111111 : node3601;
													assign node3601 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3605 = (inp[4]) ? node3617 : node3606;
											assign node3606 = (inp[13]) ? node3612 : node3607;
												assign node3607 = (inp[7]) ? node3609 : 15'b000001111111111;
													assign node3609 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3612 = (inp[7]) ? 15'b000000001111111 : node3613;
													assign node3613 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3617 = (inp[0]) ? node3625 : node3618;
												assign node3618 = (inp[1]) ? node3622 : node3619;
													assign node3619 = (inp[13]) ? 15'b000000111111111 : 15'b000000011111111;
													assign node3622 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3625 = (inp[6]) ? node3629 : node3626;
													assign node3626 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3629 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3632 = (inp[0]) ? node3644 : node3633;
										assign node3633 = (inp[7]) ? node3639 : node3634;
											assign node3634 = (inp[13]) ? 15'b000000111111111 : node3635;
												assign node3635 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3639 = (inp[10]) ? node3641 : 15'b000000011111111;
												assign node3641 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3644 = (inp[13]) ? node3652 : node3645;
											assign node3645 = (inp[10]) ? node3647 : 15'b000000011111111;
												assign node3647 = (inp[1]) ? 15'b000000001111111 : node3648;
													assign node3648 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3652 = (inp[4]) ? node3656 : node3653;
												assign node3653 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3656 = (inp[6]) ? node3660 : node3657;
													assign node3657 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3660 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3663 = (inp[13]) ? node3701 : node3664;
									assign node3664 = (inp[4]) ? node3686 : node3665;
										assign node3665 = (inp[7]) ? node3677 : node3666;
											assign node3666 = (inp[6]) ? node3672 : node3667;
												assign node3667 = (inp[8]) ? node3669 : 15'b000000111111111;
													assign node3669 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3672 = (inp[10]) ? node3674 : 15'b000000111111111;
													assign node3674 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3677 = (inp[6]) ? node3681 : node3678;
												assign node3678 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3681 = (inp[1]) ? node3683 : 15'b000000001111111;
													assign node3683 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3686 = (inp[1]) ? node3694 : node3687;
											assign node3687 = (inp[6]) ? 15'b000000001111111 : node3688;
												assign node3688 = (inp[7]) ? 15'b000000000111111 : node3689;
													assign node3689 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node3694 = (inp[0]) ? 15'b000000000111111 : node3695;
												assign node3695 = (inp[6]) ? node3697 : 15'b000000001111111;
													assign node3697 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3701 = (inp[7]) ? node3717 : node3702;
										assign node3702 = (inp[0]) ? node3710 : node3703;
											assign node3703 = (inp[8]) ? node3705 : 15'b000000011111111;
												assign node3705 = (inp[10]) ? node3707 : 15'b000000001111111;
													assign node3707 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3710 = (inp[10]) ? 15'b000000000111111 : node3711;
												assign node3711 = (inp[6]) ? node3713 : 15'b000000001111111;
													assign node3713 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3717 = (inp[1]) ? node3727 : node3718;
											assign node3718 = (inp[8]) ? node3722 : node3719;
												assign node3719 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3722 = (inp[6]) ? node3724 : 15'b000000000111111;
													assign node3724 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node3727 = (inp[8]) ? node3733 : node3728;
												assign node3728 = (inp[10]) ? node3730 : 15'b000000000111111;
													assign node3730 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3733 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3736 = (inp[10]) ? node3818 : node3737;
								assign node3737 = (inp[0]) ? node3779 : node3738;
									assign node3738 = (inp[6]) ? node3760 : node3739;
										assign node3739 = (inp[9]) ? node3747 : node3740;
											assign node3740 = (inp[8]) ? node3742 : 15'b000000111111111;
												assign node3742 = (inp[13]) ? 15'b000000011111111 : node3743;
													assign node3743 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3747 = (inp[1]) ? node3755 : node3748;
												assign node3748 = (inp[7]) ? node3752 : node3749;
													assign node3749 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3752 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3755 = (inp[13]) ? node3757 : 15'b000000001111111;
													assign node3757 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3760 = (inp[1]) ? node3768 : node3761;
											assign node3761 = (inp[13]) ? 15'b000000001111111 : node3762;
												assign node3762 = (inp[9]) ? node3764 : 15'b000000011111111;
													assign node3764 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3768 = (inp[4]) ? node3774 : node3769;
												assign node3769 = (inp[7]) ? 15'b000000001111111 : node3770;
													assign node3770 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3774 = (inp[7]) ? 15'b000000000111111 : node3775;
													assign node3775 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3779 = (inp[13]) ? node3795 : node3780;
										assign node3780 = (inp[7]) ? node3792 : node3781;
											assign node3781 = (inp[6]) ? node3787 : node3782;
												assign node3782 = (inp[4]) ? 15'b000000011111111 : node3783;
													assign node3783 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3787 = (inp[9]) ? 15'b000000001111111 : node3788;
													assign node3788 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node3792 = (inp[8]) ? 15'b000000000001111 : 15'b000000001111111;
										assign node3795 = (inp[1]) ? node3807 : node3796;
											assign node3796 = (inp[4]) ? node3800 : node3797;
												assign node3797 = (inp[7]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node3800 = (inp[6]) ? node3804 : node3801;
													assign node3801 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3804 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node3807 = (inp[4]) ? node3813 : node3808;
												assign node3808 = (inp[7]) ? node3810 : 15'b000000000111111;
													assign node3810 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3813 = (inp[9]) ? node3815 : 15'b000000000001111;
													assign node3815 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node3818 = (inp[8]) ? node3854 : node3819;
									assign node3819 = (inp[13]) ? node3833 : node3820;
										assign node3820 = (inp[1]) ? node3828 : node3821;
											assign node3821 = (inp[0]) ? 15'b000000001111111 : node3822;
												assign node3822 = (inp[7]) ? node3824 : 15'b000000011111111;
													assign node3824 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node3828 = (inp[7]) ? node3830 : 15'b000000000111111;
												assign node3830 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node3833 = (inp[7]) ? node3841 : node3834;
											assign node3834 = (inp[6]) ? 15'b000000000111111 : node3835;
												assign node3835 = (inp[9]) ? 15'b000000000111111 : node3836;
													assign node3836 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3841 = (inp[6]) ? node3849 : node3842;
												assign node3842 = (inp[4]) ? node3846 : node3843;
													assign node3843 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3846 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3849 = (inp[0]) ? node3851 : 15'b000000000011111;
													assign node3851 = (inp[4]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node3854 = (inp[6]) ? node3880 : node3855;
										assign node3855 = (inp[0]) ? node3869 : node3856;
											assign node3856 = (inp[13]) ? node3862 : node3857;
												assign node3857 = (inp[4]) ? 15'b000000000111111 : node3858;
													assign node3858 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3862 = (inp[1]) ? node3866 : node3863;
													assign node3863 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3866 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3869 = (inp[7]) ? node3875 : node3870;
												assign node3870 = (inp[13]) ? node3872 : 15'b000000000111111;
													assign node3872 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3875 = (inp[1]) ? node3877 : 15'b000000000011111;
													assign node3877 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node3880 = (inp[1]) ? node3892 : node3881;
											assign node3881 = (inp[4]) ? node3885 : node3882;
												assign node3882 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3885 = (inp[9]) ? node3889 : node3886;
													assign node3886 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3889 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node3892 = (inp[9]) ? node3896 : node3893;
												assign node3893 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node3896 = (inp[7]) ? node3900 : node3897;
													assign node3897 = (inp[13]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node3900 = (inp[4]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node3903 = (inp[2]) ? node4583 : node3904;
					assign node3904 = (inp[13]) ? node4258 : node3905;
						assign node3905 = (inp[1]) ? node4085 : node3906;
							assign node3906 = (inp[10]) ? node3996 : node3907;
								assign node3907 = (inp[8]) ? node3953 : node3908;
									assign node3908 = (inp[7]) ? node3932 : node3909;
										assign node3909 = (inp[6]) ? node3925 : node3910;
											assign node3910 = (inp[3]) ? node3918 : node3911;
												assign node3911 = (inp[5]) ? node3915 : node3912;
													assign node3912 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node3915 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3918 = (inp[9]) ? node3922 : node3919;
													assign node3919 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3922 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3925 = (inp[0]) ? node3929 : node3926;
												assign node3926 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3929 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node3932 = (inp[0]) ? node3944 : node3933;
											assign node3933 = (inp[3]) ? node3939 : node3934;
												assign node3934 = (inp[5]) ? node3936 : 15'b000011111111111;
													assign node3936 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node3939 = (inp[5]) ? 15'b000000111111111 : node3940;
													assign node3940 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3944 = (inp[6]) ? 15'b000000011111111 : node3945;
												assign node3945 = (inp[5]) ? node3949 : node3946;
													assign node3946 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3949 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3953 = (inp[5]) ? node3977 : node3954;
										assign node3954 = (inp[9]) ? node3966 : node3955;
											assign node3955 = (inp[7]) ? node3961 : node3956;
												assign node3956 = (inp[0]) ? 15'b000001111111111 : node3957;
													assign node3957 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3961 = (inp[6]) ? 15'b000000011111111 : node3962;
													assign node3962 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node3966 = (inp[0]) ? node3970 : node3967;
												assign node3967 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3970 = (inp[3]) ? node3974 : node3971;
													assign node3971 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3974 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3977 = (inp[4]) ? node3985 : node3978;
											assign node3978 = (inp[9]) ? 15'b000000011111111 : node3979;
												assign node3979 = (inp[6]) ? node3981 : 15'b000000111111111;
													assign node3981 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3985 = (inp[7]) ? node3989 : node3986;
												assign node3986 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3989 = (inp[3]) ? node3993 : node3990;
													assign node3990 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3993 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3996 = (inp[6]) ? node4042 : node3997;
									assign node3997 = (inp[3]) ? node4027 : node3998;
										assign node3998 = (inp[8]) ? node4014 : node3999;
											assign node3999 = (inp[7]) ? node4007 : node4000;
												assign node4000 = (inp[5]) ? node4004 : node4001;
													assign node4001 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4004 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4007 = (inp[9]) ? node4011 : node4008;
													assign node4008 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4011 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4014 = (inp[4]) ? node4022 : node4015;
												assign node4015 = (inp[0]) ? node4019 : node4016;
													assign node4016 = (inp[5]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node4019 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4022 = (inp[0]) ? 15'b000000001111111 : node4023;
													assign node4023 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4027 = (inp[5]) ? node4035 : node4028;
											assign node4028 = (inp[9]) ? node4030 : 15'b000000111111111;
												assign node4030 = (inp[7]) ? node4032 : 15'b000000111111111;
													assign node4032 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4035 = (inp[4]) ? node4037 : 15'b000000011111111;
												assign node4037 = (inp[9]) ? 15'b000000001111111 : node4038;
													assign node4038 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4042 = (inp[5]) ? node4064 : node4043;
										assign node4043 = (inp[3]) ? node4051 : node4044;
											assign node4044 = (inp[9]) ? 15'b000000011111111 : node4045;
												assign node4045 = (inp[4]) ? node4047 : 15'b000000111111111;
													assign node4047 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4051 = (inp[7]) ? node4057 : node4052;
												assign node4052 = (inp[4]) ? node4054 : 15'b000000011111111;
													assign node4054 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4057 = (inp[4]) ? node4061 : node4058;
													assign node4058 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4061 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4064 = (inp[4]) ? node4076 : node4065;
											assign node4065 = (inp[0]) ? node4071 : node4066;
												assign node4066 = (inp[7]) ? node4068 : 15'b000000011111111;
													assign node4068 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4071 = (inp[8]) ? node4073 : 15'b000000011111111;
													assign node4073 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4076 = (inp[7]) ? node4078 : 15'b000000001111111;
												assign node4078 = (inp[8]) ? node4082 : node4079;
													assign node4079 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node4082 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
							assign node4085 = (inp[5]) ? node4175 : node4086;
								assign node4086 = (inp[0]) ? node4134 : node4087;
									assign node4087 = (inp[4]) ? node4115 : node4088;
										assign node4088 = (inp[3]) ? node4102 : node4089;
											assign node4089 = (inp[9]) ? node4097 : node4090;
												assign node4090 = (inp[8]) ? node4094 : node4091;
													assign node4091 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4094 = (inp[10]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node4097 = (inp[7]) ? 15'b000000111111111 : node4098;
													assign node4098 = (inp[6]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node4102 = (inp[8]) ? node4110 : node4103;
												assign node4103 = (inp[10]) ? node4107 : node4104;
													assign node4104 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4107 = (inp[9]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node4110 = (inp[7]) ? node4112 : 15'b000000111111111;
													assign node4112 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4115 = (inp[7]) ? node4123 : node4116;
											assign node4116 = (inp[6]) ? 15'b000000011111111 : node4117;
												assign node4117 = (inp[3]) ? node4119 : 15'b000001111111111;
													assign node4119 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4123 = (inp[8]) ? node4129 : node4124;
												assign node4124 = (inp[6]) ? node4126 : 15'b000000111111111;
													assign node4126 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4129 = (inp[9]) ? node4131 : 15'b000000011111111;
													assign node4131 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4134 = (inp[9]) ? node4156 : node4135;
										assign node4135 = (inp[4]) ? node4145 : node4136;
											assign node4136 = (inp[7]) ? node4138 : 15'b000000111111111;
												assign node4138 = (inp[8]) ? node4142 : node4139;
													assign node4139 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4142 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4145 = (inp[7]) ? node4151 : node4146;
												assign node4146 = (inp[8]) ? node4148 : 15'b000000011111111;
													assign node4148 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4151 = (inp[10]) ? node4153 : 15'b000000011111111;
													assign node4153 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4156 = (inp[4]) ? node4170 : node4157;
											assign node4157 = (inp[8]) ? node4163 : node4158;
												assign node4158 = (inp[6]) ? 15'b000000001111111 : node4159;
													assign node4159 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node4163 = (inp[7]) ? node4167 : node4164;
													assign node4164 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4167 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4170 = (inp[8]) ? 15'b000000000111111 : node4171;
												assign node4171 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node4175 = (inp[9]) ? node4209 : node4176;
									assign node4176 = (inp[10]) ? node4194 : node4177;
										assign node4177 = (inp[0]) ? node4187 : node4178;
											assign node4178 = (inp[7]) ? node4180 : 15'b000000111111111;
												assign node4180 = (inp[6]) ? node4184 : node4181;
													assign node4181 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4184 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4187 = (inp[7]) ? node4191 : node4188;
												assign node4188 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4191 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4194 = (inp[6]) ? node4202 : node4195;
											assign node4195 = (inp[4]) ? node4197 : 15'b000000011111111;
												assign node4197 = (inp[0]) ? 15'b000000001111111 : node4198;
													assign node4198 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4202 = (inp[7]) ? node4204 : 15'b000000001111111;
												assign node4204 = (inp[0]) ? 15'b000000000111111 : node4205;
													assign node4205 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
									assign node4209 = (inp[7]) ? node4237 : node4210;
										assign node4210 = (inp[8]) ? node4222 : node4211;
											assign node4211 = (inp[10]) ? node4215 : node4212;
												assign node4212 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4215 = (inp[0]) ? node4219 : node4216;
													assign node4216 = (inp[6]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4219 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4222 = (inp[3]) ? node4230 : node4223;
												assign node4223 = (inp[6]) ? node4227 : node4224;
													assign node4224 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4227 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4230 = (inp[10]) ? node4234 : node4231;
													assign node4231 = (inp[6]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node4234 = (inp[4]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node4237 = (inp[3]) ? node4247 : node4238;
											assign node4238 = (inp[4]) ? node4242 : node4239;
												assign node4239 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4242 = (inp[0]) ? 15'b000000000011111 : node4243;
													assign node4243 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node4247 = (inp[4]) ? node4253 : node4248;
												assign node4248 = (inp[6]) ? node4250 : 15'b000000000111111;
													assign node4250 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4253 = (inp[6]) ? 15'b000000000001111 : node4254;
													assign node4254 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node4258 = (inp[7]) ? node4414 : node4259;
							assign node4259 = (inp[8]) ? node4331 : node4260;
								assign node4260 = (inp[9]) ? node4294 : node4261;
									assign node4261 = (inp[4]) ? node4279 : node4262;
										assign node4262 = (inp[6]) ? node4274 : node4263;
											assign node4263 = (inp[0]) ? node4269 : node4264;
												assign node4264 = (inp[3]) ? 15'b000001111111111 : node4265;
													assign node4265 = (inp[5]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node4269 = (inp[1]) ? 15'b000000011111111 : node4270;
													assign node4270 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4274 = (inp[10]) ? 15'b000000111111111 : node4275;
												assign node4275 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4279 = (inp[10]) ? node4287 : node4280;
											assign node4280 = (inp[5]) ? 15'b000000011111111 : node4281;
												assign node4281 = (inp[0]) ? node4283 : 15'b000011111111111;
													assign node4283 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4287 = (inp[1]) ? node4289 : 15'b000000011111111;
												assign node4289 = (inp[0]) ? 15'b000000001111111 : node4290;
													assign node4290 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4294 = (inp[10]) ? node4312 : node4295;
										assign node4295 = (inp[5]) ? node4307 : node4296;
											assign node4296 = (inp[3]) ? node4302 : node4297;
												assign node4297 = (inp[4]) ? 15'b000000111111111 : node4298;
													assign node4298 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4302 = (inp[0]) ? 15'b000000000111111 : node4303;
													assign node4303 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4307 = (inp[6]) ? node4309 : 15'b000000011111111;
												assign node4309 = (inp[1]) ? 15'b000000011111111 : 15'b000000000111111;
										assign node4312 = (inp[3]) ? node4320 : node4313;
											assign node4313 = (inp[4]) ? node4315 : 15'b000000011111111;
												assign node4315 = (inp[5]) ? node4317 : 15'b000000001111111;
													assign node4317 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4320 = (inp[5]) ? node4326 : node4321;
												assign node4321 = (inp[0]) ? 15'b000000000111111 : node4322;
													assign node4322 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4326 = (inp[1]) ? 15'b000000000011111 : node4327;
													assign node4327 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node4331 = (inp[5]) ? node4379 : node4332;
									assign node4332 = (inp[10]) ? node4358 : node4333;
										assign node4333 = (inp[1]) ? node4347 : node4334;
											assign node4334 = (inp[9]) ? node4342 : node4335;
												assign node4335 = (inp[6]) ? node4339 : node4336;
													assign node4336 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4339 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node4342 = (inp[0]) ? node4344 : 15'b000000011111111;
													assign node4344 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4347 = (inp[9]) ? node4353 : node4348;
												assign node4348 = (inp[3]) ? node4350 : 15'b000000011111111;
													assign node4350 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4353 = (inp[3]) ? 15'b000000001111111 : node4354;
													assign node4354 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4358 = (inp[4]) ? node4372 : node4359;
											assign node4359 = (inp[9]) ? node4365 : node4360;
												assign node4360 = (inp[3]) ? 15'b000000011111111 : node4361;
													assign node4361 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4365 = (inp[3]) ? node4369 : node4366;
													assign node4366 = (inp[6]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node4369 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4372 = (inp[9]) ? 15'b000000000011111 : node4373;
												assign node4373 = (inp[6]) ? node4375 : 15'b000000001111111;
													assign node4375 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4379 = (inp[9]) ? node4399 : node4380;
										assign node4380 = (inp[10]) ? node4392 : node4381;
											assign node4381 = (inp[1]) ? node4389 : node4382;
												assign node4382 = (inp[6]) ? node4386 : node4383;
													assign node4383 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node4386 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4389 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node4392 = (inp[1]) ? 15'b000000001111111 : node4393;
												assign node4393 = (inp[0]) ? 15'b000000000111111 : node4394;
													assign node4394 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4399 = (inp[1]) ? node4405 : node4400;
											assign node4400 = (inp[4]) ? 15'b000000000111111 : node4401;
												assign node4401 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4405 = (inp[10]) ? node4411 : node4406;
												assign node4406 = (inp[0]) ? node4408 : 15'b000000000111111;
													assign node4408 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4411 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node4414 = (inp[4]) ? node4492 : node4415;
								assign node4415 = (inp[10]) ? node4449 : node4416;
									assign node4416 = (inp[3]) ? node4438 : node4417;
										assign node4417 = (inp[5]) ? node4431 : node4418;
											assign node4418 = (inp[9]) ? node4426 : node4419;
												assign node4419 = (inp[0]) ? node4423 : node4420;
													assign node4420 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4423 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4426 = (inp[1]) ? 15'b000000011111111 : node4427;
													assign node4427 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node4431 = (inp[1]) ? 15'b000000001111111 : node4432;
												assign node4432 = (inp[9]) ? node4434 : 15'b000000111111111;
													assign node4434 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4438 = (inp[9]) ? node4446 : node4439;
											assign node4439 = (inp[8]) ? node4443 : node4440;
												assign node4440 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4443 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4446 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4449 = (inp[6]) ? node4463 : node4450;
										assign node4450 = (inp[8]) ? node4456 : node4451;
											assign node4451 = (inp[9]) ? 15'b000000011111111 : node4452;
												assign node4452 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4456 = (inp[0]) ? node4458 : 15'b000000001111111;
												assign node4458 = (inp[5]) ? 15'b000000000111111 : node4459;
													assign node4459 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node4463 = (inp[0]) ? node4479 : node4464;
											assign node4464 = (inp[9]) ? node4472 : node4465;
												assign node4465 = (inp[8]) ? node4469 : node4466;
													assign node4466 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node4469 = (inp[5]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node4472 = (inp[5]) ? node4476 : node4473;
													assign node4473 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4476 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4479 = (inp[1]) ? node4487 : node4480;
												assign node4480 = (inp[8]) ? node4484 : node4481;
													assign node4481 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4484 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4487 = (inp[3]) ? node4489 : 15'b000000000011111;
													assign node4489 = (inp[5]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node4492 = (inp[0]) ? node4536 : node4493;
									assign node4493 = (inp[5]) ? node4513 : node4494;
										assign node4494 = (inp[1]) ? node4500 : node4495;
											assign node4495 = (inp[9]) ? 15'b000000000111111 : node4496;
												assign node4496 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4500 = (inp[10]) ? node4508 : node4501;
												assign node4501 = (inp[8]) ? node4505 : node4502;
													assign node4502 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4505 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4508 = (inp[6]) ? node4510 : 15'b000000001111111;
													assign node4510 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4513 = (inp[1]) ? node4521 : node4514;
											assign node4514 = (inp[6]) ? node4516 : 15'b000000001111111;
												assign node4516 = (inp[3]) ? 15'b000000000011111 : node4517;
													assign node4517 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4521 = (inp[10]) ? node4529 : node4522;
												assign node4522 = (inp[9]) ? node4526 : node4523;
													assign node4523 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4526 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4529 = (inp[8]) ? node4533 : node4530;
													assign node4530 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4533 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node4536 = (inp[9]) ? node4558 : node4537;
										assign node4537 = (inp[8]) ? node4549 : node4538;
											assign node4538 = (inp[3]) ? node4546 : node4539;
												assign node4539 = (inp[10]) ? node4543 : node4540;
													assign node4540 = (inp[1]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4543 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node4546 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node4549 = (inp[1]) ? 15'b000000000011111 : node4550;
												assign node4550 = (inp[3]) ? node4554 : node4551;
													assign node4551 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4554 = (inp[6]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node4558 = (inp[5]) ? node4572 : node4559;
											assign node4559 = (inp[10]) ? node4565 : node4560;
												assign node4560 = (inp[6]) ? node4562 : 15'b000000000111111;
													assign node4562 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4565 = (inp[8]) ? node4569 : node4566;
													assign node4566 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4569 = (inp[3]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node4572 = (inp[1]) ? node4578 : node4573;
												assign node4573 = (inp[6]) ? node4575 : 15'b000000001111111;
													assign node4575 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node4578 = (inp[3]) ? node4580 : 15'b000000000001111;
													assign node4580 = (inp[8]) ? 15'b000000000000111 : 15'b000000000000111;
					assign node4583 = (inp[3]) ? node4879 : node4584;
						assign node4584 = (inp[9]) ? node4716 : node4585;
							assign node4585 = (inp[1]) ? node4649 : node4586;
								assign node4586 = (inp[10]) ? node4612 : node4587;
									assign node4587 = (inp[7]) ? node4605 : node4588;
										assign node4588 = (inp[4]) ? node4598 : node4589;
											assign node4589 = (inp[13]) ? node4595 : node4590;
												assign node4590 = (inp[0]) ? 15'b000001111111111 : node4591;
													assign node4591 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4595 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node4598 = (inp[8]) ? node4600 : 15'b000000111111111;
												assign node4600 = (inp[0]) ? 15'b000000001111111 : node4601;
													assign node4601 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4605 = (inp[4]) ? node4609 : node4606;
											assign node4606 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4609 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4612 = (inp[6]) ? node4632 : node4613;
										assign node4613 = (inp[13]) ? node4625 : node4614;
											assign node4614 = (inp[8]) ? node4620 : node4615;
												assign node4615 = (inp[4]) ? 15'b000000111111111 : node4616;
													assign node4616 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4620 = (inp[0]) ? 15'b000000011111111 : node4621;
													assign node4621 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node4625 = (inp[4]) ? node4627 : 15'b000000011111111;
												assign node4627 = (inp[0]) ? 15'b000000000111111 : node4628;
													assign node4628 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4632 = (inp[0]) ? node4640 : node4633;
											assign node4633 = (inp[4]) ? 15'b000000001111111 : node4634;
												assign node4634 = (inp[8]) ? node4636 : 15'b000000011111111;
													assign node4636 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4640 = (inp[8]) ? node4646 : node4641;
												assign node4641 = (inp[5]) ? node4643 : 15'b000000001111111;
													assign node4643 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node4646 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node4649 = (inp[5]) ? node4689 : node4650;
									assign node4650 = (inp[13]) ? node4668 : node4651;
										assign node4651 = (inp[10]) ? node4661 : node4652;
											assign node4652 = (inp[8]) ? node4658 : node4653;
												assign node4653 = (inp[7]) ? 15'b000000011111111 : node4654;
													assign node4654 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4658 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4661 = (inp[7]) ? 15'b000000001111111 : node4662;
												assign node4662 = (inp[6]) ? node4664 : 15'b000000011111111;
													assign node4664 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4668 = (inp[6]) ? node4682 : node4669;
											assign node4669 = (inp[10]) ? node4675 : node4670;
												assign node4670 = (inp[7]) ? 15'b000000011111111 : node4671;
													assign node4671 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4675 = (inp[7]) ? node4679 : node4676;
													assign node4676 = (inp[4]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4679 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4682 = (inp[4]) ? node4684 : 15'b000000001111111;
												assign node4684 = (inp[0]) ? 15'b000000000011111 : node4685;
													assign node4685 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4689 = (inp[0]) ? node4701 : node4690;
										assign node4690 = (inp[6]) ? node4694 : node4691;
											assign node4691 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4694 = (inp[13]) ? 15'b000000000111111 : node4695;
												assign node4695 = (inp[4]) ? node4697 : 15'b000000001111111;
													assign node4697 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4701 = (inp[7]) ? node4705 : node4702;
											assign node4702 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4705 = (inp[13]) ? node4711 : node4706;
												assign node4706 = (inp[6]) ? 15'b000000000111111 : node4707;
													assign node4707 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node4711 = (inp[8]) ? node4713 : 15'b000000000111111;
													assign node4713 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node4716 = (inp[5]) ? node4796 : node4717;
								assign node4717 = (inp[13]) ? node4755 : node4718;
									assign node4718 = (inp[1]) ? node4742 : node4719;
										assign node4719 = (inp[7]) ? node4733 : node4720;
											assign node4720 = (inp[8]) ? node4726 : node4721;
												assign node4721 = (inp[4]) ? node4723 : 15'b000000111111111;
													assign node4723 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node4726 = (inp[10]) ? node4730 : node4727;
													assign node4727 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4730 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4733 = (inp[8]) ? node4739 : node4734;
												assign node4734 = (inp[4]) ? node4736 : 15'b000000011111111;
													assign node4736 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4739 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4742 = (inp[10]) ? node4748 : node4743;
											assign node4743 = (inp[0]) ? 15'b000000001111111 : node4744;
												assign node4744 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4748 = (inp[6]) ? node4750 : 15'b000000001111111;
												assign node4750 = (inp[8]) ? node4752 : 15'b000000000111111;
													assign node4752 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4755 = (inp[0]) ? node4773 : node4756;
										assign node4756 = (inp[4]) ? node4762 : node4757;
											assign node4757 = (inp[10]) ? node4759 : 15'b000000011111111;
												assign node4759 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4762 = (inp[1]) ? node4768 : node4763;
												assign node4763 = (inp[8]) ? node4765 : 15'b000000011111111;
													assign node4765 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4768 = (inp[10]) ? 15'b000000000011111 : node4769;
													assign node4769 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node4773 = (inp[8]) ? node4783 : node4774;
											assign node4774 = (inp[4]) ? node4778 : node4775;
												assign node4775 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4778 = (inp[10]) ? node4780 : 15'b000000000111111;
													assign node4780 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4783 = (inp[4]) ? node4791 : node4784;
												assign node4784 = (inp[1]) ? node4788 : node4785;
													assign node4785 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4788 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4791 = (inp[10]) ? node4793 : 15'b000000000011111;
													assign node4793 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node4796 = (inp[13]) ? node4838 : node4797;
									assign node4797 = (inp[4]) ? node4815 : node4798;
										assign node4798 = (inp[1]) ? node4808 : node4799;
											assign node4799 = (inp[7]) ? node4805 : node4800;
												assign node4800 = (inp[8]) ? 15'b000000011111111 : node4801;
													assign node4801 = (inp[6]) ? 15'b000000111111111 : 15'b000000111111111;
												assign node4805 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node4808 = (inp[8]) ? node4810 : 15'b000000001111111;
												assign node4810 = (inp[0]) ? 15'b000000000011111 : node4811;
													assign node4811 = (inp[6]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node4815 = (inp[8]) ? node4827 : node4816;
											assign node4816 = (inp[1]) ? node4822 : node4817;
												assign node4817 = (inp[6]) ? 15'b000000000111111 : node4818;
													assign node4818 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node4822 = (inp[0]) ? 15'b000000000011111 : node4823;
													assign node4823 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4827 = (inp[7]) ? node4833 : node4828;
												assign node4828 = (inp[1]) ? node4830 : 15'b000000000111111;
													assign node4830 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4833 = (inp[10]) ? node4835 : 15'b000000000111111;
													assign node4835 = (inp[6]) ? 15'b000000000001111 : 15'b000000000001111;
									assign node4838 = (inp[6]) ? node4858 : node4839;
										assign node4839 = (inp[4]) ? node4851 : node4840;
											assign node4840 = (inp[8]) ? node4846 : node4841;
												assign node4841 = (inp[0]) ? node4843 : 15'b000000001111111;
													assign node4843 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4846 = (inp[10]) ? 15'b000000000111111 : node4847;
													assign node4847 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4851 = (inp[10]) ? node4855 : node4852;
												assign node4852 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4855 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4858 = (inp[7]) ? node4868 : node4859;
											assign node4859 = (inp[0]) ? node4861 : 15'b000000000111111;
												assign node4861 = (inp[4]) ? node4865 : node4862;
													assign node4862 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4865 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4868 = (inp[4]) ? node4874 : node4869;
												assign node4869 = (inp[1]) ? 15'b000000000001111 : node4870;
													assign node4870 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node4874 = (inp[0]) ? node4876 : 15'b000000000001111;
													assign node4876 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node4879 = (inp[1]) ? node5041 : node4880;
							assign node4880 = (inp[8]) ? node4952 : node4881;
								assign node4881 = (inp[10]) ? node4917 : node4882;
									assign node4882 = (inp[6]) ? node4898 : node4883;
										assign node4883 = (inp[7]) ? node4891 : node4884;
											assign node4884 = (inp[0]) ? 15'b000000011111111 : node4885;
												assign node4885 = (inp[5]) ? 15'b000000111111111 : node4886;
													assign node4886 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4891 = (inp[13]) ? node4893 : 15'b000000011111111;
												assign node4893 = (inp[9]) ? node4895 : 15'b000000011111111;
													assign node4895 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node4898 = (inp[0]) ? node4908 : node4899;
											assign node4899 = (inp[9]) ? node4901 : 15'b000000011111111;
												assign node4901 = (inp[4]) ? node4905 : node4902;
													assign node4902 = (inp[5]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node4905 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4908 = (inp[5]) ? node4910 : 15'b000000001111111;
												assign node4910 = (inp[13]) ? node4914 : node4911;
													assign node4911 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4914 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4917 = (inp[7]) ? node4935 : node4918;
										assign node4918 = (inp[9]) ? node4926 : node4919;
											assign node4919 = (inp[0]) ? node4923 : node4920;
												assign node4920 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4923 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node4926 = (inp[4]) ? node4928 : 15'b000000001111111;
												assign node4928 = (inp[5]) ? node4932 : node4929;
													assign node4929 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4932 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4935 = (inp[13]) ? node4943 : node4936;
											assign node4936 = (inp[5]) ? 15'b000000000111111 : node4937;
												assign node4937 = (inp[4]) ? node4939 : 15'b000000011111111;
													assign node4939 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4943 = (inp[9]) ? node4945 : 15'b000000000111111;
												assign node4945 = (inp[0]) ? node4949 : node4946;
													assign node4946 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node4949 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node4952 = (inp[4]) ? node4998 : node4953;
									assign node4953 = (inp[9]) ? node4973 : node4954;
										assign node4954 = (inp[0]) ? node4960 : node4955;
											assign node4955 = (inp[6]) ? node4957 : 15'b000000011111111;
												assign node4957 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4960 = (inp[5]) ? node4968 : node4961;
												assign node4961 = (inp[7]) ? node4965 : node4962;
													assign node4962 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4965 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4968 = (inp[10]) ? 15'b000000000111111 : node4969;
													assign node4969 = (inp[6]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node4973 = (inp[0]) ? node4987 : node4974;
											assign node4974 = (inp[6]) ? node4980 : node4975;
												assign node4975 = (inp[13]) ? node4977 : 15'b000000001111111;
													assign node4977 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4980 = (inp[13]) ? node4984 : node4981;
													assign node4981 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4984 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4987 = (inp[6]) ? node4993 : node4988;
												assign node4988 = (inp[5]) ? node4990 : 15'b000000000111111;
													assign node4990 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4993 = (inp[7]) ? node4995 : 15'b000000000011111;
													assign node4995 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node4998 = (inp[7]) ? node5016 : node4999;
										assign node4999 = (inp[0]) ? node5011 : node5000;
											assign node5000 = (inp[13]) ? node5006 : node5001;
												assign node5001 = (inp[5]) ? node5003 : 15'b000000001111111;
													assign node5003 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5006 = (inp[5]) ? 15'b000000000011111 : node5007;
													assign node5007 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5011 = (inp[9]) ? 15'b000000000011111 : node5012;
												assign node5012 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5016 = (inp[13]) ? node5032 : node5017;
											assign node5017 = (inp[10]) ? node5025 : node5018;
												assign node5018 = (inp[9]) ? node5022 : node5019;
													assign node5019 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node5022 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5025 = (inp[9]) ? node5029 : node5026;
													assign node5026 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5029 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5032 = (inp[6]) ? node5036 : node5033;
												assign node5033 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5036 = (inp[9]) ? node5038 : 15'b000000000001111;
													assign node5038 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node5041 = (inp[4]) ? node5127 : node5042;
								assign node5042 = (inp[5]) ? node5084 : node5043;
									assign node5043 = (inp[9]) ? node5065 : node5044;
										assign node5044 = (inp[13]) ? node5054 : node5045;
											assign node5045 = (inp[7]) ? node5051 : node5046;
												assign node5046 = (inp[6]) ? 15'b000000011111111 : node5047;
													assign node5047 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5051 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5054 = (inp[6]) ? node5060 : node5055;
												assign node5055 = (inp[0]) ? node5057 : 15'b000000001111111;
													assign node5057 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5060 = (inp[8]) ? 15'b000000000111111 : node5061;
													assign node5061 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5065 = (inp[8]) ? node5073 : node5066;
											assign node5066 = (inp[0]) ? 15'b000000000111111 : node5067;
												assign node5067 = (inp[10]) ? 15'b000000001111111 : node5068;
													assign node5068 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node5073 = (inp[0]) ? node5079 : node5074;
												assign node5074 = (inp[10]) ? node5076 : 15'b000000000111111;
													assign node5076 = (inp[7]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node5079 = (inp[7]) ? 15'b000000000011111 : node5080;
													assign node5080 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node5084 = (inp[9]) ? node5110 : node5085;
										assign node5085 = (inp[10]) ? node5097 : node5086;
											assign node5086 = (inp[13]) ? node5090 : node5087;
												assign node5087 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5090 = (inp[8]) ? node5094 : node5091;
													assign node5091 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5094 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5097 = (inp[13]) ? node5103 : node5098;
												assign node5098 = (inp[8]) ? node5100 : 15'b000000000111111;
													assign node5100 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node5103 = (inp[7]) ? node5107 : node5104;
													assign node5104 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node5107 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5110 = (inp[6]) ? node5122 : node5111;
											assign node5111 = (inp[7]) ? node5117 : node5112;
												assign node5112 = (inp[13]) ? node5114 : 15'b000000000111111;
													assign node5114 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5117 = (inp[10]) ? node5119 : 15'b000000000011111;
													assign node5119 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5122 = (inp[8]) ? 15'b000000000001111 : node5123;
												assign node5123 = (inp[7]) ? 15'b000000000011111 : 15'b000000000001111;
								assign node5127 = (inp[8]) ? node5177 : node5128;
									assign node5128 = (inp[6]) ? node5150 : node5129;
										assign node5129 = (inp[10]) ? node5137 : node5130;
											assign node5130 = (inp[7]) ? 15'b000000000011111 : node5131;
												assign node5131 = (inp[0]) ? 15'b000000001111111 : node5132;
													assign node5132 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node5137 = (inp[13]) ? node5145 : node5138;
												assign node5138 = (inp[0]) ? node5142 : node5139;
													assign node5139 = (inp[7]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node5142 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5145 = (inp[7]) ? node5147 : 15'b000000000011111;
													assign node5147 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5150 = (inp[10]) ? node5164 : node5151;
											assign node5151 = (inp[5]) ? node5157 : node5152;
												assign node5152 = (inp[0]) ? 15'b000000000011111 : node5153;
													assign node5153 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5157 = (inp[9]) ? node5161 : node5158;
													assign node5158 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5161 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5164 = (inp[13]) ? node5170 : node5165;
												assign node5165 = (inp[5]) ? node5167 : 15'b000000000011111;
													assign node5167 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node5170 = (inp[5]) ? node5174 : node5171;
													assign node5171 = (inp[0]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node5174 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node5177 = (inp[13]) ? node5197 : node5178;
										assign node5178 = (inp[7]) ? node5188 : node5179;
											assign node5179 = (inp[9]) ? node5185 : node5180;
												assign node5180 = (inp[6]) ? node5182 : 15'b000000001111111;
													assign node5182 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5185 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node5188 = (inp[6]) ? node5190 : 15'b000000000011111;
												assign node5190 = (inp[0]) ? node5194 : node5191;
													assign node5191 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node5194 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node5197 = (inp[0]) ? node5203 : node5198;
											assign node5198 = (inp[10]) ? 15'b000000000001111 : node5199;
												assign node5199 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5203 = (inp[10]) ? node5209 : node5204;
												assign node5204 = (inp[6]) ? 15'b000000000001111 : node5205;
													assign node5205 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node5209 = (inp[6]) ? 15'b000000000000011 : node5210;
													assign node5210 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
		assign node5214 = (inp[3]) ? node7892 : node5215;
			assign node5215 = (inp[5]) ? node6567 : node5216;
				assign node5216 = (inp[4]) ? node5906 : node5217;
					assign node5217 = (inp[9]) ? node5541 : node5218;
						assign node5218 = (inp[12]) ? node5378 : node5219;
							assign node5219 = (inp[13]) ? node5303 : node5220;
								assign node5220 = (inp[1]) ? node5262 : node5221;
									assign node5221 = (inp[14]) ? node5245 : node5222;
										assign node5222 = (inp[2]) ? node5232 : node5223;
											assign node5223 = (inp[10]) ? 15'b000111111111111 : node5224;
												assign node5224 = (inp[7]) ? node5228 : node5225;
													assign node5225 = (inp[6]) ? 15'b001111111111111 : 15'b011111111111111;
													assign node5228 = (inp[6]) ? 15'b000111111111111 : 15'b001111111111111;
											assign node5232 = (inp[10]) ? node5238 : node5233;
												assign node5233 = (inp[7]) ? 15'b000011111111111 : node5234;
													assign node5234 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node5238 = (inp[6]) ? node5242 : node5239;
													assign node5239 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5242 = (inp[8]) ? 15'b000000111111111 : 15'b000000111111111;
										assign node5245 = (inp[7]) ? node5255 : node5246;
											assign node5246 = (inp[6]) ? node5248 : 15'b000011111111111;
												assign node5248 = (inp[2]) ? node5252 : node5249;
													assign node5249 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5252 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5255 = (inp[2]) ? node5257 : 15'b000001111111111;
												assign node5257 = (inp[8]) ? node5259 : 15'b000001111111111;
													assign node5259 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node5262 = (inp[14]) ? node5286 : node5263;
										assign node5263 = (inp[2]) ? node5273 : node5264;
											assign node5264 = (inp[0]) ? node5268 : node5265;
												assign node5265 = (inp[10]) ? 15'b000011111111111 : 15'b001111111111111;
												assign node5268 = (inp[10]) ? 15'b000001111111111 : node5269;
													assign node5269 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node5273 = (inp[6]) ? node5279 : node5274;
												assign node5274 = (inp[10]) ? node5276 : 15'b000001111111111;
													assign node5276 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5279 = (inp[7]) ? node5283 : node5280;
													assign node5280 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5283 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5286 = (inp[0]) ? node5294 : node5287;
											assign node5287 = (inp[7]) ? 15'b000000111111111 : node5288;
												assign node5288 = (inp[10]) ? node5290 : 15'b000001111111111;
													assign node5290 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5294 = (inp[8]) ? 15'b000000011111111 : node5295;
												assign node5295 = (inp[2]) ? node5299 : node5296;
													assign node5296 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5299 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
								assign node5303 = (inp[10]) ? node5345 : node5304;
									assign node5304 = (inp[7]) ? node5320 : node5305;
										assign node5305 = (inp[2]) ? node5313 : node5306;
											assign node5306 = (inp[14]) ? node5308 : 15'b000111111111111;
												assign node5308 = (inp[6]) ? 15'b000001111111111 : node5309;
													assign node5309 = (inp[1]) ? 15'b000001111111111 : 15'b000001111111111;
											assign node5313 = (inp[14]) ? 15'b000001111111111 : node5314;
												assign node5314 = (inp[1]) ? node5316 : 15'b000001111111111;
													assign node5316 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node5320 = (inp[2]) ? node5334 : node5321;
											assign node5321 = (inp[1]) ? node5327 : node5322;
												assign node5322 = (inp[8]) ? 15'b000001111111111 : node5323;
													assign node5323 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5327 = (inp[0]) ? node5331 : node5328;
													assign node5328 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5331 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5334 = (inp[14]) ? node5340 : node5335;
												assign node5335 = (inp[6]) ? node5337 : 15'b000000111111111;
													assign node5337 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5340 = (inp[0]) ? 15'b000000011111111 : node5341;
													assign node5341 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
									assign node5345 = (inp[8]) ? node5361 : node5346;
										assign node5346 = (inp[14]) ? node5356 : node5347;
											assign node5347 = (inp[2]) ? node5353 : node5348;
												assign node5348 = (inp[7]) ? node5350 : 15'b000011111111111;
													assign node5350 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5353 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5356 = (inp[6]) ? node5358 : 15'b000000111111111;
												assign node5358 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5361 = (inp[6]) ? node5371 : node5362;
											assign node5362 = (inp[14]) ? node5368 : node5363;
												assign node5363 = (inp[2]) ? node5365 : 15'b000000111111111;
													assign node5365 = (inp[7]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node5368 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5371 = (inp[2]) ? node5373 : 15'b000000011111111;
												assign node5373 = (inp[1]) ? 15'b000000000111111 : node5374;
													assign node5374 = (inp[0]) ? 15'b000000011111111 : 15'b000000001111111;
							assign node5378 = (inp[0]) ? node5470 : node5379;
								assign node5379 = (inp[1]) ? node5431 : node5380;
									assign node5380 = (inp[7]) ? node5404 : node5381;
										assign node5381 = (inp[14]) ? node5395 : node5382;
											assign node5382 = (inp[6]) ? node5388 : node5383;
												assign node5383 = (inp[13]) ? node5385 : 15'b000111111111111;
													assign node5385 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node5388 = (inp[10]) ? node5392 : node5389;
													assign node5389 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5392 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5395 = (inp[8]) ? 15'b000000111111111 : node5396;
												assign node5396 = (inp[10]) ? node5400 : node5397;
													assign node5397 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5400 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node5404 = (inp[6]) ? node5418 : node5405;
											assign node5405 = (inp[2]) ? node5411 : node5406;
												assign node5406 = (inp[10]) ? 15'b000001111111111 : node5407;
													assign node5407 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5411 = (inp[10]) ? node5415 : node5412;
													assign node5412 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5415 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node5418 = (inp[13]) ? node5426 : node5419;
												assign node5419 = (inp[2]) ? node5423 : node5420;
													assign node5420 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node5423 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5426 = (inp[14]) ? 15'b000000011111111 : node5427;
													assign node5427 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node5431 = (inp[7]) ? node5453 : node5432;
										assign node5432 = (inp[8]) ? node5440 : node5433;
											assign node5433 = (inp[10]) ? node5435 : 15'b000011111111111;
												assign node5435 = (inp[14]) ? node5437 : 15'b000001111111111;
													assign node5437 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5440 = (inp[6]) ? node5448 : node5441;
												assign node5441 = (inp[13]) ? node5445 : node5442;
													assign node5442 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node5445 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5448 = (inp[10]) ? node5450 : 15'b000000011111111;
													assign node5450 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5453 = (inp[2]) ? node5465 : node5454;
											assign node5454 = (inp[10]) ? node5458 : node5455;
												assign node5455 = (inp[13]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node5458 = (inp[8]) ? node5462 : node5459;
													assign node5459 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5462 = (inp[14]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node5465 = (inp[10]) ? node5467 : 15'b000000011111111;
												assign node5467 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5470 = (inp[1]) ? node5508 : node5471;
									assign node5471 = (inp[14]) ? node5487 : node5472;
										assign node5472 = (inp[7]) ? node5480 : node5473;
											assign node5473 = (inp[8]) ? 15'b000000111111111 : node5474;
												assign node5474 = (inp[10]) ? node5476 : 15'b000001111111111;
													assign node5476 = (inp[6]) ? 15'b000000111111111 : 15'b000000111111111;
											assign node5480 = (inp[6]) ? 15'b000000011111111 : node5481;
												assign node5481 = (inp[2]) ? 15'b000000011111111 : node5482;
													assign node5482 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node5487 = (inp[13]) ? node5497 : node5488;
											assign node5488 = (inp[6]) ? node5492 : node5489;
												assign node5489 = (inp[10]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node5492 = (inp[2]) ? 15'b000000011111111 : node5493;
													assign node5493 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5497 = (inp[10]) ? node5503 : node5498;
												assign node5498 = (inp[2]) ? 15'b000000011111111 : node5499;
													assign node5499 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5503 = (inp[2]) ? 15'b000000000111111 : node5504;
													assign node5504 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node5508 = (inp[13]) ? node5526 : node5509;
										assign node5509 = (inp[8]) ? node5517 : node5510;
											assign node5510 = (inp[7]) ? node5512 : 15'b000000111111111;
												assign node5512 = (inp[2]) ? 15'b000000111111111 : node5513;
													assign node5513 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5517 = (inp[10]) ? 15'b000000001111111 : node5518;
												assign node5518 = (inp[14]) ? node5522 : node5519;
													assign node5519 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5522 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5526 = (inp[7]) ? node5530 : node5527;
											assign node5527 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node5530 = (inp[2]) ? node5536 : node5531;
												assign node5531 = (inp[8]) ? node5533 : 15'b000000111111111;
													assign node5533 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5536 = (inp[10]) ? node5538 : 15'b000000000111111;
													assign node5538 = (inp[14]) ? 15'b000000000011111 : 15'b000000000011111;
						assign node5541 = (inp[6]) ? node5723 : node5542;
							assign node5542 = (inp[8]) ? node5642 : node5543;
								assign node5543 = (inp[7]) ? node5591 : node5544;
									assign node5544 = (inp[10]) ? node5570 : node5545;
										assign node5545 = (inp[12]) ? node5559 : node5546;
											assign node5546 = (inp[2]) ? node5554 : node5547;
												assign node5547 = (inp[1]) ? node5551 : node5548;
													assign node5548 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node5551 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5554 = (inp[1]) ? 15'b000001111111111 : node5555;
													assign node5555 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node5559 = (inp[1]) ? node5563 : node5560;
												assign node5560 = (inp[0]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node5563 = (inp[2]) ? node5567 : node5564;
													assign node5564 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5567 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5570 = (inp[14]) ? node5586 : node5571;
											assign node5571 = (inp[13]) ? node5579 : node5572;
												assign node5572 = (inp[1]) ? node5576 : node5573;
													assign node5573 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5576 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5579 = (inp[12]) ? node5583 : node5580;
													assign node5580 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5583 = (inp[1]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node5586 = (inp[13]) ? node5588 : 15'b000000011111111;
												assign node5588 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node5591 = (inp[0]) ? node5619 : node5592;
										assign node5592 = (inp[12]) ? node5606 : node5593;
											assign node5593 = (inp[1]) ? node5601 : node5594;
												assign node5594 = (inp[10]) ? node5598 : node5595;
													assign node5595 = (inp[2]) ? 15'b000011111111111 : 15'b000001111111111;
													assign node5598 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5601 = (inp[10]) ? 15'b000000111111111 : node5602;
													assign node5602 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5606 = (inp[13]) ? node5614 : node5607;
												assign node5607 = (inp[2]) ? node5611 : node5608;
													assign node5608 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5611 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5614 = (inp[10]) ? 15'b000000011111111 : node5615;
													assign node5615 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5619 = (inp[13]) ? node5633 : node5620;
											assign node5620 = (inp[1]) ? node5628 : node5621;
												assign node5621 = (inp[2]) ? node5625 : node5622;
													assign node5622 = (inp[14]) ? 15'b000000111111111 : 15'b000000111111111;
													assign node5625 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5628 = (inp[14]) ? node5630 : 15'b000000001111111;
													assign node5630 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node5633 = (inp[14]) ? node5635 : 15'b000000011111111;
												assign node5635 = (inp[1]) ? node5639 : node5636;
													assign node5636 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5639 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5642 = (inp[10]) ? node5690 : node5643;
									assign node5643 = (inp[0]) ? node5665 : node5644;
										assign node5644 = (inp[7]) ? node5658 : node5645;
											assign node5645 = (inp[12]) ? node5653 : node5646;
												assign node5646 = (inp[13]) ? node5650 : node5647;
													assign node5647 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5650 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5653 = (inp[1]) ? 15'b000000011111111 : node5654;
													assign node5654 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5658 = (inp[2]) ? node5660 : 15'b000000111111111;
												assign node5660 = (inp[1]) ? 15'b000000011111111 : node5661;
													assign node5661 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5665 = (inp[14]) ? node5679 : node5666;
											assign node5666 = (inp[13]) ? node5672 : node5667;
												assign node5667 = (inp[1]) ? node5669 : 15'b000011111111111;
													assign node5669 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5672 = (inp[12]) ? node5676 : node5673;
													assign node5673 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5676 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5679 = (inp[12]) ? node5685 : node5680;
												assign node5680 = (inp[7]) ? node5682 : 15'b000000011111111;
													assign node5682 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5685 = (inp[7]) ? 15'b000000001111111 : node5686;
													assign node5686 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5690 = (inp[2]) ? node5704 : node5691;
										assign node5691 = (inp[12]) ? node5699 : node5692;
											assign node5692 = (inp[1]) ? 15'b000000011111111 : node5693;
												assign node5693 = (inp[14]) ? node5695 : 15'b000000111111111;
													assign node5695 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node5699 = (inp[13]) ? 15'b000000001111111 : node5700;
												assign node5700 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5704 = (inp[12]) ? node5718 : node5705;
											assign node5705 = (inp[13]) ? node5711 : node5706;
												assign node5706 = (inp[7]) ? node5708 : 15'b000000111111111;
													assign node5708 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5711 = (inp[7]) ? node5715 : node5712;
													assign node5712 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5715 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node5718 = (inp[0]) ? node5720 : 15'b000000000111111;
												assign node5720 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
							assign node5723 = (inp[7]) ? node5813 : node5724;
								assign node5724 = (inp[13]) ? node5772 : node5725;
									assign node5725 = (inp[0]) ? node5751 : node5726;
										assign node5726 = (inp[8]) ? node5738 : node5727;
											assign node5727 = (inp[1]) ? node5733 : node5728;
												assign node5728 = (inp[12]) ? node5730 : 15'b000001111111111;
													assign node5730 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5733 = (inp[2]) ? 15'b000000011111111 : node5734;
													assign node5734 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5738 = (inp[12]) ? node5746 : node5739;
												assign node5739 = (inp[2]) ? node5743 : node5740;
													assign node5740 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5743 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5746 = (inp[14]) ? node5748 : 15'b000000111111111;
													assign node5748 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node5751 = (inp[10]) ? node5763 : node5752;
											assign node5752 = (inp[1]) ? node5758 : node5753;
												assign node5753 = (inp[2]) ? node5755 : 15'b000000111111111;
													assign node5755 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5758 = (inp[8]) ? 15'b000000001111111 : node5759;
													assign node5759 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5763 = (inp[12]) ? node5769 : node5764;
												assign node5764 = (inp[2]) ? node5766 : 15'b000000111111111;
													assign node5766 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5769 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5772 = (inp[1]) ? node5790 : node5773;
										assign node5773 = (inp[2]) ? node5781 : node5774;
											assign node5774 = (inp[8]) ? 15'b000000011111111 : node5775;
												assign node5775 = (inp[0]) ? node5777 : 15'b000000111111111;
													assign node5777 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5781 = (inp[12]) ? node5787 : node5782;
												assign node5782 = (inp[14]) ? node5784 : 15'b000000011111111;
													assign node5784 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5787 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5790 = (inp[10]) ? node5802 : node5791;
											assign node5791 = (inp[12]) ? node5795 : node5792;
												assign node5792 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5795 = (inp[14]) ? node5799 : node5796;
													assign node5796 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5799 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5802 = (inp[14]) ? node5810 : node5803;
												assign node5803 = (inp[12]) ? node5807 : node5804;
													assign node5804 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5807 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node5810 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5813 = (inp[2]) ? node5855 : node5814;
									assign node5814 = (inp[0]) ? node5836 : node5815;
										assign node5815 = (inp[10]) ? node5825 : node5816;
											assign node5816 = (inp[12]) ? node5820 : node5817;
												assign node5817 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5820 = (inp[1]) ? 15'b000000011111111 : node5821;
													assign node5821 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5825 = (inp[12]) ? node5831 : node5826;
												assign node5826 = (inp[13]) ? node5828 : 15'b000000011111111;
													assign node5828 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5831 = (inp[1]) ? node5833 : 15'b000000001111111;
													assign node5833 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node5836 = (inp[8]) ? node5844 : node5837;
											assign node5837 = (inp[12]) ? node5839 : 15'b000000011111111;
												assign node5839 = (inp[13]) ? 15'b000000001111111 : node5840;
													assign node5840 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5844 = (inp[13]) ? node5850 : node5845;
												assign node5845 = (inp[14]) ? 15'b000000001111111 : node5846;
													assign node5846 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5850 = (inp[10]) ? 15'b000000000111111 : node5851;
													assign node5851 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5855 = (inp[8]) ? node5881 : node5856;
										assign node5856 = (inp[0]) ? node5868 : node5857;
											assign node5857 = (inp[12]) ? node5863 : node5858;
												assign node5858 = (inp[1]) ? 15'b000000001111111 : node5859;
													assign node5859 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5863 = (inp[13]) ? node5865 : 15'b000000001111111;
													assign node5865 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node5868 = (inp[14]) ? node5874 : node5869;
												assign node5869 = (inp[10]) ? node5871 : 15'b000000001111111;
													assign node5871 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5874 = (inp[12]) ? node5878 : node5875;
													assign node5875 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5878 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5881 = (inp[14]) ? node5893 : node5882;
											assign node5882 = (inp[1]) ? node5888 : node5883;
												assign node5883 = (inp[12]) ? node5885 : 15'b000000001111111;
													assign node5885 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5888 = (inp[13]) ? node5890 : 15'b000000000111111;
													assign node5890 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5893 = (inp[12]) ? node5901 : node5894;
												assign node5894 = (inp[10]) ? node5898 : node5895;
													assign node5895 = (inp[13]) ? 15'b000000001111111 : 15'b000000000111111;
													assign node5898 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5901 = (inp[1]) ? 15'b000000000001111 : node5902;
													assign node5902 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node5906 = (inp[2]) ? node6222 : node5907;
						assign node5907 = (inp[7]) ? node6069 : node5908;
							assign node5908 = (inp[14]) ? node5994 : node5909;
								assign node5909 = (inp[10]) ? node5947 : node5910;
									assign node5910 = (inp[6]) ? node5930 : node5911;
										assign node5911 = (inp[13]) ? node5921 : node5912;
											assign node5912 = (inp[0]) ? 15'b000000111111111 : node5913;
												assign node5913 = (inp[9]) ? node5917 : node5914;
													assign node5914 = (inp[12]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node5917 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node5921 = (inp[12]) ? node5927 : node5922;
												assign node5922 = (inp[8]) ? 15'b000000111111111 : node5923;
													assign node5923 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5927 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node5930 = (inp[9]) ? node5940 : node5931;
											assign node5931 = (inp[12]) ? node5935 : node5932;
												assign node5932 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5935 = (inp[8]) ? node5937 : 15'b000000111111111;
													assign node5937 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5940 = (inp[12]) ? 15'b000000000111111 : node5941;
												assign node5941 = (inp[13]) ? node5943 : 15'b000000111111111;
													assign node5943 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node5947 = (inp[8]) ? node5967 : node5948;
										assign node5948 = (inp[12]) ? node5954 : node5949;
											assign node5949 = (inp[0]) ? 15'b000000111111111 : node5950;
												assign node5950 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5954 = (inp[9]) ? node5962 : node5955;
												assign node5955 = (inp[6]) ? node5959 : node5956;
													assign node5956 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5959 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5962 = (inp[6]) ? 15'b000000011111111 : node5963;
													assign node5963 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
										assign node5967 = (inp[0]) ? node5981 : node5968;
											assign node5968 = (inp[6]) ? node5976 : node5969;
												assign node5969 = (inp[1]) ? node5973 : node5970;
													assign node5970 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5973 = (inp[9]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node5976 = (inp[1]) ? node5978 : 15'b000000011111111;
													assign node5978 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5981 = (inp[9]) ? node5987 : node5982;
												assign node5982 = (inp[1]) ? node5984 : 15'b000000011111111;
													assign node5984 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5987 = (inp[1]) ? node5991 : node5988;
													assign node5988 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5991 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5994 = (inp[0]) ? node6034 : node5995;
									assign node5995 = (inp[8]) ? node6017 : node5996;
										assign node5996 = (inp[12]) ? node6006 : node5997;
											assign node5997 = (inp[9]) ? node6001 : node5998;
												assign node5998 = (inp[10]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node6001 = (inp[6]) ? 15'b000000111111111 : node6002;
													assign node6002 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6006 = (inp[1]) ? node6014 : node6007;
												assign node6007 = (inp[10]) ? node6011 : node6008;
													assign node6008 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6011 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6014 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6017 = (inp[6]) ? node6029 : node6018;
											assign node6018 = (inp[12]) ? node6024 : node6019;
												assign node6019 = (inp[1]) ? node6021 : 15'b000000111111111;
													assign node6021 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6024 = (inp[1]) ? node6026 : 15'b000000001111111;
													assign node6026 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node6029 = (inp[13]) ? 15'b000000001111111 : node6030;
												assign node6030 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6034 = (inp[12]) ? node6054 : node6035;
										assign node6035 = (inp[10]) ? node6043 : node6036;
											assign node6036 = (inp[13]) ? 15'b000000011111111 : node6037;
												assign node6037 = (inp[6]) ? node6039 : 15'b000000111111111;
													assign node6039 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6043 = (inp[8]) ? node6051 : node6044;
												assign node6044 = (inp[9]) ? node6048 : node6045;
													assign node6045 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6048 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6051 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6054 = (inp[9]) ? node6064 : node6055;
											assign node6055 = (inp[10]) ? node6057 : 15'b000000011111111;
												assign node6057 = (inp[1]) ? node6061 : node6058;
													assign node6058 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6061 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6064 = (inp[13]) ? node6066 : 15'b000000001111111;
												assign node6066 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
							assign node6069 = (inp[6]) ? node6139 : node6070;
								assign node6070 = (inp[13]) ? node6108 : node6071;
									assign node6071 = (inp[0]) ? node6091 : node6072;
										assign node6072 = (inp[1]) ? node6086 : node6073;
											assign node6073 = (inp[14]) ? node6081 : node6074;
												assign node6074 = (inp[10]) ? node6078 : node6075;
													assign node6075 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6078 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6081 = (inp[10]) ? 15'b000000111111111 : node6082;
													assign node6082 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6086 = (inp[12]) ? 15'b000000011111111 : node6087;
												assign node6087 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6091 = (inp[10]) ? node6097 : node6092;
											assign node6092 = (inp[8]) ? node6094 : 15'b000000111111111;
												assign node6094 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node6097 = (inp[9]) ? node6103 : node6098;
												assign node6098 = (inp[14]) ? 15'b000000011111111 : node6099;
													assign node6099 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6103 = (inp[12]) ? 15'b000000001111111 : node6104;
													assign node6104 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6108 = (inp[9]) ? node6124 : node6109;
										assign node6109 = (inp[12]) ? node6115 : node6110;
											assign node6110 = (inp[1]) ? 15'b000000011111111 : node6111;
												assign node6111 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6115 = (inp[8]) ? node6119 : node6116;
												assign node6116 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node6119 = (inp[14]) ? 15'b000000001111111 : node6120;
													assign node6120 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6124 = (inp[8]) ? node6132 : node6125;
											assign node6125 = (inp[1]) ? 15'b000000001111111 : node6126;
												assign node6126 = (inp[0]) ? node6128 : 15'b000000011111111;
													assign node6128 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6132 = (inp[12]) ? 15'b000000000111111 : node6133;
												assign node6133 = (inp[1]) ? node6135 : 15'b000000001111111;
													assign node6135 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node6139 = (inp[10]) ? node6185 : node6140;
									assign node6140 = (inp[9]) ? node6160 : node6141;
										assign node6141 = (inp[0]) ? node6151 : node6142;
											assign node6142 = (inp[1]) ? node6146 : node6143;
												assign node6143 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node6146 = (inp[8]) ? node6148 : 15'b000000111111111;
													assign node6148 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6151 = (inp[14]) ? 15'b000000001111111 : node6152;
												assign node6152 = (inp[12]) ? node6156 : node6153;
													assign node6153 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6156 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6160 = (inp[14]) ? node6174 : node6161;
											assign node6161 = (inp[12]) ? node6167 : node6162;
												assign node6162 = (inp[13]) ? node6164 : 15'b000000011111111;
													assign node6164 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6167 = (inp[8]) ? node6171 : node6168;
													assign node6168 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node6171 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6174 = (inp[0]) ? node6180 : node6175;
												assign node6175 = (inp[13]) ? 15'b000000001111111 : node6176;
													assign node6176 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node6180 = (inp[13]) ? node6182 : 15'b000000001111111;
													assign node6182 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node6185 = (inp[12]) ? node6207 : node6186;
										assign node6186 = (inp[8]) ? node6194 : node6187;
											assign node6187 = (inp[13]) ? node6189 : 15'b000000011111111;
												assign node6189 = (inp[1]) ? 15'b000000001111111 : node6190;
													assign node6190 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6194 = (inp[9]) ? node6202 : node6195;
												assign node6195 = (inp[14]) ? node6199 : node6196;
													assign node6196 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6199 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6202 = (inp[13]) ? 15'b000000000111111 : node6203;
													assign node6203 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6207 = (inp[13]) ? node6215 : node6208;
											assign node6208 = (inp[14]) ? 15'b000000000111111 : node6209;
												assign node6209 = (inp[9]) ? node6211 : 15'b000000001111111;
													assign node6211 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6215 = (inp[1]) ? 15'b000000000111111 : node6216;
												assign node6216 = (inp[0]) ? node6218 : 15'b000000000011111;
													assign node6218 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node6222 = (inp[13]) ? node6398 : node6223;
							assign node6223 = (inp[12]) ? node6317 : node6224;
								assign node6224 = (inp[6]) ? node6272 : node6225;
									assign node6225 = (inp[0]) ? node6249 : node6226;
										assign node6226 = (inp[8]) ? node6238 : node6227;
											assign node6227 = (inp[14]) ? node6233 : node6228;
												assign node6228 = (inp[10]) ? 15'b000001111111111 : node6229;
													assign node6229 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node6233 = (inp[10]) ? 15'b000000111111111 : node6234;
													assign node6234 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6238 = (inp[1]) ? node6244 : node6239;
												assign node6239 = (inp[9]) ? 15'b000000111111111 : node6240;
													assign node6240 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6244 = (inp[10]) ? 15'b000000011111111 : node6245;
													assign node6245 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6249 = (inp[7]) ? node6261 : node6250;
											assign node6250 = (inp[1]) ? node6256 : node6251;
												assign node6251 = (inp[10]) ? 15'b000000111111111 : node6252;
													assign node6252 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6256 = (inp[10]) ? node6258 : 15'b000000111111111;
													assign node6258 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6261 = (inp[14]) ? node6267 : node6262;
												assign node6262 = (inp[9]) ? 15'b000000011111111 : node6263;
													assign node6263 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node6267 = (inp[1]) ? 15'b000000001111111 : node6268;
													assign node6268 = (inp[9]) ? 15'b000000001111111 : 15'b000000001111111;
									assign node6272 = (inp[10]) ? node6296 : node6273;
										assign node6273 = (inp[9]) ? node6281 : node6274;
											assign node6274 = (inp[0]) ? node6276 : 15'b000000111111111;
												assign node6276 = (inp[7]) ? 15'b000000011111111 : node6277;
													assign node6277 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6281 = (inp[1]) ? node6289 : node6282;
												assign node6282 = (inp[7]) ? node6286 : node6283;
													assign node6283 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6286 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6289 = (inp[0]) ? node6293 : node6290;
													assign node6290 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6293 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
										assign node6296 = (inp[9]) ? node6308 : node6297;
											assign node6297 = (inp[14]) ? node6303 : node6298;
												assign node6298 = (inp[8]) ? node6300 : 15'b000000011111111;
													assign node6300 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6303 = (inp[1]) ? node6305 : 15'b000000011111111;
													assign node6305 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6308 = (inp[7]) ? 15'b000000000111111 : node6309;
												assign node6309 = (inp[8]) ? node6313 : node6310;
													assign node6310 = (inp[14]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node6313 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node6317 = (inp[14]) ? node6361 : node6318;
									assign node6318 = (inp[9]) ? node6342 : node6319;
										assign node6319 = (inp[7]) ? node6333 : node6320;
											assign node6320 = (inp[6]) ? node6328 : node6321;
												assign node6321 = (inp[10]) ? node6325 : node6322;
													assign node6322 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6325 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6328 = (inp[8]) ? 15'b000000011111111 : node6329;
													assign node6329 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6333 = (inp[0]) ? node6337 : node6334;
												assign node6334 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node6337 = (inp[6]) ? 15'b000000001111111 : node6338;
													assign node6338 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6342 = (inp[0]) ? node6354 : node6343;
											assign node6343 = (inp[10]) ? node6349 : node6344;
												assign node6344 = (inp[6]) ? node6346 : 15'b000000111111111;
													assign node6346 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6349 = (inp[8]) ? 15'b000000000111111 : node6350;
													assign node6350 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6354 = (inp[1]) ? node6356 : 15'b000000001111111;
												assign node6356 = (inp[10]) ? 15'b000000000111111 : node6357;
													assign node6357 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node6361 = (inp[0]) ? node6381 : node6362;
										assign node6362 = (inp[8]) ? node6370 : node6363;
											assign node6363 = (inp[1]) ? 15'b000000000111111 : node6364;
												assign node6364 = (inp[6]) ? node6366 : 15'b000000111111111;
													assign node6366 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6370 = (inp[7]) ? node6374 : node6371;
												assign node6371 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6374 = (inp[6]) ? node6378 : node6375;
													assign node6375 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node6378 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6381 = (inp[7]) ? node6389 : node6382;
											assign node6382 = (inp[9]) ? 15'b000000000111111 : node6383;
												assign node6383 = (inp[1]) ? 15'b000000000111111 : node6384;
													assign node6384 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6389 = (inp[6]) ? 15'b000000000011111 : node6390;
												assign node6390 = (inp[9]) ? node6394 : node6391;
													assign node6391 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6394 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node6398 = (inp[1]) ? node6480 : node6399;
								assign node6399 = (inp[12]) ? node6439 : node6400;
									assign node6400 = (inp[14]) ? node6416 : node6401;
										assign node6401 = (inp[9]) ? node6407 : node6402;
											assign node6402 = (inp[10]) ? node6404 : 15'b000000111111111;
												assign node6404 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6407 = (inp[10]) ? node6413 : node6408;
												assign node6408 = (inp[7]) ? 15'b000000011111111 : node6409;
													assign node6409 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node6413 = (inp[6]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node6416 = (inp[6]) ? node6428 : node6417;
											assign node6417 = (inp[9]) ? node6423 : node6418;
												assign node6418 = (inp[0]) ? node6420 : 15'b000000011111111;
													assign node6420 = (inp[10]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node6423 = (inp[0]) ? 15'b000000001111111 : node6424;
													assign node6424 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6428 = (inp[0]) ? node6434 : node6429;
												assign node6429 = (inp[8]) ? 15'b000000001111111 : node6430;
													assign node6430 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6434 = (inp[10]) ? 15'b000000000111111 : node6435;
													assign node6435 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node6439 = (inp[6]) ? node6465 : node6440;
										assign node6440 = (inp[14]) ? node6454 : node6441;
											assign node6441 = (inp[10]) ? node6449 : node6442;
												assign node6442 = (inp[8]) ? node6446 : node6443;
													assign node6443 = (inp[7]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node6446 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6449 = (inp[7]) ? node6451 : 15'b000000011111111;
													assign node6451 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6454 = (inp[0]) ? node6460 : node6455;
												assign node6455 = (inp[7]) ? node6457 : 15'b000000001111111;
													assign node6457 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6460 = (inp[8]) ? node6462 : 15'b000000000111111;
													assign node6462 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6465 = (inp[0]) ? node6471 : node6466;
											assign node6466 = (inp[14]) ? 15'b000000000111111 : node6467;
												assign node6467 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6471 = (inp[10]) ? node6475 : node6472;
												assign node6472 = (inp[8]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node6475 = (inp[14]) ? 15'b000000000001111 : node6476;
													assign node6476 = (inp[7]) ? 15'b000000000001111 : 15'b000000000111111;
								assign node6480 = (inp[9]) ? node6524 : node6481;
									assign node6481 = (inp[14]) ? node6501 : node6482;
										assign node6482 = (inp[6]) ? node6490 : node6483;
											assign node6483 = (inp[7]) ? 15'b000000001111111 : node6484;
												assign node6484 = (inp[8]) ? 15'b000000011111111 : node6485;
													assign node6485 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node6490 = (inp[0]) ? node6496 : node6491;
												assign node6491 = (inp[8]) ? 15'b000000001111111 : node6492;
													assign node6492 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6496 = (inp[8]) ? node6498 : 15'b000000001111111;
													assign node6498 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6501 = (inp[0]) ? node6511 : node6502;
											assign node6502 = (inp[12]) ? node6506 : node6503;
												assign node6503 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6506 = (inp[6]) ? 15'b000000000111111 : node6507;
													assign node6507 = (inp[10]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node6511 = (inp[8]) ? node6517 : node6512;
												assign node6512 = (inp[6]) ? node6514 : 15'b000000000111111;
													assign node6514 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6517 = (inp[7]) ? node6521 : node6518;
													assign node6518 = (inp[6]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node6521 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node6524 = (inp[12]) ? node6540 : node6525;
										assign node6525 = (inp[8]) ? node6533 : node6526;
											assign node6526 = (inp[6]) ? node6528 : 15'b000000001111111;
												assign node6528 = (inp[0]) ? 15'b000000000011111 : node6529;
													assign node6529 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6533 = (inp[10]) ? node6535 : 15'b000000000111111;
												assign node6535 = (inp[0]) ? node6537 : 15'b000000000111111;
													assign node6537 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node6540 = (inp[8]) ? node6556 : node6541;
											assign node6541 = (inp[0]) ? node6549 : node6542;
												assign node6542 = (inp[6]) ? node6546 : node6543;
													assign node6543 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node6546 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6549 = (inp[10]) ? node6553 : node6550;
													assign node6550 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6553 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node6556 = (inp[14]) ? node6562 : node6557;
												assign node6557 = (inp[7]) ? node6559 : 15'b000000000011111;
													assign node6559 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node6562 = (inp[10]) ? 15'b000000000000111 : node6563;
													assign node6563 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node6567 = (inp[13]) ? node7245 : node6568;
					assign node6568 = (inp[9]) ? node6904 : node6569;
						assign node6569 = (inp[10]) ? node6755 : node6570;
							assign node6570 = (inp[14]) ? node6662 : node6571;
								assign node6571 = (inp[4]) ? node6619 : node6572;
									assign node6572 = (inp[1]) ? node6598 : node6573;
										assign node6573 = (inp[0]) ? node6587 : node6574;
											assign node6574 = (inp[6]) ? node6582 : node6575;
												assign node6575 = (inp[12]) ? node6579 : node6576;
													assign node6576 = (inp[7]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node6579 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node6582 = (inp[8]) ? 15'b000001111111111 : node6583;
													assign node6583 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node6587 = (inp[7]) ? node6595 : node6588;
												assign node6588 = (inp[6]) ? node6592 : node6589;
													assign node6589 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6592 = (inp[8]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node6595 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node6598 = (inp[7]) ? node6610 : node6599;
											assign node6599 = (inp[2]) ? node6605 : node6600;
												assign node6600 = (inp[12]) ? node6602 : 15'b000001111111111;
													assign node6602 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node6605 = (inp[6]) ? node6607 : 15'b000001111111111;
													assign node6607 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6610 = (inp[8]) ? node6612 : 15'b000000111111111;
												assign node6612 = (inp[12]) ? node6616 : node6613;
													assign node6613 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6616 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6619 = (inp[7]) ? node6639 : node6620;
										assign node6620 = (inp[6]) ? node6632 : node6621;
											assign node6621 = (inp[2]) ? node6627 : node6622;
												assign node6622 = (inp[0]) ? node6624 : 15'b000011111111111;
													assign node6624 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6627 = (inp[1]) ? 15'b000000011111111 : node6628;
													assign node6628 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6632 = (inp[12]) ? node6634 : 15'b000000111111111;
												assign node6634 = (inp[0]) ? 15'b000000011111111 : node6635;
													assign node6635 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6639 = (inp[12]) ? node6653 : node6640;
											assign node6640 = (inp[6]) ? node6648 : node6641;
												assign node6641 = (inp[0]) ? node6645 : node6642;
													assign node6642 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6645 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6648 = (inp[2]) ? 15'b000000001111111 : node6649;
													assign node6649 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6653 = (inp[1]) ? node6655 : 15'b000000011111111;
												assign node6655 = (inp[2]) ? node6659 : node6656;
													assign node6656 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6659 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6662 = (inp[0]) ? node6708 : node6663;
									assign node6663 = (inp[7]) ? node6689 : node6664;
										assign node6664 = (inp[4]) ? node6676 : node6665;
											assign node6665 = (inp[1]) ? node6669 : node6666;
												assign node6666 = (inp[6]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node6669 = (inp[6]) ? node6673 : node6670;
													assign node6670 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6673 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6676 = (inp[12]) ? node6682 : node6677;
												assign node6677 = (inp[2]) ? node6679 : 15'b000000111111111;
													assign node6679 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6682 = (inp[2]) ? node6686 : node6683;
													assign node6683 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6686 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6689 = (inp[2]) ? node6697 : node6690;
											assign node6690 = (inp[6]) ? node6692 : 15'b000000111111111;
												assign node6692 = (inp[12]) ? 15'b000000011111111 : node6693;
													assign node6693 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node6697 = (inp[8]) ? node6705 : node6698;
												assign node6698 = (inp[4]) ? node6702 : node6699;
													assign node6699 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node6702 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6705 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6708 = (inp[4]) ? node6734 : node6709;
										assign node6709 = (inp[2]) ? node6721 : node6710;
											assign node6710 = (inp[6]) ? node6716 : node6711;
												assign node6711 = (inp[8]) ? node6713 : 15'b000000111111111;
													assign node6713 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node6716 = (inp[1]) ? 15'b000000001111111 : node6717;
													assign node6717 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6721 = (inp[12]) ? node6729 : node6722;
												assign node6722 = (inp[8]) ? node6726 : node6723;
													assign node6723 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6726 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6729 = (inp[7]) ? 15'b000000001111111 : node6730;
													assign node6730 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node6734 = (inp[8]) ? node6744 : node6735;
											assign node6735 = (inp[1]) ? node6739 : node6736;
												assign node6736 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6739 = (inp[2]) ? node6741 : 15'b000000011111111;
													assign node6741 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node6744 = (inp[12]) ? node6748 : node6745;
												assign node6745 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6748 = (inp[2]) ? node6752 : node6749;
													assign node6749 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6752 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node6755 = (inp[6]) ? node6831 : node6756;
								assign node6756 = (inp[4]) ? node6792 : node6757;
									assign node6757 = (inp[1]) ? node6775 : node6758;
										assign node6758 = (inp[0]) ? node6768 : node6759;
											assign node6759 = (inp[7]) ? node6761 : 15'b000001111111111;
												assign node6761 = (inp[8]) ? node6765 : node6762;
													assign node6762 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node6765 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node6768 = (inp[8]) ? node6770 : 15'b000000111111111;
												assign node6770 = (inp[14]) ? node6772 : 15'b000000011111111;
													assign node6772 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6775 = (inp[12]) ? node6783 : node6776;
											assign node6776 = (inp[0]) ? node6778 : 15'b000000111111111;
												assign node6778 = (inp[7]) ? 15'b000000011111111 : node6779;
													assign node6779 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6783 = (inp[2]) ? node6789 : node6784;
												assign node6784 = (inp[7]) ? node6786 : 15'b000000011111111;
													assign node6786 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node6789 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node6792 = (inp[12]) ? node6812 : node6793;
										assign node6793 = (inp[14]) ? node6805 : node6794;
											assign node6794 = (inp[8]) ? node6800 : node6795;
												assign node6795 = (inp[2]) ? 15'b000000111111111 : node6796;
													assign node6796 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node6800 = (inp[7]) ? node6802 : 15'b000000111111111;
													assign node6802 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6805 = (inp[8]) ? 15'b000000000111111 : node6806;
												assign node6806 = (inp[2]) ? node6808 : 15'b000000001111111;
													assign node6808 = (inp[0]) ? 15'b000000011111111 : 15'b000000011111111;
										assign node6812 = (inp[14]) ? node6822 : node6813;
											assign node6813 = (inp[1]) ? 15'b000000001111111 : node6814;
												assign node6814 = (inp[7]) ? node6818 : node6815;
													assign node6815 = (inp[2]) ? 15'b000000111111111 : 15'b000000011111111;
													assign node6818 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6822 = (inp[2]) ? node6828 : node6823;
												assign node6823 = (inp[7]) ? node6825 : 15'b000000001111111;
													assign node6825 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6828 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node6831 = (inp[1]) ? node6873 : node6832;
									assign node6832 = (inp[7]) ? node6852 : node6833;
										assign node6833 = (inp[8]) ? node6841 : node6834;
											assign node6834 = (inp[14]) ? 15'b000000011111111 : node6835;
												assign node6835 = (inp[4]) ? 15'b000000111111111 : node6836;
													assign node6836 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6841 = (inp[4]) ? node6847 : node6842;
												assign node6842 = (inp[14]) ? 15'b000000011111111 : node6843;
													assign node6843 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6847 = (inp[0]) ? node6849 : 15'b000000001111111;
													assign node6849 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6852 = (inp[0]) ? node6866 : node6853;
											assign node6853 = (inp[14]) ? node6861 : node6854;
												assign node6854 = (inp[12]) ? node6858 : node6855;
													assign node6855 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6858 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node6861 = (inp[4]) ? node6863 : 15'b000000001111111;
													assign node6863 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node6866 = (inp[12]) ? node6868 : 15'b000000001111111;
												assign node6868 = (inp[14]) ? node6870 : 15'b000000000111111;
													assign node6870 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node6873 = (inp[0]) ? node6887 : node6874;
										assign node6874 = (inp[8]) ? node6876 : 15'b000000001111111;
											assign node6876 = (inp[14]) ? node6882 : node6877;
												assign node6877 = (inp[2]) ? node6879 : 15'b000000011111111;
													assign node6879 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6882 = (inp[4]) ? 15'b000000000111111 : node6883;
													assign node6883 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6887 = (inp[2]) ? node6895 : node6888;
											assign node6888 = (inp[8]) ? 15'b000000000111111 : node6889;
												assign node6889 = (inp[14]) ? node6891 : 15'b000000001111111;
													assign node6891 = (inp[4]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node6895 = (inp[12]) ? 15'b000000000011111 : node6896;
												assign node6896 = (inp[8]) ? node6900 : node6897;
													assign node6897 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node6900 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node6904 = (inp[1]) ? node7074 : node6905;
							assign node6905 = (inp[0]) ? node6991 : node6906;
								assign node6906 = (inp[12]) ? node6952 : node6907;
									assign node6907 = (inp[7]) ? node6933 : node6908;
										assign node6908 = (inp[6]) ? node6924 : node6909;
											assign node6909 = (inp[14]) ? node6917 : node6910;
												assign node6910 = (inp[10]) ? node6914 : node6911;
													assign node6911 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6914 = (inp[2]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node6917 = (inp[10]) ? node6921 : node6918;
													assign node6918 = (inp[8]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node6921 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6924 = (inp[8]) ? node6930 : node6925;
												assign node6925 = (inp[2]) ? 15'b000000111111111 : node6926;
													assign node6926 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6930 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6933 = (inp[10]) ? node6945 : node6934;
											assign node6934 = (inp[6]) ? node6938 : node6935;
												assign node6935 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6938 = (inp[14]) ? node6942 : node6939;
													assign node6939 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node6942 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node6945 = (inp[4]) ? 15'b000000001111111 : node6946;
												assign node6946 = (inp[6]) ? node6948 : 15'b000000011111111;
													assign node6948 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6952 = (inp[2]) ? node6970 : node6953;
										assign node6953 = (inp[6]) ? node6963 : node6954;
											assign node6954 = (inp[14]) ? node6960 : node6955;
												assign node6955 = (inp[7]) ? 15'b000000111111111 : node6956;
													assign node6956 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6960 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6963 = (inp[8]) ? 15'b000000001111111 : node6964;
												assign node6964 = (inp[14]) ? node6966 : 15'b000000111111111;
													assign node6966 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node6970 = (inp[8]) ? node6982 : node6971;
											assign node6971 = (inp[4]) ? node6977 : node6972;
												assign node6972 = (inp[14]) ? 15'b000000011111111 : node6973;
													assign node6973 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6977 = (inp[7]) ? 15'b000000000111111 : node6978;
													assign node6978 = (inp[6]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node6982 = (inp[10]) ? node6988 : node6983;
												assign node6983 = (inp[6]) ? 15'b000000000111111 : node6984;
													assign node6984 = (inp[4]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node6988 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6991 = (inp[4]) ? node7039 : node6992;
									assign node6992 = (inp[2]) ? node7014 : node6993;
										assign node6993 = (inp[6]) ? node7001 : node6994;
											assign node6994 = (inp[10]) ? node6996 : 15'b000000111111111;
												assign node6996 = (inp[7]) ? node6998 : 15'b000000111111111;
													assign node6998 = (inp[8]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node7001 = (inp[10]) ? node7009 : node7002;
												assign node7002 = (inp[7]) ? node7006 : node7003;
													assign node7003 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7006 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7009 = (inp[14]) ? node7011 : 15'b000000001111111;
													assign node7011 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7014 = (inp[7]) ? node7028 : node7015;
											assign node7015 = (inp[12]) ? node7021 : node7016;
												assign node7016 = (inp[8]) ? node7018 : 15'b000000111111111;
													assign node7018 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7021 = (inp[8]) ? node7025 : node7022;
													assign node7022 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7025 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7028 = (inp[14]) ? node7034 : node7029;
												assign node7029 = (inp[12]) ? 15'b000000000111111 : node7030;
													assign node7030 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7034 = (inp[8]) ? node7036 : 15'b000000000111111;
													assign node7036 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7039 = (inp[10]) ? node7053 : node7040;
										assign node7040 = (inp[12]) ? node7046 : node7041;
											assign node7041 = (inp[6]) ? node7043 : 15'b000000011111111;
												assign node7043 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7046 = (inp[14]) ? node7048 : 15'b000000001111111;
												assign node7048 = (inp[7]) ? 15'b000000000111111 : node7049;
													assign node7049 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7053 = (inp[7]) ? node7067 : node7054;
											assign node7054 = (inp[14]) ? node7060 : node7055;
												assign node7055 = (inp[6]) ? node7057 : 15'b000000001111111;
													assign node7057 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7060 = (inp[2]) ? node7064 : node7061;
													assign node7061 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7064 = (inp[12]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node7067 = (inp[12]) ? node7069 : 15'b000000000111111;
												assign node7069 = (inp[6]) ? node7071 : 15'b000000000011111;
													assign node7071 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node7074 = (inp[8]) ? node7162 : node7075;
								assign node7075 = (inp[12]) ? node7123 : node7076;
									assign node7076 = (inp[4]) ? node7096 : node7077;
										assign node7077 = (inp[10]) ? node7089 : node7078;
											assign node7078 = (inp[7]) ? node7084 : node7079;
												assign node7079 = (inp[6]) ? 15'b000000111111111 : node7080;
													assign node7080 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7084 = (inp[0]) ? 15'b000000011111111 : node7085;
													assign node7085 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7089 = (inp[0]) ? node7091 : 15'b000000011111111;
												assign node7091 = (inp[7]) ? node7093 : 15'b000000111111111;
													assign node7093 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7096 = (inp[7]) ? node7110 : node7097;
											assign node7097 = (inp[14]) ? node7105 : node7098;
												assign node7098 = (inp[6]) ? node7102 : node7099;
													assign node7099 = (inp[10]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node7102 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7105 = (inp[6]) ? 15'b000000001111111 : node7106;
													assign node7106 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7110 = (inp[0]) ? node7116 : node7111;
												assign node7111 = (inp[6]) ? node7113 : 15'b000000111111111;
													assign node7113 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7116 = (inp[10]) ? node7120 : node7117;
													assign node7117 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7120 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7123 = (inp[14]) ? node7149 : node7124;
										assign node7124 = (inp[7]) ? node7138 : node7125;
											assign node7125 = (inp[4]) ? node7131 : node7126;
												assign node7126 = (inp[10]) ? node7128 : 15'b000000111111111;
													assign node7128 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7131 = (inp[10]) ? node7135 : node7132;
													assign node7132 = (inp[6]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node7135 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7138 = (inp[4]) ? node7144 : node7139;
												assign node7139 = (inp[6]) ? node7141 : 15'b000000001111111;
													assign node7141 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7144 = (inp[10]) ? 15'b000000000011111 : node7145;
													assign node7145 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7149 = (inp[6]) ? node7155 : node7150;
											assign node7150 = (inp[10]) ? 15'b000000000011111 : node7151;
												assign node7151 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node7155 = (inp[0]) ? node7157 : 15'b000000000111111;
												assign node7157 = (inp[10]) ? 15'b000000000011111 : node7158;
													assign node7158 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node7162 = (inp[6]) ? node7202 : node7163;
									assign node7163 = (inp[14]) ? node7185 : node7164;
										assign node7164 = (inp[7]) ? node7176 : node7165;
											assign node7165 = (inp[12]) ? node7171 : node7166;
												assign node7166 = (inp[0]) ? 15'b000000011111111 : node7167;
													assign node7167 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7171 = (inp[0]) ? 15'b000000000111111 : node7172;
													assign node7172 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node7176 = (inp[10]) ? node7180 : node7177;
												assign node7177 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7180 = (inp[12]) ? node7182 : 15'b000000000111111;
													assign node7182 = (inp[2]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node7185 = (inp[0]) ? node7193 : node7186;
											assign node7186 = (inp[7]) ? 15'b000000000111111 : node7187;
												assign node7187 = (inp[2]) ? node7189 : 15'b000000001111111;
													assign node7189 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7193 = (inp[7]) ? 15'b000000000011111 : node7194;
												assign node7194 = (inp[10]) ? node7198 : node7195;
													assign node7195 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7198 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7202 = (inp[14]) ? node7226 : node7203;
										assign node7203 = (inp[12]) ? node7211 : node7204;
											assign node7204 = (inp[0]) ? 15'b000000000111111 : node7205;
												assign node7205 = (inp[2]) ? node7207 : 15'b000000001111111;
													assign node7207 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7211 = (inp[2]) ? node7219 : node7212;
												assign node7212 = (inp[4]) ? node7216 : node7213;
													assign node7213 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7216 = (inp[10]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node7219 = (inp[4]) ? node7223 : node7220;
													assign node7220 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7223 = (inp[0]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node7226 = (inp[4]) ? node7236 : node7227;
											assign node7227 = (inp[0]) ? 15'b000000000011111 : node7228;
												assign node7228 = (inp[2]) ? node7232 : node7229;
													assign node7229 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7232 = (inp[10]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node7236 = (inp[10]) ? node7240 : node7237;
												assign node7237 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7240 = (inp[2]) ? 15'b000000000001111 : node7241;
													assign node7241 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node7245 = (inp[2]) ? node7569 : node7246;
						assign node7246 = (inp[10]) ? node7398 : node7247;
							assign node7247 = (inp[7]) ? node7323 : node7248;
								assign node7248 = (inp[4]) ? node7294 : node7249;
									assign node7249 = (inp[12]) ? node7275 : node7250;
										assign node7250 = (inp[0]) ? node7262 : node7251;
											assign node7251 = (inp[1]) ? node7259 : node7252;
												assign node7252 = (inp[14]) ? node7256 : node7253;
													assign node7253 = (inp[8]) ? 15'b000001111111111 : 15'b000001111111111;
													assign node7256 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7259 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node7262 = (inp[6]) ? node7268 : node7263;
												assign node7263 = (inp[9]) ? 15'b000000011111111 : node7264;
													assign node7264 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7268 = (inp[14]) ? node7272 : node7269;
													assign node7269 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7272 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node7275 = (inp[14]) ? node7283 : node7276;
											assign node7276 = (inp[6]) ? node7278 : 15'b000000111111111;
												assign node7278 = (inp[0]) ? 15'b000000011111111 : node7279;
													assign node7279 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7283 = (inp[6]) ? node7289 : node7284;
												assign node7284 = (inp[0]) ? 15'b000000011111111 : node7285;
													assign node7285 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7289 = (inp[1]) ? node7291 : 15'b000000011111111;
													assign node7291 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7294 = (inp[1]) ? node7310 : node7295;
										assign node7295 = (inp[6]) ? node7303 : node7296;
											assign node7296 = (inp[0]) ? 15'b000000011111111 : node7297;
												assign node7297 = (inp[9]) ? 15'b000000111111111 : node7298;
													assign node7298 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node7303 = (inp[9]) ? node7305 : 15'b000000011111111;
												assign node7305 = (inp[14]) ? 15'b000000001111111 : node7306;
													assign node7306 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node7310 = (inp[8]) ? node7314 : node7311;
											assign node7311 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7314 = (inp[14]) ? node7320 : node7315;
												assign node7315 = (inp[0]) ? node7317 : 15'b000000001111111;
													assign node7317 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7320 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node7323 = (inp[12]) ? node7355 : node7324;
									assign node7324 = (inp[1]) ? node7336 : node7325;
										assign node7325 = (inp[6]) ? node7331 : node7326;
											assign node7326 = (inp[14]) ? 15'b000000011111111 : node7327;
												assign node7327 = (inp[9]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node7331 = (inp[14]) ? node7333 : 15'b000000011111111;
												assign node7333 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7336 = (inp[8]) ? node7346 : node7337;
											assign node7337 = (inp[6]) ? node7339 : 15'b000000011111111;
												assign node7339 = (inp[14]) ? node7343 : node7340;
													assign node7340 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7343 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7346 = (inp[4]) ? node7352 : node7347;
												assign node7347 = (inp[9]) ? 15'b000000001111111 : node7348;
													assign node7348 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7352 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node7355 = (inp[6]) ? node7379 : node7356;
										assign node7356 = (inp[1]) ? node7368 : node7357;
											assign node7357 = (inp[8]) ? node7363 : node7358;
												assign node7358 = (inp[9]) ? node7360 : 15'b000000111111111;
													assign node7360 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node7363 = (inp[0]) ? 15'b000000000111111 : node7364;
													assign node7364 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7368 = (inp[9]) ? node7374 : node7369;
												assign node7369 = (inp[14]) ? node7371 : 15'b000000001111111;
													assign node7371 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7374 = (inp[14]) ? 15'b000000000111111 : node7375;
													assign node7375 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node7379 = (inp[4]) ? node7387 : node7380;
											assign node7380 = (inp[1]) ? node7382 : 15'b000000001111111;
												assign node7382 = (inp[0]) ? 15'b000000000111111 : node7383;
													assign node7383 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7387 = (inp[8]) ? node7391 : node7388;
												assign node7388 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7391 = (inp[1]) ? node7395 : node7392;
													assign node7392 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7395 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node7398 = (inp[9]) ? node7478 : node7399;
								assign node7399 = (inp[8]) ? node7433 : node7400;
									assign node7400 = (inp[0]) ? node7420 : node7401;
										assign node7401 = (inp[14]) ? node7415 : node7402;
											assign node7402 = (inp[6]) ? node7410 : node7403;
												assign node7403 = (inp[7]) ? node7407 : node7404;
													assign node7404 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7407 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7410 = (inp[7]) ? node7412 : 15'b000000011111111;
													assign node7412 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7415 = (inp[7]) ? node7417 : 15'b000000011111111;
												assign node7417 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node7420 = (inp[12]) ? node7428 : node7421;
											assign node7421 = (inp[6]) ? 15'b000000001111111 : node7422;
												assign node7422 = (inp[14]) ? 15'b000000001111111 : node7423;
													assign node7423 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7428 = (inp[4]) ? node7430 : 15'b000000001111111;
												assign node7430 = (inp[6]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node7433 = (inp[1]) ? node7455 : node7434;
										assign node7434 = (inp[12]) ? node7446 : node7435;
											assign node7435 = (inp[14]) ? node7441 : node7436;
												assign node7436 = (inp[4]) ? 15'b000000011111111 : node7437;
													assign node7437 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7441 = (inp[4]) ? 15'b000000001111111 : node7442;
													assign node7442 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7446 = (inp[0]) ? node7452 : node7447;
												assign node7447 = (inp[4]) ? node7449 : 15'b000000011111111;
													assign node7449 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7452 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7455 = (inp[4]) ? node7469 : node7456;
											assign node7456 = (inp[14]) ? node7462 : node7457;
												assign node7457 = (inp[6]) ? node7459 : 15'b000000001111111;
													assign node7459 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7462 = (inp[12]) ? node7466 : node7463;
													assign node7463 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7466 = (inp[7]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node7469 = (inp[12]) ? node7473 : node7470;
												assign node7470 = (inp[0]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node7473 = (inp[0]) ? node7475 : 15'b000000000011111;
													assign node7475 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node7478 = (inp[12]) ? node7526 : node7479;
									assign node7479 = (inp[4]) ? node7503 : node7480;
										assign node7480 = (inp[0]) ? node7494 : node7481;
											assign node7481 = (inp[1]) ? node7489 : node7482;
												assign node7482 = (inp[6]) ? node7486 : node7483;
													assign node7483 = (inp[7]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node7486 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7489 = (inp[8]) ? node7491 : 15'b000000001111111;
													assign node7491 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7494 = (inp[1]) ? node7498 : node7495;
												assign node7495 = (inp[8]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node7498 = (inp[7]) ? node7500 : 15'b000000000111111;
													assign node7500 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7503 = (inp[1]) ? node7517 : node7504;
											assign node7504 = (inp[0]) ? node7510 : node7505;
												assign node7505 = (inp[6]) ? node7507 : 15'b000000001111111;
													assign node7507 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7510 = (inp[7]) ? node7514 : node7511;
													assign node7511 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7514 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7517 = (inp[6]) ? node7519 : 15'b000000000111111;
												assign node7519 = (inp[7]) ? node7523 : node7520;
													assign node7520 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7523 = (inp[8]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node7526 = (inp[7]) ? node7544 : node7527;
										assign node7527 = (inp[4]) ? node7539 : node7528;
											assign node7528 = (inp[8]) ? node7534 : node7529;
												assign node7529 = (inp[14]) ? 15'b000000000111111 : node7530;
													assign node7530 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7534 = (inp[14]) ? node7536 : 15'b000000000111111;
													assign node7536 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7539 = (inp[0]) ? node7541 : 15'b000000001111111;
												assign node7541 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7544 = (inp[1]) ? node7556 : node7545;
											assign node7545 = (inp[14]) ? node7551 : node7546;
												assign node7546 = (inp[6]) ? node7548 : 15'b000000000111111;
													assign node7548 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7551 = (inp[4]) ? node7553 : 15'b000000000111111;
													assign node7553 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7556 = (inp[4]) ? node7564 : node7557;
												assign node7557 = (inp[6]) ? node7561 : node7558;
													assign node7558 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node7561 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7564 = (inp[14]) ? node7566 : 15'b000000000011111;
													assign node7566 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node7569 = (inp[4]) ? node7699 : node7570;
							assign node7570 = (inp[9]) ? node7634 : node7571;
								assign node7571 = (inp[1]) ? node7597 : node7572;
									assign node7572 = (inp[14]) ? node7592 : node7573;
										assign node7573 = (inp[7]) ? node7585 : node7574;
											assign node7574 = (inp[0]) ? node7580 : node7575;
												assign node7575 = (inp[10]) ? node7577 : 15'b000011111111111;
													assign node7577 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7580 = (inp[10]) ? node7582 : 15'b000000111111111;
													assign node7582 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7585 = (inp[10]) ? 15'b000000001111111 : node7586;
												assign node7586 = (inp[0]) ? 15'b000000001111111 : node7587;
													assign node7587 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node7592 = (inp[7]) ? node7594 : 15'b000000001111111;
											assign node7594 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node7597 = (inp[8]) ? node7617 : node7598;
										assign node7598 = (inp[6]) ? node7608 : node7599;
											assign node7599 = (inp[10]) ? node7605 : node7600;
												assign node7600 = (inp[7]) ? node7602 : 15'b000000011111111;
													assign node7602 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7605 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node7608 = (inp[12]) ? node7614 : node7609;
												assign node7609 = (inp[0]) ? node7611 : 15'b000000001111111;
													assign node7611 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7614 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7617 = (inp[10]) ? node7627 : node7618;
											assign node7618 = (inp[12]) ? node7620 : 15'b000000001111111;
												assign node7620 = (inp[6]) ? node7624 : node7621;
													assign node7621 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node7624 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7627 = (inp[7]) ? node7629 : 15'b000000000111111;
												assign node7629 = (inp[12]) ? 15'b000000000011111 : node7630;
													assign node7630 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node7634 = (inp[6]) ? node7660 : node7635;
									assign node7635 = (inp[0]) ? node7645 : node7636;
										assign node7636 = (inp[10]) ? node7642 : node7637;
											assign node7637 = (inp[12]) ? 15'b000000001111111 : node7638;
												assign node7638 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node7642 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7645 = (inp[12]) ? node7653 : node7646;
											assign node7646 = (inp[7]) ? node7648 : 15'b000000011111111;
												assign node7648 = (inp[8]) ? 15'b000000000111111 : node7649;
													assign node7649 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7653 = (inp[14]) ? node7655 : 15'b000000000111111;
												assign node7655 = (inp[8]) ? 15'b000000000001111 : node7656;
													assign node7656 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7660 = (inp[7]) ? node7678 : node7661;
										assign node7661 = (inp[8]) ? node7669 : node7662;
											assign node7662 = (inp[10]) ? node7666 : node7663;
												assign node7663 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7666 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7669 = (inp[0]) ? node7671 : 15'b000000000111111;
												assign node7671 = (inp[10]) ? node7675 : node7672;
													assign node7672 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7675 = (inp[14]) ? 15'b000000000000111 : 15'b000000000011111;
										assign node7678 = (inp[12]) ? node7684 : node7679;
											assign node7679 = (inp[10]) ? 15'b000000000011111 : node7680;
												assign node7680 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node7684 = (inp[8]) ? node7692 : node7685;
												assign node7685 = (inp[10]) ? node7689 : node7686;
													assign node7686 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7689 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7692 = (inp[14]) ? node7696 : node7693;
													assign node7693 = (inp[0]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node7696 = (inp[0]) ? 15'b000000000000011 : 15'b000000000001111;
							assign node7699 = (inp[6]) ? node7793 : node7700;
								assign node7700 = (inp[0]) ? node7746 : node7701;
									assign node7701 = (inp[7]) ? node7723 : node7702;
										assign node7702 = (inp[10]) ? node7714 : node7703;
											assign node7703 = (inp[9]) ? node7711 : node7704;
												assign node7704 = (inp[14]) ? node7708 : node7705;
													assign node7705 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7708 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7711 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7714 = (inp[12]) ? node7718 : node7715;
												assign node7715 = (inp[9]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node7718 = (inp[9]) ? 15'b000000000111111 : node7719;
													assign node7719 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7723 = (inp[12]) ? node7735 : node7724;
											assign node7724 = (inp[1]) ? node7732 : node7725;
												assign node7725 = (inp[14]) ? node7729 : node7726;
													assign node7726 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7729 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7732 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7735 = (inp[1]) ? node7741 : node7736;
												assign node7736 = (inp[10]) ? 15'b000000000011111 : node7737;
													assign node7737 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7741 = (inp[14]) ? node7743 : 15'b000000000011111;
													assign node7743 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7746 = (inp[14]) ? node7766 : node7747;
										assign node7747 = (inp[12]) ? node7755 : node7748;
											assign node7748 = (inp[8]) ? 15'b000000000111111 : node7749;
												assign node7749 = (inp[7]) ? 15'b000000001111111 : node7750;
													assign node7750 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7755 = (inp[8]) ? node7759 : node7756;
												assign node7756 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7759 = (inp[9]) ? node7763 : node7760;
													assign node7760 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7763 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7766 = (inp[8]) ? node7778 : node7767;
											assign node7767 = (inp[7]) ? node7773 : node7768;
												assign node7768 = (inp[9]) ? node7770 : 15'b000000000111111;
													assign node7770 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7773 = (inp[10]) ? node7775 : 15'b000000000111111;
													assign node7775 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7778 = (inp[12]) ? node7786 : node7779;
												assign node7779 = (inp[10]) ? node7783 : node7780;
													assign node7780 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7783 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7786 = (inp[1]) ? node7790 : node7787;
													assign node7787 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7790 = (inp[7]) ? 15'b000000000000111 : 15'b000000000000111;
								assign node7793 = (inp[8]) ? node7841 : node7794;
									assign node7794 = (inp[10]) ? node7820 : node7795;
										assign node7795 = (inp[7]) ? node7809 : node7796;
											assign node7796 = (inp[0]) ? node7804 : node7797;
												assign node7797 = (inp[12]) ? node7801 : node7798;
													assign node7798 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7801 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7804 = (inp[1]) ? 15'b000000000111111 : node7805;
													assign node7805 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7809 = (inp[14]) ? node7815 : node7810;
												assign node7810 = (inp[0]) ? 15'b000000000011111 : node7811;
													assign node7811 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node7815 = (inp[9]) ? node7817 : 15'b000000000011111;
													assign node7817 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7820 = (inp[9]) ? node7832 : node7821;
											assign node7821 = (inp[7]) ? node7827 : node7822;
												assign node7822 = (inp[1]) ? node7824 : 15'b000000000111111;
													assign node7824 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7827 = (inp[12]) ? node7829 : 15'b000000000011111;
													assign node7829 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7832 = (inp[1]) ? node7838 : node7833;
												assign node7833 = (inp[14]) ? 15'b000000000001111 : node7834;
													assign node7834 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node7838 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node7841 = (inp[9]) ? node7871 : node7842;
										assign node7842 = (inp[1]) ? node7858 : node7843;
											assign node7843 = (inp[14]) ? node7851 : node7844;
												assign node7844 = (inp[7]) ? node7848 : node7845;
													assign node7845 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7848 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7851 = (inp[7]) ? node7855 : node7852;
													assign node7852 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7855 = (inp[0]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node7858 = (inp[14]) ? node7864 : node7859;
												assign node7859 = (inp[0]) ? node7861 : 15'b000000000011111;
													assign node7861 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7864 = (inp[0]) ? node7868 : node7865;
													assign node7865 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7868 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node7871 = (inp[1]) ? node7883 : node7872;
											assign node7872 = (inp[7]) ? node7878 : node7873;
												assign node7873 = (inp[14]) ? node7875 : 15'b000000000011111;
													assign node7875 = (inp[10]) ? 15'b000000000001111 : 15'b000000000001111;
												assign node7878 = (inp[10]) ? 15'b000000000001111 : node7879;
													assign node7879 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node7883 = (inp[14]) ? node7887 : node7884;
												assign node7884 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node7887 = (inp[0]) ? node7889 : 15'b000000000000111;
													assign node7889 = (inp[10]) ? 15'b000000000000001 : 15'b000000000000111;
			assign node7892 = (inp[4]) ? node9196 : node7893;
				assign node7893 = (inp[5]) ? node8507 : node7894;
					assign node7894 = (inp[8]) ? node8196 : node7895;
						assign node7895 = (inp[0]) ? node8049 : node7896;
							assign node7896 = (inp[10]) ? node7984 : node7897;
								assign node7897 = (inp[1]) ? node7943 : node7898;
									assign node7898 = (inp[6]) ? node7922 : node7899;
										assign node7899 = (inp[13]) ? node7911 : node7900;
											assign node7900 = (inp[12]) ? node7906 : node7901;
												assign node7901 = (inp[9]) ? 15'b000011111111111 : node7902;
													assign node7902 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node7906 = (inp[9]) ? 15'b000001111111111 : node7907;
													assign node7907 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node7911 = (inp[12]) ? node7917 : node7912;
												assign node7912 = (inp[9]) ? 15'b000001111111111 : node7913;
													assign node7913 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7917 = (inp[7]) ? 15'b000000111111111 : node7918;
													assign node7918 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node7922 = (inp[14]) ? node7938 : node7923;
											assign node7923 = (inp[13]) ? node7931 : node7924;
												assign node7924 = (inp[7]) ? node7928 : node7925;
													assign node7925 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7928 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7931 = (inp[2]) ? node7935 : node7932;
													assign node7932 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7935 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7938 = (inp[2]) ? 15'b000000011111111 : node7939;
												assign node7939 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node7943 = (inp[12]) ? node7967 : node7944;
										assign node7944 = (inp[2]) ? node7956 : node7945;
											assign node7945 = (inp[14]) ? node7951 : node7946;
												assign node7946 = (inp[7]) ? 15'b000001111111111 : node7947;
													assign node7947 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7951 = (inp[7]) ? node7953 : 15'b000001111111111;
													assign node7953 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7956 = (inp[9]) ? node7960 : node7957;
												assign node7957 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7960 = (inp[7]) ? node7964 : node7961;
													assign node7961 = (inp[13]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node7964 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node7967 = (inp[6]) ? node7977 : node7968;
											assign node7968 = (inp[14]) ? node7974 : node7969;
												assign node7969 = (inp[2]) ? 15'b000000011111111 : node7970;
													assign node7970 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7974 = (inp[13]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node7977 = (inp[9]) ? node7979 : 15'b000000011111111;
												assign node7979 = (inp[2]) ? 15'b000000000111111 : node7980;
													assign node7980 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node7984 = (inp[12]) ? node8024 : node7985;
									assign node7985 = (inp[1]) ? node8009 : node7986;
										assign node7986 = (inp[2]) ? node8000 : node7987;
											assign node7987 = (inp[13]) ? node7993 : node7988;
												assign node7988 = (inp[7]) ? 15'b000001111111111 : node7989;
													assign node7989 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7993 = (inp[14]) ? node7997 : node7994;
													assign node7994 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7997 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8000 = (inp[7]) ? node8002 : 15'b000000111111111;
												assign node8002 = (inp[13]) ? node8006 : node8003;
													assign node8003 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8006 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8009 = (inp[14]) ? node8017 : node8010;
											assign node8010 = (inp[13]) ? node8012 : 15'b000000111111111;
												assign node8012 = (inp[2]) ? node8014 : 15'b000000111111111;
													assign node8014 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8017 = (inp[6]) ? node8021 : node8018;
												assign node8018 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8021 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node8024 = (inp[9]) ? node8038 : node8025;
										assign node8025 = (inp[14]) ? node8031 : node8026;
											assign node8026 = (inp[7]) ? 15'b000000011111111 : node8027;
												assign node8027 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8031 = (inp[13]) ? 15'b000000001111111 : node8032;
												assign node8032 = (inp[6]) ? 15'b000000011111111 : node8033;
													assign node8033 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node8038 = (inp[7]) ? node8044 : node8039;
											assign node8039 = (inp[2]) ? 15'b000000001111111 : node8040;
												assign node8040 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8044 = (inp[1]) ? node8046 : 15'b000000001111111;
												assign node8046 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node8049 = (inp[13]) ? node8125 : node8050;
								assign node8050 = (inp[2]) ? node8092 : node8051;
									assign node8051 = (inp[7]) ? node8071 : node8052;
										assign node8052 = (inp[10]) ? node8058 : node8053;
											assign node8053 = (inp[1]) ? 15'b000000111111111 : node8054;
												assign node8054 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node8058 = (inp[6]) ? node8066 : node8059;
												assign node8059 = (inp[12]) ? node8063 : node8060;
													assign node8060 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8063 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8066 = (inp[1]) ? 15'b000000011111111 : node8067;
													assign node8067 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node8071 = (inp[1]) ? node8079 : node8072;
											assign node8072 = (inp[14]) ? node8074 : 15'b000000111111111;
												assign node8074 = (inp[9]) ? 15'b000000001111111 : node8075;
													assign node8075 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node8079 = (inp[6]) ? node8085 : node8080;
												assign node8080 = (inp[12]) ? 15'b000000011111111 : node8081;
													assign node8081 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8085 = (inp[9]) ? node8089 : node8086;
													assign node8086 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8089 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8092 = (inp[10]) ? node8110 : node8093;
										assign node8093 = (inp[7]) ? node8099 : node8094;
											assign node8094 = (inp[12]) ? 15'b000000011111111 : node8095;
												assign node8095 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node8099 = (inp[6]) ? node8105 : node8100;
												assign node8100 = (inp[9]) ? 15'b000000011111111 : node8101;
													assign node8101 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8105 = (inp[12]) ? node8107 : 15'b000000001111111;
													assign node8107 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8110 = (inp[9]) ? node8118 : node8111;
											assign node8111 = (inp[1]) ? node8113 : 15'b000000111111111;
												assign node8113 = (inp[12]) ? 15'b000000001111111 : node8114;
													assign node8114 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8118 = (inp[7]) ? 15'b000000000111111 : node8119;
												assign node8119 = (inp[14]) ? node8121 : 15'b000000001111111;
													assign node8121 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node8125 = (inp[7]) ? node8157 : node8126;
									assign node8126 = (inp[10]) ? node8138 : node8127;
										assign node8127 = (inp[14]) ? node8131 : node8128;
											assign node8128 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8131 = (inp[1]) ? node8135 : node8132;
												assign node8132 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8135 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8138 = (inp[2]) ? node8150 : node8139;
											assign node8139 = (inp[1]) ? node8143 : node8140;
												assign node8140 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8143 = (inp[6]) ? node8147 : node8144;
													assign node8144 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8147 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8150 = (inp[9]) ? node8154 : node8151;
												assign node8151 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8154 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node8157 = (inp[14]) ? node8177 : node8158;
										assign node8158 = (inp[1]) ? node8172 : node8159;
											assign node8159 = (inp[2]) ? node8167 : node8160;
												assign node8160 = (inp[12]) ? node8164 : node8161;
													assign node8161 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8164 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8167 = (inp[6]) ? node8169 : 15'b000000001111111;
													assign node8169 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node8172 = (inp[9]) ? 15'b000000000111111 : node8173;
												assign node8173 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8177 = (inp[12]) ? node8183 : node8178;
											assign node8178 = (inp[9]) ? 15'b000000000111111 : node8179;
												assign node8179 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8183 = (inp[6]) ? node8189 : node8184;
												assign node8184 = (inp[9]) ? node8186 : 15'b000000000111111;
													assign node8186 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8189 = (inp[2]) ? node8193 : node8190;
													assign node8190 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8193 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node8196 = (inp[13]) ? node8350 : node8197;
							assign node8197 = (inp[2]) ? node8267 : node8198;
								assign node8198 = (inp[6]) ? node8236 : node8199;
									assign node8199 = (inp[9]) ? node8217 : node8200;
										assign node8200 = (inp[7]) ? node8210 : node8201;
											assign node8201 = (inp[10]) ? node8205 : node8202;
												assign node8202 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8205 = (inp[1]) ? 15'b000000111111111 : node8206;
													assign node8206 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8210 = (inp[10]) ? 15'b000000011111111 : node8211;
												assign node8211 = (inp[12]) ? node8213 : 15'b000000111111111;
													assign node8213 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node8217 = (inp[1]) ? node8227 : node8218;
											assign node8218 = (inp[12]) ? node8220 : 15'b000000111111111;
												assign node8220 = (inp[10]) ? node8224 : node8221;
													assign node8221 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8224 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8227 = (inp[0]) ? node8233 : node8228;
												assign node8228 = (inp[10]) ? 15'b000000001111111 : node8229;
													assign node8229 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8233 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8236 = (inp[7]) ? node8250 : node8237;
										assign node8237 = (inp[0]) ? node8243 : node8238;
											assign node8238 = (inp[1]) ? node8240 : 15'b000000111111111;
												assign node8240 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8243 = (inp[14]) ? node8245 : 15'b000000011111111;
												assign node8245 = (inp[9]) ? 15'b000000001111111 : node8246;
													assign node8246 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8250 = (inp[10]) ? node8260 : node8251;
											assign node8251 = (inp[14]) ? 15'b000000001111111 : node8252;
												assign node8252 = (inp[0]) ? node8256 : node8253;
													assign node8253 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8256 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8260 = (inp[14]) ? 15'b000000000111111 : node8261;
												assign node8261 = (inp[1]) ? 15'b000000001111111 : node8262;
													assign node8262 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node8267 = (inp[14]) ? node8311 : node8268;
									assign node8268 = (inp[1]) ? node8292 : node8269;
										assign node8269 = (inp[7]) ? node8283 : node8270;
											assign node8270 = (inp[6]) ? node8276 : node8271;
												assign node8271 = (inp[10]) ? node8273 : 15'b000001111111111;
													assign node8273 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8276 = (inp[12]) ? node8280 : node8277;
													assign node8277 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8280 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8283 = (inp[6]) ? node8287 : node8284;
												assign node8284 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node8287 = (inp[9]) ? 15'b000000001111111 : node8288;
													assign node8288 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8292 = (inp[10]) ? node8304 : node8293;
											assign node8293 = (inp[7]) ? node8299 : node8294;
												assign node8294 = (inp[0]) ? 15'b000000001111111 : node8295;
													assign node8295 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8299 = (inp[9]) ? 15'b000000000111111 : node8300;
													assign node8300 = (inp[6]) ? 15'b000000001111111 : 15'b000000001111111;
											assign node8304 = (inp[0]) ? node8306 : 15'b000000001111111;
												assign node8306 = (inp[12]) ? 15'b000000000111111 : node8307;
													assign node8307 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8311 = (inp[1]) ? node8331 : node8312;
										assign node8312 = (inp[0]) ? node8320 : node8313;
											assign node8313 = (inp[7]) ? node8315 : 15'b000000111111111;
												assign node8315 = (inp[6]) ? 15'b000000001111111 : node8316;
													assign node8316 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8320 = (inp[9]) ? node8326 : node8321;
												assign node8321 = (inp[12]) ? node8323 : 15'b000000011111111;
													assign node8323 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8326 = (inp[12]) ? node8328 : 15'b000000000111111;
													assign node8328 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node8331 = (inp[0]) ? node8343 : node8332;
											assign node8332 = (inp[10]) ? node8338 : node8333;
												assign node8333 = (inp[7]) ? node8335 : 15'b000000001111111;
													assign node8335 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8338 = (inp[9]) ? 15'b000000000001111 : node8339;
													assign node8339 = (inp[6]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node8343 = (inp[6]) ? 15'b000000000011111 : node8344;
												assign node8344 = (inp[10]) ? node8346 : 15'b000000000111111;
													assign node8346 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
							assign node8350 = (inp[9]) ? node8428 : node8351;
								assign node8351 = (inp[2]) ? node8389 : node8352;
									assign node8352 = (inp[14]) ? node8374 : node8353;
										assign node8353 = (inp[6]) ? node8361 : node8354;
											assign node8354 = (inp[12]) ? 15'b000000111111111 : node8355;
												assign node8355 = (inp[7]) ? 15'b000001111111111 : node8356;
													assign node8356 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node8361 = (inp[0]) ? node8369 : node8362;
												assign node8362 = (inp[1]) ? node8366 : node8363;
													assign node8363 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8366 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8369 = (inp[12]) ? 15'b000000000111111 : node8370;
													assign node8370 = (inp[7]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node8374 = (inp[6]) ? node8386 : node8375;
											assign node8375 = (inp[7]) ? node8383 : node8376;
												assign node8376 = (inp[12]) ? node8380 : node8377;
													assign node8377 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8380 = (inp[10]) ? 15'b000000001111111 : 15'b000000001111111;
												assign node8383 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8386 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8389 = (inp[10]) ? node8411 : node8390;
										assign node8390 = (inp[1]) ? node8398 : node8391;
											assign node8391 = (inp[7]) ? node8395 : node8392;
												assign node8392 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node8395 = (inp[0]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node8398 = (inp[14]) ? node8406 : node8399;
												assign node8399 = (inp[0]) ? node8403 : node8400;
													assign node8400 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8403 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8406 = (inp[6]) ? node8408 : 15'b000000001111111;
													assign node8408 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8411 = (inp[6]) ? node8421 : node8412;
											assign node8412 = (inp[12]) ? node8418 : node8413;
												assign node8413 = (inp[0]) ? node8415 : 15'b000000011111111;
													assign node8415 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8418 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node8421 = (inp[1]) ? 15'b000000000011111 : node8422;
												assign node8422 = (inp[12]) ? node8424 : 15'b000000000111111;
													assign node8424 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node8428 = (inp[6]) ? node8460 : node8429;
									assign node8429 = (inp[7]) ? node8447 : node8430;
										assign node8430 = (inp[14]) ? node8440 : node8431;
											assign node8431 = (inp[0]) ? node8435 : node8432;
												assign node8432 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8435 = (inp[2]) ? node8437 : 15'b000000011111111;
													assign node8437 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8440 = (inp[2]) ? node8442 : 15'b000000001111111;
												assign node8442 = (inp[1]) ? node8444 : 15'b000000000111111;
													assign node8444 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8447 = (inp[12]) ? node8453 : node8448;
											assign node8448 = (inp[14]) ? 15'b000000000111111 : node8449;
												assign node8449 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8453 = (inp[0]) ? node8455 : 15'b000000000111111;
												assign node8455 = (inp[2]) ? 15'b000000000001111 : node8456;
													assign node8456 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node8460 = (inp[0]) ? node8484 : node8461;
										assign node8461 = (inp[2]) ? node8473 : node8462;
											assign node8462 = (inp[1]) ? node8468 : node8463;
												assign node8463 = (inp[14]) ? 15'b000000001111111 : node8464;
													assign node8464 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8468 = (inp[10]) ? node8470 : 15'b000000000111111;
													assign node8470 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8473 = (inp[12]) ? node8479 : node8474;
												assign node8474 = (inp[14]) ? node8476 : 15'b000000000111111;
													assign node8476 = (inp[10]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node8479 = (inp[1]) ? 15'b000000000001111 : node8480;
													assign node8480 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8484 = (inp[10]) ? node8494 : node8485;
											assign node8485 = (inp[1]) ? node8489 : node8486;
												assign node8486 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8489 = (inp[7]) ? node8491 : 15'b000000000111111;
													assign node8491 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node8494 = (inp[14]) ? node8500 : node8495;
												assign node8495 = (inp[1]) ? node8497 : 15'b000000000011111;
													assign node8497 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node8500 = (inp[7]) ? node8504 : node8501;
													assign node8501 = (inp[12]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node8504 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node8507 = (inp[8]) ? node8833 : node8508;
						assign node8508 = (inp[9]) ? node8678 : node8509;
							assign node8509 = (inp[14]) ? node8593 : node8510;
								assign node8510 = (inp[7]) ? node8556 : node8511;
									assign node8511 = (inp[13]) ? node8529 : node8512;
										assign node8512 = (inp[1]) ? node8522 : node8513;
											assign node8513 = (inp[0]) ? node8517 : node8514;
												assign node8514 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8517 = (inp[10]) ? node8519 : 15'b000000111111111;
													assign node8519 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8522 = (inp[2]) ? 15'b000000011111111 : node8523;
												assign node8523 = (inp[0]) ? 15'b000000111111111 : node8524;
													assign node8524 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node8529 = (inp[6]) ? node8541 : node8530;
											assign node8530 = (inp[1]) ? node8538 : node8531;
												assign node8531 = (inp[2]) ? node8535 : node8532;
													assign node8532 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8535 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8538 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8541 = (inp[10]) ? node8549 : node8542;
												assign node8542 = (inp[0]) ? node8546 : node8543;
													assign node8543 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8546 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8549 = (inp[0]) ? node8553 : node8550;
													assign node8550 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8553 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8556 = (inp[2]) ? node8576 : node8557;
										assign node8557 = (inp[0]) ? node8567 : node8558;
											assign node8558 = (inp[1]) ? node8564 : node8559;
												assign node8559 = (inp[13]) ? 15'b000000111111111 : node8560;
													assign node8560 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8564 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8567 = (inp[12]) ? node8569 : 15'b000000011111111;
												assign node8569 = (inp[1]) ? node8573 : node8570;
													assign node8570 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8573 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8576 = (inp[6]) ? node8584 : node8577;
											assign node8577 = (inp[0]) ? 15'b000000001111111 : node8578;
												assign node8578 = (inp[13]) ? node8580 : 15'b000000011111111;
													assign node8580 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8584 = (inp[10]) ? node8590 : node8585;
												assign node8585 = (inp[0]) ? node8587 : 15'b000000001111111;
													assign node8587 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8590 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node8593 = (inp[10]) ? node8639 : node8594;
									assign node8594 = (inp[0]) ? node8620 : node8595;
										assign node8595 = (inp[6]) ? node8609 : node8596;
											assign node8596 = (inp[7]) ? node8602 : node8597;
												assign node8597 = (inp[2]) ? node8599 : 15'b000000111111111;
													assign node8599 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8602 = (inp[13]) ? node8606 : node8603;
													assign node8603 = (inp[2]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node8606 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node8609 = (inp[7]) ? node8615 : node8610;
												assign node8610 = (inp[2]) ? node8612 : 15'b000000011111111;
													assign node8612 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8615 = (inp[2]) ? 15'b000000000111111 : node8616;
													assign node8616 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8620 = (inp[1]) ? node8632 : node8621;
											assign node8621 = (inp[12]) ? node8627 : node8622;
												assign node8622 = (inp[6]) ? 15'b000000001111111 : node8623;
													assign node8623 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8627 = (inp[6]) ? node8629 : 15'b000000001111111;
													assign node8629 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node8632 = (inp[2]) ? node8634 : 15'b000000001111111;
												assign node8634 = (inp[6]) ? 15'b000000000111111 : node8635;
													assign node8635 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8639 = (inp[13]) ? node8659 : node8640;
										assign node8640 = (inp[1]) ? node8646 : node8641;
											assign node8641 = (inp[2]) ? node8643 : 15'b000000011111111;
												assign node8643 = (inp[6]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node8646 = (inp[0]) ? node8652 : node8647;
												assign node8647 = (inp[7]) ? node8649 : 15'b000000001111111;
													assign node8649 = (inp[12]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node8652 = (inp[2]) ? node8656 : node8653;
													assign node8653 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8656 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8659 = (inp[0]) ? node8671 : node8660;
											assign node8660 = (inp[2]) ? node8666 : node8661;
												assign node8661 = (inp[1]) ? 15'b000000000111111 : node8662;
													assign node8662 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8666 = (inp[6]) ? node8668 : 15'b000000000111111;
													assign node8668 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8671 = (inp[1]) ? node8673 : 15'b000000000011111;
												assign node8673 = (inp[12]) ? node8675 : 15'b000000000001111;
													assign node8675 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node8678 = (inp[0]) ? node8744 : node8679;
								assign node8679 = (inp[7]) ? node8705 : node8680;
									assign node8680 = (inp[13]) ? node8696 : node8681;
										assign node8681 = (inp[6]) ? node8693 : node8682;
											assign node8682 = (inp[12]) ? node8688 : node8683;
												assign node8683 = (inp[10]) ? 15'b000000111111111 : node8684;
													assign node8684 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8688 = (inp[2]) ? 15'b000000011111111 : node8689;
													assign node8689 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8693 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8696 = (inp[1]) ? node8700 : node8697;
											assign node8697 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8700 = (inp[6]) ? node8702 : 15'b000000001111111;
												assign node8702 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node8705 = (inp[2]) ? node8727 : node8706;
										assign node8706 = (inp[12]) ? node8718 : node8707;
											assign node8707 = (inp[6]) ? node8713 : node8708;
												assign node8708 = (inp[14]) ? node8710 : 15'b000000011111111;
													assign node8710 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8713 = (inp[14]) ? 15'b000000001111111 : node8714;
													assign node8714 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8718 = (inp[1]) ? 15'b000000000111111 : node8719;
												assign node8719 = (inp[13]) ? node8723 : node8720;
													assign node8720 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8723 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node8727 = (inp[14]) ? node8733 : node8728;
											assign node8728 = (inp[13]) ? 15'b000000000111111 : node8729;
												assign node8729 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8733 = (inp[13]) ? node8739 : node8734;
												assign node8734 = (inp[1]) ? 15'b000000000011111 : node8735;
													assign node8735 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8739 = (inp[10]) ? node8741 : 15'b000000000011111;
													assign node8741 = (inp[6]) ? 15'b000000000001111 : 15'b000000000001111;
								assign node8744 = (inp[1]) ? node8780 : node8745;
									assign node8745 = (inp[12]) ? node8761 : node8746;
										assign node8746 = (inp[6]) ? node8754 : node8747;
											assign node8747 = (inp[10]) ? node8749 : 15'b000000011111111;
												assign node8749 = (inp[14]) ? 15'b000000001111111 : node8750;
													assign node8750 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8754 = (inp[14]) ? 15'b000000000111111 : node8755;
												assign node8755 = (inp[7]) ? node8757 : 15'b000000001111111;
													assign node8757 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8761 = (inp[7]) ? node8769 : node8762;
											assign node8762 = (inp[14]) ? node8764 : 15'b000000001111111;
												assign node8764 = (inp[2]) ? node8766 : 15'b000000000111111;
													assign node8766 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8769 = (inp[10]) ? node8775 : node8770;
												assign node8770 = (inp[6]) ? 15'b000000000111111 : node8771;
													assign node8771 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8775 = (inp[13]) ? node8777 : 15'b000000000111111;
													assign node8777 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node8780 = (inp[10]) ? node8808 : node8781;
										assign node8781 = (inp[2]) ? node8793 : node8782;
											assign node8782 = (inp[12]) ? node8788 : node8783;
												assign node8783 = (inp[7]) ? node8785 : 15'b000000001111111;
													assign node8785 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8788 = (inp[14]) ? 15'b000000000111111 : node8789;
													assign node8789 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8793 = (inp[14]) ? node8801 : node8794;
												assign node8794 = (inp[13]) ? node8798 : node8795;
													assign node8795 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8798 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8801 = (inp[7]) ? node8805 : node8802;
													assign node8802 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node8805 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node8808 = (inp[14]) ? node8820 : node8809;
											assign node8809 = (inp[13]) ? node8815 : node8810;
												assign node8810 = (inp[2]) ? node8812 : 15'b000000000111111;
													assign node8812 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8815 = (inp[7]) ? 15'b000000000011111 : node8816;
													assign node8816 = (inp[6]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node8820 = (inp[12]) ? node8828 : node8821;
												assign node8821 = (inp[6]) ? node8825 : node8822;
													assign node8822 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8825 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node8828 = (inp[6]) ? 15'b000000000000111 : node8829;
													assign node8829 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node8833 = (inp[7]) ? node8995 : node8834;
							assign node8834 = (inp[0]) ? node8920 : node8835;
								assign node8835 = (inp[2]) ? node8871 : node8836;
									assign node8836 = (inp[10]) ? node8850 : node8837;
										assign node8837 = (inp[6]) ? node8847 : node8838;
											assign node8838 = (inp[12]) ? 15'b000000011111111 : node8839;
												assign node8839 = (inp[14]) ? node8843 : node8840;
													assign node8840 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8843 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8847 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8850 = (inp[1]) ? node8858 : node8851;
											assign node8851 = (inp[13]) ? 15'b000000001111111 : node8852;
												assign node8852 = (inp[6]) ? 15'b000000011111111 : node8853;
													assign node8853 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8858 = (inp[6]) ? node8866 : node8859;
												assign node8859 = (inp[14]) ? node8863 : node8860;
													assign node8860 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8863 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8866 = (inp[9]) ? node8868 : 15'b000000001111111;
													assign node8868 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node8871 = (inp[12]) ? node8891 : node8872;
										assign node8872 = (inp[13]) ? node8884 : node8873;
											assign node8873 = (inp[10]) ? node8877 : node8874;
												assign node8874 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8877 = (inp[14]) ? node8881 : node8878;
													assign node8878 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8881 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8884 = (inp[9]) ? node8886 : 15'b000000001111111;
												assign node8886 = (inp[6]) ? 15'b000000000111111 : node8887;
													assign node8887 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8891 = (inp[9]) ? node8905 : node8892;
											assign node8892 = (inp[10]) ? node8898 : node8893;
												assign node8893 = (inp[14]) ? 15'b000000001111111 : node8894;
													assign node8894 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8898 = (inp[1]) ? node8902 : node8899;
													assign node8899 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node8902 = (inp[14]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node8905 = (inp[14]) ? node8913 : node8906;
												assign node8906 = (inp[13]) ? node8910 : node8907;
													assign node8907 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8910 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8913 = (inp[13]) ? node8917 : node8914;
													assign node8914 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8917 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node8920 = (inp[14]) ? node8962 : node8921;
									assign node8921 = (inp[6]) ? node8939 : node8922;
										assign node8922 = (inp[9]) ? node8932 : node8923;
											assign node8923 = (inp[1]) ? 15'b000000001111111 : node8924;
												assign node8924 = (inp[2]) ? node8928 : node8925;
													assign node8925 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8928 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8932 = (inp[10]) ? 15'b000000000111111 : node8933;
												assign node8933 = (inp[13]) ? node8935 : 15'b000000001111111;
													assign node8935 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8939 = (inp[9]) ? node8951 : node8940;
											assign node8940 = (inp[10]) ? node8946 : node8941;
												assign node8941 = (inp[13]) ? node8943 : 15'b000000011111111;
													assign node8943 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8946 = (inp[2]) ? 15'b000000000011111 : node8947;
													assign node8947 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node8951 = (inp[13]) ? node8957 : node8952;
												assign node8952 = (inp[1]) ? node8954 : 15'b000000000111111;
													assign node8954 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8957 = (inp[12]) ? 15'b000000000001111 : node8958;
													assign node8958 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node8962 = (inp[2]) ? node8978 : node8963;
										assign node8963 = (inp[6]) ? node8969 : node8964;
											assign node8964 = (inp[13]) ? 15'b000000000111111 : node8965;
												assign node8965 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8969 = (inp[13]) ? node8973 : node8970;
												assign node8970 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8973 = (inp[12]) ? 15'b000000000011111 : node8974;
													assign node8974 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node8978 = (inp[12]) ? node8986 : node8979;
											assign node8979 = (inp[9]) ? 15'b000000000011111 : node8980;
												assign node8980 = (inp[1]) ? node8982 : 15'b000000000111111;
													assign node8982 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8986 = (inp[1]) ? node8988 : 15'b000000000011111;
												assign node8988 = (inp[13]) ? node8992 : node8989;
													assign node8989 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node8992 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node8995 = (inp[1]) ? node9097 : node8996;
								assign node8996 = (inp[9]) ? node9044 : node8997;
									assign node8997 = (inp[14]) ? node9021 : node8998;
										assign node8998 = (inp[0]) ? node9008 : node8999;
											assign node8999 = (inp[12]) ? node9003 : node9000;
												assign node9000 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9003 = (inp[13]) ? node9005 : 15'b000000011111111;
													assign node9005 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9008 = (inp[13]) ? node9016 : node9009;
												assign node9009 = (inp[2]) ? node9013 : node9010;
													assign node9010 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9013 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9016 = (inp[10]) ? 15'b000000000111111 : node9017;
													assign node9017 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node9021 = (inp[6]) ? node9031 : node9022;
											assign node9022 = (inp[12]) ? node9026 : node9023;
												assign node9023 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9026 = (inp[10]) ? node9028 : 15'b000000001111111;
													assign node9028 = (inp[0]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node9031 = (inp[0]) ? node9039 : node9032;
												assign node9032 = (inp[13]) ? node9036 : node9033;
													assign node9033 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node9036 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9039 = (inp[2]) ? 15'b000000000001111 : node9040;
													assign node9040 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node9044 = (inp[10]) ? node9070 : node9045;
										assign node9045 = (inp[2]) ? node9055 : node9046;
											assign node9046 = (inp[6]) ? node9052 : node9047;
												assign node9047 = (inp[13]) ? 15'b000000001111111 : node9048;
													assign node9048 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9052 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9055 = (inp[14]) ? node9063 : node9056;
												assign node9056 = (inp[6]) ? node9060 : node9057;
													assign node9057 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9060 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9063 = (inp[13]) ? node9067 : node9064;
													assign node9064 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9067 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node9070 = (inp[14]) ? node9084 : node9071;
											assign node9071 = (inp[2]) ? node9079 : node9072;
												assign node9072 = (inp[12]) ? node9076 : node9073;
													assign node9073 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9076 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9079 = (inp[0]) ? node9081 : 15'b000000000011111;
													assign node9081 = (inp[13]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node9084 = (inp[0]) ? node9092 : node9085;
												assign node9085 = (inp[6]) ? node9089 : node9086;
													assign node9086 = (inp[12]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node9089 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9092 = (inp[13]) ? 15'b000000000001111 : node9093;
													assign node9093 = (inp[6]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node9097 = (inp[10]) ? node9147 : node9098;
									assign node9098 = (inp[6]) ? node9120 : node9099;
										assign node9099 = (inp[12]) ? node9109 : node9100;
											assign node9100 = (inp[0]) ? node9106 : node9101;
												assign node9101 = (inp[13]) ? node9103 : 15'b000000011111111;
													assign node9103 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9106 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9109 = (inp[14]) ? node9115 : node9110;
												assign node9110 = (inp[9]) ? node9112 : 15'b000000001111111;
													assign node9112 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9115 = (inp[2]) ? node9117 : 15'b000000000011111;
													assign node9117 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
										assign node9120 = (inp[2]) ? node9132 : node9121;
											assign node9121 = (inp[13]) ? node9125 : node9122;
												assign node9122 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9125 = (inp[9]) ? node9129 : node9126;
													assign node9126 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9129 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node9132 = (inp[0]) ? node9140 : node9133;
												assign node9133 = (inp[14]) ? node9137 : node9134;
													assign node9134 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node9137 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9140 = (inp[14]) ? node9144 : node9141;
													assign node9141 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node9144 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node9147 = (inp[2]) ? node9169 : node9148;
										assign node9148 = (inp[6]) ? node9158 : node9149;
											assign node9149 = (inp[14]) ? node9153 : node9150;
												assign node9150 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node9153 = (inp[0]) ? node9155 : 15'b000000000011111;
													assign node9155 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node9158 = (inp[13]) ? node9164 : node9159;
												assign node9159 = (inp[0]) ? node9161 : 15'b000000000011111;
													assign node9161 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9164 = (inp[9]) ? 15'b000000000001111 : node9165;
													assign node9165 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node9169 = (inp[9]) ? node9185 : node9170;
											assign node9170 = (inp[12]) ? node9178 : node9171;
												assign node9171 = (inp[6]) ? node9175 : node9172;
													assign node9172 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9175 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9178 = (inp[0]) ? node9182 : node9179;
													assign node9179 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node9182 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node9185 = (inp[13]) ? node9191 : node9186;
												assign node9186 = (inp[6]) ? 15'b000000000001111 : node9187;
													assign node9187 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9191 = (inp[6]) ? node9193 : 15'b000000000000111;
													assign node9193 = (inp[12]) ? 15'b000000000000011 : 15'b000000000000111;
				assign node9196 = (inp[2]) ? node9866 : node9197;
					assign node9197 = (inp[7]) ? node9527 : node9198;
						assign node9198 = (inp[1]) ? node9384 : node9199;
							assign node9199 = (inp[10]) ? node9293 : node9200;
								assign node9200 = (inp[0]) ? node9244 : node9201;
									assign node9201 = (inp[12]) ? node9227 : node9202;
										assign node9202 = (inp[8]) ? node9214 : node9203;
											assign node9203 = (inp[13]) ? node9209 : node9204;
												assign node9204 = (inp[5]) ? 15'b000001111111111 : node9205;
													assign node9205 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9209 = (inp[5]) ? 15'b000000111111111 : node9210;
													assign node9210 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node9214 = (inp[13]) ? node9222 : node9215;
												assign node9215 = (inp[9]) ? node9219 : node9216;
													assign node9216 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9219 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9222 = (inp[6]) ? node9224 : 15'b000000111111111;
													assign node9224 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9227 = (inp[8]) ? node9233 : node9228;
											assign node9228 = (inp[9]) ? node9230 : 15'b000001111111111;
												assign node9230 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node9233 = (inp[9]) ? node9239 : node9234;
												assign node9234 = (inp[13]) ? node9236 : 15'b000000011111111;
													assign node9236 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9239 = (inp[13]) ? 15'b000000000111111 : node9240;
													assign node9240 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node9244 = (inp[8]) ? node9270 : node9245;
										assign node9245 = (inp[5]) ? node9261 : node9246;
											assign node9246 = (inp[13]) ? node9254 : node9247;
												assign node9247 = (inp[9]) ? node9251 : node9248;
													assign node9248 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9251 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9254 = (inp[9]) ? node9258 : node9255;
													assign node9255 = (inp[12]) ? 15'b000000011111111 : 15'b000000011111111;
													assign node9258 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9261 = (inp[9]) ? 15'b000000001111111 : node9262;
												assign node9262 = (inp[14]) ? node9266 : node9263;
													assign node9263 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9266 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node9270 = (inp[14]) ? node9282 : node9271;
											assign node9271 = (inp[5]) ? node9277 : node9272;
												assign node9272 = (inp[6]) ? node9274 : 15'b000000011111111;
													assign node9274 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9277 = (inp[6]) ? node9279 : 15'b000000001111111;
													assign node9279 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9282 = (inp[6]) ? node9290 : node9283;
												assign node9283 = (inp[5]) ? node9287 : node9284;
													assign node9284 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9287 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9290 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9293 = (inp[9]) ? node9333 : node9294;
									assign node9294 = (inp[8]) ? node9314 : node9295;
										assign node9295 = (inp[0]) ? node9303 : node9296;
											assign node9296 = (inp[14]) ? 15'b000000011111111 : node9297;
												assign node9297 = (inp[13]) ? node9299 : 15'b000001111111111;
													assign node9299 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9303 = (inp[12]) ? node9309 : node9304;
												assign node9304 = (inp[13]) ? node9306 : 15'b000000011111111;
													assign node9306 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9309 = (inp[5]) ? 15'b000000001111111 : node9310;
													assign node9310 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9314 = (inp[12]) ? node9322 : node9315;
											assign node9315 = (inp[5]) ? node9317 : 15'b000000011111111;
												assign node9317 = (inp[14]) ? 15'b000000001111111 : node9318;
													assign node9318 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9322 = (inp[0]) ? node9328 : node9323;
												assign node9323 = (inp[13]) ? 15'b000000001111111 : node9324;
													assign node9324 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9328 = (inp[13]) ? node9330 : 15'b000000000111111;
													assign node9330 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9333 = (inp[5]) ? node9361 : node9334;
										assign node9334 = (inp[13]) ? node9346 : node9335;
											assign node9335 = (inp[8]) ? node9339 : node9336;
												assign node9336 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9339 = (inp[12]) ? node9343 : node9340;
													assign node9340 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9343 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9346 = (inp[12]) ? node9354 : node9347;
												assign node9347 = (inp[0]) ? node9351 : node9348;
													assign node9348 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node9351 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9354 = (inp[14]) ? node9358 : node9355;
													assign node9355 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9358 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9361 = (inp[14]) ? node9371 : node9362;
											assign node9362 = (inp[6]) ? node9366 : node9363;
												assign node9363 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9366 = (inp[13]) ? 15'b000000000011111 : node9367;
													assign node9367 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9371 = (inp[8]) ? node9377 : node9372;
												assign node9372 = (inp[0]) ? node9374 : 15'b000000000111111;
													assign node9374 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9377 = (inp[0]) ? node9381 : node9378;
													assign node9378 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9381 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node9384 = (inp[0]) ? node9450 : node9385;
								assign node9385 = (inp[14]) ? node9415 : node9386;
									assign node9386 = (inp[9]) ? node9402 : node9387;
										assign node9387 = (inp[12]) ? node9395 : node9388;
											assign node9388 = (inp[13]) ? node9390 : 15'b000001111111111;
												assign node9390 = (inp[5]) ? 15'b000000001111111 : node9391;
													assign node9391 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9395 = (inp[8]) ? node9397 : 15'b000000011111111;
												assign node9397 = (inp[6]) ? 15'b000000001111111 : node9398;
													assign node9398 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9402 = (inp[12]) ? node9410 : node9403;
											assign node9403 = (inp[5]) ? 15'b000000001111111 : node9404;
												assign node9404 = (inp[6]) ? 15'b000000011111111 : node9405;
													assign node9405 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9410 = (inp[8]) ? 15'b000000000111111 : node9411;
												assign node9411 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9415 = (inp[10]) ? node9429 : node9416;
										assign node9416 = (inp[13]) ? node9424 : node9417;
											assign node9417 = (inp[12]) ? 15'b000000001111111 : node9418;
												assign node9418 = (inp[8]) ? node9420 : 15'b000000011111111;
													assign node9420 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9424 = (inp[6]) ? node9426 : 15'b000000001111111;
												assign node9426 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9429 = (inp[9]) ? node9443 : node9430;
											assign node9430 = (inp[13]) ? node9436 : node9431;
												assign node9431 = (inp[6]) ? node9433 : 15'b000000001111111;
													assign node9433 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9436 = (inp[8]) ? node9440 : node9437;
													assign node9437 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9440 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9443 = (inp[6]) ? node9445 : 15'b000000000111111;
												assign node9445 = (inp[5]) ? 15'b000000000001111 : node9446;
													assign node9446 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9450 = (inp[14]) ? node9496 : node9451;
									assign node9451 = (inp[5]) ? node9475 : node9452;
										assign node9452 = (inp[9]) ? node9462 : node9453;
											assign node9453 = (inp[6]) ? node9459 : node9454;
												assign node9454 = (inp[8]) ? 15'b000000011111111 : node9455;
													assign node9455 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9459 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9462 = (inp[8]) ? node9468 : node9463;
												assign node9463 = (inp[13]) ? 15'b000000001111111 : node9464;
													assign node9464 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9468 = (inp[6]) ? node9472 : node9469;
													assign node9469 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9472 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9475 = (inp[12]) ? node9485 : node9476;
											assign node9476 = (inp[6]) ? node9480 : node9477;
												assign node9477 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9480 = (inp[10]) ? node9482 : 15'b000000000111111;
													assign node9482 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9485 = (inp[8]) ? node9491 : node9486;
												assign node9486 = (inp[6]) ? node9488 : 15'b000000011111111;
													assign node9488 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9491 = (inp[9]) ? node9493 : 15'b000000000011111;
													assign node9493 = (inp[10]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node9496 = (inp[8]) ? node9506 : node9497;
										assign node9497 = (inp[5]) ? node9501 : node9498;
											assign node9498 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9501 = (inp[6]) ? 15'b000000000011111 : node9502;
												assign node9502 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9506 = (inp[6]) ? node9514 : node9507;
											assign node9507 = (inp[10]) ? 15'b000000000011111 : node9508;
												assign node9508 = (inp[5]) ? node9510 : 15'b000000000111111;
													assign node9510 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node9514 = (inp[13]) ? node9520 : node9515;
												assign node9515 = (inp[10]) ? 15'b000000000011111 : node9516;
													assign node9516 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9520 = (inp[10]) ? node9524 : node9521;
													assign node9521 = (inp[9]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node9524 = (inp[9]) ? 15'b000000000000111 : 15'b000000000000111;
						assign node9527 = (inp[13]) ? node9681 : node9528;
							assign node9528 = (inp[10]) ? node9598 : node9529;
								assign node9529 = (inp[1]) ? node9567 : node9530;
									assign node9530 = (inp[0]) ? node9552 : node9531;
										assign node9531 = (inp[8]) ? node9541 : node9532;
											assign node9532 = (inp[12]) ? node9538 : node9533;
												assign node9533 = (inp[14]) ? 15'b000000111111111 : node9534;
													assign node9534 = (inp[6]) ? 15'b000001111111111 : 15'b000001111111111;
												assign node9538 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9541 = (inp[6]) ? node9547 : node9542;
												assign node9542 = (inp[12]) ? node9544 : 15'b000000111111111;
													assign node9544 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9547 = (inp[14]) ? 15'b000000001111111 : node9548;
													assign node9548 = (inp[9]) ? 15'b000000001111111 : 15'b000000001111111;
										assign node9552 = (inp[5]) ? node9560 : node9553;
											assign node9553 = (inp[9]) ? node9555 : 15'b000000011111111;
												assign node9555 = (inp[12]) ? 15'b000000001111111 : node9556;
													assign node9556 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9560 = (inp[8]) ? node9564 : node9561;
												assign node9561 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9564 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9567 = (inp[8]) ? node9581 : node9568;
										assign node9568 = (inp[0]) ? node9576 : node9569;
											assign node9569 = (inp[12]) ? node9571 : 15'b000000001111111;
												assign node9571 = (inp[14]) ? 15'b000000011111111 : node9572;
													assign node9572 = (inp[6]) ? 15'b000000011111111 : 15'b000000011111111;
											assign node9576 = (inp[5]) ? 15'b000000000111111 : node9577;
												assign node9577 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9581 = (inp[6]) ? node9589 : node9582;
											assign node9582 = (inp[9]) ? node9584 : 15'b000000011111111;
												assign node9584 = (inp[14]) ? node9586 : 15'b000000001111111;
													assign node9586 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9589 = (inp[9]) ? node9595 : node9590;
												assign node9590 = (inp[12]) ? node9592 : 15'b000000000111111;
													assign node9592 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9595 = (inp[12]) ? 15'b000000000011111 : 15'b000000000001111;
								assign node9598 = (inp[14]) ? node9642 : node9599;
									assign node9599 = (inp[0]) ? node9619 : node9600;
										assign node9600 = (inp[6]) ? node9610 : node9601;
											assign node9601 = (inp[9]) ? node9607 : node9602;
												assign node9602 = (inp[5]) ? node9604 : 15'b000000111111111;
													assign node9604 = (inp[12]) ? 15'b000000011111111 : 15'b000000011111111;
												assign node9607 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9610 = (inp[8]) ? node9614 : node9611;
												assign node9611 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9614 = (inp[12]) ? node9616 : 15'b000000000111111;
													assign node9616 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9619 = (inp[12]) ? node9631 : node9620;
											assign node9620 = (inp[9]) ? node9626 : node9621;
												assign node9621 = (inp[1]) ? node9623 : 15'b000000001111111;
													assign node9623 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9626 = (inp[1]) ? node9628 : 15'b000000000111111;
													assign node9628 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9631 = (inp[6]) ? node9637 : node9632;
												assign node9632 = (inp[1]) ? node9634 : 15'b000000000111111;
													assign node9634 = (inp[9]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node9637 = (inp[5]) ? node9639 : 15'b000000000011111;
													assign node9639 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node9642 = (inp[8]) ? node9658 : node9643;
										assign node9643 = (inp[9]) ? node9647 : node9644;
											assign node9644 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9647 = (inp[6]) ? node9653 : node9648;
												assign node9648 = (inp[12]) ? node9650 : 15'b000000000111111;
													assign node9650 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9653 = (inp[0]) ? 15'b000000000011111 : node9654;
													assign node9654 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9658 = (inp[6]) ? node9668 : node9659;
											assign node9659 = (inp[9]) ? node9663 : node9660;
												assign node9660 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node9663 = (inp[12]) ? node9665 : 15'b000000000011111;
													assign node9665 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node9668 = (inp[1]) ? node9676 : node9669;
												assign node9669 = (inp[9]) ? node9673 : node9670;
													assign node9670 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9673 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9676 = (inp[5]) ? 15'b000000000001111 : node9677;
													assign node9677 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node9681 = (inp[9]) ? node9773 : node9682;
								assign node9682 = (inp[6]) ? node9724 : node9683;
									assign node9683 = (inp[14]) ? node9703 : node9684;
										assign node9684 = (inp[1]) ? node9690 : node9685;
											assign node9685 = (inp[10]) ? node9687 : 15'b000000011111111;
												assign node9687 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9690 = (inp[0]) ? node9696 : node9691;
												assign node9691 = (inp[8]) ? 15'b000000001111111 : node9692;
													assign node9692 = (inp[12]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node9696 = (inp[12]) ? node9700 : node9697;
													assign node9697 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9700 = (inp[10]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node9703 = (inp[5]) ? node9713 : node9704;
											assign node9704 = (inp[1]) ? node9706 : 15'b000000011111111;
												assign node9706 = (inp[10]) ? node9710 : node9707;
													assign node9707 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9710 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9713 = (inp[0]) ? node9719 : node9714;
												assign node9714 = (inp[1]) ? node9716 : 15'b000000000111111;
													assign node9716 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9719 = (inp[12]) ? node9721 : 15'b000000001111111;
													assign node9721 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node9724 = (inp[12]) ? node9754 : node9725;
										assign node9725 = (inp[1]) ? node9739 : node9726;
											assign node9726 = (inp[14]) ? node9734 : node9727;
												assign node9727 = (inp[0]) ? node9731 : node9728;
													assign node9728 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9731 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node9734 = (inp[8]) ? node9736 : 15'b000000000111111;
													assign node9736 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9739 = (inp[5]) ? node9747 : node9740;
												assign node9740 = (inp[10]) ? node9744 : node9741;
													assign node9741 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9744 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9747 = (inp[8]) ? node9751 : node9748;
													assign node9748 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
													assign node9751 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node9754 = (inp[0]) ? node9760 : node9755;
											assign node9755 = (inp[14]) ? 15'b000000000011111 : node9756;
												assign node9756 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node9760 = (inp[8]) ? node9766 : node9761;
												assign node9761 = (inp[10]) ? 15'b000000000011111 : node9762;
													assign node9762 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9766 = (inp[5]) ? node9770 : node9767;
													assign node9767 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node9770 = (inp[1]) ? 15'b000000000000011 : 15'b000000000001111;
								assign node9773 = (inp[14]) ? node9815 : node9774;
									assign node9774 = (inp[5]) ? node9794 : node9775;
										assign node9775 = (inp[12]) ? node9785 : node9776;
											assign node9776 = (inp[0]) ? node9780 : node9777;
												assign node9777 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9780 = (inp[6]) ? 15'b000000000011111 : node9781;
													assign node9781 = (inp[10]) ? 15'b000000000111111 : 15'b000000000111111;
											assign node9785 = (inp[10]) ? node9787 : 15'b000000000111111;
												assign node9787 = (inp[0]) ? node9791 : node9788;
													assign node9788 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9791 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node9794 = (inp[0]) ? node9802 : node9795;
											assign node9795 = (inp[10]) ? 15'b000000000011111 : node9796;
												assign node9796 = (inp[1]) ? node9798 : 15'b000000000111111;
													assign node9798 = (inp[8]) ? 15'b000000000011111 : 15'b000000000011111;
											assign node9802 = (inp[1]) ? node9808 : node9803;
												assign node9803 = (inp[12]) ? 15'b000000000011111 : node9804;
													assign node9804 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node9808 = (inp[6]) ? node9812 : node9809;
													assign node9809 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node9812 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node9815 = (inp[6]) ? node9843 : node9816;
										assign node9816 = (inp[0]) ? node9830 : node9817;
											assign node9817 = (inp[5]) ? node9825 : node9818;
												assign node9818 = (inp[1]) ? node9822 : node9819;
													assign node9819 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9822 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node9825 = (inp[10]) ? 15'b000000000011111 : node9826;
													assign node9826 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9830 = (inp[8]) ? node9836 : node9831;
												assign node9831 = (inp[12]) ? node9833 : 15'b000000001111111;
													assign node9833 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9836 = (inp[1]) ? node9840 : node9837;
													assign node9837 = (inp[12]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node9840 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node9843 = (inp[10]) ? node9857 : node9844;
											assign node9844 = (inp[12]) ? node9850 : node9845;
												assign node9845 = (inp[1]) ? node9847 : 15'b000000000011111;
													assign node9847 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node9850 = (inp[1]) ? node9854 : node9851;
													assign node9851 = (inp[0]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node9854 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node9857 = (inp[5]) ? node9859 : 15'b000000000001111;
												assign node9859 = (inp[8]) ? node9863 : node9860;
													assign node9860 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node9863 = (inp[1]) ? 15'b000000000000011 : 15'b000000000000111;
					assign node9866 = (inp[9]) ? node10212 : node9867;
						assign node9867 = (inp[13]) ? node10031 : node9868;
							assign node9868 = (inp[1]) ? node9940 : node9869;
								assign node9869 = (inp[14]) ? node9911 : node9870;
									assign node9870 = (inp[6]) ? node9890 : node9871;
										assign node9871 = (inp[12]) ? node9879 : node9872;
											assign node9872 = (inp[7]) ? node9876 : node9873;
												assign node9873 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9876 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9879 = (inp[7]) ? node9885 : node9880;
												assign node9880 = (inp[8]) ? 15'b000000011111111 : node9881;
													assign node9881 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9885 = (inp[10]) ? node9887 : 15'b000000011111111;
													assign node9887 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9890 = (inp[0]) ? node9904 : node9891;
											assign node9891 = (inp[5]) ? node9897 : node9892;
												assign node9892 = (inp[8]) ? node9894 : 15'b000000011111111;
													assign node9894 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9897 = (inp[7]) ? node9901 : node9898;
													assign node9898 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9901 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9904 = (inp[8]) ? node9906 : 15'b000000001111111;
												assign node9906 = (inp[7]) ? 15'b000000000111111 : node9907;
													assign node9907 = (inp[10]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node9911 = (inp[10]) ? node9921 : node9912;
										assign node9912 = (inp[12]) ? node9916 : node9913;
											assign node9913 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9916 = (inp[7]) ? 15'b000000000111111 : node9917;
												assign node9917 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9921 = (inp[5]) ? node9931 : node9922;
											assign node9922 = (inp[6]) ? node9928 : node9923;
												assign node9923 = (inp[12]) ? node9925 : 15'b000000001111111;
													assign node9925 = (inp[8]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node9928 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9931 = (inp[0]) ? node9935 : node9932;
												assign node9932 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9935 = (inp[6]) ? node9937 : 15'b000000000011111;
													assign node9937 = (inp[7]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node9940 = (inp[8]) ? node9984 : node9941;
									assign node9941 = (inp[5]) ? node9965 : node9942;
										assign node9942 = (inp[10]) ? node9954 : node9943;
											assign node9943 = (inp[0]) ? node9947 : node9944;
												assign node9944 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9947 = (inp[12]) ? node9951 : node9948;
													assign node9948 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9951 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9954 = (inp[6]) ? node9958 : node9955;
												assign node9955 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9958 = (inp[7]) ? node9962 : node9959;
													assign node9959 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9962 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9965 = (inp[0]) ? node9977 : node9966;
											assign node9966 = (inp[12]) ? node9972 : node9967;
												assign node9967 = (inp[14]) ? node9969 : 15'b000000001111111;
													assign node9969 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node9972 = (inp[7]) ? 15'b000000000111111 : node9973;
													assign node9973 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9977 = (inp[12]) ? 15'b000000000011111 : node9978;
												assign node9978 = (inp[7]) ? 15'b000000000111111 : node9979;
													assign node9979 = (inp[6]) ? 15'b000000001111111 : 15'b000000000111111;
									assign node9984 = (inp[6]) ? node10008 : node9985;
										assign node9985 = (inp[14]) ? node9997 : node9986;
											assign node9986 = (inp[5]) ? node9992 : node9987;
												assign node9987 = (inp[0]) ? node9989 : 15'b000000011111111;
													assign node9989 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9992 = (inp[0]) ? 15'b000000000011111 : node9993;
													assign node9993 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9997 = (inp[0]) ? node10003 : node9998;
												assign node9998 = (inp[10]) ? node10000 : 15'b000000001111111;
													assign node10000 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10003 = (inp[10]) ? 15'b000000000001111 : node10004;
													assign node10004 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10008 = (inp[0]) ? node10020 : node10009;
											assign node10009 = (inp[5]) ? node10015 : node10010;
												assign node10010 = (inp[12]) ? 15'b000000000011111 : node10011;
													assign node10011 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10015 = (inp[7]) ? node10017 : 15'b000000000011111;
													assign node10017 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10020 = (inp[5]) ? node10026 : node10021;
												assign node10021 = (inp[12]) ? node10023 : 15'b000000000011111;
													assign node10023 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10026 = (inp[7]) ? node10028 : 15'b000000000011111;
													assign node10028 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node10031 = (inp[6]) ? node10129 : node10032;
								assign node10032 = (inp[12]) ? node10074 : node10033;
									assign node10033 = (inp[10]) ? node10055 : node10034;
										assign node10034 = (inp[1]) ? node10046 : node10035;
											assign node10035 = (inp[0]) ? node10041 : node10036;
												assign node10036 = (inp[5]) ? 15'b000000001111111 : node10037;
													assign node10037 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10041 = (inp[7]) ? node10043 : 15'b000000011111111;
													assign node10043 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10046 = (inp[0]) ? 15'b000000000011111 : node10047;
												assign node10047 = (inp[5]) ? node10051 : node10048;
													assign node10048 = (inp[8]) ? 15'b000000001111111 : 15'b000000001111111;
													assign node10051 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10055 = (inp[7]) ? node10063 : node10056;
											assign node10056 = (inp[1]) ? node10058 : 15'b000000001111111;
												assign node10058 = (inp[14]) ? 15'b000000000111111 : node10059;
													assign node10059 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10063 = (inp[0]) ? node10069 : node10064;
												assign node10064 = (inp[5]) ? 15'b000000000111111 : node10065;
													assign node10065 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10069 = (inp[8]) ? node10071 : 15'b000000000011111;
													assign node10071 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node10074 = (inp[0]) ? node10102 : node10075;
										assign node10075 = (inp[14]) ? node10087 : node10076;
											assign node10076 = (inp[8]) ? node10082 : node10077;
												assign node10077 = (inp[10]) ? node10079 : 15'b000000011111111;
													assign node10079 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10082 = (inp[1]) ? node10084 : 15'b000000000111111;
													assign node10084 = (inp[7]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node10087 = (inp[7]) ? node10095 : node10088;
												assign node10088 = (inp[8]) ? node10092 : node10089;
													assign node10089 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10092 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10095 = (inp[10]) ? node10099 : node10096;
													assign node10096 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10099 = (inp[5]) ? 15'b000000000001111 : 15'b000000000001111;
										assign node10102 = (inp[10]) ? node10114 : node10103;
											assign node10103 = (inp[1]) ? node10109 : node10104;
												assign node10104 = (inp[7]) ? node10106 : 15'b000000000111111;
													assign node10106 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10109 = (inp[5]) ? 15'b000000000011111 : node10110;
													assign node10110 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10114 = (inp[5]) ? node10122 : node10115;
												assign node10115 = (inp[7]) ? node10119 : node10116;
													assign node10116 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10119 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10122 = (inp[14]) ? node10126 : node10123;
													assign node10123 = (inp[7]) ? 15'b000000000011111 : 15'b000000000001111;
													assign node10126 = (inp[7]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node10129 = (inp[14]) ? node10173 : node10130;
									assign node10130 = (inp[5]) ? node10152 : node10131;
										assign node10131 = (inp[7]) ? node10141 : node10132;
											assign node10132 = (inp[0]) ? node10136 : node10133;
												assign node10133 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10136 = (inp[1]) ? node10138 : 15'b000000000111111;
													assign node10138 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10141 = (inp[10]) ? node10147 : node10142;
												assign node10142 = (inp[0]) ? node10144 : 15'b000000000111111;
													assign node10144 = (inp[1]) ? 15'b000000000011111 : 15'b000000000011111;
												assign node10147 = (inp[0]) ? 15'b000000000011111 : node10148;
													assign node10148 = (inp[1]) ? 15'b000000000011111 : 15'b000000000011111;
										assign node10152 = (inp[10]) ? node10164 : node10153;
											assign node10153 = (inp[7]) ? node10159 : node10154;
												assign node10154 = (inp[1]) ? 15'b000000000111111 : node10155;
													assign node10155 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10159 = (inp[8]) ? 15'b000000000000111 : node10160;
													assign node10160 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10164 = (inp[8]) ? node10168 : node10165;
												assign node10165 = (inp[7]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10168 = (inp[12]) ? node10170 : 15'b000000000001111;
													assign node10170 = (inp[1]) ? 15'b000000000000011 : 15'b000000000000111;
									assign node10173 = (inp[7]) ? node10193 : node10174;
										assign node10174 = (inp[8]) ? node10184 : node10175;
											assign node10175 = (inp[12]) ? 15'b000000000011111 : node10176;
												assign node10176 = (inp[1]) ? node10180 : node10177;
													assign node10177 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10180 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10184 = (inp[12]) ? node10190 : node10185;
												assign node10185 = (inp[5]) ? node10187 : 15'b000000000011111;
													assign node10187 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10190 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node10193 = (inp[10]) ? node10205 : node10194;
											assign node10194 = (inp[0]) ? node10200 : node10195;
												assign node10195 = (inp[8]) ? node10197 : 15'b000000000011111;
													assign node10197 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10200 = (inp[1]) ? node10202 : 15'b000000000001111;
													assign node10202 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node10205 = (inp[5]) ? node10207 : 15'b000000000001111;
												assign node10207 = (inp[1]) ? node10209 : 15'b000000000000111;
													assign node10209 = (inp[0]) ? 15'b000000000000011 : 15'b000000000000111;
						assign node10212 = (inp[8]) ? node10378 : node10213;
							assign node10213 = (inp[6]) ? node10291 : node10214;
								assign node10214 = (inp[5]) ? node10250 : node10215;
									assign node10215 = (inp[13]) ? node10235 : node10216;
										assign node10216 = (inp[0]) ? node10226 : node10217;
											assign node10217 = (inp[10]) ? node10221 : node10218;
												assign node10218 = (inp[14]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node10221 = (inp[14]) ? 15'b000000000111111 : node10222;
													assign node10222 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10226 = (inp[7]) ? node10228 : 15'b000000001111111;
												assign node10228 = (inp[10]) ? node10232 : node10229;
													assign node10229 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10232 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10235 = (inp[12]) ? node10243 : node10236;
											assign node10236 = (inp[7]) ? node10240 : node10237;
												assign node10237 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10240 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10243 = (inp[14]) ? node10245 : 15'b000000000111111;
												assign node10245 = (inp[10]) ? 15'b000000000011111 : node10246;
													assign node10246 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10250 = (inp[12]) ? node10274 : node10251;
										assign node10251 = (inp[10]) ? node10263 : node10252;
											assign node10252 = (inp[0]) ? node10258 : node10253;
												assign node10253 = (inp[13]) ? node10255 : 15'b000000001111111;
													assign node10255 = (inp[14]) ? 15'b000000000111111 : 15'b000000000111111;
												assign node10258 = (inp[14]) ? 15'b000000000111111 : node10259;
													assign node10259 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10263 = (inp[7]) ? node10267 : node10264;
												assign node10264 = (inp[0]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node10267 = (inp[14]) ? node10271 : node10268;
													assign node10268 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10271 = (inp[13]) ? 15'b000000000011111 : 15'b000000000001111;
										assign node10274 = (inp[0]) ? node10282 : node10275;
											assign node10275 = (inp[13]) ? node10277 : 15'b000000000111111;
												assign node10277 = (inp[14]) ? 15'b000000000011111 : node10278;
													assign node10278 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10282 = (inp[14]) ? node10288 : node10283;
												assign node10283 = (inp[10]) ? 15'b000000000001111 : node10284;
													assign node10284 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10288 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node10291 = (inp[5]) ? node10337 : node10292;
									assign node10292 = (inp[0]) ? node10320 : node10293;
										assign node10293 = (inp[7]) ? node10305 : node10294;
											assign node10294 = (inp[13]) ? node10300 : node10295;
												assign node10295 = (inp[10]) ? 15'b000000001111111 : node10296;
													assign node10296 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10300 = (inp[14]) ? 15'b000000000111111 : node10301;
													assign node10301 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10305 = (inp[13]) ? node10313 : node10306;
												assign node10306 = (inp[12]) ? node10310 : node10307;
													assign node10307 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10310 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10313 = (inp[12]) ? node10317 : node10314;
													assign node10314 = (inp[10]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node10317 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node10320 = (inp[10]) ? node10332 : node10321;
											assign node10321 = (inp[13]) ? node10327 : node10322;
												assign node10322 = (inp[7]) ? 15'b000000000111111 : node10323;
													assign node10323 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10327 = (inp[1]) ? node10329 : 15'b000000000011111;
													assign node10329 = (inp[7]) ? 15'b000000000001111 : 15'b000000000001111;
											assign node10332 = (inp[14]) ? 15'b000000000000111 : node10333;
												assign node10333 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node10337 = (inp[7]) ? node10359 : node10338;
										assign node10338 = (inp[13]) ? node10350 : node10339;
											assign node10339 = (inp[12]) ? node10345 : node10340;
												assign node10340 = (inp[10]) ? 15'b000000000011111 : node10341;
													assign node10341 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node10345 = (inp[0]) ? 15'b000000000001111 : node10346;
													assign node10346 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10350 = (inp[12]) ? node10356 : node10351;
												assign node10351 = (inp[10]) ? node10353 : 15'b000000000011111;
													assign node10353 = (inp[1]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node10356 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node10359 = (inp[0]) ? node10365 : node10360;
											assign node10360 = (inp[14]) ? 15'b000000000001111 : node10361;
												assign node10361 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10365 = (inp[14]) ? node10371 : node10366;
												assign node10366 = (inp[12]) ? node10368 : 15'b000000000001111;
													assign node10368 = (inp[1]) ? 15'b000000000000111 : 15'b000000000000111;
												assign node10371 = (inp[10]) ? node10375 : node10372;
													assign node10372 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node10375 = (inp[12]) ? 15'b000000000000001 : 15'b000000000000111;
							assign node10378 = (inp[7]) ? node10462 : node10379;
								assign node10379 = (inp[1]) ? node10419 : node10380;
									assign node10380 = (inp[10]) ? node10394 : node10381;
										assign node10381 = (inp[0]) ? node10389 : node10382;
											assign node10382 = (inp[6]) ? node10384 : 15'b000000001111111;
												assign node10384 = (inp[14]) ? 15'b000000000111111 : node10385;
													assign node10385 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10389 = (inp[14]) ? node10391 : 15'b000000000111111;
												assign node10391 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10394 = (inp[13]) ? node10410 : node10395;
											assign node10395 = (inp[5]) ? node10403 : node10396;
												assign node10396 = (inp[0]) ? node10400 : node10397;
													assign node10397 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10400 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10403 = (inp[0]) ? node10407 : node10404;
													assign node10404 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10407 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10410 = (inp[14]) ? node10414 : node10411;
												assign node10411 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10414 = (inp[12]) ? node10416 : 15'b000000000001111;
													assign node10416 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node10419 = (inp[0]) ? node10445 : node10420;
										assign node10420 = (inp[14]) ? node10430 : node10421;
											assign node10421 = (inp[10]) ? node10425 : node10422;
												assign node10422 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10425 = (inp[6]) ? node10427 : 15'b000000000011111;
													assign node10427 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10430 = (inp[5]) ? node10438 : node10431;
												assign node10431 = (inp[12]) ? node10435 : node10432;
													assign node10432 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10435 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10438 = (inp[6]) ? node10442 : node10439;
													assign node10439 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node10442 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node10445 = (inp[13]) ? node10457 : node10446;
											assign node10446 = (inp[10]) ? node10452 : node10447;
												assign node10447 = (inp[5]) ? 15'b000000000011111 : node10448;
													assign node10448 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10452 = (inp[12]) ? 15'b000000000000111 : node10453;
													assign node10453 = (inp[5]) ? 15'b000000000000111 : 15'b000000000011111;
											assign node10457 = (inp[12]) ? 15'b000000000000111 : node10458;
												assign node10458 = (inp[14]) ? 15'b000000000000011 : 15'b000000000001111;
								assign node10462 = (inp[12]) ? node10506 : node10463;
									assign node10463 = (inp[13]) ? node10485 : node10464;
										assign node10464 = (inp[5]) ? node10474 : node10465;
											assign node10465 = (inp[6]) ? 15'b000000000011111 : node10466;
												assign node10466 = (inp[14]) ? node10470 : node10467;
													assign node10467 = (inp[1]) ? 15'b000000000111111 : 15'b000000000111111;
													assign node10470 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10474 = (inp[0]) ? node10480 : node10475;
												assign node10475 = (inp[10]) ? node10477 : 15'b000000000011111;
													assign node10477 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10480 = (inp[14]) ? node10482 : 15'b000000000011111;
													assign node10482 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node10485 = (inp[10]) ? node10499 : node10486;
											assign node10486 = (inp[1]) ? node10492 : node10487;
												assign node10487 = (inp[14]) ? node10489 : 15'b000000000111111;
													assign node10489 = (inp[6]) ? 15'b000000000001111 : 15'b000000000001111;
												assign node10492 = (inp[0]) ? node10496 : node10493;
													assign node10493 = (inp[6]) ? 15'b000000000001111 : 15'b000000000001111;
													assign node10496 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node10499 = (inp[6]) ? node10501 : 15'b000000000000111;
												assign node10501 = (inp[1]) ? 15'b000000000000111 : node10502;
													assign node10502 = (inp[5]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node10506 = (inp[1]) ? node10526 : node10507;
										assign node10507 = (inp[0]) ? node10517 : node10508;
											assign node10508 = (inp[10]) ? node10512 : node10509;
												assign node10509 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10512 = (inp[13]) ? 15'b000000000001111 : node10513;
													assign node10513 = (inp[6]) ? 15'b000000000011111 : 15'b000000000001111;
											assign node10517 = (inp[5]) ? 15'b000000000000111 : node10518;
												assign node10518 = (inp[13]) ? node10522 : node10519;
													assign node10519 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node10522 = (inp[10]) ? 15'b000000000000011 : 15'b000000000001111;
										assign node10526 = (inp[6]) ? node10540 : node10527;
											assign node10527 = (inp[5]) ? node10535 : node10528;
												assign node10528 = (inp[13]) ? node10532 : node10529;
													assign node10529 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node10532 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node10535 = (inp[0]) ? node10537 : 15'b000000000001111;
													assign node10537 = (inp[13]) ? 15'b000000000000001 : 15'b000000000000011;
											assign node10540 = (inp[13]) ? node10548 : node10541;
												assign node10541 = (inp[0]) ? node10545 : node10542;
													assign node10542 = (inp[14]) ? 15'b000000000000011 : 15'b000000000000111;
													assign node10545 = (inp[14]) ? 15'b000000000000001 : 15'b000000000000011;
												assign node10548 = (inp[14]) ? node10550 : 15'b000000000000011;
													assign node10550 = (inp[5]) ? 15'b000000000000000 : 15'b000000000000001;

endmodule