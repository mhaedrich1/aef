module dtc_split66_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node701;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node980;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1099;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1110;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1121;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1191;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1200;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1224;
	wire [3-1:0] node1226;
	wire [3-1:0] node1228;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1238;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1244;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1299;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1318;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1337;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1355;
	wire [3-1:0] node1356;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1388;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1414;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1425;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1441;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1461;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1468;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1474;
	wire [3-1:0] node1477;
	wire [3-1:0] node1479;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1491;
	wire [3-1:0] node1494;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1500;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1514;
	wire [3-1:0] node1516;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1521;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1535;
	wire [3-1:0] node1536;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1548;
	wire [3-1:0] node1549;
	wire [3-1:0] node1552;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1560;
	wire [3-1:0] node1563;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1570;
	wire [3-1:0] node1571;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1581;
	wire [3-1:0] node1584;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1591;
	wire [3-1:0] node1593;
	wire [3-1:0] node1594;
	wire [3-1:0] node1598;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1609;
	wire [3-1:0] node1610;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1615;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1622;
	wire [3-1:0] node1625;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1631;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1638;
	wire [3-1:0] node1640;
	wire [3-1:0] node1643;
	wire [3-1:0] node1645;
	wire [3-1:0] node1648;
	wire [3-1:0] node1649;
	wire [3-1:0] node1650;
	wire [3-1:0] node1653;
	wire [3-1:0] node1657;
	wire [3-1:0] node1658;
	wire [3-1:0] node1659;
	wire [3-1:0] node1660;
	wire [3-1:0] node1663;
	wire [3-1:0] node1666;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1676;
	wire [3-1:0] node1679;
	wire [3-1:0] node1680;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1686;
	wire [3-1:0] node1687;
	wire [3-1:0] node1688;
	wire [3-1:0] node1691;
	wire [3-1:0] node1694;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1701;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1712;
	wire [3-1:0] node1713;
	wire [3-1:0] node1714;
	wire [3-1:0] node1716;
	wire [3-1:0] node1719;
	wire [3-1:0] node1720;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1727;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1737;
	wire [3-1:0] node1739;
	wire [3-1:0] node1742;
	wire [3-1:0] node1743;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1750;
	wire [3-1:0] node1754;
	wire [3-1:0] node1755;
	wire [3-1:0] node1759;
	wire [3-1:0] node1760;
	wire [3-1:0] node1762;
	wire [3-1:0] node1765;
	wire [3-1:0] node1766;
	wire [3-1:0] node1769;
	wire [3-1:0] node1772;
	wire [3-1:0] node1773;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1776;
	wire [3-1:0] node1779;
	wire [3-1:0] node1782;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1787;
	wire [3-1:0] node1791;
	wire [3-1:0] node1793;
	wire [3-1:0] node1796;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1800;
	wire [3-1:0] node1803;
	wire [3-1:0] node1804;
	wire [3-1:0] node1807;
	wire [3-1:0] node1810;
	wire [3-1:0] node1811;
	wire [3-1:0] node1813;
	wire [3-1:0] node1816;
	wire [3-1:0] node1817;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1825;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1828;
	wire [3-1:0] node1832;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1838;
	wire [3-1:0] node1841;
	wire [3-1:0] node1842;
	wire [3-1:0] node1846;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1853;
	wire [3-1:0] node1854;
	wire [3-1:0] node1858;
	wire [3-1:0] node1859;
	wire [3-1:0] node1861;
	wire [3-1:0] node1864;
	wire [3-1:0] node1865;
	wire [3-1:0] node1869;
	wire [3-1:0] node1870;
	wire [3-1:0] node1871;
	wire [3-1:0] node1872;
	wire [3-1:0] node1875;
	wire [3-1:0] node1877;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1884;
	wire [3-1:0] node1887;
	wire [3-1:0] node1888;
	wire [3-1:0] node1890;
	wire [3-1:0] node1893;
	wire [3-1:0] node1894;
	wire [3-1:0] node1895;
	wire [3-1:0] node1898;
	wire [3-1:0] node1901;
	wire [3-1:0] node1903;
	wire [3-1:0] node1906;
	wire [3-1:0] node1907;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1910;
	wire [3-1:0] node1911;
	wire [3-1:0] node1912;
	wire [3-1:0] node1913;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1921;
	wire [3-1:0] node1924;
	wire [3-1:0] node1925;
	wire [3-1:0] node1929;
	wire [3-1:0] node1930;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1936;
	wire [3-1:0] node1937;
	wire [3-1:0] node1940;
	wire [3-1:0] node1943;
	wire [3-1:0] node1944;
	wire [3-1:0] node1947;
	wire [3-1:0] node1950;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1953;
	wire [3-1:0] node1955;
	wire [3-1:0] node1959;
	wire [3-1:0] node1960;
	wire [3-1:0] node1962;
	wire [3-1:0] node1965;
	wire [3-1:0] node1966;
	wire [3-1:0] node1969;
	wire [3-1:0] node1972;
	wire [3-1:0] node1973;
	wire [3-1:0] node1974;
	wire [3-1:0] node1976;
	wire [3-1:0] node1979;
	wire [3-1:0] node1981;
	wire [3-1:0] node1984;
	wire [3-1:0] node1985;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1991;
	wire [3-1:0] node1992;
	wire [3-1:0] node1993;
	wire [3-1:0] node1994;
	wire [3-1:0] node1997;
	wire [3-1:0] node2000;
	wire [3-1:0] node2001;
	wire [3-1:0] node2005;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2010;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2017;
	wire [3-1:0] node2020;
	wire [3-1:0] node2021;
	wire [3-1:0] node2022;
	wire [3-1:0] node2023;
	wire [3-1:0] node2028;
	wire [3-1:0] node2029;
	wire [3-1:0] node2030;
	wire [3-1:0] node2033;
	wire [3-1:0] node2036;
	wire [3-1:0] node2039;
	wire [3-1:0] node2040;
	wire [3-1:0] node2041;
	wire [3-1:0] node2042;
	wire [3-1:0] node2043;
	wire [3-1:0] node2047;
	wire [3-1:0] node2049;
	wire [3-1:0] node2052;
	wire [3-1:0] node2053;
	wire [3-1:0] node2054;
	wire [3-1:0] node2057;
	wire [3-1:0] node2060;
	wire [3-1:0] node2062;
	wire [3-1:0] node2065;
	wire [3-1:0] node2066;
	wire [3-1:0] node2067;
	wire [3-1:0] node2068;
	wire [3-1:0] node2071;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2081;
	wire [3-1:0] node2084;
	wire [3-1:0] node2087;
	wire [3-1:0] node2088;
	wire [3-1:0] node2091;
	wire [3-1:0] node2094;
	wire [3-1:0] node2095;
	wire [3-1:0] node2096;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2100;
	wire [3-1:0] node2104;
	wire [3-1:0] node2106;
	wire [3-1:0] node2109;
	wire [3-1:0] node2111;
	wire [3-1:0] node2113;
	wire [3-1:0] node2116;
	wire [3-1:0] node2117;
	wire [3-1:0] node2118;
	wire [3-1:0] node2119;
	wire [3-1:0] node2126;
	wire [3-1:0] node2127;
	wire [3-1:0] node2128;
	wire [3-1:0] node2129;
	wire [3-1:0] node2130;
	wire [3-1:0] node2131;
	wire [3-1:0] node2135;
	wire [3-1:0] node2137;
	wire [3-1:0] node2140;
	wire [3-1:0] node2141;
	wire [3-1:0] node2144;
	wire [3-1:0] node2145;
	wire [3-1:0] node2148;
	wire [3-1:0] node2151;
	wire [3-1:0] node2152;
	wire [3-1:0] node2153;
	wire [3-1:0] node2154;
	wire [3-1:0] node2157;
	wire [3-1:0] node2160;
	wire [3-1:0] node2161;
	wire [3-1:0] node2165;
	wire [3-1:0] node2166;
	wire [3-1:0] node2167;
	wire [3-1:0] node2170;
	wire [3-1:0] node2173;
	wire [3-1:0] node2175;
	wire [3-1:0] node2178;
	wire [3-1:0] node2179;
	wire [3-1:0] node2180;
	wire [3-1:0] node2181;
	wire [3-1:0] node2184;
	wire [3-1:0] node2185;
	wire [3-1:0] node2189;
	wire [3-1:0] node2190;
	wire [3-1:0] node2192;
	wire [3-1:0] node2195;
	wire [3-1:0] node2196;
	wire [3-1:0] node2199;
	wire [3-1:0] node2202;
	wire [3-1:0] node2203;
	wire [3-1:0] node2204;
	wire [3-1:0] node2205;
	wire [3-1:0] node2209;
	wire [3-1:0] node2210;

	assign outp = (inp[6]) ? node898 : node1;
		assign node1 = (inp[3]) ? node643 : node2;
			assign node2 = (inp[9]) ? node364 : node3;
				assign node3 = (inp[4]) ? node187 : node4;
					assign node4 = (inp[0]) ? node98 : node5;
						assign node5 = (inp[1]) ? node53 : node6;
							assign node6 = (inp[7]) ? node36 : node7;
								assign node7 = (inp[10]) ? node23 : node8;
									assign node8 = (inp[5]) ? node16 : node9;
										assign node9 = (inp[8]) ? node13 : node10;
											assign node10 = (inp[2]) ? 3'b101 : 3'b011;
											assign node13 = (inp[11]) ? 3'b011 : 3'b011;
										assign node16 = (inp[11]) ? node20 : node17;
											assign node17 = (inp[8]) ? 3'b011 : 3'b101;
											assign node20 = (inp[2]) ? 3'b001 : 3'b001;
									assign node23 = (inp[2]) ? node29 : node24;
										assign node24 = (inp[8]) ? 3'b001 : node25;
											assign node25 = (inp[5]) ? 3'b001 : 3'b101;
										assign node29 = (inp[11]) ? node33 : node30;
											assign node30 = (inp[5]) ? 3'b001 : 3'b101;
											assign node33 = (inp[5]) ? 3'b110 : 3'b001;
								assign node36 = (inp[2]) ? node46 : node37;
									assign node37 = (inp[5]) ? node43 : node38;
										assign node38 = (inp[8]) ? node40 : 3'b001;
											assign node40 = (inp[10]) ? 3'b001 : 3'b000;
										assign node43 = (inp[8]) ? 3'b001 : 3'b000;
									assign node46 = (inp[8]) ? 3'b001 : node47;
										assign node47 = (inp[5]) ? node49 : 3'b001;
											assign node49 = (inp[10]) ? 3'b000 : 3'b001;
							assign node53 = (inp[7]) ? node75 : node54;
								assign node54 = (inp[10]) ? node64 : node55;
									assign node55 = (inp[5]) ? node59 : node56;
										assign node56 = (inp[8]) ? 3'b101 : 3'b001;
										assign node59 = (inp[8]) ? 3'b001 : node60;
											assign node60 = (inp[11]) ? 3'b110 : 3'b001;
									assign node64 = (inp[8]) ? node70 : node65;
										assign node65 = (inp[11]) ? node67 : 3'b110;
											assign node67 = (inp[2]) ? 3'b010 : 3'b110;
										assign node70 = (inp[2]) ? 3'b110 : node71;
											assign node71 = (inp[5]) ? 3'b000 : 3'b001;
								assign node75 = (inp[8]) ? node87 : node76;
									assign node76 = (inp[11]) ? node82 : node77;
										assign node77 = (inp[5]) ? 3'b101 : node78;
											assign node78 = (inp[2]) ? 3'b011 : 3'b101;
										assign node82 = (inp[2]) ? node84 : 3'b001;
											assign node84 = (inp[10]) ? 3'b001 : 3'b101;
									assign node87 = (inp[10]) ? node95 : node88;
										assign node88 = (inp[5]) ? node92 : node89;
											assign node89 = (inp[2]) ? 3'b011 : 3'b111;
											assign node92 = (inp[11]) ? 3'b001 : 3'b011;
										assign node95 = (inp[11]) ? 3'b001 : 3'b011;
						assign node98 = (inp[7]) ? node144 : node99;
							assign node99 = (inp[10]) ? node121 : node100;
								assign node100 = (inp[11]) ? node114 : node101;
									assign node101 = (inp[1]) ? node107 : node102;
										assign node102 = (inp[2]) ? 3'b001 : node103;
											assign node103 = (inp[8]) ? 3'b001 : 3'b110;
										assign node107 = (inp[2]) ? node111 : node108;
											assign node108 = (inp[5]) ? 3'b110 : 3'b001;
											assign node111 = (inp[5]) ? 3'b010 : 3'b110;
									assign node114 = (inp[5]) ? node118 : node115;
										assign node115 = (inp[8]) ? 3'b110 : 3'b010;
										assign node118 = (inp[1]) ? 3'b100 : 3'b110;
								assign node121 = (inp[11]) ? node135 : node122;
									assign node122 = (inp[1]) ? node130 : node123;
										assign node123 = (inp[5]) ? node127 : node124;
											assign node124 = (inp[8]) ? 3'b010 : 3'b110;
											assign node127 = (inp[2]) ? 3'b010 : 3'b110;
										assign node130 = (inp[5]) ? node132 : 3'b010;
											assign node132 = (inp[8]) ? 3'b010 : 3'b100;
									assign node135 = (inp[1]) ? node141 : node136;
										assign node136 = (inp[2]) ? 3'b100 : node137;
											assign node137 = (inp[8]) ? 3'b010 : 3'b000;
										assign node141 = (inp[5]) ? 3'b100 : 3'b110;
							assign node144 = (inp[1]) ? node164 : node145;
								assign node145 = (inp[10]) ? node157 : node146;
									assign node146 = (inp[8]) ? node152 : node147;
										assign node147 = (inp[5]) ? 3'b001 : node148;
											assign node148 = (inp[11]) ? 3'b101 : 3'b001;
										assign node152 = (inp[5]) ? 3'b101 : node153;
											assign node153 = (inp[2]) ? 3'b101 : 3'b010;
									assign node157 = (inp[8]) ? node161 : node158;
										assign node158 = (inp[5]) ? 3'b110 : 3'b001;
										assign node161 = (inp[5]) ? 3'b001 : 3'b101;
								assign node164 = (inp[10]) ? node176 : node165;
									assign node165 = (inp[8]) ? node171 : node166;
										assign node166 = (inp[5]) ? 3'b110 : node167;
											assign node167 = (inp[2]) ? 3'b001 : 3'b001;
										assign node171 = (inp[5]) ? 3'b001 : node172;
											assign node172 = (inp[11]) ? 3'b001 : 3'b101;
									assign node176 = (inp[5]) ? node182 : node177;
										assign node177 = (inp[8]) ? node179 : 3'b110;
											assign node179 = (inp[11]) ? 3'b010 : 3'b001;
										assign node182 = (inp[8]) ? 3'b110 : node183;
											assign node183 = (inp[11]) ? 3'b010 : 3'b010;
					assign node187 = (inp[7]) ? node273 : node188;
						assign node188 = (inp[0]) ? node240 : node189;
							assign node189 = (inp[1]) ? node217 : node190;
								assign node190 = (inp[10]) ? node204 : node191;
									assign node191 = (inp[8]) ? node197 : node192;
										assign node192 = (inp[5]) ? 3'b110 : node193;
											assign node193 = (inp[11]) ? 3'b010 : 3'b000;
										assign node197 = (inp[5]) ? node201 : node198;
											assign node198 = (inp[11]) ? 3'b000 : 3'b100;
											assign node201 = (inp[2]) ? 3'b000 : 3'b000;
									assign node204 = (inp[11]) ? node212 : node205;
										assign node205 = (inp[2]) ? node209 : node206;
											assign node206 = (inp[8]) ? 3'b110 : 3'b100;
											assign node209 = (inp[5]) ? 3'b000 : 3'b000;
										assign node212 = (inp[2]) ? 3'b110 : node213;
											assign node213 = (inp[8]) ? 3'b000 : 3'b010;
								assign node217 = (inp[2]) ? node227 : node218;
									assign node218 = (inp[8]) ? node224 : node219;
										assign node219 = (inp[11]) ? node221 : 3'b010;
											assign node221 = (inp[10]) ? 3'b010 : 3'b010;
										assign node224 = (inp[5]) ? 3'b010 : 3'b000;
									assign node227 = (inp[10]) ? node233 : node228;
										assign node228 = (inp[8]) ? 3'b110 : node229;
											assign node229 = (inp[5]) ? 3'b010 : 3'b110;
										assign node233 = (inp[8]) ? node237 : node234;
											assign node234 = (inp[5]) ? 3'b100 : 3'b010;
											assign node237 = (inp[11]) ? 3'b010 : 3'b010;
							assign node240 = (inp[10]) ? node256 : node241;
								assign node241 = (inp[1]) ? node249 : node242;
									assign node242 = (inp[5]) ? node246 : node243;
										assign node243 = (inp[11]) ? 3'b010 : 3'b110;
										assign node246 = (inp[8]) ? 3'b010 : 3'b100;
									assign node249 = (inp[5]) ? node251 : 3'b100;
										assign node251 = (inp[11]) ? node253 : 3'b100;
											assign node253 = (inp[8]) ? 3'b100 : 3'b000;
								assign node256 = (inp[1]) ? node266 : node257;
									assign node257 = (inp[2]) ? node263 : node258;
										assign node258 = (inp[5]) ? 3'b100 : node259;
											assign node259 = (inp[8]) ? 3'b000 : 3'b100;
										assign node263 = (inp[5]) ? 3'b000 : 3'b100;
									assign node266 = (inp[11]) ? 3'b000 : node267;
										assign node267 = (inp[8]) ? node269 : 3'b000;
											assign node269 = (inp[2]) ? 3'b000 : 3'b000;
						assign node273 = (inp[0]) ? node317 : node274;
							assign node274 = (inp[5]) ? node294 : node275;
								assign node275 = (inp[11]) ? node285 : node276;
									assign node276 = (inp[1]) ? node280 : node277;
										assign node277 = (inp[10]) ? 3'b001 : 3'b111;
										assign node280 = (inp[10]) ? node282 : 3'b001;
											assign node282 = (inp[8]) ? 3'b001 : 3'b110;
									assign node285 = (inp[10]) ? 3'b001 : node286;
										assign node286 = (inp[1]) ? node290 : node287;
											assign node287 = (inp[8]) ? 3'b011 : 3'b001;
											assign node290 = (inp[8]) ? 3'b101 : 3'b001;
								assign node294 = (inp[1]) ? node306 : node295;
									assign node295 = (inp[10]) ? node299 : node296;
										assign node296 = (inp[11]) ? 3'b101 : 3'b111;
										assign node299 = (inp[11]) ? node303 : node300;
											assign node300 = (inp[2]) ? 3'b001 : 3'b001;
											assign node303 = (inp[2]) ? 3'b000 : 3'b001;
									assign node306 = (inp[10]) ? node312 : node307;
										assign node307 = (inp[8]) ? node309 : 3'b110;
											assign node309 = (inp[2]) ? 3'b001 : 3'b101;
										assign node312 = (inp[2]) ? node314 : 3'b110;
											assign node314 = (inp[8]) ? 3'b110 : 3'b010;
							assign node317 = (inp[1]) ? node345 : node318;
								assign node318 = (inp[10]) ? node334 : node319;
									assign node319 = (inp[8]) ? node327 : node320;
										assign node320 = (inp[11]) ? node324 : node321;
											assign node321 = (inp[5]) ? 3'b110 : 3'b001;
											assign node324 = (inp[2]) ? 3'b010 : 3'b010;
										assign node327 = (inp[11]) ? node331 : node328;
											assign node328 = (inp[2]) ? 3'b001 : 3'b001;
											assign node331 = (inp[5]) ? 3'b110 : 3'b000;
									assign node334 = (inp[5]) ? node340 : node335;
										assign node335 = (inp[11]) ? 3'b010 : node336;
											assign node336 = (inp[8]) ? 3'b010 : 3'b110;
										assign node340 = (inp[11]) ? node342 : 3'b010;
											assign node342 = (inp[8]) ? 3'b010 : 3'b000;
								assign node345 = (inp[8]) ? node357 : node346;
									assign node346 = (inp[10]) ? node352 : node347;
										assign node347 = (inp[5]) ? 3'b010 : node348;
											assign node348 = (inp[11]) ? 3'b010 : 3'b111;
										assign node352 = (inp[5]) ? node354 : 3'b010;
											assign node354 = (inp[11]) ? 3'b000 : 3'b100;
									assign node357 = (inp[2]) ? node359 : 3'b110;
										assign node359 = (inp[10]) ? 3'b010 : node360;
											assign node360 = (inp[5]) ? 3'b010 : 3'b110;
				assign node364 = (inp[4]) ? node546 : node365;
					assign node365 = (inp[7]) ? node451 : node366;
						assign node366 = (inp[10]) ? node416 : node367;
							assign node367 = (inp[11]) ? node391 : node368;
								assign node368 = (inp[0]) ? node380 : node369;
									assign node369 = (inp[1]) ? node375 : node370;
										assign node370 = (inp[8]) ? 3'b010 : node371;
											assign node371 = (inp[5]) ? 3'b100 : 3'b010;
										assign node375 = (inp[5]) ? 3'b010 : node376;
											assign node376 = (inp[2]) ? 3'b010 : 3'b011;
									assign node380 = (inp[1]) ? node386 : node381;
										assign node381 = (inp[5]) ? node383 : 3'b010;
											assign node383 = (inp[8]) ? 3'b010 : 3'b100;
										assign node386 = (inp[8]) ? 3'b100 : node387;
											assign node387 = (inp[5]) ? 3'b000 : 3'b100;
								assign node391 = (inp[5]) ? node405 : node392;
									assign node392 = (inp[0]) ? node400 : node393;
										assign node393 = (inp[1]) ? node397 : node394;
											assign node394 = (inp[8]) ? 3'b010 : 3'b000;
											assign node397 = (inp[2]) ? 3'b010 : 3'b110;
										assign node400 = (inp[2]) ? node402 : 3'b000;
											assign node402 = (inp[1]) ? 3'b100 : 3'b010;
									assign node405 = (inp[0]) ? node411 : node406;
										assign node406 = (inp[1]) ? 3'b100 : node407;
											assign node407 = (inp[8]) ? 3'b000 : 3'b000;
										assign node411 = (inp[2]) ? node413 : 3'b000;
											assign node413 = (inp[8]) ? 3'b100 : 3'b000;
							assign node416 = (inp[0]) ? node438 : node417;
								assign node417 = (inp[1]) ? node431 : node418;
									assign node418 = (inp[5]) ? node426 : node419;
										assign node419 = (inp[2]) ? node423 : node420;
											assign node420 = (inp[11]) ? 3'b100 : 3'b000;
											assign node423 = (inp[11]) ? 3'b000 : 3'b100;
										assign node426 = (inp[8]) ? node428 : 3'b000;
											assign node428 = (inp[11]) ? 3'b000 : 3'b100;
									assign node431 = (inp[5]) ? node433 : 3'b010;
										assign node433 = (inp[11]) ? 3'b100 : node434;
											assign node434 = (inp[2]) ? 3'b100 : 3'b110;
								assign node438 = (inp[1]) ? 3'b000 : node439;
									assign node439 = (inp[2]) ? node445 : node440;
										assign node440 = (inp[8]) ? 3'b100 : node441;
											assign node441 = (inp[5]) ? 3'b000 : 3'b100;
										assign node445 = (inp[5]) ? 3'b000 : node446;
											assign node446 = (inp[11]) ? 3'b000 : 3'b000;
						assign node451 = (inp[0]) ? node499 : node452;
							assign node452 = (inp[1]) ? node474 : node453;
								assign node453 = (inp[5]) ? node467 : node454;
									assign node454 = (inp[8]) ? node462 : node455;
										assign node455 = (inp[10]) ? node459 : node456;
											assign node456 = (inp[11]) ? 3'b000 : 3'b001;
											assign node459 = (inp[11]) ? 3'b100 : 3'b000;
										assign node462 = (inp[11]) ? node464 : 3'b101;
											assign node464 = (inp[10]) ? 3'b000 : 3'b101;
									assign node467 = (inp[11]) ? node469 : 3'b000;
										assign node469 = (inp[10]) ? 3'b100 : node470;
											assign node470 = (inp[8]) ? 3'b101 : 3'b000;
								assign node474 = (inp[8]) ? node488 : node475;
									assign node475 = (inp[11]) ? node483 : node476;
										assign node476 = (inp[5]) ? node480 : node477;
											assign node477 = (inp[10]) ? 3'b110 : 3'b001;
											assign node480 = (inp[10]) ? 3'b101 : 3'b110;
										assign node483 = (inp[10]) ? node485 : 3'b110;
											assign node485 = (inp[2]) ? 3'b010 : 3'b110;
									assign node488 = (inp[5]) ? node494 : node489;
										assign node489 = (inp[10]) ? 3'b001 : node490;
											assign node490 = (inp[11]) ? 3'b001 : 3'b101;
										assign node494 = (inp[10]) ? node496 : 3'b001;
											assign node496 = (inp[2]) ? 3'b010 : 3'b110;
							assign node499 = (inp[1]) ? node525 : node500;
								assign node500 = (inp[2]) ? node514 : node501;
									assign node501 = (inp[8]) ? node507 : node502;
										assign node502 = (inp[10]) ? node504 : 3'b010;
											assign node504 = (inp[11]) ? 3'b100 : 3'b000;
										assign node507 = (inp[10]) ? node511 : node508;
											assign node508 = (inp[5]) ? 3'b110 : 3'b000;
											assign node511 = (inp[5]) ? 3'b010 : 3'b110;
									assign node514 = (inp[10]) ? node520 : node515;
										assign node515 = (inp[8]) ? 3'b110 : node516;
											assign node516 = (inp[5]) ? 3'b010 : 3'b110;
										assign node520 = (inp[11]) ? 3'b010 : node521;
											assign node521 = (inp[5]) ? 3'b010 : 3'b010;
								assign node525 = (inp[10]) ? node537 : node526;
									assign node526 = (inp[11]) ? node532 : node527;
										assign node527 = (inp[5]) ? node529 : 3'b110;
											assign node529 = (inp[8]) ? 3'b010 : 3'b100;
										assign node532 = (inp[5]) ? node534 : 3'b010;
											assign node534 = (inp[8]) ? 3'b010 : 3'b100;
									assign node537 = (inp[8]) ? node541 : node538;
										assign node538 = (inp[5]) ? 3'b000 : 3'b100;
										assign node541 = (inp[11]) ? node543 : 3'b010;
											assign node543 = (inp[2]) ? 3'b100 : 3'b000;
					assign node546 = (inp[0]) ? node610 : node547;
						assign node547 = (inp[1]) ? node575 : node548;
							assign node548 = (inp[7]) ? node554 : node549;
								assign node549 = (inp[5]) ? node551 : 3'b010;
									assign node551 = (inp[10]) ? 3'b000 : 3'b010;
								assign node554 = (inp[5]) ? node568 : node555;
									assign node555 = (inp[10]) ? node561 : node556;
										assign node556 = (inp[11]) ? node558 : 3'b010;
											assign node558 = (inp[8]) ? 3'b000 : 3'b100;
										assign node561 = (inp[8]) ? node565 : node562;
											assign node562 = (inp[11]) ? 3'b000 : 3'b100;
											assign node565 = (inp[11]) ? 3'b100 : 3'b000;
									assign node568 = (inp[8]) ? node570 : 3'b000;
										assign node570 = (inp[11]) ? node572 : 3'b100;
											assign node572 = (inp[10]) ? 3'b000 : 3'b100;
							assign node575 = (inp[7]) ? node589 : node576;
								assign node576 = (inp[8]) ? node582 : node577;
									assign node577 = (inp[5]) ? 3'b000 : node578;
										assign node578 = (inp[10]) ? 3'b000 : 3'b100;
									assign node582 = (inp[10]) ? node586 : node583;
										assign node583 = (inp[5]) ? 3'b100 : 3'b000;
										assign node586 = (inp[5]) ? 3'b000 : 3'b100;
								assign node589 = (inp[10]) ? node603 : node590;
									assign node590 = (inp[11]) ? node598 : node591;
										assign node591 = (inp[8]) ? node595 : node592;
											assign node592 = (inp[5]) ? 3'b010 : 3'b010;
											assign node595 = (inp[2]) ? 3'b010 : 3'b110;
										assign node598 = (inp[8]) ? node600 : 3'b100;
											assign node600 = (inp[5]) ? 3'b010 : 3'b110;
									assign node603 = (inp[8]) ? node605 : 3'b100;
										assign node605 = (inp[2]) ? 3'b010 : node606;
											assign node606 = (inp[11]) ? 3'b100 : 3'b110;
						assign node610 = (inp[7]) ? node612 : 3'b000;
							assign node612 = (inp[1]) ? node636 : node613;
								assign node613 = (inp[10]) ? node625 : node614;
									assign node614 = (inp[11]) ? node620 : node615;
										assign node615 = (inp[5]) ? node617 : 3'b010;
											assign node617 = (inp[8]) ? 3'b110 : 3'b100;
										assign node620 = (inp[8]) ? node622 : 3'b100;
											assign node622 = (inp[5]) ? 3'b100 : 3'b000;
									assign node625 = (inp[11]) ? node631 : node626;
										assign node626 = (inp[2]) ? 3'b100 : node627;
											assign node627 = (inp[8]) ? 3'b000 : 3'b100;
										assign node631 = (inp[8]) ? node633 : 3'b000;
											assign node633 = (inp[5]) ? 3'b000 : 3'b100;
								assign node636 = (inp[10]) ? 3'b000 : node637;
									assign node637 = (inp[8]) ? node639 : 3'b000;
										assign node639 = (inp[11]) ? 3'b000 : 3'b100;
			assign node643 = (inp[9]) ? node861 : node644;
				assign node644 = (inp[7]) ? node712 : node645;
					assign node645 = (inp[4]) ? node701 : node646;
						assign node646 = (inp[0]) ? node686 : node647;
							assign node647 = (inp[1]) ? node661 : node648;
								assign node648 = (inp[10]) ? 3'b000 : node649;
									assign node649 = (inp[11]) ? node655 : node650;
										assign node650 = (inp[5]) ? node652 : 3'b100;
											assign node652 = (inp[8]) ? 3'b100 : 3'b000;
										assign node655 = (inp[8]) ? node657 : 3'b000;
											assign node657 = (inp[5]) ? 3'b000 : 3'b000;
								assign node661 = (inp[10]) ? node673 : node662;
									assign node662 = (inp[11]) ? node666 : node663;
										assign node663 = (inp[2]) ? 3'b010 : 3'b110;
										assign node666 = (inp[8]) ? node670 : node667;
											assign node667 = (inp[5]) ? 3'b000 : 3'b100;
											assign node670 = (inp[2]) ? 3'b010 : 3'b000;
									assign node673 = (inp[8]) ? node679 : node674;
										assign node674 = (inp[5]) ? 3'b000 : node675;
											assign node675 = (inp[11]) ? 3'b000 : 3'b100;
										assign node679 = (inp[11]) ? node683 : node680;
											assign node680 = (inp[2]) ? 3'b100 : 3'b000;
											assign node683 = (inp[5]) ? 3'b000 : 3'b100;
							assign node686 = (inp[10]) ? 3'b000 : node687;
								assign node687 = (inp[1]) ? 3'b000 : node688;
									assign node688 = (inp[8]) ? node694 : node689;
										assign node689 = (inp[11]) ? 3'b000 : node690;
											assign node690 = (inp[5]) ? 3'b000 : 3'b100;
										assign node694 = (inp[11]) ? node696 : 3'b100;
											assign node696 = (inp[5]) ? 3'b000 : 3'b100;
						assign node701 = (inp[2]) ? node703 : 3'b000;
							assign node703 = (inp[11]) ? 3'b000 : node704;
								assign node704 = (inp[10]) ? 3'b000 : node705;
									assign node705 = (inp[8]) ? node707 : 3'b000;
										assign node707 = (inp[1]) ? 3'b100 : 3'b000;
					assign node712 = (inp[4]) ? node806 : node713;
						assign node713 = (inp[0]) ? node765 : node714;
							assign node714 = (inp[1]) ? node738 : node715;
								assign node715 = (inp[10]) ? node727 : node716;
									assign node716 = (inp[5]) ? node722 : node717;
										assign node717 = (inp[8]) ? node719 : 3'b000;
											assign node719 = (inp[11]) ? 3'b000 : 3'b100;
										assign node722 = (inp[8]) ? node724 : 3'b110;
											assign node724 = (inp[2]) ? 3'b010 : 3'b000;
									assign node727 = (inp[5]) ? node733 : node728;
										assign node728 = (inp[8]) ? node730 : 3'b110;
											assign node730 = (inp[2]) ? 3'b000 : 3'b000;
										assign node733 = (inp[8]) ? 3'b110 : node734;
											assign node734 = (inp[11]) ? 3'b010 : 3'b100;
								assign node738 = (inp[8]) ? node752 : node739;
									assign node739 = (inp[5]) ? node747 : node740;
										assign node740 = (inp[11]) ? node744 : node741;
											assign node741 = (inp[10]) ? 3'b010 : 3'b110;
											assign node744 = (inp[10]) ? 3'b110 : 3'b000;
										assign node747 = (inp[10]) ? node749 : 3'b010;
											assign node749 = (inp[11]) ? 3'b100 : 3'b000;
									assign node752 = (inp[2]) ? node758 : node753;
										assign node753 = (inp[10]) ? node755 : 3'b110;
											assign node755 = (inp[11]) ? 3'b010 : 3'b110;
										assign node758 = (inp[11]) ? node762 : node759;
											assign node759 = (inp[5]) ? 3'b010 : 3'b001;
											assign node762 = (inp[5]) ? 3'b010 : 3'b010;
							assign node765 = (inp[1]) ? node787 : node766;
								assign node766 = (inp[10]) ? node774 : node767;
									assign node767 = (inp[5]) ? 3'b100 : node768;
										assign node768 = (inp[11]) ? node770 : 3'b110;
											assign node770 = (inp[2]) ? 3'b010 : 3'b110;
									assign node774 = (inp[11]) ? node782 : node775;
										assign node775 = (inp[5]) ? node779 : node776;
											assign node776 = (inp[8]) ? 3'b010 : 3'b100;
											assign node779 = (inp[2]) ? 3'b000 : 3'b100;
										assign node782 = (inp[5]) ? node784 : 3'b100;
											assign node784 = (inp[8]) ? 3'b100 : 3'b000;
								assign node787 = (inp[8]) ? node795 : node788;
									assign node788 = (inp[5]) ? 3'b000 : node789;
										assign node789 = (inp[2]) ? 3'b000 : node790;
											assign node790 = (inp[10]) ? 3'b000 : 3'b000;
									assign node795 = (inp[10]) ? node801 : node796;
										assign node796 = (inp[11]) ? 3'b100 : node797;
											assign node797 = (inp[5]) ? 3'b000 : 3'b010;
										assign node801 = (inp[11]) ? 3'b000 : node802;
											assign node802 = (inp[5]) ? 3'b000 : 3'b100;
						assign node806 = (inp[0]) ? node846 : node807;
							assign node807 = (inp[1]) ? node821 : node808;
								assign node808 = (inp[10]) ? 3'b000 : node809;
									assign node809 = (inp[11]) ? node815 : node810;
										assign node810 = (inp[8]) ? 3'b100 : node811;
											assign node811 = (inp[5]) ? 3'b000 : 3'b100;
										assign node815 = (inp[8]) ? node817 : 3'b000;
											assign node817 = (inp[2]) ? 3'b100 : 3'b000;
								assign node821 = (inp[10]) ? node835 : node822;
									assign node822 = (inp[5]) ? node828 : node823;
										assign node823 = (inp[2]) ? 3'b010 : node824;
											assign node824 = (inp[11]) ? 3'b100 : 3'b010;
										assign node828 = (inp[2]) ? node832 : node829;
											assign node829 = (inp[11]) ? 3'b100 : 3'b010;
											assign node832 = (inp[11]) ? 3'b000 : 3'b100;
									assign node835 = (inp[11]) ? node841 : node836;
										assign node836 = (inp[2]) ? 3'b100 : node837;
											assign node837 = (inp[5]) ? 3'b000 : 3'b000;
										assign node841 = (inp[8]) ? node843 : 3'b000;
											assign node843 = (inp[5]) ? 3'b000 : 3'b100;
							assign node846 = (inp[1]) ? 3'b000 : node847;
								assign node847 = (inp[10]) ? 3'b000 : node848;
									assign node848 = (inp[11]) ? node854 : node849;
										assign node849 = (inp[5]) ? node851 : 3'b100;
											assign node851 = (inp[8]) ? 3'b100 : 3'b000;
										assign node854 = (inp[5]) ? 3'b000 : node855;
											assign node855 = (inp[2]) ? 3'b100 : 3'b000;
				assign node861 = (inp[7]) ? node863 : 3'b000;
					assign node863 = (inp[4]) ? 3'b000 : node864;
						assign node864 = (inp[0]) ? node888 : node865;
							assign node865 = (inp[1]) ? node871 : node866;
								assign node866 = (inp[10]) ? node868 : 3'b010;
									assign node868 = (inp[5]) ? 3'b000 : 3'b010;
								assign node871 = (inp[5]) ? node883 : node872;
									assign node872 = (inp[2]) ? node878 : node873;
										assign node873 = (inp[11]) ? 3'b100 : node874;
											assign node874 = (inp[8]) ? 3'b000 : 3'b100;
										assign node878 = (inp[10]) ? 3'b000 : node879;
											assign node879 = (inp[11]) ? 3'b100 : 3'b000;
									assign node883 = (inp[8]) ? node885 : 3'b000;
										assign node885 = (inp[11]) ? 3'b000 : 3'b100;
							assign node888 = (inp[1]) ? 3'b000 : node889;
								assign node889 = (inp[2]) ? node891 : 3'b000;
									assign node891 = (inp[8]) ? node893 : 3'b000;
										assign node893 = (inp[11]) ? 3'b000 : 3'b100;
		assign node898 = (inp[3]) ? node1540 : node899;
			assign node899 = (inp[0]) ? node1169 : node900;
				assign node900 = (inp[9]) ? node998 : node901;
					assign node901 = (inp[7]) ? node969 : node902;
						assign node902 = (inp[1]) ? node922 : node903;
							assign node903 = (inp[4]) ? node905 : 3'b111;
								assign node905 = (inp[10]) ? node913 : node906;
									assign node906 = (inp[5]) ? node908 : 3'b111;
										assign node908 = (inp[8]) ? node910 : 3'b011;
											assign node910 = (inp[2]) ? 3'b011 : 3'b111;
									assign node913 = (inp[5]) ? node917 : node914;
										assign node914 = (inp[11]) ? 3'b011 : 3'b111;
										assign node917 = (inp[11]) ? node919 : 3'b011;
											assign node919 = (inp[2]) ? 3'b111 : 3'b011;
							assign node922 = (inp[4]) ? node946 : node923;
								assign node923 = (inp[11]) ? node933 : node924;
									assign node924 = (inp[10]) ? node928 : node925;
										assign node925 = (inp[8]) ? 3'b011 : 3'b111;
										assign node928 = (inp[8]) ? node930 : 3'b011;
											assign node930 = (inp[2]) ? 3'b011 : 3'b011;
									assign node933 = (inp[8]) ? node939 : node934;
										assign node934 = (inp[10]) ? node936 : 3'b011;
											assign node936 = (inp[5]) ? 3'b010 : 3'b011;
										assign node939 = (inp[2]) ? node943 : node940;
											assign node940 = (inp[10]) ? 3'b111 : 3'b010;
											assign node943 = (inp[5]) ? 3'b011 : 3'b011;
								assign node946 = (inp[10]) ? node960 : node947;
									assign node947 = (inp[8]) ? node953 : node948;
										assign node948 = (inp[5]) ? 3'b101 : node949;
											assign node949 = (inp[11]) ? 3'b101 : 3'b011;
										assign node953 = (inp[2]) ? node957 : node954;
											assign node954 = (inp[5]) ? 3'b011 : 3'b111;
											assign node957 = (inp[5]) ? 3'b101 : 3'b011;
									assign node960 = (inp[5]) ? 3'b101 : node961;
										assign node961 = (inp[8]) ? node965 : node962;
											assign node962 = (inp[11]) ? 3'b001 : 3'b101;
											assign node965 = (inp[11]) ? 3'b101 : 3'b011;
						assign node969 = (inp[1]) ? node971 : 3'b111;
							assign node971 = (inp[4]) ? node973 : 3'b111;
								assign node973 = (inp[10]) ? node985 : node974;
									assign node974 = (inp[5]) ? node980 : node975;
										assign node975 = (inp[8]) ? 3'b111 : node976;
											assign node976 = (inp[11]) ? 3'b101 : 3'b111;
										assign node980 = (inp[11]) ? node982 : 3'b111;
											assign node982 = (inp[8]) ? 3'b111 : 3'b011;
									assign node985 = (inp[11]) ? node991 : node986;
										assign node986 = (inp[8]) ? node988 : 3'b011;
											assign node988 = (inp[5]) ? 3'b011 : 3'b111;
										assign node991 = (inp[5]) ? node995 : node992;
											assign node992 = (inp[8]) ? 3'b111 : 3'b011;
											assign node995 = (inp[8]) ? 3'b011 : 3'b101;
					assign node998 = (inp[7]) ? node1088 : node999;
						assign node999 = (inp[4]) ? node1055 : node1000;
							assign node1000 = (inp[1]) ? node1028 : node1001;
								assign node1001 = (inp[8]) ? node1015 : node1002;
									assign node1002 = (inp[5]) ? node1010 : node1003;
										assign node1003 = (inp[10]) ? node1007 : node1004;
											assign node1004 = (inp[2]) ? 3'b011 : 3'b001;
											assign node1007 = (inp[11]) ? 3'b101 : 3'b001;
										assign node1010 = (inp[2]) ? 3'b101 : node1011;
											assign node1011 = (inp[10]) ? 3'b001 : 3'b011;
									assign node1015 = (inp[5]) ? node1023 : node1016;
										assign node1016 = (inp[10]) ? node1020 : node1017;
											assign node1017 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1020 = (inp[2]) ? 3'b011 : 3'b011;
										assign node1023 = (inp[2]) ? node1025 : 3'b011;
											assign node1025 = (inp[10]) ? 3'b111 : 3'b011;
								assign node1028 = (inp[10]) ? node1042 : node1029;
									assign node1029 = (inp[11]) ? node1037 : node1030;
										assign node1030 = (inp[8]) ? node1034 : node1031;
											assign node1031 = (inp[2]) ? 3'b101 : 3'b111;
											assign node1034 = (inp[5]) ? 3'b001 : 3'b011;
										assign node1037 = (inp[8]) ? 3'b011 : node1038;
											assign node1038 = (inp[2]) ? 3'b001 : 3'b001;
									assign node1042 = (inp[8]) ? node1050 : node1043;
										assign node1043 = (inp[11]) ? node1047 : node1044;
											assign node1044 = (inp[5]) ? 3'b001 : 3'b001;
											assign node1047 = (inp[5]) ? 3'b001 : 3'b001;
										assign node1050 = (inp[2]) ? 3'b101 : node1051;
											assign node1051 = (inp[5]) ? 3'b001 : 3'b001;
							assign node1055 = (inp[10]) ? node1073 : node1056;
								assign node1056 = (inp[1]) ? node1064 : node1057;
									assign node1057 = (inp[11]) ? 3'b101 : node1058;
										assign node1058 = (inp[8]) ? node1060 : 3'b001;
											assign node1060 = (inp[5]) ? 3'b101 : 3'b001;
									assign node1064 = (inp[8]) ? node1066 : 3'b110;
										assign node1066 = (inp[2]) ? node1070 : node1067;
											assign node1067 = (inp[11]) ? 3'b001 : 3'b001;
											assign node1070 = (inp[5]) ? 3'b110 : 3'b001;
								assign node1073 = (inp[8]) ? node1079 : node1074;
									assign node1074 = (inp[11]) ? node1076 : 3'b110;
										assign node1076 = (inp[1]) ? 3'b010 : 3'b000;
									assign node1079 = (inp[5]) ? node1085 : node1080;
										assign node1080 = (inp[1]) ? 3'b001 : node1081;
											assign node1081 = (inp[11]) ? 3'b001 : 3'b011;
										assign node1085 = (inp[1]) ? 3'b110 : 3'b001;
						assign node1088 = (inp[4]) ? node1126 : node1089;
							assign node1089 = (inp[10]) ? node1103 : node1090;
								assign node1090 = (inp[8]) ? 3'b111 : node1091;
									assign node1091 = (inp[1]) ? node1097 : node1092;
										assign node1092 = (inp[11]) ? node1094 : 3'b111;
											assign node1094 = (inp[5]) ? 3'b111 : 3'b011;
										assign node1097 = (inp[5]) ? node1099 : 3'b111;
											assign node1099 = (inp[11]) ? 3'b111 : 3'b011;
								assign node1103 = (inp[1]) ? node1115 : node1104;
									assign node1104 = (inp[5]) ? node1110 : node1105;
										assign node1105 = (inp[8]) ? 3'b111 : node1106;
											assign node1106 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1110 = (inp[11]) ? node1112 : 3'b011;
											assign node1112 = (inp[2]) ? 3'b111 : 3'b011;
									assign node1115 = (inp[8]) ? node1121 : node1116;
										assign node1116 = (inp[5]) ? 3'b101 : node1117;
											assign node1117 = (inp[2]) ? 3'b001 : 3'b011;
										assign node1121 = (inp[2]) ? node1123 : 3'b011;
											assign node1123 = (inp[11]) ? 3'b011 : 3'b001;
							assign node1126 = (inp[10]) ? node1150 : node1127;
								assign node1127 = (inp[1]) ? node1139 : node1128;
									assign node1128 = (inp[8]) ? node1134 : node1129;
										assign node1129 = (inp[5]) ? node1131 : 3'b011;
											assign node1131 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1134 = (inp[5]) ? node1136 : 3'b111;
											assign node1136 = (inp[2]) ? 3'b011 : 3'b011;
									assign node1139 = (inp[5]) ? node1145 : node1140;
										assign node1140 = (inp[8]) ? 3'b011 : node1141;
											assign node1141 = (inp[11]) ? 3'b001 : 3'b011;
										assign node1145 = (inp[2]) ? node1147 : 3'b001;
											assign node1147 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1150 = (inp[2]) ? node1160 : node1151;
									assign node1151 = (inp[1]) ? node1157 : node1152;
										assign node1152 = (inp[8]) ? node1154 : 3'b101;
											assign node1154 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1157 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1160 = (inp[1]) ? node1166 : node1161;
										assign node1161 = (inp[11]) ? node1163 : 3'b111;
											assign node1163 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1166 = (inp[11]) ? 3'b110 : 3'b101;
				assign node1169 = (inp[9]) ? node1355 : node1170;
					assign node1170 = (inp[1]) ? node1248 : node1171;
						assign node1171 = (inp[7]) ? node1221 : node1172;
							assign node1172 = (inp[10]) ? node1194 : node1173;
								assign node1173 = (inp[4]) ? node1185 : node1174;
									assign node1174 = (inp[5]) ? node1180 : node1175;
										assign node1175 = (inp[8]) ? 3'b111 : node1176;
											assign node1176 = (inp[11]) ? 3'b011 : 3'b011;
										assign node1180 = (inp[2]) ? 3'b011 : node1181;
											assign node1181 = (inp[8]) ? 3'b011 : 3'b001;
									assign node1185 = (inp[5]) ? node1191 : node1186;
										assign node1186 = (inp[2]) ? 3'b101 : node1187;
											assign node1187 = (inp[8]) ? 3'b011 : 3'b111;
										assign node1191 = (inp[8]) ? 3'b101 : 3'b001;
								assign node1194 = (inp[4]) ? node1208 : node1195;
									assign node1195 = (inp[11]) ? node1203 : node1196;
										assign node1196 = (inp[2]) ? node1200 : node1197;
											assign node1197 = (inp[5]) ? 3'b011 : 3'b111;
											assign node1200 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1203 = (inp[5]) ? node1205 : 3'b101;
											assign node1205 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1208 = (inp[8]) ? node1214 : node1209;
										assign node1209 = (inp[2]) ? 3'b110 : node1210;
											assign node1210 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1214 = (inp[11]) ? node1218 : node1215;
											assign node1215 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1218 = (inp[5]) ? 3'b110 : 3'b101;
							assign node1221 = (inp[4]) ? node1231 : node1222;
								assign node1222 = (inp[11]) ? node1224 : 3'b111;
									assign node1224 = (inp[5]) ? node1226 : 3'b111;
										assign node1226 = (inp[10]) ? node1228 : 3'b111;
											assign node1228 = (inp[8]) ? 3'b011 : 3'b011;
								assign node1231 = (inp[5]) ? node1241 : node1232;
									assign node1232 = (inp[2]) ? node1234 : 3'b111;
										assign node1234 = (inp[8]) ? node1238 : node1235;
											assign node1235 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1238 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1241 = (inp[11]) ? 3'b101 : node1242;
										assign node1242 = (inp[8]) ? node1244 : 3'b111;
											assign node1244 = (inp[10]) ? 3'b001 : 3'b011;
						assign node1248 = (inp[4]) ? node1302 : node1249;
							assign node1249 = (inp[7]) ? node1281 : node1250;
								assign node1250 = (inp[10]) ? node1266 : node1251;
									assign node1251 = (inp[8]) ? node1259 : node1252;
										assign node1252 = (inp[5]) ? node1256 : node1253;
											assign node1253 = (inp[11]) ? 3'b001 : 3'b011;
											assign node1256 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1259 = (inp[11]) ? node1263 : node1260;
											assign node1260 = (inp[2]) ? 3'b011 : 3'b011;
											assign node1263 = (inp[5]) ? 3'b001 : 3'b010;
									assign node1266 = (inp[5]) ? node1274 : node1267;
										assign node1267 = (inp[8]) ? node1271 : node1268;
											assign node1268 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1271 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1274 = (inp[11]) ? node1278 : node1275;
											assign node1275 = (inp[8]) ? 3'b101 : 3'b001;
											assign node1278 = (inp[8]) ? 3'b001 : 3'b010;
								assign node1281 = (inp[2]) ? node1291 : node1282;
									assign node1282 = (inp[10]) ? node1288 : node1283;
										assign node1283 = (inp[11]) ? node1285 : 3'b111;
											assign node1285 = (inp[5]) ? 3'b111 : 3'b011;
										assign node1288 = (inp[5]) ? 3'b101 : 3'b111;
									assign node1291 = (inp[10]) ? node1295 : node1292;
										assign node1292 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1295 = (inp[5]) ? node1299 : node1296;
											assign node1296 = (inp[11]) ? 3'b011 : 3'b011;
											assign node1299 = (inp[8]) ? 3'b001 : 3'b101;
							assign node1302 = (inp[7]) ? node1326 : node1303;
								assign node1303 = (inp[10]) ? node1315 : node1304;
									assign node1304 = (inp[8]) ? node1310 : node1305;
										assign node1305 = (inp[5]) ? 3'b110 : node1306;
											assign node1306 = (inp[11]) ? 3'b001 : 3'b001;
										assign node1310 = (inp[5]) ? 3'b001 : node1311;
											assign node1311 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1315 = (inp[8]) ? node1321 : node1316;
										assign node1316 = (inp[2]) ? node1318 : 3'b110;
											assign node1318 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1321 = (inp[2]) ? 3'b110 : node1322;
											assign node1322 = (inp[5]) ? 3'b110 : 3'b000;
								assign node1326 = (inp[11]) ? node1340 : node1327;
									assign node1327 = (inp[2]) ? node1333 : node1328;
										assign node1328 = (inp[10]) ? node1330 : 3'b101;
											assign node1330 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1333 = (inp[5]) ? node1337 : node1334;
											assign node1334 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1337 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1340 = (inp[2]) ? node1348 : node1341;
										assign node1341 = (inp[8]) ? node1345 : node1342;
											assign node1342 = (inp[5]) ? 3'b000 : 3'b001;
											assign node1345 = (inp[5]) ? 3'b001 : 3'b000;
										assign node1348 = (inp[10]) ? node1352 : node1349;
											assign node1349 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1352 = (inp[5]) ? 3'b110 : 3'b001;
					assign node1355 = (inp[4]) ? node1455 : node1356;
						assign node1356 = (inp[10]) ? node1406 : node1357;
							assign node1357 = (inp[11]) ? node1381 : node1358;
								assign node1358 = (inp[8]) ? node1368 : node1359;
									assign node1359 = (inp[7]) ? node1361 : 3'b001;
										assign node1361 = (inp[1]) ? node1365 : node1362;
											assign node1362 = (inp[5]) ? 3'b101 : 3'b011;
											assign node1365 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1368 = (inp[7]) ? node1374 : node1369;
										assign node1369 = (inp[2]) ? 3'b001 : node1370;
											assign node1370 = (inp[1]) ? 3'b101 : 3'b001;
										assign node1374 = (inp[5]) ? node1378 : node1375;
											assign node1375 = (inp[1]) ? 3'b011 : 3'b111;
											assign node1378 = (inp[1]) ? 3'b101 : 3'b011;
								assign node1381 = (inp[7]) ? node1393 : node1382;
									assign node1382 = (inp[5]) ? node1388 : node1383;
										assign node1383 = (inp[2]) ? 3'b001 : node1384;
											assign node1384 = (inp[1]) ? 3'b000 : 3'b101;
										assign node1388 = (inp[1]) ? node1390 : 3'b110;
											assign node1390 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1393 = (inp[2]) ? node1401 : node1394;
										assign node1394 = (inp[5]) ? node1398 : node1395;
											assign node1395 = (inp[8]) ? 3'b111 : 3'b011;
											assign node1398 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1401 = (inp[1]) ? node1403 : 3'b011;
											assign node1403 = (inp[8]) ? 3'b101 : 3'b001;
							assign node1406 = (inp[7]) ? node1430 : node1407;
								assign node1407 = (inp[8]) ? node1417 : node1408;
									assign node1408 = (inp[5]) ? node1410 : 3'b110;
										assign node1410 = (inp[2]) ? node1414 : node1411;
											assign node1411 = (inp[1]) ? 3'b010 : 3'b110;
											assign node1414 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1417 = (inp[1]) ? node1425 : node1418;
										assign node1418 = (inp[5]) ? node1422 : node1419;
											assign node1419 = (inp[11]) ? 3'b001 : 3'b001;
											assign node1422 = (inp[2]) ? 3'b110 : 3'b000;
										assign node1425 = (inp[2]) ? node1427 : 3'b010;
											assign node1427 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1430 = (inp[1]) ? node1444 : node1431;
									assign node1431 = (inp[11]) ? node1437 : node1432;
										assign node1432 = (inp[8]) ? 3'b011 : node1433;
											assign node1433 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1437 = (inp[5]) ? node1441 : node1438;
											assign node1438 = (inp[2]) ? 3'b101 : 3'b011;
											assign node1441 = (inp[2]) ? 3'b001 : 3'b001;
									assign node1444 = (inp[8]) ? node1450 : node1445;
										assign node1445 = (inp[11]) ? node1447 : 3'b010;
											assign node1447 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1450 = (inp[11]) ? node1452 : 3'b101;
											assign node1452 = (inp[2]) ? 3'b000 : 3'b001;
						assign node1455 = (inp[7]) ? node1503 : node1456;
							assign node1456 = (inp[1]) ? node1482 : node1457;
								assign node1457 = (inp[2]) ? node1471 : node1458;
									assign node1458 = (inp[10]) ? node1464 : node1459;
										assign node1459 = (inp[5]) ? node1461 : 3'b001;
											assign node1461 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1464 = (inp[5]) ? node1468 : node1465;
											assign node1465 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1468 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1471 = (inp[10]) ? node1477 : node1472;
										assign node1472 = (inp[11]) ? node1474 : 3'b110;
											assign node1474 = (inp[8]) ? 3'b010 : 3'b010;
										assign node1477 = (inp[11]) ? node1479 : 3'b010;
											assign node1479 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1482 = (inp[5]) ? node1494 : node1483;
									assign node1483 = (inp[10]) ? node1489 : node1484;
										assign node1484 = (inp[8]) ? node1486 : 3'b010;
											assign node1486 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1489 = (inp[11]) ? node1491 : 3'b010;
											assign node1491 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1494 = (inp[2]) ? node1496 : 3'b100;
										assign node1496 = (inp[10]) ? node1500 : node1497;
											assign node1497 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1500 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1503 = (inp[10]) ? node1519 : node1504;
								assign node1504 = (inp[1]) ? node1508 : node1505;
									assign node1505 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1508 = (inp[5]) ? node1514 : node1509;
										assign node1509 = (inp[11]) ? 3'b000 : node1510;
											assign node1510 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1514 = (inp[8]) ? node1516 : 3'b110;
											assign node1516 = (inp[11]) ? 3'b010 : 3'b001;
								assign node1519 = (inp[1]) ? node1531 : node1520;
									assign node1520 = (inp[8]) ? node1526 : node1521;
										assign node1521 = (inp[11]) ? node1523 : 3'b110;
											assign node1523 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1526 = (inp[5]) ? 3'b110 : node1527;
											assign node1527 = (inp[2]) ? 3'b011 : 3'b001;
									assign node1531 = (inp[5]) ? node1535 : node1532;
										assign node1532 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1535 = (inp[8]) ? 3'b010 : node1536;
											assign node1536 = (inp[11]) ? 3'b000 : 3'b010;
			assign node1540 = (inp[9]) ? node1906 : node1541;
				assign node1541 = (inp[7]) ? node1731 : node1542;
					assign node1542 = (inp[4]) ? node1634 : node1543;
						assign node1543 = (inp[10]) ? node1589 : node1544;
							assign node1544 = (inp[5]) ? node1570 : node1545;
								assign node1545 = (inp[0]) ? node1555 : node1546;
									assign node1546 = (inp[1]) ? node1548 : 3'b101;
										assign node1548 = (inp[11]) ? node1552 : node1549;
											assign node1549 = (inp[2]) ? 3'b001 : 3'b011;
											assign node1552 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1555 = (inp[1]) ? node1563 : node1556;
										assign node1556 = (inp[11]) ? node1560 : node1557;
											assign node1557 = (inp[8]) ? 3'b001 : 3'b001;
											assign node1560 = (inp[2]) ? 3'b001 : 3'b001;
										assign node1563 = (inp[11]) ? node1567 : node1564;
											assign node1564 = (inp[2]) ? 3'b110 : 3'b001;
											assign node1567 = (inp[8]) ? 3'b110 : 3'b100;
								assign node1570 = (inp[1]) ? node1578 : node1571;
									assign node1571 = (inp[2]) ? 3'b110 : node1572;
										assign node1572 = (inp[8]) ? 3'b100 : node1573;
											assign node1573 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1578 = (inp[0]) ? node1584 : node1579;
										assign node1579 = (inp[11]) ? node1581 : 3'b001;
											assign node1581 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1584 = (inp[8]) ? node1586 : 3'b010;
											assign node1586 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1589 = (inp[0]) ? node1609 : node1590;
								assign node1590 = (inp[2]) ? node1598 : node1591;
									assign node1591 = (inp[8]) ? node1593 : 3'b110;
										assign node1593 = (inp[5]) ? 3'b110 : node1594;
											assign node1594 = (inp[1]) ? 3'b001 : 3'b100;
									assign node1598 = (inp[11]) ? node1604 : node1599;
										assign node1599 = (inp[1]) ? 3'b110 : node1600;
											assign node1600 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1604 = (inp[8]) ? 3'b110 : node1605;
											assign node1605 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1609 = (inp[5]) ? node1625 : node1610;
									assign node1610 = (inp[8]) ? node1618 : node1611;
										assign node1611 = (inp[11]) ? node1615 : node1612;
											assign node1612 = (inp[1]) ? 3'b010 : 3'b110;
											assign node1615 = (inp[1]) ? 3'b000 : 3'b010;
										assign node1618 = (inp[1]) ? node1622 : node1619;
											assign node1619 = (inp[2]) ? 3'b110 : 3'b100;
											assign node1622 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1625 = (inp[8]) ? node1627 : 3'b100;
										assign node1627 = (inp[11]) ? node1631 : node1628;
											assign node1628 = (inp[1]) ? 3'b010 : 3'b110;
											assign node1631 = (inp[1]) ? 3'b100 : 3'b010;
						assign node1634 = (inp[10]) ? node1684 : node1635;
							assign node1635 = (inp[2]) ? node1657 : node1636;
								assign node1636 = (inp[0]) ? node1648 : node1637;
									assign node1637 = (inp[8]) ? node1643 : node1638;
										assign node1638 = (inp[1]) ? node1640 : 3'b110;
											assign node1640 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1643 = (inp[1]) ? node1645 : 3'b000;
											assign node1645 = (inp[5]) ? 3'b110 : 3'b000;
									assign node1648 = (inp[1]) ? 3'b100 : node1649;
										assign node1649 = (inp[5]) ? node1653 : node1650;
											assign node1650 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1653 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1657 = (inp[11]) ? node1671 : node1658;
									assign node1658 = (inp[1]) ? node1666 : node1659;
										assign node1659 = (inp[0]) ? node1663 : node1660;
											assign node1660 = (inp[8]) ? 3'b000 : 3'b110;
											assign node1663 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1666 = (inp[0]) ? node1668 : 3'b110;
											assign node1668 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1671 = (inp[0]) ? node1679 : node1672;
										assign node1672 = (inp[1]) ? node1676 : node1673;
											assign node1673 = (inp[8]) ? 3'b000 : 3'b110;
											assign node1676 = (inp[8]) ? 3'b010 : 3'b010;
										assign node1679 = (inp[8]) ? 3'b010 : node1680;
											assign node1680 = (inp[5]) ? 3'b000 : 3'b010;
							assign node1684 = (inp[0]) ? node1712 : node1685;
								assign node1685 = (inp[5]) ? node1701 : node1686;
									assign node1686 = (inp[8]) ? node1694 : node1687;
										assign node1687 = (inp[1]) ? node1691 : node1688;
											assign node1688 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1691 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1694 = (inp[1]) ? node1698 : node1695;
											assign node1695 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1698 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1701 = (inp[8]) ? node1707 : node1702;
										assign node1702 = (inp[11]) ? 3'b100 : node1703;
											assign node1703 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1707 = (inp[1]) ? 3'b100 : node1708;
											assign node1708 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1712 = (inp[1]) ? node1724 : node1713;
									assign node1713 = (inp[5]) ? node1719 : node1714;
										assign node1714 = (inp[8]) ? node1716 : 3'b100;
											assign node1716 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1719 = (inp[8]) ? 3'b100 : node1720;
											assign node1720 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1724 = (inp[11]) ? 3'b000 : node1725;
										assign node1725 = (inp[8]) ? node1727 : 3'b000;
											assign node1727 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1731 = (inp[0]) ? node1823 : node1732;
						assign node1732 = (inp[4]) ? node1772 : node1733;
							assign node1733 = (inp[1]) ? node1747 : node1734;
								assign node1734 = (inp[10]) ? node1742 : node1735;
									assign node1735 = (inp[11]) ? node1737 : 3'b111;
										assign node1737 = (inp[2]) ? node1739 : 3'b111;
											assign node1739 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1742 = (inp[11]) ? 3'b011 : node1743;
										assign node1743 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1747 = (inp[10]) ? node1759 : node1748;
									assign node1748 = (inp[8]) ? node1754 : node1749;
										assign node1749 = (inp[5]) ? 3'b101 : node1750;
											assign node1750 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1754 = (inp[11]) ? 3'b011 : node1755;
											assign node1755 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1759 = (inp[2]) ? node1765 : node1760;
										assign node1760 = (inp[11]) ? node1762 : 3'b101;
											assign node1762 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1765 = (inp[8]) ? node1769 : node1766;
											assign node1766 = (inp[5]) ? 3'b001 : 3'b001;
											assign node1769 = (inp[5]) ? 3'b001 : 3'b011;
							assign node1772 = (inp[8]) ? node1796 : node1773;
								assign node1773 = (inp[11]) ? node1785 : node1774;
									assign node1774 = (inp[1]) ? node1782 : node1775;
										assign node1775 = (inp[5]) ? node1779 : node1776;
											assign node1776 = (inp[2]) ? 3'b011 : 3'b101;
											assign node1779 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1782 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1785 = (inp[10]) ? node1791 : node1786;
										assign node1786 = (inp[1]) ? 3'b110 : node1787;
											assign node1787 = (inp[5]) ? 3'b001 : 3'b100;
										assign node1791 = (inp[5]) ? node1793 : 3'b110;
											assign node1793 = (inp[1]) ? 3'b010 : 3'b110;
								assign node1796 = (inp[2]) ? node1810 : node1797;
									assign node1797 = (inp[10]) ? node1803 : node1798;
										assign node1798 = (inp[5]) ? node1800 : 3'b011;
											assign node1800 = (inp[11]) ? 3'b001 : 3'b011;
										assign node1803 = (inp[11]) ? node1807 : node1804;
											assign node1804 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1807 = (inp[5]) ? 3'b000 : 3'b001;
									assign node1810 = (inp[10]) ? node1816 : node1811;
										assign node1811 = (inp[5]) ? node1813 : 3'b101;
											assign node1813 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1816 = (inp[1]) ? node1820 : node1817;
											assign node1817 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1820 = (inp[5]) ? 3'b110 : 3'b001;
						assign node1823 = (inp[4]) ? node1869 : node1824;
							assign node1824 = (inp[10]) ? node1846 : node1825;
								assign node1825 = (inp[8]) ? node1835 : node1826;
									assign node1826 = (inp[5]) ? node1832 : node1827;
										assign node1827 = (inp[11]) ? 3'b001 : node1828;
											assign node1828 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1832 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1835 = (inp[5]) ? node1841 : node1836;
										assign node1836 = (inp[1]) ? node1838 : 3'b011;
											assign node1838 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1841 = (inp[1]) ? 3'b001 : node1842;
											assign node1842 = (inp[2]) ? 3'b001 : 3'b101;
								assign node1846 = (inp[8]) ? node1858 : node1847;
									assign node1847 = (inp[5]) ? node1853 : node1848;
										assign node1848 = (inp[1]) ? 3'b110 : node1849;
											assign node1849 = (inp[11]) ? 3'b000 : 3'b001;
										assign node1853 = (inp[2]) ? 3'b110 : node1854;
											assign node1854 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1858 = (inp[5]) ? node1864 : node1859;
										assign node1859 = (inp[1]) ? node1861 : 3'b101;
											assign node1861 = (inp[11]) ? 3'b010 : 3'b001;
										assign node1864 = (inp[1]) ? 3'b110 : node1865;
											assign node1865 = (inp[2]) ? 3'b000 : 3'b001;
							assign node1869 = (inp[8]) ? node1887 : node1870;
								assign node1870 = (inp[10]) ? node1880 : node1871;
									assign node1871 = (inp[5]) ? node1875 : node1872;
										assign node1872 = (inp[1]) ? 3'b100 : 3'b110;
										assign node1875 = (inp[2]) ? node1877 : 3'b010;
											assign node1877 = (inp[1]) ? 3'b000 : 3'b010;
									assign node1880 = (inp[5]) ? node1884 : node1881;
										assign node1881 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1884 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1887 = (inp[11]) ? node1893 : node1888;
									assign node1888 = (inp[1]) ? node1890 : 3'b110;
										assign node1890 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1893 = (inp[1]) ? node1901 : node1894;
										assign node1894 = (inp[5]) ? node1898 : node1895;
											assign node1895 = (inp[10]) ? 3'b110 : 3'b001;
											assign node1898 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1901 = (inp[5]) ? node1903 : 3'b110;
											assign node1903 = (inp[2]) ? 3'b100 : 3'b110;
				assign node1906 = (inp[0]) ? node2094 : node1907;
					assign node1907 = (inp[1]) ? node1989 : node1908;
						assign node1908 = (inp[7]) ? node1950 : node1909;
							assign node1909 = (inp[4]) ? node1929 : node1910;
								assign node1910 = (inp[10]) ? node1924 : node1911;
									assign node1911 = (inp[2]) ? node1919 : node1912;
										assign node1912 = (inp[11]) ? node1916 : node1913;
											assign node1913 = (inp[5]) ? 3'b000 : 3'b001;
											assign node1916 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1919 = (inp[5]) ? node1921 : 3'b111;
											assign node1921 = (inp[8]) ? 3'b110 : 3'b110;
									assign node1924 = (inp[11]) ? 3'b010 : node1925;
										assign node1925 = (inp[5]) ? 3'b110 : 3'b011;
								assign node1929 = (inp[5]) ? node1943 : node1930;
									assign node1930 = (inp[8]) ? node1936 : node1931;
										assign node1931 = (inp[10]) ? 3'b110 : node1932;
											assign node1932 = (inp[11]) ? 3'b010 : 3'b010;
										assign node1936 = (inp[10]) ? node1940 : node1937;
											assign node1937 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1940 = (inp[2]) ? 3'b010 : 3'b010;
									assign node1943 = (inp[10]) ? node1947 : node1944;
										assign node1944 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1947 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1950 = (inp[10]) ? node1972 : node1951;
								assign node1951 = (inp[4]) ? node1959 : node1952;
									assign node1952 = (inp[11]) ? 3'b101 : node1953;
										assign node1953 = (inp[8]) ? node1955 : 3'b001;
											assign node1955 = (inp[5]) ? 3'b101 : 3'b011;
									assign node1959 = (inp[5]) ? node1965 : node1960;
										assign node1960 = (inp[11]) ? node1962 : 3'b001;
											assign node1962 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1965 = (inp[8]) ? node1969 : node1966;
											assign node1966 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1969 = (inp[2]) ? 3'b110 : 3'b001;
								assign node1972 = (inp[11]) ? node1984 : node1973;
									assign node1973 = (inp[4]) ? node1979 : node1974;
										assign node1974 = (inp[8]) ? node1976 : 3'b110;
											assign node1976 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1979 = (inp[5]) ? node1981 : 3'b110;
											assign node1981 = (inp[2]) ? 3'b010 : 3'b010;
									assign node1984 = (inp[4]) ? 3'b010 : node1985;
										assign node1985 = (inp[8]) ? 3'b001 : 3'b000;
						assign node1989 = (inp[7]) ? node2039 : node1990;
							assign node1990 = (inp[4]) ? node2020 : node1991;
								assign node1991 = (inp[2]) ? node2005 : node1992;
									assign node1992 = (inp[11]) ? node2000 : node1993;
										assign node1993 = (inp[5]) ? node1997 : node1994;
											assign node1994 = (inp[10]) ? 3'b000 : 3'b111;
											assign node1997 = (inp[10]) ? 3'b100 : 3'b000;
										assign node2000 = (inp[10]) ? 3'b100 : node2001;
											assign node2001 = (inp[5]) ? 3'b100 : 3'b110;
									assign node2005 = (inp[11]) ? node2013 : node2006;
										assign node2006 = (inp[10]) ? node2010 : node2007;
											assign node2007 = (inp[5]) ? 3'b000 : 3'b100;
											assign node2010 = (inp[5]) ? 3'b110 : 3'b010;
										assign node2013 = (inp[10]) ? node2017 : node2014;
											assign node2014 = (inp[5]) ? 3'b010 : 3'b000;
											assign node2017 = (inp[8]) ? 3'b000 : 3'b000;
								assign node2020 = (inp[8]) ? node2028 : node2021;
									assign node2021 = (inp[5]) ? 3'b000 : node2022;
										assign node2022 = (inp[10]) ? 3'b000 : node2023;
											assign node2023 = (inp[11]) ? 3'b000 : 3'b100;
									assign node2028 = (inp[10]) ? node2036 : node2029;
										assign node2029 = (inp[5]) ? node2033 : node2030;
											assign node2030 = (inp[11]) ? 3'b100 : 3'b000;
											assign node2033 = (inp[11]) ? 3'b000 : 3'b100;
										assign node2036 = (inp[5]) ? 3'b000 : 3'b100;
							assign node2039 = (inp[11]) ? node2065 : node2040;
								assign node2040 = (inp[10]) ? node2052 : node2041;
									assign node2041 = (inp[2]) ? node2047 : node2042;
										assign node2042 = (inp[8]) ? 3'b001 : node2043;
											assign node2043 = (inp[5]) ? 3'b010 : 3'b011;
										assign node2047 = (inp[4]) ? node2049 : 3'b110;
											assign node2049 = (inp[8]) ? 3'b010 : 3'b010;
									assign node2052 = (inp[4]) ? node2060 : node2053;
										assign node2053 = (inp[8]) ? node2057 : node2054;
											assign node2054 = (inp[5]) ? 3'b001 : 3'b110;
											assign node2057 = (inp[5]) ? 3'b110 : 3'b001;
										assign node2060 = (inp[8]) ? node2062 : 3'b100;
											assign node2062 = (inp[2]) ? 3'b000 : 3'b010;
								assign node2065 = (inp[4]) ? node2079 : node2066;
									assign node2066 = (inp[8]) ? node2074 : node2067;
										assign node2067 = (inp[10]) ? node2071 : node2068;
											assign node2068 = (inp[2]) ? 3'b110 : 3'b010;
											assign node2071 = (inp[5]) ? 3'b010 : 3'b010;
										assign node2074 = (inp[2]) ? 3'b110 : node2075;
											assign node2075 = (inp[10]) ? 3'b000 : 3'b001;
									assign node2079 = (inp[8]) ? node2087 : node2080;
										assign node2080 = (inp[2]) ? node2084 : node2081;
											assign node2081 = (inp[5]) ? 3'b100 : 3'b100;
											assign node2084 = (inp[5]) ? 3'b000 : 3'b010;
										assign node2087 = (inp[10]) ? node2091 : node2088;
											assign node2088 = (inp[5]) ? 3'b010 : 3'b110;
											assign node2091 = (inp[5]) ? 3'b100 : 3'b010;
					assign node2094 = (inp[7]) ? node2126 : node2095;
						assign node2095 = (inp[4]) ? 3'b000 : node2096;
							assign node2096 = (inp[10]) ? node2116 : node2097;
								assign node2097 = (inp[5]) ? node2109 : node2098;
									assign node2098 = (inp[1]) ? node2104 : node2099;
										assign node2099 = (inp[11]) ? 3'b100 : node2100;
											assign node2100 = (inp[2]) ? 3'b010 : 3'b010;
										assign node2104 = (inp[11]) ? node2106 : 3'b100;
											assign node2106 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2109 = (inp[8]) ? node2111 : 3'b000;
										assign node2111 = (inp[11]) ? node2113 : 3'b100;
											assign node2113 = (inp[1]) ? 3'b000 : 3'b100;
								assign node2116 = (inp[1]) ? 3'b000 : node2117;
									assign node2117 = (inp[5]) ? 3'b000 : node2118;
										assign node2118 = (inp[2]) ? 3'b100 : node2119;
											assign node2119 = (inp[11]) ? 3'b000 : 3'b010;
						assign node2126 = (inp[1]) ? node2178 : node2127;
							assign node2127 = (inp[4]) ? node2151 : node2128;
								assign node2128 = (inp[8]) ? node2140 : node2129;
									assign node2129 = (inp[10]) ? node2135 : node2130;
										assign node2130 = (inp[5]) ? 3'b010 : node2131;
											assign node2131 = (inp[11]) ? 3'b010 : 3'b010;
										assign node2135 = (inp[5]) ? node2137 : 3'b010;
											assign node2137 = (inp[2]) ? 3'b100 : 3'b000;
									assign node2140 = (inp[5]) ? node2144 : node2141;
										assign node2141 = (inp[10]) ? 3'b110 : 3'b001;
										assign node2144 = (inp[10]) ? node2148 : node2145;
											assign node2145 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2148 = (inp[2]) ? 3'b100 : 3'b010;
								assign node2151 = (inp[11]) ? node2165 : node2152;
									assign node2152 = (inp[2]) ? node2160 : node2153;
										assign node2153 = (inp[8]) ? node2157 : node2154;
											assign node2154 = (inp[10]) ? 3'b110 : 3'b010;
											assign node2157 = (inp[5]) ? 3'b010 : 3'b010;
										assign node2160 = (inp[10]) ? 3'b100 : node2161;
											assign node2161 = (inp[5]) ? 3'b100 : 3'b010;
									assign node2165 = (inp[5]) ? node2173 : node2166;
										assign node2166 = (inp[8]) ? node2170 : node2167;
											assign node2167 = (inp[10]) ? 3'b000 : 3'b100;
											assign node2170 = (inp[10]) ? 3'b100 : 3'b010;
										assign node2173 = (inp[8]) ? node2175 : 3'b000;
											assign node2175 = (inp[10]) ? 3'b000 : 3'b100;
							assign node2178 = (inp[4]) ? node2202 : node2179;
								assign node2179 = (inp[10]) ? node2189 : node2180;
									assign node2180 = (inp[8]) ? node2184 : node2181;
										assign node2181 = (inp[5]) ? 3'b100 : 3'b010;
										assign node2184 = (inp[5]) ? 3'b010 : node2185;
											assign node2185 = (inp[2]) ? 3'b010 : 3'b110;
									assign node2189 = (inp[11]) ? node2195 : node2190;
										assign node2190 = (inp[8]) ? node2192 : 3'b100;
											assign node2192 = (inp[5]) ? 3'b100 : 3'b010;
										assign node2195 = (inp[8]) ? node2199 : node2196;
											assign node2196 = (inp[5]) ? 3'b000 : 3'b100;
											assign node2199 = (inp[2]) ? 3'b100 : 3'b000;
								assign node2202 = (inp[10]) ? 3'b000 : node2203;
									assign node2203 = (inp[11]) ? node2209 : node2204;
										assign node2204 = (inp[8]) ? 3'b100 : node2205;
											assign node2205 = (inp[5]) ? 3'b000 : 3'b100;
										assign node2209 = (inp[5]) ? 3'b000 : node2210;
											assign node2210 = (inp[8]) ? 3'b100 : 3'b000;

endmodule