module dtc_split05_bm23 (
	input  wire [12-1:0] inp,
	output wire [12-1:0] outp
);

	wire [12-1:0] node1;
	wire [12-1:0] node2;
	wire [12-1:0] node3;
	wire [12-1:0] node4;
	wire [12-1:0] node5;
	wire [12-1:0] node7;
	wire [12-1:0] node8;
	wire [12-1:0] node11;
	wire [12-1:0] node14;
	wire [12-1:0] node15;
	wire [12-1:0] node16;
	wire [12-1:0] node20;
	wire [12-1:0] node23;
	wire [12-1:0] node24;
	wire [12-1:0] node26;
	wire [12-1:0] node27;
	wire [12-1:0] node31;
	wire [12-1:0] node33;
	wire [12-1:0] node36;
	wire [12-1:0] node37;
	wire [12-1:0] node38;
	wire [12-1:0] node39;
	wire [12-1:0] node40;
	wire [12-1:0] node44;
	wire [12-1:0] node45;
	wire [12-1:0] node48;
	wire [12-1:0] node52;
	wire [12-1:0] node53;
	wire [12-1:0] node54;
	wire [12-1:0] node58;
	wire [12-1:0] node60;
	wire [12-1:0] node63;
	wire [12-1:0] node64;
	wire [12-1:0] node65;
	wire [12-1:0] node66;
	wire [12-1:0] node67;
	wire [12-1:0] node69;
	wire [12-1:0] node72;
	wire [12-1:0] node73;
	wire [12-1:0] node76;
	wire [12-1:0] node80;
	wire [12-1:0] node81;
	wire [12-1:0] node82;
	wire [12-1:0] node85;
	wire [12-1:0] node86;
	wire [12-1:0] node89;
	wire [12-1:0] node92;
	wire [12-1:0] node93;
	wire [12-1:0] node97;
	wire [12-1:0] node98;
	wire [12-1:0] node99;
	wire [12-1:0] node100;
	wire [12-1:0] node103;
	wire [12-1:0] node106;
	wire [12-1:0] node108;
	wire [12-1:0] node111;
	wire [12-1:0] node112;
	wire [12-1:0] node113;
	wire [12-1:0] node115;
	wire [12-1:0] node118;
	wire [12-1:0] node120;
	wire [12-1:0] node123;
	wire [12-1:0] node124;
	wire [12-1:0] node125;
	wire [12-1:0] node130;
	wire [12-1:0] node131;
	wire [12-1:0] node132;
	wire [12-1:0] node133;
	wire [12-1:0] node134;
	wire [12-1:0] node137;
	wire [12-1:0] node140;
	wire [12-1:0] node141;
	wire [12-1:0] node143;
	wire [12-1:0] node144;
	wire [12-1:0] node148;
	wire [12-1:0] node149;
	wire [12-1:0] node151;
	wire [12-1:0] node155;
	wire [12-1:0] node156;
	wire [12-1:0] node157;
	wire [12-1:0] node158;
	wire [12-1:0] node161;
	wire [12-1:0] node162;
	wire [12-1:0] node165;
	wire [12-1:0] node168;
	wire [12-1:0] node170;
	wire [12-1:0] node172;
	wire [12-1:0] node175;
	wire [12-1:0] node176;
	wire [12-1:0] node179;
	wire [12-1:0] node180;
	wire [12-1:0] node183;
	wire [12-1:0] node186;
	wire [12-1:0] node187;
	wire [12-1:0] node188;
	wire [12-1:0] node189;
	wire [12-1:0] node190;
	wire [12-1:0] node193;
	wire [12-1:0] node196;
	wire [12-1:0] node198;
	wire [12-1:0] node199;
	wire [12-1:0] node202;
	wire [12-1:0] node205;
	wire [12-1:0] node206;
	wire [12-1:0] node208;
	wire [12-1:0] node209;
	wire [12-1:0] node212;
	wire [12-1:0] node215;
	wire [12-1:0] node216;
	wire [12-1:0] node217;
	wire [12-1:0] node221;
	wire [12-1:0] node224;
	wire [12-1:0] node225;
	wire [12-1:0] node226;
	wire [12-1:0] node227;
	wire [12-1:0] node229;
	wire [12-1:0] node232;
	wire [12-1:0] node234;
	wire [12-1:0] node237;
	wire [12-1:0] node238;
	wire [12-1:0] node241;
	wire [12-1:0] node244;
	wire [12-1:0] node245;
	wire [12-1:0] node246;
	wire [12-1:0] node249;
	wire [12-1:0] node252;
	wire [12-1:0] node253;
	wire [12-1:0] node256;
	wire [12-1:0] node258;

	assign outp = (inp[11]) ? node130 : node1;
		assign node1 = (inp[5]) ? node63 : node2;
			assign node2 = (inp[9]) ? node36 : node3;
				assign node3 = (inp[10]) ? node23 : node4;
					assign node4 = (inp[4]) ? node14 : node5;
						assign node5 = (inp[8]) ? node7 : 12'b001111111111;
							assign node7 = (inp[0]) ? node11 : node8;
								assign node8 = (inp[7]) ? 12'b001111111111 : 12'b000111111111;
								assign node11 = (inp[6]) ? 12'b000001111111 : 12'b000111111111;
						assign node14 = (inp[1]) ? node20 : node15;
							assign node15 = (inp[6]) ? 12'b000011111111 : node16;
								assign node16 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
							assign node20 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
					assign node23 = (inp[7]) ? node31 : node24;
						assign node24 = (inp[0]) ? node26 : 12'b000111111111;
							assign node26 = (inp[3]) ? 12'b000001111111 : node27;
								assign node27 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
						assign node31 = (inp[6]) ? node33 : 12'b000001111111;
							assign node33 = (inp[3]) ? 12'b000000111111 : 12'b000011111111;
				assign node36 = (inp[0]) ? node52 : node37;
					assign node37 = (inp[3]) ? 12'b000001111111 : node38;
						assign node38 = (inp[10]) ? node44 : node39;
							assign node39 = (inp[6]) ? 12'b000001111111 : node40;
								assign node40 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
							assign node44 = (inp[7]) ? node48 : node45;
								assign node45 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
								assign node48 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
					assign node52 = (inp[1]) ? node58 : node53;
						assign node53 = (inp[10]) ? 12'b000000111111 : node54;
							assign node54 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
						assign node58 = (inp[8]) ? node60 : 12'b000000111111;
							assign node60 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
			assign node63 = (inp[3]) ? node97 : node64;
				assign node64 = (inp[8]) ? node80 : node65;
					assign node65 = (inp[1]) ? 12'b000000011111 : node66;
						assign node66 = (inp[10]) ? node72 : node67;
							assign node67 = (inp[7]) ? node69 : 12'b000111111111;
								assign node69 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
							assign node72 = (inp[7]) ? node76 : node73;
								assign node73 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node76 = (inp[9]) ? 12'b000001111111 : 12'b000000111111;
					assign node80 = (inp[0]) ? node92 : node81;
						assign node81 = (inp[6]) ? node85 : node82;
							assign node82 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
							assign node85 = (inp[4]) ? node89 : node86;
								assign node86 = (inp[1]) ? 12'b000000111111 : 12'b000011111111;
								assign node89 = (inp[10]) ? 12'b000000111111 : 12'b000000011111;
						assign node92 = (inp[1]) ? 12'b000000000011 : node93;
							assign node93 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
				assign node97 = (inp[2]) ? node111 : node98;
					assign node98 = (inp[7]) ? node106 : node99;
						assign node99 = (inp[6]) ? node103 : node100;
							assign node100 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
							assign node103 = (inp[4]) ? 12'b000001111111 : 12'b000000111111;
						assign node106 = (inp[4]) ? node108 : 12'b000000111111;
							assign node108 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
					assign node111 = (inp[0]) ? node123 : node112;
						assign node112 = (inp[10]) ? node118 : node113;
							assign node113 = (inp[4]) ? node115 : 12'b000001111111;
								assign node115 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
							assign node118 = (inp[1]) ? node120 : 12'b000000111111;
								assign node120 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
						assign node123 = (inp[8]) ? 12'b000000001111 : node124;
							assign node124 = (inp[6]) ? 12'b000000011111 : node125;
								assign node125 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
		assign node130 = (inp[7]) ? node186 : node131;
			assign node131 = (inp[10]) ? node155 : node132;
				assign node132 = (inp[4]) ? node140 : node133;
					assign node133 = (inp[1]) ? node137 : node134;
						assign node134 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
						assign node137 = (inp[6]) ? 12'b000011111111 : 12'b000001111111;
					assign node140 = (inp[5]) ? node148 : node141;
						assign node141 = (inp[2]) ? node143 : 12'b000001111111;
							assign node143 = (inp[1]) ? 12'b000000011111 : node144;
								assign node144 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
						assign node148 = (inp[6]) ? 12'b000000011111 : node149;
							assign node149 = (inp[3]) ? node151 : 12'b000000111111;
								assign node151 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
				assign node155 = (inp[0]) ? node175 : node156;
					assign node156 = (inp[2]) ? node168 : node157;
						assign node157 = (inp[3]) ? node161 : node158;
							assign node158 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
							assign node161 = (inp[9]) ? node165 : node162;
								assign node162 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
								assign node165 = (inp[4]) ? 12'b000000111111 : 12'b000000011111;
						assign node168 = (inp[8]) ? node170 : 12'b000000111111;
							assign node170 = (inp[5]) ? node172 : 12'b000000111111;
								assign node172 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
					assign node175 = (inp[3]) ? node179 : node176;
						assign node176 = (inp[4]) ? 12'b000000011111 : 12'b000001111111;
						assign node179 = (inp[4]) ? node183 : node180;
							assign node180 = (inp[1]) ? 12'b000000001111 : 12'b000000111111;
							assign node183 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
			assign node186 = (inp[4]) ? node224 : node187;
				assign node187 = (inp[3]) ? node205 : node188;
					assign node188 = (inp[10]) ? node196 : node189;
						assign node189 = (inp[0]) ? node193 : node190;
							assign node190 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
							assign node193 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
						assign node196 = (inp[5]) ? node198 : 12'b000000111111;
							assign node198 = (inp[6]) ? node202 : node199;
								assign node199 = (inp[2]) ? 12'b000000011111 : 12'b000000011111;
								assign node202 = (inp[0]) ? 12'b000000000011 : 12'b000000001111;
					assign node205 = (inp[1]) ? node215 : node206;
						assign node206 = (inp[0]) ? node208 : 12'b000000001111;
							assign node208 = (inp[8]) ? node212 : node209;
								assign node209 = (inp[9]) ? 12'b000000011111 : 12'b000001111111;
								assign node212 = (inp[5]) ? 12'b000000011111 : 12'b000000011111;
						assign node215 = (inp[5]) ? node221 : node216;
							assign node216 = (inp[0]) ? 12'b000000001111 : node217;
								assign node217 = (inp[8]) ? 12'b000000111111 : 12'b000000011111;
							assign node221 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
				assign node224 = (inp[1]) ? node244 : node225;
					assign node225 = (inp[5]) ? node237 : node226;
						assign node226 = (inp[8]) ? node232 : node227;
							assign node227 = (inp[10]) ? node229 : 12'b000001111111;
								assign node229 = (inp[0]) ? 12'b000000111111 : 12'b000000011111;
							assign node232 = (inp[2]) ? node234 : 12'b000000011111;
								assign node234 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
						assign node237 = (inp[10]) ? node241 : node238;
							assign node238 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
							assign node241 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
					assign node244 = (inp[9]) ? node252 : node245;
						assign node245 = (inp[5]) ? node249 : node246;
							assign node246 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
							assign node249 = (inp[8]) ? 12'b000000000111 : 12'b000000001111;
						assign node252 = (inp[10]) ? node256 : node253;
							assign node253 = (inp[2]) ? 12'b000000000011 : 12'b000000001111;
							assign node256 = (inp[6]) ? node258 : 12'b000000000111;
								assign node258 = (inp[2]) ? 12'b000000000011 : 12'b000000000011;

endmodule