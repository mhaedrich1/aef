module dtc_split875_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node13;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node69;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node78;
	wire [1-1:0] node80;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node100;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node122;
	wire [1-1:0] node125;
	wire [1-1:0] node127;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node153;
	wire [1-1:0] node155;
	wire [1-1:0] node158;
	wire [1-1:0] node159;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node171;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node179;
	wire [1-1:0] node182;
	wire [1-1:0] node184;
	wire [1-1:0] node187;
	wire [1-1:0] node189;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node198;
	wire [1-1:0] node201;
	wire [1-1:0] node203;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node211;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node220;
	wire [1-1:0] node222;
	wire [1-1:0] node225;
	wire [1-1:0] node227;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node233;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node245;
	wire [1-1:0] node247;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node258;
	wire [1-1:0] node261;
	wire [1-1:0] node262;
	wire [1-1:0] node264;
	wire [1-1:0] node267;
	wire [1-1:0] node269;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node277;
	wire [1-1:0] node278;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node285;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node294;
	wire [1-1:0] node295;
	wire [1-1:0] node296;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node302;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node311;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node316;
	wire [1-1:0] node317;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node326;
	wire [1-1:0] node328;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node360;
	wire [1-1:0] node363;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node374;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node381;
	wire [1-1:0] node383;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node394;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node406;
	wire [1-1:0] node408;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node421;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node430;
	wire [1-1:0] node432;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node440;
	wire [1-1:0] node443;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node454;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node462;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node468;
	wire [1-1:0] node470;
	wire [1-1:0] node473;
	wire [1-1:0] node474;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node480;
	wire [1-1:0] node483;
	wire [1-1:0] node484;
	wire [1-1:0] node488;
	wire [1-1:0] node489;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node501;
	wire [1-1:0] node504;
	wire [1-1:0] node505;
	wire [1-1:0] node507;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node516;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node519;
	wire [1-1:0] node521;
	wire [1-1:0] node524;
	wire [1-1:0] node525;
	wire [1-1:0] node527;
	wire [1-1:0] node530;
	wire [1-1:0] node531;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node538;
	wire [1-1:0] node539;
	wire [1-1:0] node540;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node550;
	wire [1-1:0] node551;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node556;
	wire [1-1:0] node559;
	wire [1-1:0] node560;
	wire [1-1:0] node562;
	wire [1-1:0] node565;
	wire [1-1:0] node569;
	wire [1-1:0] node570;
	wire [1-1:0] node571;
	wire [1-1:0] node572;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node579;
	wire [1-1:0] node582;
	wire [1-1:0] node584;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node593;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node601;
	wire [1-1:0] node602;
	wire [1-1:0] node604;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node618;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node631;
	wire [1-1:0] node632;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node638;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node646;
	wire [1-1:0] node648;
	wire [1-1:0] node652;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node657;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node661;
	wire [1-1:0] node664;
	wire [1-1:0] node666;
	wire [1-1:0] node669;
	wire [1-1:0] node671;
	wire [1-1:0] node675;
	wire [1-1:0] node676;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node684;
	wire [1-1:0] node686;
	wire [1-1:0] node689;
	wire [1-1:0] node691;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node698;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node704;
	wire [1-1:0] node707;
	wire [1-1:0] node708;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node721;
	wire [1-1:0] node722;
	wire [1-1:0] node723;
	wire [1-1:0] node727;
	wire [1-1:0] node729;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node735;
	wire [1-1:0] node736;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node742;
	wire [1-1:0] node745;
	wire [1-1:0] node746;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node756;
	wire [1-1:0] node757;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node761;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node769;
	wire [1-1:0] node770;
	wire [1-1:0] node774;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node782;
	wire [1-1:0] node783;
	wire [1-1:0] node785;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node793;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node797;
	wire [1-1:0] node799;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node805;
	wire [1-1:0] node808;
	wire [1-1:0] node810;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node818;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node825;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node831;
	wire [1-1:0] node832;
	wire [1-1:0] node837;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node860;
	wire [1-1:0] node863;
	wire [1-1:0] node864;
	wire [1-1:0] node865;
	wire [1-1:0] node869;
	wire [1-1:0] node870;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node880;
	wire [1-1:0] node883;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node895;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node898;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node904;
	wire [1-1:0] node905;
	wire [1-1:0] node906;
	wire [1-1:0] node907;
	wire [1-1:0] node908;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node917;
	wire [1-1:0] node919;
	wire [1-1:0] node923;
	wire [1-1:0] node924;
	wire [1-1:0] node925;
	wire [1-1:0] node926;
	wire [1-1:0] node928;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node933;
	wire [1-1:0] node937;
	wire [1-1:0] node939;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node945;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node955;
	wire [1-1:0] node957;
	wire [1-1:0] node960;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node966;
	wire [1-1:0] node969;
	wire [1-1:0] node970;
	wire [1-1:0] node972;
	wire [1-1:0] node975;
	wire [1-1:0] node977;
	wire [1-1:0] node981;
	wire [1-1:0] node982;
	wire [1-1:0] node983;
	wire [1-1:0] node984;
	wire [1-1:0] node985;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node994;
	wire [1-1:0] node996;
	wire [1-1:0] node999;
	wire [1-1:0] node1001;
	wire [1-1:0] node1005;
	wire [1-1:0] node1006;
	wire [1-1:0] node1007;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1013;
	wire [1-1:0] node1014;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1023;
	wire [1-1:0] node1025;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1031;
	wire [1-1:0] node1032;
	wire [1-1:0] node1033;
	wire [1-1:0] node1037;
	wire [1-1:0] node1039;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1045;
	wire [1-1:0] node1046;
	wire [1-1:0] node1047;
	wire [1-1:0] node1049;
	wire [1-1:0] node1052;
	wire [1-1:0] node1054;
	wire [1-1:0] node1057;
	wire [1-1:0] node1058;
	wire [1-1:0] node1063;
	wire [1-1:0] node1064;
	wire [1-1:0] node1065;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1075;
	wire [1-1:0] node1077;
	wire [1-1:0] node1080;
	wire [1-1:0] node1082;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1088;
	wire [1-1:0] node1090;
	wire [1-1:0] node1091;
	wire [1-1:0] node1093;
	wire [1-1:0] node1096;
	wire [1-1:0] node1098;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1106;
	wire [1-1:0] node1109;
	wire [1-1:0] node1110;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1119;
	wire [1-1:0] node1120;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1129;
	wire [1-1:0] node1131;
	wire [1-1:0] node1134;
	wire [1-1:0] node1136;
	wire [1-1:0] node1140;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1143;
	wire [1-1:0] node1144;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1151;
	wire [1-1:0] node1154;
	wire [1-1:0] node1155;
	wire [1-1:0] node1159;
	wire [1-1:0] node1161;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1167;
	wire [1-1:0] node1168;
	wire [1-1:0] node1172;
	wire [1-1:0] node1173;
	wire [1-1:0] node1175;
	wire [1-1:0] node1178;
	wire [1-1:0] node1180;
	wire [1-1:0] node1182;
	wire [1-1:0] node1185;
	wire [1-1:0] node1187;
	wire [1-1:0] node1189;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1196;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1200;
	wire [1-1:0] node1202;
	wire [1-1:0] node1205;
	wire [1-1:0] node1206;
	wire [1-1:0] node1208;
	wire [1-1:0] node1211;
	wire [1-1:0] node1213;
	wire [1-1:0] node1217;
	wire [1-1:0] node1218;
	wire [1-1:0] node1219;
	wire [1-1:0] node1221;
	wire [1-1:0] node1222;
	wire [1-1:0] node1223;
	wire [1-1:0] node1225;
	wire [1-1:0] node1228;
	wire [1-1:0] node1229;
	wire [1-1:0] node1231;
	wire [1-1:0] node1234;
	wire [1-1:0] node1235;
	wire [1-1:0] node1240;
	wire [1-1:0] node1241;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1245;
	wire [1-1:0] node1248;
	wire [1-1:0] node1249;
	wire [1-1:0] node1251;
	wire [1-1:0] node1254;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1265;
	wire [1-1:0] node1266;
	wire [1-1:0] node1270;
	wire [1-1:0] node1272;
	wire [1-1:0] node1275;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1287;
	wire [1-1:0] node1290;
	wire [1-1:0] node1291;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1300;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1304;
	wire [1-1:0] node1307;
	wire [1-1:0] node1309;
	wire [1-1:0] node1312;
	wire [1-1:0] node1313;
	wire [1-1:0] node1318;
	wire [1-1:0] node1319;
	wire [1-1:0] node1320;
	wire [1-1:0] node1321;
	wire [1-1:0] node1322;
	wire [1-1:0] node1323;
	wire [1-1:0] node1325;
	wire [1-1:0] node1328;
	wire [1-1:0] node1329;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1347;
	wire [1-1:0] node1351;
	wire [1-1:0] node1352;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1359;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1371;
	wire [1-1:0] node1373;
	wire [1-1:0] node1377;
	wire [1-1:0] node1378;
	wire [1-1:0] node1379;
	wire [1-1:0] node1380;
	wire [1-1:0] node1381;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1385;
	wire [1-1:0] node1386;
	wire [1-1:0] node1390;
	wire [1-1:0] node1392;
	wire [1-1:0] node1395;
	wire [1-1:0] node1397;
	wire [1-1:0] node1401;
	wire [1-1:0] node1402;
	wire [1-1:0] node1403;
	wire [1-1:0] node1405;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1410;
	wire [1-1:0] node1414;
	wire [1-1:0] node1416;
	wire [1-1:0] node1419;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1424;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1433;
	wire [1-1:0] node1435;
	wire [1-1:0] node1438;
	wire [1-1:0] node1440;
	wire [1-1:0] node1441;
	wire [1-1:0] node1442;
	wire [1-1:0] node1443;
	wire [1-1:0] node1445;
	wire [1-1:0] node1448;
	wire [1-1:0] node1449;
	wire [1-1:0] node1453;
	wire [1-1:0] node1455;
	wire [1-1:0] node1459;
	wire [1-1:0] node1460;
	wire [1-1:0] node1461;
	wire [1-1:0] node1462;
	wire [1-1:0] node1463;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1468;
	wire [1-1:0] node1471;
	wire [1-1:0] node1472;
	wire [1-1:0] node1474;
	wire [1-1:0] node1477;
	wire [1-1:0] node1479;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1486;
	wire [1-1:0] node1490;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1501;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1505;
	wire [1-1:0] node1507;
	wire [1-1:0] node1510;
	wire [1-1:0] node1511;
	wire [1-1:0] node1515;
	wire [1-1:0] node1516;
	wire [1-1:0] node1520;
	wire [1-1:0] node1521;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1525;
	wire [1-1:0] node1527;
	wire [1-1:0] node1530;
	wire [1-1:0] node1532;
	wire [1-1:0] node1535;
	wire [1-1:0] node1537;
	wire [1-1:0] node1541;
	wire [1-1:0] node1542;
	wire [1-1:0] node1543;
	wire [1-1:0] node1544;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1550;
	wire [1-1:0] node1553;
	wire [1-1:0] node1554;
	wire [1-1:0] node1558;
	wire [1-1:0] node1559;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1568;
	wire [1-1:0] node1570;
	wire [1-1:0] node1573;
	wire [1-1:0] node1574;
	wire [1-1:0] node1578;
	wire [1-1:0] node1580;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1586;
	wire [1-1:0] node1587;
	wire [1-1:0] node1591;
	wire [1-1:0] node1592;
	wire [1-1:0] node1596;
	wire [1-1:0] node1598;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1604;
	wire [1-1:0] node1605;
	wire [1-1:0] node1606;
	wire [1-1:0] node1607;
	wire [1-1:0] node1611;
	wire [1-1:0] node1613;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1622;
	wire [1-1:0] node1623;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1627;
	wire [1-1:0] node1629;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1634;
	wire [1-1:0] node1638;
	wire [1-1:0] node1639;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1652;
	wire [1-1:0] node1653;
	wire [1-1:0] node1655;
	wire [1-1:0] node1658;
	wire [1-1:0] node1659;
	wire [1-1:0] node1663;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1667;
	wire [1-1:0] node1669;
	wire [1-1:0] node1672;
	wire [1-1:0] node1674;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1682;
	wire [1-1:0] node1684;
	wire [1-1:0] node1685;
	wire [1-1:0] node1686;
	wire [1-1:0] node1687;
	wire [1-1:0] node1689;
	wire [1-1:0] node1692;
	wire [1-1:0] node1693;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1706;
	wire [1-1:0] node1707;
	wire [1-1:0] node1708;
	wire [1-1:0] node1709;
	wire [1-1:0] node1711;
	wire [1-1:0] node1712;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1719;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1731;
	wire [1-1:0] node1732;
	wire [1-1:0] node1733;
	wire [1-1:0] node1734;
	wire [1-1:0] node1735;
	wire [1-1:0] node1739;
	wire [1-1:0] node1741;
	wire [1-1:0] node1744;
	wire [1-1:0] node1746;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1754;
	wire [1-1:0] node1757;
	wire [1-1:0] node1759;
	wire [1-1:0] node1762;
	wire [1-1:0] node1763;
	wire [1-1:0] node1767;
	wire [1-1:0] node1769;
	wire [1-1:0] node1770;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1776;
	wire [1-1:0] node1777;
	wire [1-1:0] node1779;
	wire [1-1:0] node1782;
	wire [1-1:0] node1783;
	wire [1-1:0] node1788;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1791;
	wire [1-1:0] node1793;
	wire [1-1:0] node1794;
	wire [1-1:0] node1795;
	wire [1-1:0] node1796;
	wire [1-1:0] node1800;
	wire [1-1:0] node1802;
	wire [1-1:0] node1805;
	wire [1-1:0] node1807;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1813;
	wire [1-1:0] node1814;
	wire [1-1:0] node1815;
	wire [1-1:0] node1817;
	wire [1-1:0] node1820;
	wire [1-1:0] node1822;
	wire [1-1:0] node1825;
	wire [1-1:0] node1826;
	wire [1-1:0] node1831;
	wire [1-1:0] node1832;
	wire [1-1:0] node1834;
	wire [1-1:0] node1837;
	wire [1-1:0] node1838;
	wire [1-1:0] node1840;
	wire [1-1:0] node1843;
	wire [1-1:0] node1845;
	wire [1-1:0] node1848;
	wire [1-1:0] node1850;
	wire [1-1:0] node1851;
	wire [1-1:0] node1852;
	wire [1-1:0] node1853;
	wire [1-1:0] node1855;
	wire [1-1:0] node1858;
	wire [1-1:0] node1860;
	wire [1-1:0] node1863;
	wire [1-1:0] node1865;
	wire [1-1:0] node1869;
	wire [1-1:0] node1870;
	wire [1-1:0] node1871;
	wire [1-1:0] node1873;
	wire [1-1:0] node1874;
	wire [1-1:0] node1875;
	wire [1-1:0] node1879;
	wire [1-1:0] node1880;
	wire [1-1:0] node1882;
	wire [1-1:0] node1885;
	wire [1-1:0] node1886;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1893;
	wire [1-1:0] node1894;
	wire [1-1:0] node1895;
	wire [1-1:0] node1897;
	wire [1-1:0] node1900;
	wire [1-1:0] node1901;
	wire [1-1:0] node1902;
	wire [1-1:0] node1906;
	wire [1-1:0] node1907;
	wire [1-1:0] node1912;
	wire [1-1:0] node1913;
	wire [1-1:0] node1915;
	wire [1-1:0] node1918;
	wire [1-1:0] node1919;
	wire [1-1:0] node1920;
	wire [1-1:0] node1924;
	wire [1-1:0] node1925;
	wire [1-1:0] node1929;
	wire [1-1:0] node1930;
	wire [1-1:0] node1932;
	wire [1-1:0] node1933;
	wire [1-1:0] node1934;
	wire [1-1:0] node1935;
	wire [1-1:0] node1939;
	wire [1-1:0] node1941;
	wire [1-1:0] node1944;
	wire [1-1:0] node1946;
	wire [1-1:0] node1950;
	wire [1-1:0] node1951;
	wire [1-1:0] node1952;
	wire [1-1:0] node1953;
	wire [1-1:0] node1955;
	wire [1-1:0] node1956;
	wire [1-1:0] node1957;
	wire [1-1:0] node1958;
	wire [1-1:0] node1962;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1968;
	wire [1-1:0] node1969;
	wire [1-1:0] node1974;
	wire [1-1:0] node1975;
	wire [1-1:0] node1976;
	wire [1-1:0] node1977;
	wire [1-1:0] node1978;
	wire [1-1:0] node1982;
	wire [1-1:0] node1984;
	wire [1-1:0] node1987;
	wire [1-1:0] node1989;
	wire [1-1:0] node1992;
	wire [1-1:0] node1994;
	wire [1-1:0] node1995;
	wire [1-1:0] node1996;
	wire [1-1:0] node1998;
	wire [1-1:0] node2001;
	wire [1-1:0] node2002;
	wire [1-1:0] node2006;
	wire [1-1:0] node2008;
	wire [1-1:0] node2011;
	wire [1-1:0] node2013;
	wire [1-1:0] node2014;
	wire [1-1:0] node2015;
	wire [1-1:0] node2016;
	wire [1-1:0] node2020;
	wire [1-1:0] node2021;
	wire [1-1:0] node2022;
	wire [1-1:0] node2026;
	wire [1-1:0] node2028;
	wire [1-1:0] node2032;
	wire [1-1:0] node2033;
	wire [1-1:0] node2034;
	wire [1-1:0] node2035;
	wire [1-1:0] node2037;
	wire [1-1:0] node2038;
	wire [1-1:0] node2039;
	wire [1-1:0] node2040;
	wire [1-1:0] node2042;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2050;
	wire [1-1:0] node2051;
	wire [1-1:0] node2056;
	wire [1-1:0] node2057;
	wire [1-1:0] node2058;
	wire [1-1:0] node2059;
	wire [1-1:0] node2060;
	wire [1-1:0] node2064;
	wire [1-1:0] node2066;
	wire [1-1:0] node2069;
	wire [1-1:0] node2071;
	wire [1-1:0] node2074;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2079;
	wire [1-1:0] node2082;
	wire [1-1:0] node2083;
	wire [1-1:0] node2085;
	wire [1-1:0] node2088;
	wire [1-1:0] node2089;
	wire [1-1:0] node2093;
	wire [1-1:0] node2094;
	wire [1-1:0] node2096;
	wire [1-1:0] node2097;
	wire [1-1:0] node2098;
	wire [1-1:0] node2100;
	wire [1-1:0] node2103;
	wire [1-1:0] node2105;
	wire [1-1:0] node2108;
	wire [1-1:0] node2109;
	wire [1-1:0] node2114;
	wire [1-1:0] node2115;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2119;
	wire [1-1:0] node2120;
	wire [1-1:0] node2122;
	wire [1-1:0] node2125;
	wire [1-1:0] node2127;
	wire [1-1:0] node2130;
	wire [1-1:0] node2131;
	wire [1-1:0] node2136;
	wire [1-1:0] node2137;
	wire [1-1:0] node2138;
	wire [1-1:0] node2139;
	wire [1-1:0] node2140;
	wire [1-1:0] node2142;
	wire [1-1:0] node2145;
	wire [1-1:0] node2146;
	wire [1-1:0] node2148;
	wire [1-1:0] node2151;
	wire [1-1:0] node2153;
	wire [1-1:0] node2157;
	wire [1-1:0] node2158;
	wire [1-1:0] node2159;
	wire [1-1:0] node2161;
	wire [1-1:0] node2164;
	wire [1-1:0] node2165;
	wire [1-1:0] node2169;
	wire [1-1:0] node2171;
	wire [1-1:0] node2174;
	wire [1-1:0] node2176;
	wire [1-1:0] node2177;
	wire [1-1:0] node2178;
	wire [1-1:0] node2179;
	wire [1-1:0] node2180;
	wire [1-1:0] node2184;
	wire [1-1:0] node2185;
	wire [1-1:0] node2189;
	wire [1-1:0] node2191;
	wire [1-1:0] node2195;
	wire [1-1:0] node2196;
	wire [1-1:0] node2197;
	wire [1-1:0] node2199;
	wire [1-1:0] node2200;
	wire [1-1:0] node2201;
	wire [1-1:0] node2202;
	wire [1-1:0] node2203;
	wire [1-1:0] node2207;
	wire [1-1:0] node2209;
	wire [1-1:0] node2212;
	wire [1-1:0] node2214;
	wire [1-1:0] node2218;
	wire [1-1:0] node2219;
	wire [1-1:0] node2220;
	wire [1-1:0] node2221;
	wire [1-1:0] node2222;
	wire [1-1:0] node2223;
	wire [1-1:0] node2227;
	wire [1-1:0] node2229;
	wire [1-1:0] node2232;
	wire [1-1:0] node2234;
	wire [1-1:0] node2237;
	wire [1-1:0] node2239;
	wire [1-1:0] node2240;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2246;
	wire [1-1:0] node2247;
	wire [1-1:0] node2251;
	wire [1-1:0] node2253;
	wire [1-1:0] node2256;
	wire [1-1:0] node2258;
	wire [1-1:0] node2259;
	wire [1-1:0] node2260;
	wire [1-1:0] node2261;
	wire [1-1:0] node2265;
	wire [1-1:0] node2266;
	wire [1-1:0] node2268;
	wire [1-1:0] node2271;
	wire [1-1:0] node2272;
	wire [1-1:0] node2277;
	wire [1-1:0] node2278;
	wire [1-1:0] node2279;
	wire [1-1:0] node2280;
	wire [1-1:0] node2282;
	wire [1-1:0] node2283;
	wire [1-1:0] node2284;
	wire [1-1:0] node2285;
	wire [1-1:0] node2289;
	wire [1-1:0] node2290;
	wire [1-1:0] node2294;
	wire [1-1:0] node2296;
	wire [1-1:0] node2300;
	wire [1-1:0] node2301;
	wire [1-1:0] node2302;
	wire [1-1:0] node2303;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2309;
	wire [1-1:0] node2310;
	wire [1-1:0] node2312;
	wire [1-1:0] node2315;
	wire [1-1:0] node2317;
	wire [1-1:0] node2321;
	wire [1-1:0] node2322;
	wire [1-1:0] node2323;
	wire [1-1:0] node2327;
	wire [1-1:0] node2328;
	wire [1-1:0] node2329;
	wire [1-1:0] node2333;
	wire [1-1:0] node2334;
	wire [1-1:0] node2338;
	wire [1-1:0] node2340;
	wire [1-1:0] node2341;
	wire [1-1:0] node2342;
	wire [1-1:0] node2343;
	wire [1-1:0] node2347;
	wire [1-1:0] node2348;
	wire [1-1:0] node2349;
	wire [1-1:0] node2353;
	wire [1-1:0] node2355;
	wire [1-1:0] node2359;
	wire [1-1:0] node2360;
	wire [1-1:0] node2361;
	wire [1-1:0] node2363;
	wire [1-1:0] node2364;
	wire [1-1:0] node2365;
	wire [1-1:0] node2366;
	wire [1-1:0] node2370;
	wire [1-1:0] node2371;
	wire [1-1:0] node2373;
	wire [1-1:0] node2376;
	wire [1-1:0] node2377;
	wire [1-1:0] node2382;
	wire [1-1:0] node2383;
	wire [1-1:0] node2384;
	wire [1-1:0] node2385;
	wire [1-1:0] node2387;
	wire [1-1:0] node2390;
	wire [1-1:0] node2391;
	wire [1-1:0] node2393;
	wire [1-1:0] node2396;
	wire [1-1:0] node2398;
	wire [1-1:0] node2402;
	wire [1-1:0] node2403;
	wire [1-1:0] node2404;
	wire [1-1:0] node2408;
	wire [1-1:0] node2409;
	wire [1-1:0] node2411;
	wire [1-1:0] node2414;
	wire [1-1:0] node2416;
	wire [1-1:0] node2419;
	wire [1-1:0] node2421;
	wire [1-1:0] node2422;
	wire [1-1:0] node2423;
	wire [1-1:0] node2424;
	wire [1-1:0] node2428;
	wire [1-1:0] node2429;
	wire [1-1:0] node2430;
	wire [1-1:0] node2434;
	wire [1-1:0] node2436;
	wire [1-1:0] node2440;
	wire [1-1:0] node2441;
	wire [1-1:0] node2442;
	wire [1-1:0] node2443;
	wire [1-1:0] node2444;
	wire [1-1:0] node2446;
	wire [1-1:0] node2447;
	wire [1-1:0] node2448;
	wire [1-1:0] node2450;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2456;
	wire [1-1:0] node2459;
	wire [1-1:0] node2460;
	wire [1-1:0] node2465;
	wire [1-1:0] node2466;
	wire [1-1:0] node2467;
	wire [1-1:0] node2468;
	wire [1-1:0] node2470;
	wire [1-1:0] node2473;
	wire [1-1:0] node2475;
	wire [1-1:0] node2478;
	wire [1-1:0] node2480;
	wire [1-1:0] node2483;
	wire [1-1:0] node2485;
	wire [1-1:0] node2486;
	wire [1-1:0] node2488;
	wire [1-1:0] node2491;
	wire [1-1:0] node2492;
	wire [1-1:0] node2494;
	wire [1-1:0] node2497;
	wire [1-1:0] node2498;
	wire [1-1:0] node2502;
	wire [1-1:0] node2503;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;
	wire [1-1:0] node2508;
	wire [1-1:0] node2511;
	wire [1-1:0] node2512;
	wire [1-1:0] node2514;
	wire [1-1:0] node2517;
	wire [1-1:0] node2518;
	wire [1-1:0] node2523;
	wire [1-1:0] node2524;
	wire [1-1:0] node2525;
	wire [1-1:0] node2526;
	wire [1-1:0] node2527;
	wire [1-1:0] node2529;
	wire [1-1:0] node2530;
	wire [1-1:0] node2531;
	wire [1-1:0] node2532;
	wire [1-1:0] node2536;
	wire [1-1:0] node2537;
	wire [1-1:0] node2539;
	wire [1-1:0] node2542;
	wire [1-1:0] node2543;
	wire [1-1:0] node2548;
	wire [1-1:0] node2549;
	wire [1-1:0] node2550;
	wire [1-1:0] node2551;
	wire [1-1:0] node2552;
	wire [1-1:0] node2553;
	wire [1-1:0] node2557;
	wire [1-1:0] node2558;
	wire [1-1:0] node2560;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2569;
	wire [1-1:0] node2570;
	wire [1-1:0] node2572;
	wire [1-1:0] node2575;
	wire [1-1:0] node2576;
	wire [1-1:0] node2578;
	wire [1-1:0] node2581;
	wire [1-1:0] node2582;
	wire [1-1:0] node2586;
	wire [1-1:0] node2587;
	wire [1-1:0] node2589;
	wire [1-1:0] node2590;
	wire [1-1:0] node2591;
	wire [1-1:0] node2592;
	wire [1-1:0] node2596;
	wire [1-1:0] node2597;
	wire [1-1:0] node2601;
	wire [1-1:0] node2602;
	wire [1-1:0] node2607;
	wire [1-1:0] node2608;
	wire [1-1:0] node2609;
	wire [1-1:0] node2611;
	wire [1-1:0] node2612;
	wire [1-1:0] node2613;
	wire [1-1:0] node2614;
	wire [1-1:0] node2616;
	wire [1-1:0] node2619;
	wire [1-1:0] node2620;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2630;
	wire [1-1:0] node2631;
	wire [1-1:0] node2632;
	wire [1-1:0] node2633;
	wire [1-1:0] node2634;
	wire [1-1:0] node2636;
	wire [1-1:0] node2639;
	wire [1-1:0] node2640;
	wire [1-1:0] node2644;
	wire [1-1:0] node2646;
	wire [1-1:0] node2650;
	wire [1-1:0] node2651;
	wire [1-1:0] node2652;
	wire [1-1:0] node2656;
	wire [1-1:0] node2657;
	wire [1-1:0] node2659;
	wire [1-1:0] node2662;
	wire [1-1:0] node2663;
	wire [1-1:0] node2667;
	wire [1-1:0] node2669;
	wire [1-1:0] node2670;
	wire [1-1:0] node2671;
	wire [1-1:0] node2672;
	wire [1-1:0] node2676;
	wire [1-1:0] node2677;
	wire [1-1:0] node2679;
	wire [1-1:0] node2682;
	wire [1-1:0] node2683;
	wire [1-1:0] node2688;
	wire [1-1:0] node2689;
	wire [1-1:0] node2690;
	wire [1-1:0] node2691;
	wire [1-1:0] node2693;
	wire [1-1:0] node2694;
	wire [1-1:0] node2695;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2701;
	wire [1-1:0] node2705;
	wire [1-1:0] node2706;
	wire [1-1:0] node2711;
	wire [1-1:0] node2712;
	wire [1-1:0] node2713;
	wire [1-1:0] node2715;
	wire [1-1:0] node2718;
	wire [1-1:0] node2719;
	wire [1-1:0] node2721;
	wire [1-1:0] node2724;
	wire [1-1:0] node2726;
	wire [1-1:0] node2729;
	wire [1-1:0] node2731;
	wire [1-1:0] node2732;
	wire [1-1:0] node2733;
	wire [1-1:0] node2737;
	wire [1-1:0] node2738;
	wire [1-1:0] node2740;
	wire [1-1:0] node2743;
	wire [1-1:0] node2745;
	wire [1-1:0] node2748;
	wire [1-1:0] node2750;
	wire [1-1:0] node2751;
	wire [1-1:0] node2752;
	wire [1-1:0] node2753;
	wire [1-1:0] node2757;
	wire [1-1:0] node2758;
	wire [1-1:0] node2760;
	wire [1-1:0] node2763;
	wire [1-1:0] node2765;
	wire [1-1:0] node2769;
	wire [1-1:0] node2770;
	wire [1-1:0] node2771;
	wire [1-1:0] node2772;
	wire [1-1:0] node2773;
	wire [1-1:0] node2774;
	wire [1-1:0] node2775;
	wire [1-1:0] node2777;
	wire [1-1:0] node2778;
	wire [1-1:0] node2780;
	wire [1-1:0] node2783;
	wire [1-1:0] node2784;
	wire [1-1:0] node2785;
	wire [1-1:0] node2789;
	wire [1-1:0] node2791;
	wire [1-1:0] node2795;
	wire [1-1:0] node2796;
	wire [1-1:0] node2797;
	wire [1-1:0] node2799;
	wire [1-1:0] node2802;
	wire [1-1:0] node2803;
	wire [1-1:0] node2805;
	wire [1-1:0] node2808;
	wire [1-1:0] node2810;
	wire [1-1:0] node2813;
	wire [1-1:0] node2815;
	wire [1-1:0] node2816;
	wire [1-1:0] node2817;
	wire [1-1:0] node2821;
	wire [1-1:0] node2822;
	wire [1-1:0] node2824;
	wire [1-1:0] node2827;
	wire [1-1:0] node2829;
	wire [1-1:0] node2832;
	wire [1-1:0] node2834;
	wire [1-1:0] node2835;
	wire [1-1:0] node2836;
	wire [1-1:0] node2838;
	wire [1-1:0] node2841;
	wire [1-1:0] node2842;
	wire [1-1:0] node2843;
	wire [1-1:0] node2847;
	wire [1-1:0] node2849;
	wire [1-1:0] node2853;
	wire [1-1:0] node2854;
	wire [1-1:0] node2855;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2859;
	wire [1-1:0] node2860;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2866;
	wire [1-1:0] node2870;
	wire [1-1:0] node2872;
	wire [1-1:0] node2876;
	wire [1-1:0] node2877;
	wire [1-1:0] node2878;
	wire [1-1:0] node2879;
	wire [1-1:0] node2880;
	wire [1-1:0] node2884;
	wire [1-1:0] node2885;
	wire [1-1:0] node2889;
	wire [1-1:0] node2890;
	wire [1-1:0] node2894;
	wire [1-1:0] node2896;
	wire [1-1:0] node2897;
	wire [1-1:0] node2899;
	wire [1-1:0] node2902;
	wire [1-1:0] node2903;
	wire [1-1:0] node2904;
	wire [1-1:0] node2908;
	wire [1-1:0] node2909;
	wire [1-1:0] node2913;
	wire [1-1:0] node2914;
	wire [1-1:0] node2916;
	wire [1-1:0] node2917;
	wire [1-1:0] node2918;
	wire [1-1:0] node2919;
	wire [1-1:0] node2923;
	wire [1-1:0] node2925;
	wire [1-1:0] node2928;
	wire [1-1:0] node2930;
	wire [1-1:0] node2934;
	wire [1-1:0] node2935;
	wire [1-1:0] node2937;
	wire [1-1:0] node2938;
	wire [1-1:0] node2939;
	wire [1-1:0] node2940;
	wire [1-1:0] node2941;
	wire [1-1:0] node2945;
	wire [1-1:0] node2947;
	wire [1-1:0] node2950;
	wire [1-1:0] node2952;
	wire [1-1:0] node2956;
	wire [1-1:0] node2957;
	wire [1-1:0] node2958;
	wire [1-1:0] node2959;
	wire [1-1:0] node2960;
	wire [1-1:0] node2961;
	wire [1-1:0] node2962;
	wire [1-1:0] node2966;
	wire [1-1:0] node2968;
	wire [1-1:0] node2971;
	wire [1-1:0] node2972;
	wire [1-1:0] node2977;
	wire [1-1:0] node2978;
	wire [1-1:0] node2979;
	wire [1-1:0] node2981;
	wire [1-1:0] node2984;
	wire [1-1:0] node2986;
	wire [1-1:0] node2989;
	wire [1-1:0] node2991;
	wire [1-1:0] node2994;
	wire [1-1:0] node2995;
	wire [1-1:0] node2997;
	wire [1-1:0] node2998;
	wire [1-1:0] node3000;
	wire [1-1:0] node3003;
	wire [1-1:0] node3004;
	wire [1-1:0] node3005;
	wire [1-1:0] node3009;
	wire [1-1:0] node3010;
	wire [1-1:0] node3015;
	wire [1-1:0] node3016;
	wire [1-1:0] node3017;
	wire [1-1:0] node3018;
	wire [1-1:0] node3020;
	wire [1-1:0] node3021;
	wire [1-1:0] node3022;
	wire [1-1:0] node3023;
	wire [1-1:0] node3027;
	wire [1-1:0] node3028;
	wire [1-1:0] node3029;
	wire [1-1:0] node3033;
	wire [1-1:0] node3034;
	wire [1-1:0] node3039;
	wire [1-1:0] node3040;
	wire [1-1:0] node3041;
	wire [1-1:0] node3042;
	wire [1-1:0] node3044;
	wire [1-1:0] node3047;
	wire [1-1:0] node3048;
	wire [1-1:0] node3049;
	wire [1-1:0] node3053;
	wire [1-1:0] node3054;
	wire [1-1:0] node3058;
	wire [1-1:0] node3060;
	wire [1-1:0] node3061;
	wire [1-1:0] node3062;
	wire [1-1:0] node3063;
	wire [1-1:0] node3067;
	wire [1-1:0] node3069;
	wire [1-1:0] node3072;
	wire [1-1:0] node3073;
	wire [1-1:0] node3077;
	wire [1-1:0] node3078;
	wire [1-1:0] node3080;
	wire [1-1:0] node3081;
	wire [1-1:0] node3082;
	wire [1-1:0] node3084;
	wire [1-1:0] node3087;
	wire [1-1:0] node3089;
	wire [1-1:0] node3092;
	wire [1-1:0] node3094;
	wire [1-1:0] node3098;
	wire [1-1:0] node3099;
	wire [1-1:0] node3100;
	wire [1-1:0] node3102;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3105;
	wire [1-1:0] node3109;
	wire [1-1:0] node3110;
	wire [1-1:0] node3112;
	wire [1-1:0] node3115;
	wire [1-1:0] node3117;
	wire [1-1:0] node3121;
	wire [1-1:0] node3122;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3125;
	wire [1-1:0] node3126;
	wire [1-1:0] node3131;
	wire [1-1:0] node3133;
	wire [1-1:0] node3137;
	wire [1-1:0] node3138;
	wire [1-1:0] node3140;
	wire [1-1:0] node3143;
	wire [1-1:0] node3144;
	wire [1-1:0] node3146;
	wire [1-1:0] node3149;
	wire [1-1:0] node3151;
	wire [1-1:0] node3154;
	wire [1-1:0] node3156;
	wire [1-1:0] node3157;
	wire [1-1:0] node3158;
	wire [1-1:0] node3160;
	wire [1-1:0] node3163;
	wire [1-1:0] node3164;
	wire [1-1:0] node3165;
	wire [1-1:0] node3169;
	wire [1-1:0] node3171;
	wire [1-1:0] node3175;
	wire [1-1:0] node3176;
	wire [1-1:0] node3177;
	wire [1-1:0] node3179;
	wire [1-1:0] node3180;
	wire [1-1:0] node3181;
	wire [1-1:0] node3182;
	wire [1-1:0] node3183;
	wire [1-1:0] node3187;
	wire [1-1:0] node3189;
	wire [1-1:0] node3192;
	wire [1-1:0] node3194;
	wire [1-1:0] node3198;
	wire [1-1:0] node3199;
	wire [1-1:0] node3200;
	wire [1-1:0] node3202;
	wire [1-1:0] node3205;
	wire [1-1:0] node3206;
	wire [1-1:0] node3208;
	wire [1-1:0] node3211;
	wire [1-1:0] node3212;
	wire [1-1:0] node3216;
	wire [1-1:0] node3218;
	wire [1-1:0] node3219;
	wire [1-1:0] node3220;
	wire [1-1:0] node3222;
	wire [1-1:0] node3225;
	wire [1-1:0] node3226;
	wire [1-1:0] node3230;
	wire [1-1:0] node3232;
	wire [1-1:0] node3235;
	wire [1-1:0] node3237;
	wire [1-1:0] node3238;
	wire [1-1:0] node3239;
	wire [1-1:0] node3240;
	wire [1-1:0] node3241;
	wire [1-1:0] node3245;
	wire [1-1:0] node3246;
	wire [1-1:0] node3250;
	wire [1-1:0] node3252;
	wire [1-1:0] node3256;
	wire [1-1:0] node3257;
	wire [1-1:0] node3258;
	wire [1-1:0] node3260;
	wire [1-1:0] node3261;
	wire [1-1:0] node3262;
	wire [1-1:0] node3264;
	wire [1-1:0] node3267;
	wire [1-1:0] node3268;
	wire [1-1:0] node3270;
	wire [1-1:0] node3273;
	wire [1-1:0] node3274;
	wire [1-1:0] node3279;
	wire [1-1:0] node3280;
	wire [1-1:0] node3281;
	wire [1-1:0] node3283;
	wire [1-1:0] node3286;
	wire [1-1:0] node3287;
	wire [1-1:0] node3288;
	wire [1-1:0] node3292;
	wire [1-1:0] node3294;
	wire [1-1:0] node3297;
	wire [1-1:0] node3299;
	wire [1-1:0] node3300;
	wire [1-1:0] node3301;
	wire [1-1:0] node3305;
	wire [1-1:0] node3306;
	wire [1-1:0] node3308;
	wire [1-1:0] node3311;
	wire [1-1:0] node3312;
	wire [1-1:0] node3316;
	wire [1-1:0] node3317;
	wire [1-1:0] node3319;
	wire [1-1:0] node3320;
	wire [1-1:0] node3321;
	wire [1-1:0] node3323;
	wire [1-1:0] node3326;
	wire [1-1:0] node3327;
	wire [1-1:0] node3331;
	wire [1-1:0] node3332;

	assign outp = (inp[5]) ? node2440 : node1;
		assign node1 = (inp[6]) ? node895 : node2;
			assign node2 = (inp[12]) ? node84 : node3;
				assign node3 = (inp[1]) ? node25 : node4;
					assign node4 = (inp[0]) ? node6 : 1'b1;
						assign node6 = (inp[4]) ? 1'b1 : node7;
							assign node7 = (inp[13]) ? node13 : node8;
								assign node8 = (inp[2]) ? 1'b0 : node9;
									assign node9 = (inp[14]) ? 1'b1 : 1'b0;
								assign node13 = (inp[11]) ? node19 : node14;
									assign node14 = (inp[2]) ? 1'b1 : node15;
										assign node15 = (inp[14]) ? 1'b0 : 1'b1;
									assign node19 = (inp[14]) ? node21 : 1'b0;
										assign node21 = (inp[2]) ? 1'b0 : 1'b1;
					assign node25 = (inp[8]) ? node63 : node26;
						assign node26 = (inp[4]) ? node46 : node27;
							assign node27 = (inp[0]) ? 1'b1 : node28;
								assign node28 = (inp[14]) ? node34 : node29;
									assign node29 = (inp[11]) ? 1'b0 : node30;
										assign node30 = (inp[13]) ? 1'b1 : 1'b0;
									assign node34 = (inp[2]) ? node40 : node35;
										assign node35 = (inp[11]) ? 1'b1 : node36;
											assign node36 = (inp[13]) ? 1'b0 : 1'b1;
										assign node40 = (inp[11]) ? 1'b0 : node41;
											assign node41 = (inp[13]) ? 1'b1 : 1'b0;
							assign node46 = (inp[11]) ? node58 : node47;
								assign node47 = (inp[13]) ? node53 : node48;
									assign node48 = (inp[2]) ? 1'b0 : node49;
										assign node49 = (inp[14]) ? 1'b1 : 1'b0;
									assign node53 = (inp[2]) ? 1'b1 : node54;
										assign node54 = (inp[14]) ? 1'b0 : 1'b1;
								assign node58 = (inp[2]) ? 1'b0 : node59;
									assign node59 = (inp[14]) ? 1'b1 : 1'b0;
						assign node63 = (inp[0]) ? node65 : 1'b1;
							assign node65 = (inp[4]) ? 1'b1 : node66;
								assign node66 = (inp[14]) ? node72 : node67;
									assign node67 = (inp[13]) ? node69 : 1'b0;
										assign node69 = (inp[11]) ? 1'b0 : 1'b1;
									assign node72 = (inp[2]) ? node78 : node73;
										assign node73 = (inp[11]) ? 1'b1 : node74;
											assign node74 = (inp[13]) ? 1'b0 : 1'b1;
										assign node78 = (inp[13]) ? node80 : 1'b0;
											assign node80 = (inp[11]) ? 1'b0 : 1'b1;
				assign node84 = (inp[15]) ? node814 : node85;
					assign node85 = (inp[10]) ? node569 : node86;
						assign node86 = (inp[9]) ? node332 : node87;
							assign node87 = (inp[3]) ? node169 : node88;
								assign node88 = (inp[1]) ? node110 : node89;
									assign node89 = (inp[0]) ? node91 : 1'b0;
										assign node91 = (inp[4]) ? 1'b0 : node92;
											assign node92 = (inp[2]) ? node104 : node93;
												assign node93 = (inp[14]) ? node99 : node94;
													assign node94 = (inp[13]) ? node96 : 1'b1;
														assign node96 = (inp[11]) ? 1'b1 : 1'b0;
													assign node99 = (inp[11]) ? 1'b0 : node100;
														assign node100 = (inp[13]) ? 1'b1 : 1'b0;
												assign node104 = (inp[11]) ? 1'b1 : node105;
													assign node105 = (inp[13]) ? 1'b0 : 1'b1;
									assign node110 = (inp[8]) ? node148 : node111;
										assign node111 = (inp[4]) ? node131 : node112;
											assign node112 = (inp[0]) ? 1'b0 : node113;
												assign node113 = (inp[14]) ? node119 : node114;
													assign node114 = (inp[13]) ? node116 : 1'b1;
														assign node116 = (inp[11]) ? 1'b1 : 1'b0;
													assign node119 = (inp[2]) ? node125 : node120;
														assign node120 = (inp[13]) ? node122 : 1'b0;
															assign node122 = (inp[11]) ? 1'b0 : 1'b1;
														assign node125 = (inp[13]) ? node127 : 1'b1;
															assign node127 = (inp[11]) ? 1'b1 : 1'b0;
											assign node131 = (inp[14]) ? node137 : node132;
												assign node132 = (inp[11]) ? 1'b1 : node133;
													assign node133 = (inp[13]) ? 1'b0 : 1'b1;
												assign node137 = (inp[2]) ? node143 : node138;
													assign node138 = (inp[11]) ? 1'b0 : node139;
														assign node139 = (inp[13]) ? 1'b1 : 1'b0;
													assign node143 = (inp[11]) ? 1'b1 : node144;
														assign node144 = (inp[13]) ? 1'b0 : 1'b1;
										assign node148 = (inp[4]) ? 1'b0 : node149;
											assign node149 = (inp[0]) ? node151 : 1'b0;
												assign node151 = (inp[11]) ? node163 : node152;
													assign node152 = (inp[13]) ? node158 : node153;
														assign node153 = (inp[14]) ? node155 : 1'b1;
															assign node155 = (inp[2]) ? 1'b1 : 1'b0;
														assign node158 = (inp[2]) ? 1'b0 : node159;
															assign node159 = (inp[14]) ? 1'b1 : 1'b0;
													assign node163 = (inp[14]) ? node165 : 1'b1;
														assign node165 = (inp[2]) ? 1'b1 : 1'b0;
								assign node169 = (inp[7]) ? node251 : node170;
									assign node170 = (inp[8]) ? node230 : node171;
										assign node171 = (inp[1]) ? node193 : node172;
											assign node172 = (inp[0]) ? node174 : 1'b1;
												assign node174 = (inp[4]) ? 1'b1 : node175;
													assign node175 = (inp[2]) ? node187 : node176;
														assign node176 = (inp[14]) ? node182 : node177;
															assign node177 = (inp[13]) ? node179 : 1'b0;
																assign node179 = (inp[11]) ? 1'b0 : 1'b1;
															assign node182 = (inp[13]) ? node184 : 1'b1;
																assign node184 = (inp[11]) ? 1'b1 : 1'b0;
														assign node187 = (inp[13]) ? node189 : 1'b0;
															assign node189 = (inp[11]) ? 1'b0 : 1'b1;
											assign node193 = (inp[0]) ? node211 : node194;
												assign node194 = (inp[2]) ? node206 : node195;
													assign node195 = (inp[14]) ? node201 : node196;
														assign node196 = (inp[13]) ? node198 : 1'b0;
															assign node198 = (inp[11]) ? 1'b0 : 1'b1;
														assign node201 = (inp[13]) ? node203 : 1'b1;
															assign node203 = (inp[11]) ? 1'b1 : 1'b0;
													assign node206 = (inp[11]) ? 1'b0 : node207;
														assign node207 = (inp[13]) ? 1'b1 : 1'b0;
												assign node211 = (inp[4]) ? node213 : 1'b1;
													assign node213 = (inp[2]) ? node225 : node214;
														assign node214 = (inp[14]) ? node220 : node215;
															assign node215 = (inp[11]) ? 1'b0 : node216;
																assign node216 = (inp[13]) ? 1'b1 : 1'b0;
															assign node220 = (inp[13]) ? node222 : 1'b1;
																assign node222 = (inp[11]) ? 1'b1 : 1'b0;
														assign node225 = (inp[13]) ? node227 : 1'b0;
															assign node227 = (inp[11]) ? 1'b0 : 1'b1;
										assign node230 = (inp[4]) ? 1'b1 : node231;
											assign node231 = (inp[0]) ? node233 : 1'b1;
												assign node233 = (inp[2]) ? node245 : node234;
													assign node234 = (inp[14]) ? node240 : node235;
														assign node235 = (inp[11]) ? 1'b0 : node236;
															assign node236 = (inp[13]) ? 1'b1 : 1'b0;
														assign node240 = (inp[11]) ? 1'b1 : node241;
															assign node241 = (inp[13]) ? 1'b0 : 1'b1;
													assign node245 = (inp[13]) ? node247 : 1'b0;
														assign node247 = (inp[11]) ? 1'b0 : 1'b1;
									assign node251 = (inp[1]) ? node273 : node252;
										assign node252 = (inp[4]) ? 1'b0 : node253;
											assign node253 = (inp[0]) ? node255 : 1'b0;
												assign node255 = (inp[14]) ? node261 : node256;
													assign node256 = (inp[13]) ? node258 : 1'b1;
														assign node258 = (inp[11]) ? 1'b1 : 1'b0;
													assign node261 = (inp[2]) ? node267 : node262;
														assign node262 = (inp[13]) ? node264 : 1'b0;
															assign node264 = (inp[11]) ? 1'b0 : 1'b1;
														assign node267 = (inp[13]) ? node269 : 1'b1;
															assign node269 = (inp[11]) ? 1'b1 : 1'b0;
										assign node273 = (inp[8]) ? node311 : node274;
											assign node274 = (inp[4]) ? node294 : node275;
												assign node275 = (inp[0]) ? 1'b0 : node276;
													assign node276 = (inp[13]) ? node282 : node277;
														assign node277 = (inp[2]) ? 1'b1 : node278;
															assign node278 = (inp[14]) ? 1'b0 : 1'b1;
														assign node282 = (inp[11]) ? node288 : node283;
															assign node283 = (inp[14]) ? node285 : 1'b0;
																assign node285 = (inp[2]) ? 1'b0 : 1'b1;
															assign node288 = (inp[2]) ? 1'b1 : node289;
																assign node289 = (inp[14]) ? 1'b0 : 1'b1;
												assign node294 = (inp[14]) ? node300 : node295;
													assign node295 = (inp[11]) ? 1'b1 : node296;
														assign node296 = (inp[13]) ? 1'b0 : 1'b1;
													assign node300 = (inp[2]) ? node306 : node301;
														assign node301 = (inp[11]) ? 1'b0 : node302;
															assign node302 = (inp[13]) ? 1'b1 : 1'b0;
														assign node306 = (inp[11]) ? 1'b1 : node307;
															assign node307 = (inp[13]) ? 1'b0 : 1'b1;
											assign node311 = (inp[0]) ? node313 : 1'b0;
												assign node313 = (inp[4]) ? 1'b0 : node314;
													assign node314 = (inp[2]) ? node326 : node315;
														assign node315 = (inp[14]) ? node321 : node316;
															assign node316 = (inp[11]) ? 1'b1 : node317;
																assign node317 = (inp[13]) ? 1'b0 : 1'b1;
															assign node321 = (inp[11]) ? 1'b0 : node322;
																assign node322 = (inp[13]) ? 1'b1 : 1'b0;
														assign node326 = (inp[13]) ? node328 : 1'b1;
															assign node328 = (inp[11]) ? 1'b1 : 1'b0;
							assign node332 = (inp[3]) ? node412 : node333;
								assign node333 = (inp[8]) ? node391 : node334;
									assign node334 = (inp[1]) ? node356 : node335;
										assign node335 = (inp[0]) ? node337 : 1'b1;
											assign node337 = (inp[4]) ? 1'b1 : node338;
												assign node338 = (inp[11]) ? node350 : node339;
													assign node339 = (inp[13]) ? node345 : node340;
														assign node340 = (inp[2]) ? 1'b0 : node341;
															assign node341 = (inp[14]) ? 1'b1 : 1'b0;
														assign node345 = (inp[2]) ? 1'b1 : node346;
															assign node346 = (inp[14]) ? 1'b0 : 1'b1;
													assign node350 = (inp[2]) ? 1'b0 : node351;
														assign node351 = (inp[14]) ? 1'b1 : 1'b0;
										assign node356 = (inp[0]) ? node374 : node357;
											assign node357 = (inp[13]) ? node363 : node358;
												assign node358 = (inp[14]) ? node360 : 1'b0;
													assign node360 = (inp[2]) ? 1'b0 : 1'b1;
												assign node363 = (inp[11]) ? node369 : node364;
													assign node364 = (inp[14]) ? node366 : 1'b1;
														assign node366 = (inp[2]) ? 1'b1 : 1'b0;
													assign node369 = (inp[2]) ? 1'b0 : node370;
														assign node370 = (inp[14]) ? 1'b1 : 1'b0;
											assign node374 = (inp[4]) ? node376 : 1'b1;
												assign node376 = (inp[11]) ? node386 : node377;
													assign node377 = (inp[13]) ? node381 : node378;
														assign node378 = (inp[2]) ? 1'b0 : 1'b1;
														assign node381 = (inp[14]) ? node383 : 1'b1;
															assign node383 = (inp[2]) ? 1'b1 : 1'b0;
													assign node386 = (inp[2]) ? 1'b0 : node387;
														assign node387 = (inp[14]) ? 1'b1 : 1'b0;
									assign node391 = (inp[4]) ? 1'b1 : node392;
										assign node392 = (inp[0]) ? node394 : 1'b1;
											assign node394 = (inp[11]) ? node406 : node395;
												assign node395 = (inp[13]) ? node401 : node396;
													assign node396 = (inp[2]) ? 1'b0 : node397;
														assign node397 = (inp[14]) ? 1'b1 : 1'b0;
													assign node401 = (inp[2]) ? 1'b1 : node402;
														assign node402 = (inp[14]) ? 1'b0 : 1'b1;
												assign node406 = (inp[14]) ? node408 : 1'b0;
													assign node408 = (inp[2]) ? 1'b0 : 1'b1;
								assign node412 = (inp[7]) ? node494 : node413;
									assign node413 = (inp[8]) ? node473 : node414;
										assign node414 = (inp[1]) ? node436 : node415;
											assign node415 = (inp[4]) ? 1'b0 : node416;
												assign node416 = (inp[0]) ? node418 : 1'b0;
													assign node418 = (inp[14]) ? node424 : node419;
														assign node419 = (inp[13]) ? node421 : 1'b1;
															assign node421 = (inp[11]) ? 1'b1 : 1'b0;
														assign node424 = (inp[2]) ? node430 : node425;
															assign node425 = (inp[11]) ? 1'b0 : node426;
																assign node426 = (inp[13]) ? 1'b1 : 1'b0;
															assign node430 = (inp[13]) ? node432 : 1'b1;
																assign node432 = (inp[11]) ? 1'b1 : 1'b0;
											assign node436 = (inp[0]) ? node454 : node437;
												assign node437 = (inp[13]) ? node443 : node438;
													assign node438 = (inp[14]) ? node440 : 1'b1;
														assign node440 = (inp[2]) ? 1'b1 : 1'b0;
													assign node443 = (inp[11]) ? node449 : node444;
														assign node444 = (inp[2]) ? 1'b0 : node445;
															assign node445 = (inp[14]) ? 1'b1 : 1'b0;
														assign node449 = (inp[14]) ? node451 : 1'b1;
															assign node451 = (inp[2]) ? 1'b1 : 1'b0;
												assign node454 = (inp[4]) ? node456 : 1'b0;
													assign node456 = (inp[13]) ? node462 : node457;
														assign node457 = (inp[2]) ? 1'b1 : node458;
															assign node458 = (inp[14]) ? 1'b0 : 1'b1;
														assign node462 = (inp[11]) ? node468 : node463;
															assign node463 = (inp[2]) ? 1'b0 : node464;
																assign node464 = (inp[14]) ? 1'b1 : 1'b0;
															assign node468 = (inp[14]) ? node470 : 1'b1;
																assign node470 = (inp[2]) ? 1'b1 : 1'b0;
										assign node473 = (inp[4]) ? 1'b0 : node474;
											assign node474 = (inp[0]) ? node476 : 1'b0;
												assign node476 = (inp[2]) ? node488 : node477;
													assign node477 = (inp[14]) ? node483 : node478;
														assign node478 = (inp[13]) ? node480 : 1'b1;
															assign node480 = (inp[11]) ? 1'b1 : 1'b0;
														assign node483 = (inp[11]) ? 1'b0 : node484;
															assign node484 = (inp[13]) ? 1'b1 : 1'b0;
													assign node488 = (inp[11]) ? 1'b1 : node489;
														assign node489 = (inp[13]) ? 1'b0 : 1'b1;
									assign node494 = (inp[0]) ? node516 : node495;
										assign node495 = (inp[8]) ? 1'b1 : node496;
											assign node496 = (inp[1]) ? node498 : 1'b1;
												assign node498 = (inp[14]) ? node504 : node499;
													assign node499 = (inp[13]) ? node501 : 1'b0;
														assign node501 = (inp[11]) ? 1'b0 : 1'b1;
													assign node504 = (inp[2]) ? node510 : node505;
														assign node505 = (inp[13]) ? node507 : 1'b1;
															assign node507 = (inp[11]) ? 1'b1 : 1'b0;
														assign node510 = (inp[11]) ? 1'b0 : node511;
															assign node511 = (inp[13]) ? 1'b1 : 1'b0;
										assign node516 = (inp[4]) ? node550 : node517;
											assign node517 = (inp[1]) ? node535 : node518;
												assign node518 = (inp[14]) ? node524 : node519;
													assign node519 = (inp[13]) ? node521 : 1'b0;
														assign node521 = (inp[11]) ? 1'b0 : 1'b1;
													assign node524 = (inp[2]) ? node530 : node525;
														assign node525 = (inp[13]) ? node527 : 1'b1;
															assign node527 = (inp[11]) ? 1'b1 : 1'b0;
														assign node530 = (inp[11]) ? 1'b0 : node531;
															assign node531 = (inp[13]) ? 1'b1 : 1'b0;
												assign node535 = (inp[8]) ? node537 : 1'b1;
													assign node537 = (inp[11]) ? node545 : node538;
														assign node538 = (inp[13]) ? 1'b1 : node539;
															assign node539 = (inp[2]) ? 1'b0 : node540;
																assign node540 = (inp[14]) ? 1'b1 : 1'b0;
														assign node545 = (inp[2]) ? 1'b0 : node546;
															assign node546 = (inp[13]) ? 1'b0 : 1'b1;
											assign node550 = (inp[8]) ? 1'b1 : node551;
												assign node551 = (inp[1]) ? node553 : 1'b1;
													assign node553 = (inp[13]) ? node559 : node554;
														assign node554 = (inp[14]) ? node556 : 1'b0;
															assign node556 = (inp[2]) ? 1'b0 : 1'b1;
														assign node559 = (inp[11]) ? node565 : node560;
															assign node560 = (inp[14]) ? node562 : 1'b1;
																assign node562 = (inp[2]) ? 1'b1 : 1'b0;
															assign node565 = (inp[2]) ? 1'b0 : 1'b1;
						assign node569 = (inp[7]) ? node733 : node570;
							assign node570 = (inp[3]) ? node652 : node571;
								assign node571 = (inp[1]) ? node593 : node572;
									assign node572 = (inp[0]) ? node574 : 1'b0;
										assign node574 = (inp[4]) ? 1'b0 : node575;
											assign node575 = (inp[2]) ? node587 : node576;
												assign node576 = (inp[14]) ? node582 : node577;
													assign node577 = (inp[13]) ? node579 : 1'b1;
														assign node579 = (inp[11]) ? 1'b1 : 1'b0;
													assign node582 = (inp[13]) ? node584 : 1'b0;
														assign node584 = (inp[11]) ? 1'b0 : 1'b1;
												assign node587 = (inp[11]) ? 1'b1 : node588;
													assign node588 = (inp[13]) ? 1'b0 : 1'b1;
									assign node593 = (inp[8]) ? node631 : node594;
										assign node594 = (inp[0]) ? node612 : node595;
											assign node595 = (inp[14]) ? node601 : node596;
												assign node596 = (inp[11]) ? 1'b1 : node597;
													assign node597 = (inp[13]) ? 1'b0 : 1'b1;
												assign node601 = (inp[2]) ? node607 : node602;
													assign node602 = (inp[13]) ? node604 : 1'b0;
														assign node604 = (inp[11]) ? 1'b0 : 1'b1;
													assign node607 = (inp[11]) ? 1'b1 : node608;
														assign node608 = (inp[13]) ? 1'b0 : 1'b1;
											assign node612 = (inp[4]) ? node614 : 1'b0;
												assign node614 = (inp[2]) ? node626 : node615;
													assign node615 = (inp[14]) ? node621 : node616;
														assign node616 = (inp[13]) ? node618 : 1'b1;
															assign node618 = (inp[11]) ? 1'b1 : 1'b0;
														assign node621 = (inp[11]) ? 1'b0 : node622;
															assign node622 = (inp[13]) ? 1'b1 : 1'b0;
													assign node626 = (inp[11]) ? 1'b1 : node627;
														assign node627 = (inp[13]) ? 1'b0 : 1'b1;
										assign node631 = (inp[4]) ? 1'b0 : node632;
											assign node632 = (inp[0]) ? node634 : 1'b0;
												assign node634 = (inp[2]) ? node646 : node635;
													assign node635 = (inp[14]) ? node641 : node636;
														assign node636 = (inp[13]) ? node638 : 1'b1;
															assign node638 = (inp[11]) ? 1'b1 : 1'b0;
														assign node641 = (inp[11]) ? 1'b0 : node642;
															assign node642 = (inp[13]) ? 1'b1 : 1'b0;
													assign node646 = (inp[13]) ? node648 : 1'b1;
														assign node648 = (inp[11]) ? 1'b1 : 1'b0;
								assign node652 = (inp[4]) ? node712 : node653;
									assign node653 = (inp[0]) ? node675 : node654;
										assign node654 = (inp[8]) ? 1'b1 : node655;
											assign node655 = (inp[1]) ? node657 : 1'b1;
												assign node657 = (inp[11]) ? node669 : node658;
													assign node658 = (inp[13]) ? node664 : node659;
														assign node659 = (inp[14]) ? node661 : 1'b0;
															assign node661 = (inp[2]) ? 1'b0 : 1'b1;
														assign node664 = (inp[14]) ? node666 : 1'b1;
															assign node666 = (inp[2]) ? 1'b1 : 1'b0;
													assign node669 = (inp[14]) ? node671 : 1'b0;
														assign node671 = (inp[2]) ? 1'b0 : 1'b1;
										assign node675 = (inp[8]) ? node695 : node676;
											assign node676 = (inp[1]) ? 1'b1 : node677;
												assign node677 = (inp[2]) ? node689 : node678;
													assign node678 = (inp[14]) ? node684 : node679;
														assign node679 = (inp[11]) ? 1'b0 : node680;
															assign node680 = (inp[13]) ? 1'b1 : 1'b0;
														assign node684 = (inp[13]) ? node686 : 1'b1;
															assign node686 = (inp[11]) ? 1'b1 : 1'b0;
													assign node689 = (inp[13]) ? node691 : 1'b0;
														assign node691 = (inp[11]) ? 1'b0 : 1'b1;
											assign node695 = (inp[13]) ? node701 : node696;
												assign node696 = (inp[14]) ? node698 : 1'b0;
													assign node698 = (inp[2]) ? 1'b0 : 1'b1;
												assign node701 = (inp[11]) ? node707 : node702;
													assign node702 = (inp[14]) ? node704 : 1'b1;
														assign node704 = (inp[2]) ? 1'b1 : 1'b0;
													assign node707 = (inp[2]) ? 1'b0 : node708;
														assign node708 = (inp[14]) ? 1'b1 : 1'b0;
									assign node712 = (inp[8]) ? 1'b1 : node713;
										assign node713 = (inp[1]) ? node715 : 1'b1;
											assign node715 = (inp[13]) ? node721 : node716;
												assign node716 = (inp[2]) ? 1'b0 : node717;
													assign node717 = (inp[14]) ? 1'b1 : 1'b0;
												assign node721 = (inp[11]) ? node727 : node722;
													assign node722 = (inp[2]) ? 1'b1 : node723;
														assign node723 = (inp[14]) ? 1'b0 : 1'b1;
													assign node727 = (inp[14]) ? node729 : 1'b0;
														assign node729 = (inp[2]) ? 1'b0 : 1'b1;
							assign node733 = (inp[8]) ? node793 : node734;
								assign node734 = (inp[1]) ? node756 : node735;
									assign node735 = (inp[4]) ? 1'b0 : node736;
										assign node736 = (inp[0]) ? node738 : 1'b0;
											assign node738 = (inp[2]) ? node750 : node739;
												assign node739 = (inp[14]) ? node745 : node740;
													assign node740 = (inp[13]) ? node742 : 1'b1;
														assign node742 = (inp[11]) ? 1'b1 : 1'b0;
													assign node745 = (inp[11]) ? 1'b0 : node746;
														assign node746 = (inp[13]) ? 1'b1 : 1'b0;
												assign node750 = (inp[13]) ? node752 : 1'b1;
													assign node752 = (inp[11]) ? 1'b1 : 1'b0;
									assign node756 = (inp[0]) ? node774 : node757;
										assign node757 = (inp[2]) ? node769 : node758;
											assign node758 = (inp[14]) ? node764 : node759;
												assign node759 = (inp[13]) ? node761 : 1'b1;
													assign node761 = (inp[11]) ? 1'b1 : 1'b0;
												assign node764 = (inp[11]) ? 1'b0 : node765;
													assign node765 = (inp[13]) ? 1'b1 : 1'b0;
											assign node769 = (inp[11]) ? 1'b1 : node770;
												assign node770 = (inp[13]) ? 1'b0 : 1'b1;
										assign node774 = (inp[4]) ? node776 : 1'b0;
											assign node776 = (inp[14]) ? node782 : node777;
												assign node777 = (inp[11]) ? 1'b1 : node778;
													assign node778 = (inp[13]) ? 1'b0 : 1'b1;
												assign node782 = (inp[2]) ? node788 : node783;
													assign node783 = (inp[13]) ? node785 : 1'b0;
														assign node785 = (inp[11]) ? 1'b0 : 1'b1;
													assign node788 = (inp[11]) ? 1'b1 : node789;
														assign node789 = (inp[13]) ? 1'b0 : 1'b1;
								assign node793 = (inp[0]) ? node795 : 1'b0;
									assign node795 = (inp[4]) ? 1'b0 : node796;
										assign node796 = (inp[13]) ? node802 : node797;
											assign node797 = (inp[14]) ? node799 : 1'b1;
												assign node799 = (inp[2]) ? 1'b1 : 1'b0;
											assign node802 = (inp[11]) ? node808 : node803;
												assign node803 = (inp[14]) ? node805 : 1'b0;
													assign node805 = (inp[2]) ? 1'b0 : 1'b1;
												assign node808 = (inp[14]) ? node810 : 1'b1;
													assign node810 = (inp[2]) ? 1'b1 : 1'b0;
					assign node814 = (inp[4]) ? node874 : node815;
						assign node815 = (inp[0]) ? node837 : node816;
							assign node816 = (inp[1]) ? node818 : 1'b1;
								assign node818 = (inp[8]) ? 1'b1 : node819;
									assign node819 = (inp[14]) ? node825 : node820;
										assign node820 = (inp[11]) ? 1'b0 : node821;
											assign node821 = (inp[13]) ? 1'b1 : 1'b0;
										assign node825 = (inp[2]) ? node831 : node826;
											assign node826 = (inp[11]) ? 1'b1 : node827;
												assign node827 = (inp[13]) ? 1'b0 : 1'b1;
											assign node831 = (inp[11]) ? 1'b0 : node832;
												assign node832 = (inp[13]) ? 1'b1 : 1'b0;
							assign node837 = (inp[8]) ? node857 : node838;
								assign node838 = (inp[1]) ? 1'b1 : node839;
									assign node839 = (inp[14]) ? node845 : node840;
										assign node840 = (inp[11]) ? 1'b0 : node841;
											assign node841 = (inp[13]) ? 1'b1 : 1'b0;
										assign node845 = (inp[2]) ? node851 : node846;
											assign node846 = (inp[11]) ? 1'b1 : node847;
												assign node847 = (inp[13]) ? 1'b0 : 1'b1;
											assign node851 = (inp[13]) ? node853 : 1'b0;
												assign node853 = (inp[11]) ? 1'b0 : 1'b1;
								assign node857 = (inp[14]) ? node863 : node858;
									assign node858 = (inp[13]) ? node860 : 1'b0;
										assign node860 = (inp[11]) ? 1'b0 : 1'b1;
									assign node863 = (inp[2]) ? node869 : node864;
										assign node864 = (inp[11]) ? 1'b1 : node865;
											assign node865 = (inp[13]) ? 1'b0 : 1'b1;
										assign node869 = (inp[11]) ? 1'b0 : node870;
											assign node870 = (inp[13]) ? 1'b1 : 1'b0;
						assign node874 = (inp[8]) ? 1'b1 : node875;
							assign node875 = (inp[1]) ? node877 : 1'b1;
								assign node877 = (inp[13]) ? node883 : node878;
									assign node878 = (inp[14]) ? node880 : 1'b0;
										assign node880 = (inp[2]) ? 1'b0 : 1'b1;
									assign node883 = (inp[11]) ? node889 : node884;
										assign node884 = (inp[2]) ? 1'b1 : node885;
											assign node885 = (inp[14]) ? 1'b0 : 1'b1;
										assign node889 = (inp[2]) ? 1'b0 : node890;
											assign node890 = (inp[14]) ? 1'b1 : 1'b0;
			assign node895 = (inp[15]) ? node1703 : node896;
				assign node896 = (inp[12]) ? node1622 : node897;
					assign node897 = (inp[10]) ? node1377 : node898;
						assign node898 = (inp[9]) ? node1140 : node899;
							assign node899 = (inp[3]) ? node981 : node900;
								assign node900 = (inp[4]) ? node960 : node901;
									assign node901 = (inp[0]) ? node923 : node902;
										assign node902 = (inp[1]) ? node904 : 1'b0;
											assign node904 = (inp[8]) ? 1'b0 : node905;
												assign node905 = (inp[2]) ? node917 : node906;
													assign node906 = (inp[14]) ? node912 : node907;
														assign node907 = (inp[11]) ? 1'b1 : node908;
															assign node908 = (inp[13]) ? 1'b0 : 1'b1;
														assign node912 = (inp[11]) ? 1'b0 : node913;
															assign node913 = (inp[13]) ? 1'b1 : 1'b0;
													assign node917 = (inp[13]) ? node919 : 1'b1;
														assign node919 = (inp[11]) ? 1'b1 : 1'b0;
										assign node923 = (inp[8]) ? node943 : node924;
											assign node924 = (inp[1]) ? 1'b0 : node925;
												assign node925 = (inp[13]) ? node931 : node926;
													assign node926 = (inp[14]) ? node928 : 1'b1;
														assign node928 = (inp[2]) ? 1'b1 : 1'b0;
													assign node931 = (inp[11]) ? node937 : node932;
														assign node932 = (inp[2]) ? 1'b0 : node933;
															assign node933 = (inp[14]) ? 1'b1 : 1'b0;
														assign node937 = (inp[14]) ? node939 : 1'b1;
															assign node939 = (inp[2]) ? 1'b1 : 1'b0;
											assign node943 = (inp[14]) ? node949 : node944;
												assign node944 = (inp[11]) ? 1'b1 : node945;
													assign node945 = (inp[13]) ? 1'b0 : 1'b1;
												assign node949 = (inp[2]) ? node955 : node950;
													assign node950 = (inp[11]) ? 1'b0 : node951;
														assign node951 = (inp[13]) ? 1'b1 : 1'b0;
													assign node955 = (inp[13]) ? node957 : 1'b1;
														assign node957 = (inp[11]) ? 1'b1 : 1'b0;
									assign node960 = (inp[1]) ? node962 : 1'b0;
										assign node962 = (inp[8]) ? 1'b0 : node963;
											assign node963 = (inp[14]) ? node969 : node964;
												assign node964 = (inp[13]) ? node966 : 1'b1;
													assign node966 = (inp[11]) ? 1'b1 : 1'b0;
												assign node969 = (inp[2]) ? node975 : node970;
													assign node970 = (inp[13]) ? node972 : 1'b0;
														assign node972 = (inp[11]) ? 1'b0 : 1'b1;
													assign node975 = (inp[13]) ? node977 : 1'b1;
														assign node977 = (inp[11]) ? 1'b1 : 1'b0;
								assign node981 = (inp[7]) ? node1063 : node982;
									assign node982 = (inp[8]) ? node1042 : node983;
										assign node983 = (inp[1]) ? node1005 : node984;
											assign node984 = (inp[4]) ? 1'b1 : node985;
												assign node985 = (inp[0]) ? node987 : 1'b1;
													assign node987 = (inp[11]) ? node999 : node988;
														assign node988 = (inp[13]) ? node994 : node989;
															assign node989 = (inp[14]) ? node991 : 1'b0;
																assign node991 = (inp[2]) ? 1'b0 : 1'b1;
															assign node994 = (inp[14]) ? node996 : 1'b1;
																assign node996 = (inp[2]) ? 1'b1 : 1'b0;
														assign node999 = (inp[14]) ? node1001 : 1'b0;
															assign node1001 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1005 = (inp[0]) ? node1023 : node1006;
												assign node1006 = (inp[2]) ? node1018 : node1007;
													assign node1007 = (inp[14]) ? node1013 : node1008;
														assign node1008 = (inp[11]) ? 1'b0 : node1009;
															assign node1009 = (inp[13]) ? 1'b1 : 1'b0;
														assign node1013 = (inp[11]) ? 1'b1 : node1014;
															assign node1014 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1018 = (inp[11]) ? 1'b0 : node1019;
														assign node1019 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1023 = (inp[4]) ? node1025 : 1'b1;
													assign node1025 = (inp[14]) ? node1031 : node1026;
														assign node1026 = (inp[11]) ? 1'b0 : node1027;
															assign node1027 = (inp[13]) ? 1'b1 : 1'b0;
														assign node1031 = (inp[2]) ? node1037 : node1032;
															assign node1032 = (inp[11]) ? 1'b1 : node1033;
																assign node1033 = (inp[13]) ? 1'b0 : 1'b1;
															assign node1037 = (inp[13]) ? node1039 : 1'b0;
																assign node1039 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1042 = (inp[4]) ? 1'b1 : node1043;
											assign node1043 = (inp[0]) ? node1045 : 1'b1;
												assign node1045 = (inp[11]) ? node1057 : node1046;
													assign node1046 = (inp[13]) ? node1052 : node1047;
														assign node1047 = (inp[14]) ? node1049 : 1'b0;
															assign node1049 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1052 = (inp[14]) ? node1054 : 1'b1;
															assign node1054 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1057 = (inp[2]) ? 1'b0 : node1058;
														assign node1058 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1063 = (inp[8]) ? node1119 : node1064;
										assign node1064 = (inp[1]) ? node1086 : node1065;
											assign node1065 = (inp[0]) ? node1067 : 1'b0;
												assign node1067 = (inp[4]) ? 1'b0 : node1068;
													assign node1068 = (inp[11]) ? node1080 : node1069;
														assign node1069 = (inp[13]) ? node1075 : node1070;
															assign node1070 = (inp[2]) ? 1'b1 : node1071;
																assign node1071 = (inp[14]) ? 1'b0 : 1'b1;
															assign node1075 = (inp[14]) ? node1077 : 1'b0;
																assign node1077 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1080 = (inp[14]) ? node1082 : 1'b1;
															assign node1082 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1086 = (inp[4]) ? node1102 : node1087;
												assign node1087 = (inp[0]) ? 1'b0 : node1088;
													assign node1088 = (inp[13]) ? node1090 : 1'b1;
														assign node1090 = (inp[11]) ? node1096 : node1091;
															assign node1091 = (inp[14]) ? node1093 : 1'b0;
																assign node1093 = (inp[2]) ? 1'b0 : 1'b1;
															assign node1096 = (inp[14]) ? node1098 : 1'b1;
																assign node1098 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1102 = (inp[11]) ? node1114 : node1103;
													assign node1103 = (inp[13]) ? node1109 : node1104;
														assign node1104 = (inp[14]) ? node1106 : 1'b1;
															assign node1106 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1109 = (inp[2]) ? 1'b0 : node1110;
															assign node1110 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1114 = (inp[2]) ? 1'b1 : node1115;
														assign node1115 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1119 = (inp[4]) ? 1'b0 : node1120;
											assign node1120 = (inp[0]) ? node1122 : 1'b0;
												assign node1122 = (inp[11]) ? node1134 : node1123;
													assign node1123 = (inp[13]) ? node1129 : node1124;
														assign node1124 = (inp[2]) ? 1'b1 : node1125;
															assign node1125 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1129 = (inp[14]) ? node1131 : 1'b0;
															assign node1131 = (inp[1]) ? 1'b0 : 1'b1;
													assign node1134 = (inp[14]) ? node1136 : 1'b1;
														assign node1136 = (inp[2]) ? 1'b1 : 1'b0;
							assign node1140 = (inp[7]) ? node1296 : node1141;
								assign node1141 = (inp[3]) ? node1217 : node1142;
									assign node1142 = (inp[4]) ? node1196 : node1143;
										assign node1143 = (inp[0]) ? node1165 : node1144;
											assign node1144 = (inp[1]) ? node1146 : 1'b1;
												assign node1146 = (inp[8]) ? 1'b1 : node1147;
													assign node1147 = (inp[11]) ? node1159 : node1148;
														assign node1148 = (inp[13]) ? node1154 : node1149;
															assign node1149 = (inp[14]) ? node1151 : 1'b0;
																assign node1151 = (inp[2]) ? 1'b0 : 1'b1;
															assign node1154 = (inp[2]) ? 1'b1 : node1155;
																assign node1155 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1159 = (inp[14]) ? node1161 : 1'b0;
															assign node1161 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1165 = (inp[1]) ? node1185 : node1166;
												assign node1166 = (inp[14]) ? node1172 : node1167;
													assign node1167 = (inp[11]) ? 1'b0 : node1168;
														assign node1168 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1172 = (inp[2]) ? node1178 : node1173;
														assign node1173 = (inp[13]) ? node1175 : 1'b1;
															assign node1175 = (inp[11]) ? 1'b1 : 1'b0;
														assign node1178 = (inp[8]) ? node1180 : 1'b0;
															assign node1180 = (inp[13]) ? node1182 : 1'b0;
																assign node1182 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1185 = (inp[8]) ? node1187 : 1'b1;
													assign node1187 = (inp[13]) ? node1189 : 1'b0;
														assign node1189 = (inp[11]) ? node1191 : 1'b1;
															assign node1191 = (inp[2]) ? 1'b0 : node1192;
																assign node1192 = (inp[14]) ? 1'b1 : 1'b0;
										assign node1196 = (inp[1]) ? node1198 : 1'b1;
											assign node1198 = (inp[8]) ? 1'b1 : node1199;
												assign node1199 = (inp[13]) ? node1205 : node1200;
													assign node1200 = (inp[14]) ? node1202 : 1'b0;
														assign node1202 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1205 = (inp[11]) ? node1211 : node1206;
														assign node1206 = (inp[14]) ? node1208 : 1'b1;
															assign node1208 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1211 = (inp[14]) ? node1213 : 1'b0;
															assign node1213 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1217 = (inp[8]) ? node1275 : node1218;
										assign node1218 = (inp[1]) ? node1240 : node1219;
											assign node1219 = (inp[0]) ? node1221 : 1'b0;
												assign node1221 = (inp[4]) ? 1'b0 : node1222;
													assign node1222 = (inp[13]) ? node1228 : node1223;
														assign node1223 = (inp[14]) ? node1225 : 1'b1;
															assign node1225 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1228 = (inp[11]) ? node1234 : node1229;
															assign node1229 = (inp[14]) ? node1231 : 1'b0;
																assign node1231 = (inp[2]) ? 1'b0 : 1'b1;
															assign node1234 = (inp[2]) ? 1'b1 : node1235;
																assign node1235 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1240 = (inp[4]) ? node1258 : node1241;
												assign node1241 = (inp[0]) ? 1'b0 : node1242;
													assign node1242 = (inp[13]) ? node1248 : node1243;
														assign node1243 = (inp[14]) ? node1245 : 1'b1;
															assign node1245 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1248 = (inp[11]) ? node1254 : node1249;
															assign node1249 = (inp[14]) ? node1251 : 1'b0;
																assign node1251 = (inp[2]) ? 1'b0 : 1'b1;
															assign node1254 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1258 = (inp[11]) ? node1270 : node1259;
													assign node1259 = (inp[13]) ? node1265 : node1260;
														assign node1260 = (inp[2]) ? 1'b1 : node1261;
															assign node1261 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1265 = (inp[2]) ? 1'b0 : node1266;
															assign node1266 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1270 = (inp[14]) ? node1272 : 1'b1;
														assign node1272 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1275 = (inp[0]) ? node1277 : 1'b0;
											assign node1277 = (inp[4]) ? 1'b0 : node1278;
												assign node1278 = (inp[14]) ? node1284 : node1279;
													assign node1279 = (inp[11]) ? 1'b1 : node1280;
														assign node1280 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1284 = (inp[2]) ? node1290 : node1285;
														assign node1285 = (inp[13]) ? node1287 : 1'b0;
															assign node1287 = (inp[11]) ? 1'b0 : 1'b1;
														assign node1290 = (inp[11]) ? 1'b1 : node1291;
															assign node1291 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1296 = (inp[0]) ? node1318 : node1297;
									assign node1297 = (inp[8]) ? 1'b1 : node1298;
										assign node1298 = (inp[1]) ? node1300 : 1'b1;
											assign node1300 = (inp[2]) ? node1312 : node1301;
												assign node1301 = (inp[14]) ? node1307 : node1302;
													assign node1302 = (inp[13]) ? node1304 : 1'b0;
														assign node1304 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1307 = (inp[13]) ? node1309 : 1'b1;
														assign node1309 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1312 = (inp[11]) ? 1'b0 : node1313;
													assign node1313 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1318 = (inp[4]) ? node1356 : node1319;
										assign node1319 = (inp[8]) ? node1339 : node1320;
											assign node1320 = (inp[1]) ? 1'b1 : node1321;
												assign node1321 = (inp[11]) ? node1333 : node1322;
													assign node1322 = (inp[13]) ? node1328 : node1323;
														assign node1323 = (inp[14]) ? node1325 : 1'b0;
															assign node1325 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1328 = (inp[2]) ? 1'b1 : node1329;
															assign node1329 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1333 = (inp[2]) ? 1'b0 : node1334;
														assign node1334 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1339 = (inp[14]) ? node1345 : node1340;
												assign node1340 = (inp[11]) ? 1'b0 : node1341;
													assign node1341 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1345 = (inp[2]) ? node1351 : node1346;
													assign node1346 = (inp[11]) ? 1'b1 : node1347;
														assign node1347 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1351 = (inp[11]) ? 1'b0 : node1352;
														assign node1352 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1356 = (inp[8]) ? 1'b1 : node1357;
											assign node1357 = (inp[1]) ? node1359 : 1'b1;
												assign node1359 = (inp[14]) ? node1365 : node1360;
													assign node1360 = (inp[11]) ? 1'b0 : node1361;
														assign node1361 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1365 = (inp[2]) ? node1371 : node1366;
														assign node1366 = (inp[11]) ? 1'b1 : node1367;
															assign node1367 = (inp[13]) ? 1'b0 : 1'b1;
														assign node1371 = (inp[13]) ? node1373 : 1'b0;
															assign node1373 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1377 = (inp[3]) ? node1459 : node1378;
							assign node1378 = (inp[8]) ? node1438 : node1379;
								assign node1379 = (inp[1]) ? node1401 : node1380;
									assign node1380 = (inp[4]) ? 1'b0 : node1381;
										assign node1381 = (inp[0]) ? node1383 : 1'b0;
											assign node1383 = (inp[11]) ? node1395 : node1384;
												assign node1384 = (inp[13]) ? node1390 : node1385;
													assign node1385 = (inp[2]) ? 1'b1 : node1386;
														assign node1386 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1390 = (inp[14]) ? node1392 : 1'b0;
														assign node1392 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1395 = (inp[14]) ? node1397 : 1'b1;
													assign node1397 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1401 = (inp[0]) ? node1419 : node1402;
										assign node1402 = (inp[13]) ? node1408 : node1403;
											assign node1403 = (inp[14]) ? node1405 : 1'b1;
												assign node1405 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1408 = (inp[11]) ? node1414 : node1409;
												assign node1409 = (inp[2]) ? 1'b0 : node1410;
													assign node1410 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1414 = (inp[14]) ? node1416 : 1'b1;
													assign node1416 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1419 = (inp[4]) ? node1421 : 1'b0;
											assign node1421 = (inp[14]) ? node1427 : node1422;
												assign node1422 = (inp[13]) ? node1424 : 1'b1;
													assign node1424 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1427 = (inp[2]) ? node1433 : node1428;
													assign node1428 = (inp[11]) ? 1'b0 : node1429;
														assign node1429 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1433 = (inp[13]) ? node1435 : 1'b1;
														assign node1435 = (inp[11]) ? 1'b1 : 1'b0;
								assign node1438 = (inp[0]) ? node1440 : 1'b0;
									assign node1440 = (inp[4]) ? 1'b0 : node1441;
										assign node1441 = (inp[2]) ? node1453 : node1442;
											assign node1442 = (inp[14]) ? node1448 : node1443;
												assign node1443 = (inp[13]) ? node1445 : 1'b1;
													assign node1445 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1448 = (inp[11]) ? 1'b0 : node1449;
													assign node1449 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1453 = (inp[13]) ? node1455 : 1'b1;
												assign node1455 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1459 = (inp[7]) ? node1541 : node1460;
								assign node1460 = (inp[4]) ? node1520 : node1461;
									assign node1461 = (inp[0]) ? node1483 : node1462;
										assign node1462 = (inp[8]) ? 1'b1 : node1463;
											assign node1463 = (inp[1]) ? node1465 : 1'b1;
												assign node1465 = (inp[14]) ? node1471 : node1466;
													assign node1466 = (inp[13]) ? node1468 : 1'b0;
														assign node1468 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1471 = (inp[2]) ? node1477 : node1472;
														assign node1472 = (inp[13]) ? node1474 : 1'b1;
															assign node1474 = (inp[11]) ? 1'b1 : 1'b0;
														assign node1477 = (inp[13]) ? node1479 : 1'b0;
															assign node1479 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1483 = (inp[1]) ? node1501 : node1484;
											assign node1484 = (inp[13]) ? node1490 : node1485;
												assign node1485 = (inp[2]) ? 1'b0 : node1486;
													assign node1486 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1490 = (inp[11]) ? node1496 : node1491;
													assign node1491 = (inp[2]) ? 1'b1 : node1492;
														assign node1492 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1496 = (inp[2]) ? 1'b0 : node1497;
														assign node1497 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1501 = (inp[8]) ? node1503 : 1'b1;
												assign node1503 = (inp[11]) ? node1515 : node1504;
													assign node1504 = (inp[13]) ? node1510 : node1505;
														assign node1505 = (inp[14]) ? node1507 : 1'b0;
															assign node1507 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1510 = (inp[2]) ? 1'b1 : node1511;
															assign node1511 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1515 = (inp[2]) ? 1'b0 : node1516;
														assign node1516 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1520 = (inp[8]) ? 1'b1 : node1521;
										assign node1521 = (inp[1]) ? node1523 : 1'b1;
											assign node1523 = (inp[11]) ? node1535 : node1524;
												assign node1524 = (inp[13]) ? node1530 : node1525;
													assign node1525 = (inp[14]) ? node1527 : 1'b0;
														assign node1527 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1530 = (inp[14]) ? node1532 : 1'b1;
														assign node1532 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1535 = (inp[14]) ? node1537 : 1'b0;
													assign node1537 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1541 = (inp[8]) ? node1601 : node1542;
									assign node1542 = (inp[1]) ? node1564 : node1543;
										assign node1543 = (inp[4]) ? 1'b0 : node1544;
											assign node1544 = (inp[0]) ? node1546 : 1'b0;
												assign node1546 = (inp[2]) ? node1558 : node1547;
													assign node1547 = (inp[14]) ? node1553 : node1548;
														assign node1548 = (inp[13]) ? node1550 : 1'b1;
															assign node1550 = (inp[11]) ? 1'b1 : 1'b0;
														assign node1553 = (inp[11]) ? 1'b0 : node1554;
															assign node1554 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1558 = (inp[11]) ? 1'b1 : node1559;
														assign node1559 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1564 = (inp[4]) ? node1584 : node1565;
											assign node1565 = (inp[0]) ? 1'b0 : node1566;
												assign node1566 = (inp[11]) ? node1578 : node1567;
													assign node1567 = (inp[13]) ? node1573 : node1568;
														assign node1568 = (inp[14]) ? node1570 : 1'b1;
															assign node1570 = (inp[2]) ? 1'b1 : 1'b0;
														assign node1573 = (inp[2]) ? 1'b0 : node1574;
															assign node1574 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1578 = (inp[14]) ? node1580 : 1'b1;
														assign node1580 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1584 = (inp[11]) ? node1596 : node1585;
												assign node1585 = (inp[13]) ? node1591 : node1586;
													assign node1586 = (inp[2]) ? 1'b1 : node1587;
														assign node1587 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1591 = (inp[2]) ? 1'b0 : node1592;
														assign node1592 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1596 = (inp[14]) ? node1598 : 1'b1;
													assign node1598 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1601 = (inp[4]) ? 1'b0 : node1602;
										assign node1602 = (inp[0]) ? node1604 : 1'b0;
											assign node1604 = (inp[2]) ? node1616 : node1605;
												assign node1605 = (inp[14]) ? node1611 : node1606;
													assign node1606 = (inp[11]) ? 1'b1 : node1607;
														assign node1607 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1611 = (inp[13]) ? node1613 : 1'b0;
														assign node1613 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1616 = (inp[11]) ? 1'b1 : node1617;
													assign node1617 = (inp[13]) ? 1'b0 : 1'b1;
					assign node1622 = (inp[0]) ? node1644 : node1623;
						assign node1623 = (inp[1]) ? node1625 : 1'b1;
							assign node1625 = (inp[8]) ? 1'b1 : node1626;
								assign node1626 = (inp[13]) ? node1632 : node1627;
									assign node1627 = (inp[14]) ? node1629 : 1'b0;
										assign node1629 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1632 = (inp[11]) ? node1638 : node1633;
										assign node1633 = (inp[2]) ? 1'b1 : node1634;
											assign node1634 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1638 = (inp[2]) ? 1'b0 : node1639;
											assign node1639 = (inp[14]) ? 1'b1 : 1'b0;
						assign node1644 = (inp[4]) ? node1682 : node1645;
							assign node1645 = (inp[1]) ? node1663 : node1646;
								assign node1646 = (inp[13]) ? node1652 : node1647;
									assign node1647 = (inp[2]) ? 1'b0 : node1648;
										assign node1648 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1652 = (inp[11]) ? node1658 : node1653;
										assign node1653 = (inp[14]) ? node1655 : 1'b1;
											assign node1655 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1658 = (inp[2]) ? 1'b0 : node1659;
											assign node1659 = (inp[14]) ? 1'b1 : 1'b0;
								assign node1663 = (inp[8]) ? node1665 : 1'b1;
									assign node1665 = (inp[2]) ? node1677 : node1666;
										assign node1666 = (inp[14]) ? node1672 : node1667;
											assign node1667 = (inp[13]) ? node1669 : 1'b0;
												assign node1669 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1672 = (inp[13]) ? node1674 : 1'b1;
												assign node1674 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1677 = (inp[11]) ? 1'b0 : node1678;
											assign node1678 = (inp[13]) ? 1'b1 : 1'b0;
							assign node1682 = (inp[1]) ? node1684 : 1'b1;
								assign node1684 = (inp[8]) ? 1'b1 : node1685;
									assign node1685 = (inp[11]) ? node1697 : node1686;
										assign node1686 = (inp[13]) ? node1692 : node1687;
											assign node1687 = (inp[14]) ? node1689 : 1'b0;
												assign node1689 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1692 = (inp[2]) ? 1'b1 : node1693;
												assign node1693 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1697 = (inp[2]) ? 1'b0 : node1698;
											assign node1698 = (inp[14]) ? 1'b1 : 1'b0;
				assign node1703 = (inp[7]) ? node2195 : node1704;
					assign node1704 = (inp[3]) ? node1950 : node1705;
						assign node1705 = (inp[10]) ? node1869 : node1706;
							assign node1706 = (inp[9]) ? node1788 : node1707;
								assign node1707 = (inp[1]) ? node1729 : node1708;
									assign node1708 = (inp[4]) ? 1'b0 : node1709;
										assign node1709 = (inp[0]) ? node1711 : 1'b0;
											assign node1711 = (inp[13]) ? node1717 : node1712;
												assign node1712 = (inp[14]) ? node1714 : 1'b1;
													assign node1714 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1717 = (inp[11]) ? node1723 : node1718;
													assign node1718 = (inp[2]) ? 1'b0 : node1719;
														assign node1719 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1723 = (inp[2]) ? 1'b1 : node1724;
														assign node1724 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1729 = (inp[8]) ? node1767 : node1730;
										assign node1730 = (inp[4]) ? node1750 : node1731;
											assign node1731 = (inp[0]) ? 1'b0 : node1732;
												assign node1732 = (inp[2]) ? node1744 : node1733;
													assign node1733 = (inp[14]) ? node1739 : node1734;
														assign node1734 = (inp[11]) ? 1'b1 : node1735;
															assign node1735 = (inp[13]) ? 1'b0 : 1'b1;
														assign node1739 = (inp[13]) ? node1741 : 1'b0;
															assign node1741 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1744 = (inp[13]) ? node1746 : 1'b1;
														assign node1746 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1750 = (inp[11]) ? node1762 : node1751;
												assign node1751 = (inp[13]) ? node1757 : node1752;
													assign node1752 = (inp[14]) ? node1754 : 1'b1;
														assign node1754 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1757 = (inp[14]) ? node1759 : 1'b0;
														assign node1759 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1762 = (inp[2]) ? 1'b1 : node1763;
													assign node1763 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1767 = (inp[0]) ? node1769 : 1'b0;
											assign node1769 = (inp[4]) ? 1'b0 : node1770;
												assign node1770 = (inp[13]) ? node1776 : node1771;
													assign node1771 = (inp[2]) ? 1'b1 : node1772;
														assign node1772 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1776 = (inp[11]) ? node1782 : node1777;
														assign node1777 = (inp[14]) ? node1779 : 1'b0;
															assign node1779 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1782 = (inp[2]) ? 1'b1 : node1783;
															assign node1783 = (inp[14]) ? 1'b0 : 1'b1;
								assign node1788 = (inp[8]) ? node1848 : node1789;
									assign node1789 = (inp[1]) ? node1811 : node1790;
										assign node1790 = (inp[4]) ? 1'b1 : node1791;
											assign node1791 = (inp[0]) ? node1793 : 1'b1;
												assign node1793 = (inp[11]) ? node1805 : node1794;
													assign node1794 = (inp[13]) ? node1800 : node1795;
														assign node1795 = (inp[2]) ? 1'b0 : node1796;
															assign node1796 = (inp[14]) ? 1'b1 : 1'b0;
														assign node1800 = (inp[14]) ? node1802 : 1'b1;
															assign node1802 = (inp[12]) ? 1'b1 : 1'b0;
													assign node1805 = (inp[14]) ? node1807 : 1'b0;
														assign node1807 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1811 = (inp[4]) ? node1831 : node1812;
											assign node1812 = (inp[0]) ? 1'b1 : node1813;
												assign node1813 = (inp[2]) ? node1825 : node1814;
													assign node1814 = (inp[14]) ? node1820 : node1815;
														assign node1815 = (inp[13]) ? node1817 : 1'b0;
															assign node1817 = (inp[11]) ? 1'b0 : 1'b1;
														assign node1820 = (inp[13]) ? node1822 : 1'b1;
															assign node1822 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1825 = (inp[11]) ? 1'b0 : node1826;
														assign node1826 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1831 = (inp[13]) ? node1837 : node1832;
												assign node1832 = (inp[14]) ? node1834 : 1'b0;
													assign node1834 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1837 = (inp[11]) ? node1843 : node1838;
													assign node1838 = (inp[14]) ? node1840 : 1'b1;
														assign node1840 = (inp[2]) ? 1'b1 : 1'b0;
													assign node1843 = (inp[14]) ? node1845 : 1'b0;
														assign node1845 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1848 = (inp[0]) ? node1850 : 1'b1;
										assign node1850 = (inp[4]) ? 1'b1 : node1851;
											assign node1851 = (inp[11]) ? node1863 : node1852;
												assign node1852 = (inp[13]) ? node1858 : node1853;
													assign node1853 = (inp[14]) ? node1855 : 1'b0;
														assign node1855 = (inp[2]) ? 1'b0 : 1'b1;
													assign node1858 = (inp[14]) ? node1860 : 1'b1;
														assign node1860 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1863 = (inp[14]) ? node1865 : 1'b0;
													assign node1865 = (inp[2]) ? 1'b0 : 1'b1;
							assign node1869 = (inp[1]) ? node1891 : node1870;
								assign node1870 = (inp[4]) ? 1'b0 : node1871;
									assign node1871 = (inp[0]) ? node1873 : 1'b0;
										assign node1873 = (inp[14]) ? node1879 : node1874;
											assign node1874 = (inp[11]) ? 1'b1 : node1875;
												assign node1875 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1879 = (inp[2]) ? node1885 : node1880;
												assign node1880 = (inp[13]) ? node1882 : 1'b0;
													assign node1882 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1885 = (inp[11]) ? 1'b1 : node1886;
													assign node1886 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1891 = (inp[8]) ? node1929 : node1892;
									assign node1892 = (inp[4]) ? node1912 : node1893;
										assign node1893 = (inp[0]) ? 1'b0 : node1894;
											assign node1894 = (inp[14]) ? node1900 : node1895;
												assign node1895 = (inp[13]) ? node1897 : 1'b1;
													assign node1897 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1900 = (inp[2]) ? node1906 : node1901;
													assign node1901 = (inp[11]) ? 1'b0 : node1902;
														assign node1902 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1906 = (inp[11]) ? 1'b1 : node1907;
														assign node1907 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1912 = (inp[14]) ? node1918 : node1913;
											assign node1913 = (inp[13]) ? node1915 : 1'b1;
												assign node1915 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1918 = (inp[2]) ? node1924 : node1919;
												assign node1919 = (inp[11]) ? 1'b0 : node1920;
													assign node1920 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1924 = (inp[11]) ? 1'b1 : node1925;
													assign node1925 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1929 = (inp[4]) ? 1'b0 : node1930;
										assign node1930 = (inp[0]) ? node1932 : 1'b0;
											assign node1932 = (inp[2]) ? node1944 : node1933;
												assign node1933 = (inp[14]) ? node1939 : node1934;
													assign node1934 = (inp[11]) ? 1'b1 : node1935;
														assign node1935 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1939 = (inp[13]) ? node1941 : 1'b0;
														assign node1941 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1944 = (inp[13]) ? node1946 : 1'b1;
													assign node1946 = (inp[11]) ? 1'b1 : 1'b0;
						assign node1950 = (inp[9]) ? node2032 : node1951;
							assign node1951 = (inp[4]) ? node2011 : node1952;
								assign node1952 = (inp[0]) ? node1974 : node1953;
									assign node1953 = (inp[1]) ? node1955 : 1'b1;
										assign node1955 = (inp[8]) ? 1'b1 : node1956;
											assign node1956 = (inp[14]) ? node1962 : node1957;
												assign node1957 = (inp[11]) ? 1'b0 : node1958;
													assign node1958 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1962 = (inp[2]) ? node1968 : node1963;
													assign node1963 = (inp[11]) ? 1'b1 : node1964;
														assign node1964 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1968 = (inp[11]) ? 1'b0 : node1969;
														assign node1969 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1974 = (inp[1]) ? node1992 : node1975;
										assign node1975 = (inp[11]) ? node1987 : node1976;
											assign node1976 = (inp[13]) ? node1982 : node1977;
												assign node1977 = (inp[2]) ? 1'b0 : node1978;
													assign node1978 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1982 = (inp[14]) ? node1984 : 1'b1;
													assign node1984 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1987 = (inp[14]) ? node1989 : 1'b0;
												assign node1989 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1992 = (inp[8]) ? node1994 : 1'b1;
											assign node1994 = (inp[2]) ? node2006 : node1995;
												assign node1995 = (inp[14]) ? node2001 : node1996;
													assign node1996 = (inp[13]) ? node1998 : 1'b0;
														assign node1998 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2001 = (inp[11]) ? 1'b1 : node2002;
														assign node2002 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2006 = (inp[13]) ? node2008 : 1'b0;
													assign node2008 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2011 = (inp[1]) ? node2013 : 1'b1;
									assign node2013 = (inp[8]) ? 1'b1 : node2014;
										assign node2014 = (inp[14]) ? node2020 : node2015;
											assign node2015 = (inp[11]) ? 1'b0 : node2016;
												assign node2016 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2020 = (inp[2]) ? node2026 : node2021;
												assign node2021 = (inp[11]) ? 1'b1 : node2022;
													assign node2022 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2026 = (inp[13]) ? node2028 : 1'b0;
													assign node2028 = (inp[11]) ? 1'b0 : 1'b1;
							assign node2032 = (inp[10]) ? node2114 : node2033;
								assign node2033 = (inp[8]) ? node2093 : node2034;
									assign node2034 = (inp[1]) ? node2056 : node2035;
										assign node2035 = (inp[0]) ? node2037 : 1'b0;
											assign node2037 = (inp[4]) ? 1'b0 : node2038;
												assign node2038 = (inp[2]) ? node2050 : node2039;
													assign node2039 = (inp[14]) ? node2045 : node2040;
														assign node2040 = (inp[13]) ? node2042 : 1'b1;
															assign node2042 = (inp[11]) ? 1'b1 : 1'b0;
														assign node2045 = (inp[11]) ? 1'b0 : node2046;
															assign node2046 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2050 = (inp[11]) ? 1'b1 : node2051;
														assign node2051 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2056 = (inp[0]) ? node2074 : node2057;
											assign node2057 = (inp[11]) ? node2069 : node2058;
												assign node2058 = (inp[13]) ? node2064 : node2059;
													assign node2059 = (inp[2]) ? 1'b1 : node2060;
														assign node2060 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2064 = (inp[14]) ? node2066 : 1'b0;
														assign node2066 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2069 = (inp[14]) ? node2071 : 1'b1;
													assign node2071 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2074 = (inp[4]) ? node2076 : 1'b0;
												assign node2076 = (inp[13]) ? node2082 : node2077;
													assign node2077 = (inp[14]) ? node2079 : 1'b1;
														assign node2079 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2082 = (inp[11]) ? node2088 : node2083;
														assign node2083 = (inp[14]) ? node2085 : 1'b0;
															assign node2085 = (inp[2]) ? 1'b0 : 1'b1;
														assign node2088 = (inp[2]) ? 1'b1 : node2089;
															assign node2089 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2093 = (inp[4]) ? 1'b0 : node2094;
										assign node2094 = (inp[0]) ? node2096 : 1'b0;
											assign node2096 = (inp[11]) ? node2108 : node2097;
												assign node2097 = (inp[13]) ? node2103 : node2098;
													assign node2098 = (inp[14]) ? node2100 : 1'b1;
														assign node2100 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2103 = (inp[14]) ? node2105 : 1'b0;
														assign node2105 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2108 = (inp[2]) ? 1'b1 : node2109;
													assign node2109 = (inp[14]) ? 1'b0 : 1'b1;
								assign node2114 = (inp[0]) ? node2136 : node2115;
									assign node2115 = (inp[1]) ? node2117 : 1'b1;
										assign node2117 = (inp[8]) ? 1'b1 : node2118;
											assign node2118 = (inp[2]) ? node2130 : node2119;
												assign node2119 = (inp[14]) ? node2125 : node2120;
													assign node2120 = (inp[13]) ? node2122 : 1'b0;
														assign node2122 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2125 = (inp[13]) ? node2127 : 1'b1;
														assign node2127 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2130 = (inp[11]) ? 1'b0 : node2131;
													assign node2131 = (inp[13]) ? 1'b1 : 1'b0;
									assign node2136 = (inp[4]) ? node2174 : node2137;
										assign node2137 = (inp[8]) ? node2157 : node2138;
											assign node2138 = (inp[1]) ? 1'b1 : node2139;
												assign node2139 = (inp[13]) ? node2145 : node2140;
													assign node2140 = (inp[14]) ? node2142 : 1'b0;
														assign node2142 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2145 = (inp[11]) ? node2151 : node2146;
														assign node2146 = (inp[14]) ? node2148 : 1'b1;
															assign node2148 = (inp[2]) ? 1'b1 : 1'b0;
														assign node2151 = (inp[14]) ? node2153 : 1'b0;
															assign node2153 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2157 = (inp[2]) ? node2169 : node2158;
												assign node2158 = (inp[14]) ? node2164 : node2159;
													assign node2159 = (inp[13]) ? node2161 : 1'b0;
														assign node2161 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2164 = (inp[11]) ? 1'b1 : node2165;
														assign node2165 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2169 = (inp[13]) ? node2171 : 1'b0;
													assign node2171 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2174 = (inp[1]) ? node2176 : 1'b1;
											assign node2176 = (inp[8]) ? 1'b1 : node2177;
												assign node2177 = (inp[2]) ? node2189 : node2178;
													assign node2178 = (inp[14]) ? node2184 : node2179;
														assign node2179 = (inp[11]) ? 1'b0 : node2180;
															assign node2180 = (inp[13]) ? 1'b1 : 1'b0;
														assign node2184 = (inp[11]) ? 1'b1 : node2185;
															assign node2185 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2189 = (inp[13]) ? node2191 : 1'b0;
														assign node2191 = (inp[11]) ? 1'b0 : 1'b1;
					assign node2195 = (inp[9]) ? node2277 : node2196;
						assign node2196 = (inp[1]) ? node2218 : node2197;
							assign node2197 = (inp[0]) ? node2199 : 1'b0;
								assign node2199 = (inp[4]) ? 1'b0 : node2200;
									assign node2200 = (inp[2]) ? node2212 : node2201;
										assign node2201 = (inp[14]) ? node2207 : node2202;
											assign node2202 = (inp[11]) ? 1'b1 : node2203;
												assign node2203 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2207 = (inp[13]) ? node2209 : 1'b0;
												assign node2209 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2212 = (inp[13]) ? node2214 : 1'b1;
											assign node2214 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2218 = (inp[8]) ? node2256 : node2219;
								assign node2219 = (inp[0]) ? node2237 : node2220;
									assign node2220 = (inp[2]) ? node2232 : node2221;
										assign node2221 = (inp[14]) ? node2227 : node2222;
											assign node2222 = (inp[11]) ? 1'b1 : node2223;
												assign node2223 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2227 = (inp[13]) ? node2229 : 1'b0;
												assign node2229 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2232 = (inp[13]) ? node2234 : 1'b1;
											assign node2234 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2237 = (inp[4]) ? node2239 : 1'b0;
										assign node2239 = (inp[2]) ? node2251 : node2240;
											assign node2240 = (inp[14]) ? node2246 : node2241;
												assign node2241 = (inp[11]) ? 1'b1 : node2242;
													assign node2242 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2246 = (inp[11]) ? 1'b0 : node2247;
													assign node2247 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2251 = (inp[13]) ? node2253 : 1'b1;
												assign node2253 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2256 = (inp[0]) ? node2258 : 1'b0;
									assign node2258 = (inp[4]) ? 1'b0 : node2259;
										assign node2259 = (inp[13]) ? node2265 : node2260;
											assign node2260 = (inp[2]) ? 1'b1 : node2261;
												assign node2261 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2265 = (inp[11]) ? node2271 : node2266;
												assign node2266 = (inp[14]) ? node2268 : 1'b0;
													assign node2268 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2271 = (inp[2]) ? 1'b1 : node2272;
													assign node2272 = (inp[14]) ? 1'b0 : 1'b1;
						assign node2277 = (inp[10]) ? node2359 : node2278;
							assign node2278 = (inp[1]) ? node2300 : node2279;
								assign node2279 = (inp[4]) ? 1'b1 : node2280;
									assign node2280 = (inp[0]) ? node2282 : 1'b1;
										assign node2282 = (inp[11]) ? node2294 : node2283;
											assign node2283 = (inp[13]) ? node2289 : node2284;
												assign node2284 = (inp[2]) ? 1'b0 : node2285;
													assign node2285 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2289 = (inp[2]) ? 1'b1 : node2290;
													assign node2290 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2294 = (inp[14]) ? node2296 : 1'b0;
												assign node2296 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2300 = (inp[8]) ? node2338 : node2301;
									assign node2301 = (inp[4]) ? node2321 : node2302;
										assign node2302 = (inp[0]) ? 1'b1 : node2303;
											assign node2303 = (inp[14]) ? node2309 : node2304;
												assign node2304 = (inp[11]) ? 1'b0 : node2305;
													assign node2305 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2309 = (inp[2]) ? node2315 : node2310;
													assign node2310 = (inp[13]) ? node2312 : 1'b1;
														assign node2312 = (inp[11]) ? 1'b1 : 1'b0;
													assign node2315 = (inp[13]) ? node2317 : 1'b0;
														assign node2317 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2321 = (inp[14]) ? node2327 : node2322;
											assign node2322 = (inp[11]) ? 1'b0 : node2323;
												assign node2323 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2327 = (inp[2]) ? node2333 : node2328;
												assign node2328 = (inp[11]) ? 1'b1 : node2329;
													assign node2329 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2333 = (inp[11]) ? 1'b0 : node2334;
													assign node2334 = (inp[13]) ? 1'b1 : 1'b0;
									assign node2338 = (inp[0]) ? node2340 : 1'b1;
										assign node2340 = (inp[4]) ? 1'b1 : node2341;
											assign node2341 = (inp[13]) ? node2347 : node2342;
												assign node2342 = (inp[2]) ? 1'b0 : node2343;
													assign node2343 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2347 = (inp[11]) ? node2353 : node2348;
													assign node2348 = (inp[2]) ? 1'b1 : node2349;
														assign node2349 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2353 = (inp[14]) ? node2355 : 1'b0;
														assign node2355 = (inp[2]) ? 1'b0 : 1'b1;
							assign node2359 = (inp[8]) ? node2419 : node2360;
								assign node2360 = (inp[1]) ? node2382 : node2361;
									assign node2361 = (inp[0]) ? node2363 : 1'b0;
										assign node2363 = (inp[4]) ? 1'b0 : node2364;
											assign node2364 = (inp[14]) ? node2370 : node2365;
												assign node2365 = (inp[11]) ? 1'b1 : node2366;
													assign node2366 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2370 = (inp[2]) ? node2376 : node2371;
													assign node2371 = (inp[13]) ? node2373 : 1'b0;
														assign node2373 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2376 = (inp[11]) ? 1'b1 : node2377;
														assign node2377 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2382 = (inp[4]) ? node2402 : node2383;
										assign node2383 = (inp[0]) ? 1'b0 : node2384;
											assign node2384 = (inp[13]) ? node2390 : node2385;
												assign node2385 = (inp[14]) ? node2387 : 1'b1;
													assign node2387 = (inp[2]) ? 1'b1 : 1'b0;
												assign node2390 = (inp[11]) ? node2396 : node2391;
													assign node2391 = (inp[14]) ? node2393 : 1'b0;
														assign node2393 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2396 = (inp[14]) ? node2398 : 1'b1;
														assign node2398 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2402 = (inp[14]) ? node2408 : node2403;
											assign node2403 = (inp[11]) ? 1'b1 : node2404;
												assign node2404 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2408 = (inp[2]) ? node2414 : node2409;
												assign node2409 = (inp[13]) ? node2411 : 1'b0;
													assign node2411 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2414 = (inp[13]) ? node2416 : 1'b1;
													assign node2416 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2419 = (inp[0]) ? node2421 : 1'b0;
									assign node2421 = (inp[4]) ? 1'b0 : node2422;
										assign node2422 = (inp[13]) ? node2428 : node2423;
											assign node2423 = (inp[2]) ? 1'b1 : node2424;
												assign node2424 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2428 = (inp[11]) ? node2434 : node2429;
												assign node2429 = (inp[2]) ? 1'b0 : node2430;
													assign node2430 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2434 = (inp[14]) ? node2436 : 1'b1;
													assign node2436 = (inp[2]) ? 1'b1 : 1'b0;
		assign node2440 = (inp[15]) ? node3256 : node2441;
			assign node2441 = (inp[12]) ? node2523 : node2442;
				assign node2442 = (inp[8]) ? node2502 : node2443;
					assign node2443 = (inp[1]) ? node2465 : node2444;
						assign node2444 = (inp[0]) ? node2446 : 1'b1;
							assign node2446 = (inp[4]) ? 1'b1 : node2447;
								assign node2447 = (inp[14]) ? node2453 : node2448;
									assign node2448 = (inp[13]) ? node2450 : 1'b0;
										assign node2450 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2453 = (inp[2]) ? node2459 : node2454;
										assign node2454 = (inp[13]) ? node2456 : 1'b1;
											assign node2456 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2459 = (inp[11]) ? 1'b0 : node2460;
											assign node2460 = (inp[13]) ? 1'b1 : 1'b0;
						assign node2465 = (inp[0]) ? node2483 : node2466;
							assign node2466 = (inp[2]) ? node2478 : node2467;
								assign node2467 = (inp[14]) ? node2473 : node2468;
									assign node2468 = (inp[13]) ? node2470 : 1'b0;
										assign node2470 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2473 = (inp[13]) ? node2475 : 1'b1;
										assign node2475 = (inp[11]) ? 1'b1 : 1'b0;
								assign node2478 = (inp[13]) ? node2480 : 1'b0;
									assign node2480 = (inp[11]) ? 1'b0 : 1'b1;
							assign node2483 = (inp[4]) ? node2485 : 1'b1;
								assign node2485 = (inp[13]) ? node2491 : node2486;
									assign node2486 = (inp[14]) ? node2488 : 1'b0;
										assign node2488 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2491 = (inp[11]) ? node2497 : node2492;
										assign node2492 = (inp[14]) ? node2494 : 1'b1;
											assign node2494 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2497 = (inp[2]) ? 1'b0 : node2498;
											assign node2498 = (inp[14]) ? 1'b1 : 1'b0;
					assign node2502 = (inp[4]) ? 1'b1 : node2503;
						assign node2503 = (inp[0]) ? node2505 : 1'b1;
							assign node2505 = (inp[14]) ? node2511 : node2506;
								assign node2506 = (inp[13]) ? node2508 : 1'b0;
									assign node2508 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2511 = (inp[2]) ? node2517 : node2512;
									assign node2512 = (inp[13]) ? node2514 : 1'b1;
										assign node2514 = (inp[11]) ? 1'b1 : 1'b0;
									assign node2517 = (inp[11]) ? 1'b0 : node2518;
										assign node2518 = (inp[13]) ? 1'b1 : 1'b0;
				assign node2523 = (inp[9]) ? node2769 : node2524;
					assign node2524 = (inp[7]) ? node2688 : node2525;
						assign node2525 = (inp[3]) ? node2607 : node2526;
							assign node2526 = (inp[1]) ? node2548 : node2527;
								assign node2527 = (inp[0]) ? node2529 : 1'b0;
									assign node2529 = (inp[4]) ? 1'b0 : node2530;
										assign node2530 = (inp[13]) ? node2536 : node2531;
											assign node2531 = (inp[2]) ? 1'b1 : node2532;
												assign node2532 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2536 = (inp[11]) ? node2542 : node2537;
												assign node2537 = (inp[14]) ? node2539 : 1'b0;
													assign node2539 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2542 = (inp[2]) ? 1'b1 : node2543;
													assign node2543 = (inp[14]) ? 1'b0 : 1'b1;
								assign node2548 = (inp[8]) ? node2586 : node2549;
									assign node2549 = (inp[4]) ? node2569 : node2550;
										assign node2550 = (inp[0]) ? 1'b0 : node2551;
											assign node2551 = (inp[13]) ? node2557 : node2552;
												assign node2552 = (inp[2]) ? 1'b1 : node2553;
													assign node2553 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2557 = (inp[11]) ? node2563 : node2558;
													assign node2558 = (inp[14]) ? node2560 : 1'b0;
														assign node2560 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2563 = (inp[2]) ? 1'b1 : node2564;
														assign node2564 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2569 = (inp[13]) ? node2575 : node2570;
											assign node2570 = (inp[14]) ? node2572 : 1'b1;
												assign node2572 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2575 = (inp[11]) ? node2581 : node2576;
												assign node2576 = (inp[14]) ? node2578 : 1'b0;
													assign node2578 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2581 = (inp[2]) ? 1'b1 : node2582;
													assign node2582 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2586 = (inp[4]) ? 1'b0 : node2587;
										assign node2587 = (inp[0]) ? node2589 : 1'b0;
											assign node2589 = (inp[2]) ? node2601 : node2590;
												assign node2590 = (inp[14]) ? node2596 : node2591;
													assign node2591 = (inp[11]) ? 1'b1 : node2592;
														assign node2592 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2596 = (inp[11]) ? 1'b0 : node2597;
														assign node2597 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2601 = (inp[11]) ? 1'b1 : node2602;
													assign node2602 = (inp[13]) ? 1'b0 : 1'b1;
							assign node2607 = (inp[8]) ? node2667 : node2608;
								assign node2608 = (inp[1]) ? node2630 : node2609;
									assign node2609 = (inp[0]) ? node2611 : 1'b1;
										assign node2611 = (inp[4]) ? 1'b1 : node2612;
											assign node2612 = (inp[2]) ? node2624 : node2613;
												assign node2613 = (inp[14]) ? node2619 : node2614;
													assign node2614 = (inp[13]) ? node2616 : 1'b0;
														assign node2616 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2619 = (inp[11]) ? 1'b1 : node2620;
														assign node2620 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2624 = (inp[11]) ? 1'b0 : node2625;
													assign node2625 = (inp[13]) ? 1'b1 : 1'b0;
									assign node2630 = (inp[4]) ? node2650 : node2631;
										assign node2631 = (inp[0]) ? 1'b1 : node2632;
											assign node2632 = (inp[11]) ? node2644 : node2633;
												assign node2633 = (inp[13]) ? node2639 : node2634;
													assign node2634 = (inp[14]) ? node2636 : 1'b0;
														assign node2636 = (inp[2]) ? 1'b0 : 1'b1;
													assign node2639 = (inp[2]) ? 1'b1 : node2640;
														assign node2640 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2644 = (inp[14]) ? node2646 : 1'b0;
													assign node2646 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2650 = (inp[14]) ? node2656 : node2651;
											assign node2651 = (inp[11]) ? 1'b0 : node2652;
												assign node2652 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2656 = (inp[2]) ? node2662 : node2657;
												assign node2657 = (inp[13]) ? node2659 : 1'b1;
													assign node2659 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2662 = (inp[11]) ? 1'b0 : node2663;
													assign node2663 = (inp[13]) ? 1'b1 : 1'b0;
								assign node2667 = (inp[0]) ? node2669 : 1'b1;
									assign node2669 = (inp[4]) ? 1'b1 : node2670;
										assign node2670 = (inp[14]) ? node2676 : node2671;
											assign node2671 = (inp[11]) ? 1'b0 : node2672;
												assign node2672 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2676 = (inp[2]) ? node2682 : node2677;
												assign node2677 = (inp[13]) ? node2679 : 1'b1;
													assign node2679 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2682 = (inp[11]) ? 1'b0 : node2683;
													assign node2683 = (inp[13]) ? 1'b1 : 1'b0;
						assign node2688 = (inp[8]) ? node2748 : node2689;
							assign node2689 = (inp[1]) ? node2711 : node2690;
								assign node2690 = (inp[4]) ? 1'b0 : node2691;
									assign node2691 = (inp[0]) ? node2693 : 1'b0;
										assign node2693 = (inp[14]) ? node2699 : node2694;
											assign node2694 = (inp[11]) ? 1'b1 : node2695;
												assign node2695 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2699 = (inp[2]) ? node2705 : node2700;
												assign node2700 = (inp[11]) ? 1'b0 : node2701;
													assign node2701 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2705 = (inp[11]) ? 1'b1 : node2706;
													assign node2706 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2711 = (inp[0]) ? node2729 : node2712;
									assign node2712 = (inp[13]) ? node2718 : node2713;
										assign node2713 = (inp[14]) ? node2715 : 1'b1;
											assign node2715 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2718 = (inp[11]) ? node2724 : node2719;
											assign node2719 = (inp[14]) ? node2721 : 1'b0;
												assign node2721 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2724 = (inp[14]) ? node2726 : 1'b1;
												assign node2726 = (inp[2]) ? 1'b1 : 1'b0;
									assign node2729 = (inp[4]) ? node2731 : 1'b0;
										assign node2731 = (inp[14]) ? node2737 : node2732;
											assign node2732 = (inp[11]) ? 1'b1 : node2733;
												assign node2733 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2737 = (inp[2]) ? node2743 : node2738;
												assign node2738 = (inp[13]) ? node2740 : 1'b0;
													assign node2740 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2743 = (inp[13]) ? node2745 : 1'b1;
													assign node2745 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2748 = (inp[0]) ? node2750 : 1'b0;
								assign node2750 = (inp[4]) ? 1'b0 : node2751;
									assign node2751 = (inp[13]) ? node2757 : node2752;
										assign node2752 = (inp[2]) ? 1'b1 : node2753;
											assign node2753 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2757 = (inp[11]) ? node2763 : node2758;
											assign node2758 = (inp[14]) ? node2760 : 1'b0;
												assign node2760 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2763 = (inp[14]) ? node2765 : 1'b1;
												assign node2765 = (inp[2]) ? 1'b1 : 1'b0;
					assign node2769 = (inp[10]) ? node3015 : node2770;
						assign node2770 = (inp[7]) ? node2934 : node2771;
							assign node2771 = (inp[3]) ? node2853 : node2772;
								assign node2772 = (inp[4]) ? node2832 : node2773;
									assign node2773 = (inp[0]) ? node2795 : node2774;
										assign node2774 = (inp[8]) ? 1'b1 : node2775;
											assign node2775 = (inp[1]) ? node2777 : 1'b1;
												assign node2777 = (inp[14]) ? node2783 : node2778;
													assign node2778 = (inp[13]) ? node2780 : 1'b0;
														assign node2780 = (inp[11]) ? 1'b0 : 1'b1;
													assign node2783 = (inp[2]) ? node2789 : node2784;
														assign node2784 = (inp[11]) ? 1'b1 : node2785;
															assign node2785 = (inp[13]) ? 1'b0 : 1'b1;
														assign node2789 = (inp[13]) ? node2791 : 1'b0;
															assign node2791 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2795 = (inp[1]) ? node2813 : node2796;
											assign node2796 = (inp[13]) ? node2802 : node2797;
												assign node2797 = (inp[14]) ? node2799 : 1'b0;
													assign node2799 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2802 = (inp[11]) ? node2808 : node2803;
													assign node2803 = (inp[14]) ? node2805 : 1'b1;
														assign node2805 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2808 = (inp[14]) ? node2810 : 1'b0;
														assign node2810 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2813 = (inp[8]) ? node2815 : 1'b1;
												assign node2815 = (inp[14]) ? node2821 : node2816;
													assign node2816 = (inp[11]) ? 1'b0 : node2817;
														assign node2817 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2821 = (inp[2]) ? node2827 : node2822;
														assign node2822 = (inp[13]) ? node2824 : 1'b1;
															assign node2824 = (inp[11]) ? 1'b1 : 1'b0;
														assign node2827 = (inp[13]) ? node2829 : 1'b0;
															assign node2829 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2832 = (inp[1]) ? node2834 : 1'b1;
										assign node2834 = (inp[8]) ? 1'b1 : node2835;
											assign node2835 = (inp[14]) ? node2841 : node2836;
												assign node2836 = (inp[13]) ? node2838 : 1'b0;
													assign node2838 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2841 = (inp[2]) ? node2847 : node2842;
													assign node2842 = (inp[11]) ? 1'b1 : node2843;
														assign node2843 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2847 = (inp[13]) ? node2849 : 1'b0;
														assign node2849 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2853 = (inp[8]) ? node2913 : node2854;
									assign node2854 = (inp[1]) ? node2876 : node2855;
										assign node2855 = (inp[0]) ? node2857 : 1'b0;
											assign node2857 = (inp[4]) ? 1'b0 : node2858;
												assign node2858 = (inp[13]) ? node2864 : node2859;
													assign node2859 = (inp[2]) ? 1'b1 : node2860;
														assign node2860 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2864 = (inp[11]) ? node2870 : node2865;
														assign node2865 = (inp[2]) ? 1'b0 : node2866;
															assign node2866 = (inp[14]) ? 1'b1 : 1'b0;
														assign node2870 = (inp[14]) ? node2872 : 1'b1;
															assign node2872 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2876 = (inp[0]) ? node2894 : node2877;
											assign node2877 = (inp[11]) ? node2889 : node2878;
												assign node2878 = (inp[13]) ? node2884 : node2879;
													assign node2879 = (inp[2]) ? 1'b1 : node2880;
														assign node2880 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2884 = (inp[2]) ? 1'b0 : node2885;
														assign node2885 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2889 = (inp[2]) ? 1'b1 : node2890;
													assign node2890 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2894 = (inp[4]) ? node2896 : 1'b0;
												assign node2896 = (inp[13]) ? node2902 : node2897;
													assign node2897 = (inp[14]) ? node2899 : 1'b1;
														assign node2899 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2902 = (inp[11]) ? node2908 : node2903;
														assign node2903 = (inp[2]) ? 1'b0 : node2904;
															assign node2904 = (inp[14]) ? 1'b1 : 1'b0;
														assign node2908 = (inp[2]) ? 1'b1 : node2909;
															assign node2909 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2913 = (inp[4]) ? 1'b0 : node2914;
										assign node2914 = (inp[0]) ? node2916 : 1'b0;
											assign node2916 = (inp[2]) ? node2928 : node2917;
												assign node2917 = (inp[14]) ? node2923 : node2918;
													assign node2918 = (inp[11]) ? 1'b1 : node2919;
														assign node2919 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2923 = (inp[13]) ? node2925 : 1'b0;
														assign node2925 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2928 = (inp[13]) ? node2930 : 1'b1;
													assign node2930 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2934 = (inp[0]) ? node2956 : node2935;
								assign node2935 = (inp[1]) ? node2937 : 1'b1;
									assign node2937 = (inp[8]) ? 1'b1 : node2938;
										assign node2938 = (inp[11]) ? node2950 : node2939;
											assign node2939 = (inp[13]) ? node2945 : node2940;
												assign node2940 = (inp[2]) ? 1'b0 : node2941;
													assign node2941 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2945 = (inp[14]) ? node2947 : 1'b1;
													assign node2947 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2950 = (inp[14]) ? node2952 : 1'b0;
												assign node2952 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2956 = (inp[4]) ? node2994 : node2957;
									assign node2957 = (inp[8]) ? node2977 : node2958;
										assign node2958 = (inp[1]) ? 1'b1 : node2959;
											assign node2959 = (inp[2]) ? node2971 : node2960;
												assign node2960 = (inp[14]) ? node2966 : node2961;
													assign node2961 = (inp[11]) ? 1'b0 : node2962;
														assign node2962 = (inp[13]) ? 1'b1 : 1'b0;
													assign node2966 = (inp[13]) ? node2968 : 1'b1;
														assign node2968 = (inp[11]) ? 1'b1 : 1'b0;
												assign node2971 = (inp[11]) ? 1'b0 : node2972;
													assign node2972 = (inp[13]) ? 1'b1 : 1'b0;
										assign node2977 = (inp[2]) ? node2989 : node2978;
											assign node2978 = (inp[14]) ? node2984 : node2979;
												assign node2979 = (inp[13]) ? node2981 : 1'b0;
													assign node2981 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2984 = (inp[13]) ? node2986 : 1'b1;
													assign node2986 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2989 = (inp[13]) ? node2991 : 1'b0;
												assign node2991 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2994 = (inp[8]) ? 1'b1 : node2995;
										assign node2995 = (inp[1]) ? node2997 : 1'b1;
											assign node2997 = (inp[14]) ? node3003 : node2998;
												assign node2998 = (inp[13]) ? node3000 : 1'b0;
													assign node3000 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3003 = (inp[2]) ? node3009 : node3004;
													assign node3004 = (inp[11]) ? 1'b1 : node3005;
														assign node3005 = (inp[13]) ? 1'b0 : 1'b1;
													assign node3009 = (inp[11]) ? 1'b0 : node3010;
														assign node3010 = (inp[13]) ? 1'b1 : 1'b0;
						assign node3015 = (inp[7]) ? node3175 : node3016;
							assign node3016 = (inp[3]) ? node3098 : node3017;
								assign node3017 = (inp[0]) ? node3039 : node3018;
									assign node3018 = (inp[1]) ? node3020 : 1'b0;
										assign node3020 = (inp[8]) ? 1'b0 : node3021;
											assign node3021 = (inp[14]) ? node3027 : node3022;
												assign node3022 = (inp[11]) ? 1'b1 : node3023;
													assign node3023 = (inp[13]) ? 1'b0 : 1'b1;
												assign node3027 = (inp[2]) ? node3033 : node3028;
													assign node3028 = (inp[11]) ? 1'b0 : node3029;
														assign node3029 = (inp[13]) ? 1'b1 : 1'b0;
													assign node3033 = (inp[11]) ? 1'b1 : node3034;
														assign node3034 = (inp[13]) ? 1'b0 : 1'b1;
									assign node3039 = (inp[4]) ? node3077 : node3040;
										assign node3040 = (inp[1]) ? node3058 : node3041;
											assign node3041 = (inp[13]) ? node3047 : node3042;
												assign node3042 = (inp[14]) ? node3044 : 1'b1;
													assign node3044 = (inp[2]) ? 1'b1 : 1'b0;
												assign node3047 = (inp[11]) ? node3053 : node3048;
													assign node3048 = (inp[2]) ? 1'b0 : node3049;
														assign node3049 = (inp[14]) ? 1'b1 : 1'b0;
													assign node3053 = (inp[2]) ? 1'b1 : node3054;
														assign node3054 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3058 = (inp[8]) ? node3060 : 1'b0;
												assign node3060 = (inp[11]) ? node3072 : node3061;
													assign node3061 = (inp[13]) ? node3067 : node3062;
														assign node3062 = (inp[2]) ? 1'b1 : node3063;
															assign node3063 = (inp[14]) ? 1'b0 : 1'b1;
														assign node3067 = (inp[14]) ? node3069 : 1'b0;
															assign node3069 = (inp[2]) ? 1'b0 : 1'b1;
													assign node3072 = (inp[2]) ? 1'b1 : node3073;
														assign node3073 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3077 = (inp[8]) ? 1'b0 : node3078;
											assign node3078 = (inp[1]) ? node3080 : 1'b0;
												assign node3080 = (inp[2]) ? node3092 : node3081;
													assign node3081 = (inp[14]) ? node3087 : node3082;
														assign node3082 = (inp[13]) ? node3084 : 1'b1;
															assign node3084 = (inp[11]) ? 1'b1 : 1'b0;
														assign node3087 = (inp[13]) ? node3089 : 1'b0;
															assign node3089 = (inp[11]) ? 1'b0 : 1'b1;
													assign node3092 = (inp[13]) ? node3094 : 1'b1;
														assign node3094 = (inp[11]) ? 1'b1 : 1'b0;
								assign node3098 = (inp[8]) ? node3154 : node3099;
									assign node3099 = (inp[1]) ? node3121 : node3100;
										assign node3100 = (inp[0]) ? node3102 : 1'b1;
											assign node3102 = (inp[4]) ? 1'b1 : node3103;
												assign node3103 = (inp[13]) ? node3109 : node3104;
													assign node3104 = (inp[2]) ? 1'b0 : node3105;
														assign node3105 = (inp[14]) ? 1'b1 : 1'b0;
													assign node3109 = (inp[11]) ? node3115 : node3110;
														assign node3110 = (inp[14]) ? node3112 : 1'b1;
															assign node3112 = (inp[2]) ? 1'b1 : 1'b0;
														assign node3115 = (inp[14]) ? node3117 : 1'b0;
															assign node3117 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3121 = (inp[4]) ? node3137 : node3122;
											assign node3122 = (inp[0]) ? 1'b1 : node3123;
												assign node3123 = (inp[11]) ? node3131 : node3124;
													assign node3124 = (inp[13]) ? 1'b1 : node3125;
														assign node3125 = (inp[2]) ? 1'b0 : node3126;
															assign node3126 = (inp[14]) ? 1'b1 : 1'b0;
													assign node3131 = (inp[14]) ? node3133 : 1'b0;
														assign node3133 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3137 = (inp[13]) ? node3143 : node3138;
												assign node3138 = (inp[14]) ? node3140 : 1'b0;
													assign node3140 = (inp[2]) ? 1'b0 : 1'b1;
												assign node3143 = (inp[11]) ? node3149 : node3144;
													assign node3144 = (inp[14]) ? node3146 : 1'b1;
														assign node3146 = (inp[2]) ? 1'b1 : 1'b0;
													assign node3149 = (inp[14]) ? node3151 : 1'b0;
														assign node3151 = (inp[2]) ? 1'b0 : 1'b1;
									assign node3154 = (inp[0]) ? node3156 : 1'b1;
										assign node3156 = (inp[4]) ? 1'b1 : node3157;
											assign node3157 = (inp[13]) ? node3163 : node3158;
												assign node3158 = (inp[14]) ? node3160 : 1'b0;
													assign node3160 = (inp[2]) ? 1'b0 : 1'b1;
												assign node3163 = (inp[11]) ? node3169 : node3164;
													assign node3164 = (inp[2]) ? 1'b1 : node3165;
														assign node3165 = (inp[14]) ? 1'b0 : 1'b1;
													assign node3169 = (inp[14]) ? node3171 : 1'b0;
														assign node3171 = (inp[2]) ? 1'b0 : 1'b1;
							assign node3175 = (inp[8]) ? node3235 : node3176;
								assign node3176 = (inp[1]) ? node3198 : node3177;
									assign node3177 = (inp[0]) ? node3179 : 1'b0;
										assign node3179 = (inp[4]) ? 1'b0 : node3180;
											assign node3180 = (inp[2]) ? node3192 : node3181;
												assign node3181 = (inp[14]) ? node3187 : node3182;
													assign node3182 = (inp[11]) ? 1'b1 : node3183;
														assign node3183 = (inp[13]) ? 1'b0 : 1'b1;
													assign node3187 = (inp[13]) ? node3189 : 1'b0;
														assign node3189 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3192 = (inp[13]) ? node3194 : 1'b1;
													assign node3194 = (inp[11]) ? 1'b1 : 1'b0;
									assign node3198 = (inp[0]) ? node3216 : node3199;
										assign node3199 = (inp[14]) ? node3205 : node3200;
											assign node3200 = (inp[13]) ? node3202 : 1'b1;
												assign node3202 = (inp[11]) ? 1'b1 : 1'b0;
											assign node3205 = (inp[2]) ? node3211 : node3206;
												assign node3206 = (inp[13]) ? node3208 : 1'b0;
													assign node3208 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3211 = (inp[11]) ? 1'b1 : node3212;
													assign node3212 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3216 = (inp[4]) ? node3218 : 1'b0;
											assign node3218 = (inp[2]) ? node3230 : node3219;
												assign node3219 = (inp[14]) ? node3225 : node3220;
													assign node3220 = (inp[13]) ? node3222 : 1'b1;
														assign node3222 = (inp[11]) ? 1'b1 : 1'b0;
													assign node3225 = (inp[11]) ? 1'b0 : node3226;
														assign node3226 = (inp[13]) ? 1'b1 : 1'b0;
												assign node3230 = (inp[13]) ? node3232 : 1'b1;
													assign node3232 = (inp[11]) ? 1'b1 : 1'b0;
								assign node3235 = (inp[0]) ? node3237 : 1'b0;
									assign node3237 = (inp[4]) ? 1'b0 : node3238;
										assign node3238 = (inp[2]) ? node3250 : node3239;
											assign node3239 = (inp[14]) ? node3245 : node3240;
												assign node3240 = (inp[11]) ? 1'b1 : node3241;
													assign node3241 = (inp[13]) ? 1'b0 : 1'b1;
												assign node3245 = (inp[11]) ? 1'b0 : node3246;
													assign node3246 = (inp[13]) ? 1'b1 : 1'b0;
											assign node3250 = (inp[13]) ? node3252 : 1'b1;
												assign node3252 = (inp[11]) ? 1'b1 : 1'b0;
			assign node3256 = (inp[8]) ? node3316 : node3257;
				assign node3257 = (inp[1]) ? node3279 : node3258;
					assign node3258 = (inp[0]) ? node3260 : 1'b1;
						assign node3260 = (inp[4]) ? 1'b1 : node3261;
							assign node3261 = (inp[14]) ? node3267 : node3262;
								assign node3262 = (inp[13]) ? node3264 : 1'b0;
									assign node3264 = (inp[11]) ? 1'b0 : 1'b1;
								assign node3267 = (inp[2]) ? node3273 : node3268;
									assign node3268 = (inp[13]) ? node3270 : 1'b1;
										assign node3270 = (inp[11]) ? 1'b1 : 1'b0;
									assign node3273 = (inp[11]) ? 1'b0 : node3274;
										assign node3274 = (inp[13]) ? 1'b1 : 1'b0;
					assign node3279 = (inp[0]) ? node3297 : node3280;
						assign node3280 = (inp[13]) ? node3286 : node3281;
							assign node3281 = (inp[14]) ? node3283 : 1'b0;
								assign node3283 = (inp[2]) ? 1'b0 : 1'b1;
							assign node3286 = (inp[11]) ? node3292 : node3287;
								assign node3287 = (inp[2]) ? 1'b1 : node3288;
									assign node3288 = (inp[14]) ? 1'b0 : 1'b1;
								assign node3292 = (inp[14]) ? node3294 : 1'b0;
									assign node3294 = (inp[2]) ? 1'b0 : 1'b1;
						assign node3297 = (inp[4]) ? node3299 : 1'b1;
							assign node3299 = (inp[14]) ? node3305 : node3300;
								assign node3300 = (inp[11]) ? 1'b0 : node3301;
									assign node3301 = (inp[13]) ? 1'b1 : 1'b0;
								assign node3305 = (inp[2]) ? node3311 : node3306;
									assign node3306 = (inp[13]) ? node3308 : 1'b1;
										assign node3308 = (inp[11]) ? 1'b1 : 1'b0;
									assign node3311 = (inp[11]) ? 1'b0 : node3312;
										assign node3312 = (inp[13]) ? 1'b1 : 1'b0;
				assign node3316 = (inp[4]) ? 1'b1 : node3317;
					assign node3317 = (inp[0]) ? node3319 : 1'b1;
						assign node3319 = (inp[11]) ? node3331 : node3320;
							assign node3320 = (inp[13]) ? node3326 : node3321;
								assign node3321 = (inp[14]) ? node3323 : 1'b0;
									assign node3323 = (inp[2]) ? 1'b0 : 1'b1;
								assign node3326 = (inp[2]) ? 1'b1 : node3327;
									assign node3327 = (inp[14]) ? 1'b0 : 1'b1;
							assign node3331 = (inp[2]) ? 1'b0 : node3332;
								assign node3332 = (inp[14]) ? 1'b1 : 1'b0;

endmodule