module dtc_split25_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;

	assign outp = (inp[6]) ? node174 : node1;
		assign node1 = (inp[9]) ? node153 : node2;
			assign node2 = (inp[7]) ? node38 : node3;
				assign node3 = (inp[0]) ? 3'b000 : node4;
					assign node4 = (inp[10]) ? node30 : node5;
						assign node5 = (inp[1]) ? node21 : node6;
							assign node6 = (inp[11]) ? node14 : node7;
								assign node7 = (inp[3]) ? 3'b110 : node8;
									assign node8 = (inp[8]) ? node10 : 3'b010;
										assign node10 = (inp[4]) ? 3'b110 : 3'b010;
								assign node14 = (inp[8]) ? 3'b010 : node15;
									assign node15 = (inp[5]) ? node17 : 3'b000;
										assign node17 = (inp[3]) ? 3'b100 : 3'b110;
							assign node21 = (inp[8]) ? node23 : 3'b000;
								assign node23 = (inp[11]) ? 3'b100 : node24;
									assign node24 = (inp[2]) ? node26 : 3'b010;
										assign node26 = (inp[3]) ? 3'b100 : 3'b010;
						assign node30 = (inp[1]) ? 3'b000 : node31;
							assign node31 = (inp[11]) ? 3'b000 : node32;
								assign node32 = (inp[8]) ? 3'b100 : 3'b000;
				assign node38 = (inp[0]) ? node102 : node39;
					assign node39 = (inp[10]) ? node65 : node40;
						assign node40 = (inp[1]) ? node54 : node41;
							assign node41 = (inp[8]) ? node47 : node42;
								assign node42 = (inp[11]) ? node44 : 3'b001;
									assign node44 = (inp[4]) ? 3'b010 : 3'b110;
								assign node47 = (inp[11]) ? node49 : 3'b101;
									assign node49 = (inp[2]) ? 3'b001 : node50;
										assign node50 = (inp[3]) ? 3'b001 : 3'b101;
							assign node54 = (inp[11]) ? node62 : node55;
								assign node55 = (inp[8]) ? node57 : 3'b110;
									assign node57 = (inp[3]) ? node59 : 3'b001;
										assign node59 = (inp[2]) ? 3'b110 : 3'b001;
								assign node62 = (inp[8]) ? 3'b110 : 3'b010;
						assign node65 = (inp[1]) ? node87 : node66;
							assign node66 = (inp[5]) ? node78 : node67;
								assign node67 = (inp[2]) ? node73 : node68;
									assign node68 = (inp[8]) ? 3'b110 : node69;
										assign node69 = (inp[3]) ? 3'b010 : 3'b110;
									assign node73 = (inp[8]) ? node75 : 3'b100;
										assign node75 = (inp[4]) ? 3'b010 : 3'b110;
								assign node78 = (inp[11]) ? 3'b010 : node79;
									assign node79 = (inp[8]) ? 3'b110 : node80;
										assign node80 = (inp[4]) ? node82 : 3'b010;
											assign node82 = (inp[3]) ? 3'b100 : 3'b010;
							assign node87 = (inp[11]) ? node95 : node88;
								assign node88 = (inp[8]) ? node90 : 3'b100;
									assign node90 = (inp[3]) ? node92 : 3'b010;
										assign node92 = (inp[2]) ? 3'b100 : 3'b010;
								assign node95 = (inp[3]) ? 3'b000 : node96;
									assign node96 = (inp[8]) ? 3'b100 : node97;
										assign node97 = (inp[4]) ? 3'b000 : 3'b100;
					assign node102 = (inp[10]) ? node146 : node103;
						assign node103 = (inp[11]) ? node135 : node104;
							assign node104 = (inp[2]) ? node126 : node105;
								assign node105 = (inp[5]) ? node117 : node106;
									assign node106 = (inp[3]) ? node112 : node107;
										assign node107 = (inp[1]) ? 3'b010 : node108;
											assign node108 = (inp[8]) ? 3'b110 : 3'b010;
										assign node112 = (inp[8]) ? 3'b010 : node113;
											assign node113 = (inp[1]) ? 3'b000 : 3'b010;
									assign node117 = (inp[1]) ? node121 : node118;
										assign node118 = (inp[8]) ? 3'b110 : 3'b010;
										assign node121 = (inp[8]) ? node123 : 3'b100;
											assign node123 = (inp[4]) ? 3'b100 : 3'b010;
								assign node126 = (inp[5]) ? node128 : 3'b100;
									assign node128 = (inp[8]) ? node132 : node129;
										assign node129 = (inp[1]) ? 3'b000 : 3'b100;
										assign node132 = (inp[4]) ? 3'b010 : 3'b110;
							assign node135 = (inp[1]) ? node141 : node136;
								assign node136 = (inp[2]) ? 3'b100 : node137;
									assign node137 = (inp[8]) ? 3'b010 : 3'b100;
								assign node141 = (inp[8]) ? node143 : 3'b000;
									assign node143 = (inp[2]) ? 3'b000 : 3'b100;
						assign node146 = (inp[8]) ? node148 : 3'b000;
							assign node148 = (inp[2]) ? 3'b000 : node149;
								assign node149 = (inp[5]) ? 3'b100 : 3'b000;
			assign node153 = (inp[1]) ? 3'b000 : node154;
				assign node154 = (inp[0]) ? 3'b000 : node155;
					assign node155 = (inp[7]) ? node157 : 3'b000;
						assign node157 = (inp[3]) ? node167 : node158;
							assign node158 = (inp[10]) ? 3'b000 : node159;
								assign node159 = (inp[8]) ? 3'b100 : node160;
									assign node160 = (inp[5]) ? node162 : 3'b000;
										assign node162 = (inp[4]) ? 3'b100 : 3'b000;
							assign node167 = (inp[8]) ? node169 : 3'b000;
								assign node169 = (inp[11]) ? 3'b000 : 3'b010;
		assign node174 = (inp[9]) ? node404 : node175;
			assign node175 = (inp[0]) ? node269 : node176;
				assign node176 = (inp[1]) ? node208 : node177;
					assign node177 = (inp[10]) ? node187 : node178;
						assign node178 = (inp[11]) ? node180 : 3'b111;
							assign node180 = (inp[7]) ? 3'b111 : node181;
								assign node181 = (inp[8]) ? node183 : 3'b101;
									assign node183 = (inp[2]) ? 3'b011 : 3'b111;
						assign node187 = (inp[7]) ? node195 : node188;
							assign node188 = (inp[8]) ? node192 : node189;
								assign node189 = (inp[2]) ? 3'b110 : 3'b101;
								assign node192 = (inp[5]) ? 3'b001 : 3'b101;
							assign node195 = (inp[8]) ? 3'b111 : node196;
								assign node196 = (inp[11]) ? node204 : node197;
									assign node197 = (inp[2]) ? 3'b011 : node198;
										assign node198 = (inp[4]) ? node200 : 3'b111;
											assign node200 = (inp[5]) ? 3'b011 : 3'b111;
									assign node204 = (inp[2]) ? 3'b101 : 3'b011;
					assign node208 = (inp[10]) ? node244 : node209;
						assign node209 = (inp[7]) ? node235 : node210;
							assign node210 = (inp[11]) ? node228 : node211;
								assign node211 = (inp[8]) ? node219 : node212;
									assign node212 = (inp[3]) ? node216 : node213;
										assign node213 = (inp[2]) ? 3'b101 : 3'b011;
										assign node216 = (inp[2]) ? 3'b001 : 3'b101;
									assign node219 = (inp[4]) ? node223 : node220;
										assign node220 = (inp[2]) ? 3'b011 : 3'b111;
										assign node223 = (inp[2]) ? node225 : 3'b011;
											assign node225 = (inp[3]) ? 3'b101 : 3'b011;
								assign node228 = (inp[8]) ? 3'b101 : node229;
									assign node229 = (inp[3]) ? 3'b001 : node230;
										assign node230 = (inp[4]) ? 3'b001 : 3'b101;
							assign node235 = (inp[8]) ? 3'b111 : node236;
								assign node236 = (inp[11]) ? 3'b011 : node237;
									assign node237 = (inp[5]) ? node239 : 3'b111;
										assign node239 = (inp[4]) ? 3'b011 : 3'b111;
						assign node244 = (inp[7]) ? node260 : node245;
							assign node245 = (inp[11]) ? node255 : node246;
								assign node246 = (inp[4]) ? node248 : 3'b001;
									assign node248 = (inp[5]) ? node252 : node249;
										assign node249 = (inp[3]) ? 3'b010 : 3'b110;
										assign node252 = (inp[3]) ? 3'b110 : 3'b001;
								assign node255 = (inp[5]) ? node257 : 3'b110;
									assign node257 = (inp[8]) ? 3'b110 : 3'b010;
							assign node260 = (inp[11]) ? node266 : node261;
								assign node261 = (inp[8]) ? node263 : 3'b101;
									assign node263 = (inp[2]) ? 3'b011 : 3'b111;
								assign node266 = (inp[8]) ? 3'b101 : 3'b001;
				assign node269 = (inp[10]) ? node355 : node270;
					assign node270 = (inp[7]) ? node316 : node271;
						assign node271 = (inp[1]) ? node293 : node272;
							assign node272 = (inp[8]) ? node284 : node273;
								assign node273 = (inp[11]) ? node281 : node274;
									assign node274 = (inp[2]) ? node276 : 3'b001;
										assign node276 = (inp[4]) ? 3'b110 : node277;
											assign node277 = (inp[3]) ? 3'b110 : 3'b001;
									assign node281 = (inp[2]) ? 3'b010 : 3'b110;
								assign node284 = (inp[11]) ? node288 : node285;
									assign node285 = (inp[5]) ? 3'b001 : 3'b101;
									assign node288 = (inp[5]) ? node290 : 3'b001;
										assign node290 = (inp[2]) ? 3'b110 : 3'b001;
							assign node293 = (inp[8]) ? node305 : node294;
								assign node294 = (inp[11]) ? node298 : node295;
									assign node295 = (inp[2]) ? 3'b010 : 3'b110;
									assign node298 = (inp[2]) ? 3'b100 : node299;
										assign node299 = (inp[4]) ? node301 : 3'b010;
											assign node301 = (inp[3]) ? 3'b100 : 3'b010;
								assign node305 = (inp[11]) ? node311 : node306;
									assign node306 = (inp[5]) ? node308 : 3'b001;
										assign node308 = (inp[2]) ? 3'b110 : 3'b001;
									assign node311 = (inp[2]) ? node313 : 3'b110;
										assign node313 = (inp[4]) ? 3'b010 : 3'b110;
						assign node316 = (inp[1]) ? node328 : node317;
							assign node317 = (inp[11]) ? node325 : node318;
								assign node318 = (inp[8]) ? 3'b111 : node319;
									assign node319 = (inp[3]) ? node321 : 3'b011;
										assign node321 = (inp[2]) ? 3'b101 : 3'b011;
								assign node325 = (inp[8]) ? 3'b011 : 3'b101;
							assign node328 = (inp[4]) ? node336 : node329;
								assign node329 = (inp[8]) ? node333 : node330;
									assign node330 = (inp[3]) ? 3'b001 : 3'b101;
									assign node333 = (inp[11]) ? 3'b001 : 3'b011;
								assign node336 = (inp[5]) ? node342 : node337;
									assign node337 = (inp[11]) ? node339 : 3'b101;
										assign node339 = (inp[8]) ? 3'b101 : 3'b001;
									assign node342 = (inp[3]) ? 3'b110 : node343;
										assign node343 = (inp[8]) ? node347 : node344;
											assign node344 = (inp[2]) ? 3'b110 : 3'b001;
											assign node347 = (inp[2]) ? node351 : node348;
												assign node348 = (inp[11]) ? 3'b101 : 3'b011;
												assign node351 = (inp[11]) ? 3'b001 : 3'b101;
					assign node355 = (inp[7]) ? node379 : node356;
						assign node356 = (inp[11]) ? node366 : node357;
							assign node357 = (inp[8]) ? node361 : node358;
								assign node358 = (inp[2]) ? 3'b000 : 3'b010;
								assign node361 = (inp[1]) ? 3'b010 : node362;
									assign node362 = (inp[2]) ? 3'b010 : 3'b110;
							assign node366 = (inp[8]) ? node374 : node367;
								assign node367 = (inp[1]) ? 3'b000 : node368;
									assign node368 = (inp[2]) ? node370 : 3'b100;
										assign node370 = (inp[3]) ? 3'b000 : 3'b100;
								assign node374 = (inp[5]) ? node376 : 3'b100;
									assign node376 = (inp[1]) ? 3'b000 : 3'b100;
						assign node379 = (inp[11]) ? node393 : node380;
							assign node380 = (inp[8]) ? node390 : node381;
								assign node381 = (inp[1]) ? node387 : node382;
									assign node382 = (inp[3]) ? node384 : 3'b001;
										assign node384 = (inp[2]) ? 3'b110 : 3'b001;
									assign node387 = (inp[4]) ? 3'b010 : 3'b110;
								assign node390 = (inp[2]) ? 3'b101 : 3'b001;
							assign node393 = (inp[1]) ? node397 : node394;
								assign node394 = (inp[8]) ? 3'b101 : 3'b110;
								assign node397 = (inp[4]) ? node399 : 3'b010;
									assign node399 = (inp[3]) ? 3'b100 : node400;
										assign node400 = (inp[5]) ? 3'b110 : 3'b010;
			assign node404 = (inp[0]) ? node532 : node405;
				assign node405 = (inp[7]) ? node463 : node406;
					assign node406 = (inp[10]) ? node444 : node407;
						assign node407 = (inp[11]) ? node429 : node408;
							assign node408 = (inp[8]) ? node418 : node409;
								assign node409 = (inp[1]) ? node411 : 3'b110;
									assign node411 = (inp[4]) ? node415 : node412;
										assign node412 = (inp[3]) ? 3'b100 : 3'b010;
										assign node415 = (inp[3]) ? 3'b000 : 3'b100;
								assign node418 = (inp[4]) ? node422 : node419;
									assign node419 = (inp[1]) ? 3'b010 : 3'b001;
									assign node422 = (inp[1]) ? node424 : 3'b110;
										assign node424 = (inp[3]) ? 3'b010 : node425;
											assign node425 = (inp[2]) ? 3'b010 : 3'b110;
							assign node429 = (inp[1]) ? node439 : node430;
								assign node430 = (inp[2]) ? 3'b100 : node431;
									assign node431 = (inp[5]) ? node435 : node432;
										assign node432 = (inp[4]) ? 3'b100 : 3'b110;
										assign node435 = (inp[3]) ? 3'b010 : 3'b110;
								assign node439 = (inp[8]) ? 3'b100 : node440;
									assign node440 = (inp[4]) ? 3'b000 : 3'b100;
						assign node444 = (inp[1]) ? node456 : node445;
							assign node445 = (inp[2]) ? node451 : node446;
								assign node446 = (inp[8]) ? node448 : 3'b100;
									assign node448 = (inp[11]) ? 3'b100 : 3'b010;
								assign node451 = (inp[11]) ? 3'b000 : node452;
									assign node452 = (inp[3]) ? 3'b100 : 3'b000;
							assign node456 = (inp[2]) ? 3'b000 : node457;
								assign node457 = (inp[3]) ? 3'b000 : node458;
									assign node458 = (inp[8]) ? 3'b100 : 3'b000;
					assign node463 = (inp[10]) ? node497 : node464;
						assign node464 = (inp[8]) ? node478 : node465;
							assign node465 = (inp[3]) ? node473 : node466;
								assign node466 = (inp[2]) ? 3'b110 : node467;
									assign node467 = (inp[4]) ? node469 : 3'b001;
										assign node469 = (inp[1]) ? 3'b110 : 3'b001;
								assign node473 = (inp[11]) ? node475 : 3'b110;
									assign node475 = (inp[5]) ? 3'b010 : 3'b110;
							assign node478 = (inp[4]) ? node486 : node479;
								assign node479 = (inp[3]) ? node481 : 3'b101;
									assign node481 = (inp[5]) ? 3'b001 : node482;
										assign node482 = (inp[11]) ? 3'b001 : 3'b101;
								assign node486 = (inp[1]) ? node492 : node487;
									assign node487 = (inp[2]) ? node489 : 3'b101;
										assign node489 = (inp[11]) ? 3'b001 : 3'b101;
									assign node492 = (inp[2]) ? 3'b110 : node493;
										assign node493 = (inp[5]) ? 3'b001 : 3'b110;
						assign node497 = (inp[1]) ? node513 : node498;
							assign node498 = (inp[8]) ? node508 : node499;
								assign node499 = (inp[4]) ? node501 : 3'b010;
									assign node501 = (inp[3]) ? 3'b010 : node502;
										assign node502 = (inp[2]) ? 3'b100 : node503;
											assign node503 = (inp[11]) ? 3'b010 : 3'b110;
								assign node508 = (inp[11]) ? 3'b110 : node509;
									assign node509 = (inp[3]) ? 3'b110 : 3'b001;
							assign node513 = (inp[8]) ? node527 : node514;
								assign node514 = (inp[4]) ? node520 : node515;
									assign node515 = (inp[2]) ? node517 : 3'b100;
										assign node517 = (inp[3]) ? 3'b100 : 3'b000;
									assign node520 = (inp[11]) ? node522 : 3'b010;
										assign node522 = (inp[5]) ? 3'b000 : node523;
											assign node523 = (inp[3]) ? 3'b000 : 3'b100;
								assign node527 = (inp[4]) ? 3'b100 : node528;
									assign node528 = (inp[3]) ? 3'b010 : 3'b110;
				assign node532 = (inp[10]) ? node576 : node533;
					assign node533 = (inp[7]) ? node541 : node534;
						assign node534 = (inp[11]) ? 3'b000 : node535;
							assign node535 = (inp[1]) ? 3'b000 : node536;
								assign node536 = (inp[8]) ? 3'b100 : 3'b000;
						assign node541 = (inp[2]) ? node565 : node542;
							assign node542 = (inp[11]) ? node556 : node543;
								assign node543 = (inp[3]) ? node549 : node544;
									assign node544 = (inp[1]) ? node546 : 3'b001;
										assign node546 = (inp[8]) ? 3'b010 : 3'b100;
									assign node549 = (inp[5]) ? 3'b010 : node550;
										assign node550 = (inp[1]) ? 3'b100 : node551;
											assign node551 = (inp[8]) ? 3'b110 : 3'b010;
								assign node556 = (inp[8]) ? node560 : node557;
									assign node557 = (inp[1]) ? 3'b000 : 3'b100;
									assign node560 = (inp[1]) ? 3'b100 : node561;
										assign node561 = (inp[3]) ? 3'b010 : 3'b110;
							assign node565 = (inp[1]) ? node569 : node566;
								assign node566 = (inp[8]) ? 3'b110 : 3'b100;
								assign node569 = (inp[5]) ? node573 : node570;
									assign node570 = (inp[8]) ? 3'b010 : 3'b100;
									assign node573 = (inp[8]) ? 3'b100 : 3'b000;
					assign node576 = (inp[1]) ? 3'b000 : node577;
						assign node577 = (inp[8]) ? node579 : 3'b000;
							assign node579 = (inp[7]) ? node581 : 3'b000;
								assign node581 = (inp[5]) ? 3'b100 : node582;
									assign node582 = (inp[11]) ? 3'b000 : node583;
										assign node583 = (inp[2]) ? 3'b100 : 3'b011;

endmodule