module dtc_split25_bm37 (
	input  wire [8-1:0] inp,
	output wire [63-1:0] outp
);

	wire [63-1:0] node1;
	wire [63-1:0] node2;
	wire [63-1:0] node3;
	wire [63-1:0] node4;
	wire [63-1:0] node5;
	wire [63-1:0] node9;
	wire [63-1:0] node12;
	wire [63-1:0] node13;
	wire [63-1:0] node16;
	wire [63-1:0] node18;
	wire [63-1:0] node20;
	wire [63-1:0] node23;
	wire [63-1:0] node24;
	wire [63-1:0] node25;
	wire [63-1:0] node26;
	wire [63-1:0] node30;
	wire [63-1:0] node32;
	wire [63-1:0] node35;
	wire [63-1:0] node36;
	wire [63-1:0] node39;
	wire [63-1:0] node42;
	wire [63-1:0] node43;
	wire [63-1:0] node44;
	wire [63-1:0] node47;
	wire [63-1:0] node48;
	wire [63-1:0] node51;
	wire [63-1:0] node53;
	wire [63-1:0] node55;
	wire [63-1:0] node58;
	wire [63-1:0] node59;
	wire [63-1:0] node60;
	wire [63-1:0] node61;
	wire [63-1:0] node62;
	wire [63-1:0] node67;
	wire [63-1:0] node69;
	wire [63-1:0] node72;
	wire [63-1:0] node73;
	wire [63-1:0] node74;
	wire [63-1:0] node77;
	wire [63-1:0] node80;
	wire [63-1:0] node81;
	wire [63-1:0] node84;

	assign outp = (inp[7]) ? node42 : node1;
		assign node1 = (inp[2]) ? node23 : node2;
			assign node2 = (inp[6]) ? node12 : node3;
				assign node3 = (inp[1]) ? node9 : node4;
					assign node4 = (inp[3]) ? 63'b100110101001100000110001101110110011010101001100000101001010101 : node5;
						assign node5 = (inp[0]) ? 63'b100111101001100000110001101110110010010101001101001101001010101 : 63'b100111101001100000110001101110110010010101001100001101001010101;
					assign node9 = (inp[3]) ? 63'b100001101001100000010001101110010010010101001100101101000010101 : 63'b100111101001100000010001101110010010010101001100101101000000101;
				assign node12 = (inp[3]) ? node16 : node13;
					assign node13 = (inp[4]) ? 63'b100110101001100000110001101110110001010101000101101101001010000 : 63'b100110101001100000110001101110110011010101000100001101001010001;
					assign node16 = (inp[1]) ? node18 : 63'b100110101001100000110001101110110011010001001100001101001010101;
						assign node18 = (inp[4]) ? node20 : 63'b100110101001100000110001101110100011010101001100100101001010100;
							assign node20 = (inp[0]) ? 63'b100110101001100000110001101110100011010101001100100101001010100 : 63'b100110101001100000110001101110100011010101001100100101001010100;
			assign node23 = (inp[0]) ? node35 : node24;
				assign node24 = (inp[5]) ? node30 : node25;
					assign node25 = (inp[4]) ? 63'b110111100001000000110001101100110011010101001100111101001010101 : node26;
						assign node26 = (inp[6]) ? 63'b100111101001100000111001101110110011010001001100100101001010100 : 63'b101110100001100000110001101110110011010101001100101101001010100;
					assign node30 = (inp[4]) ? node32 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node32 = (inp[1]) ? 63'b100111101001100000110101101110110011010101001100101101001010101 : 63'b100101101001110000110001101110110011010101001100101101001010101;
				assign node35 = (inp[4]) ? node39 : node36;
					assign node36 = (inp[1]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : 63'b100111101001000000110001101110110011000110001100101001001010101;
					assign node39 = (inp[5]) ? 63'b100001101001100000110001101110010010010101011101101101000010101 : 63'b100110101001100000110001101110110011010101011100000101001010101;
		assign node42 = (inp[2]) ? node58 : node43;
			assign node43 = (inp[6]) ? node47 : node44;
				assign node44 = (inp[3]) ? 63'b000111101001001000110001101010110011000101001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101000010101;
				assign node47 = (inp[3]) ? node51 : node48;
					assign node48 = (inp[4]) ? 63'b100111101001000000110001101000110111010101001100101100001010101 : 63'b100111101000000000110001100000110011010101001100101100001010101;
					assign node51 = (inp[5]) ? node53 : 63'b100111101011100000100001101110110010010101001100101101000010101;
						assign node53 = (inp[4]) ? node55 : 63'b100111101000000000110000100100110011010101101100101101001010101;
							assign node55 = (inp[0]) ? 63'b100111101001000000110000100100110011010101101101101101001010101 : 63'b100111101001000000110000100100110011010101101100101101001010101;
			assign node58 = (inp[0]) ? node72 : node59;
				assign node59 = (inp[4]) ? node67 : node60;
					assign node60 = (inp[5]) ? 63'b100111101001100100110001101110110011010101001100101101001010101 : node61;
						assign node61 = (inp[6]) ? 63'b100111101001100000110001101110110011010001001100101101001010100 : node62;
							assign node62 = (inp[3]) ? 63'b100111101001100000110001101110110011010101001100001101001010101 : 63'b100111101001100000110001101110110011010101001110101101001010101;
					assign node67 = (inp[6]) ? node69 : 63'b100111101001000000110001101110110011100100001100101001001010101;
						assign node69 = (inp[5]) ? 63'b100101101001110000110001101110110011010101001100101101001010101 : 63'b100111001001100000110001101110110011010101000100101101001000001;
				assign node72 = (inp[4]) ? node80 : node73;
					assign node73 = (inp[1]) ? node77 : node74;
						assign node74 = (inp[6]) ? 63'b100111101011000000110001101110110011000110001100101001001010101 : 63'b100001101001000000110001101110110011000110001100101001001010101;
						assign node77 = (inp[5]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node80 = (inp[6]) ? node84 : node81;
						assign node81 = (inp[5]) ? 63'b100111101000000000110001101001110011010101011101101100001010101 : 63'b100111101000000000110000101100110011010101011100101101001011101;
						assign node84 = (inp[3]) ? 63'b100111101001100000100001101110110010010101011100101101000010101 : 63'b100111101001100000110001001110110011010101011100101101000010101;

endmodule