module dtc_split875_bm76 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node396;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node422;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node460;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node632;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node711;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node764;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node806;

	assign outp = (inp[9]) ? node554 : node1;
		assign node1 = (inp[6]) ? node261 : node2;
			assign node2 = (inp[10]) ? node98 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[3]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[8]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? node13 : 3'b111;
										assign node13 = (inp[5]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node55 : node18;
						assign node18 = (inp[8]) ? node36 : node19;
							assign node19 = (inp[3]) ? node21 : 3'b111;
								assign node21 = (inp[4]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? node31 : node24;
										assign node24 = (inp[0]) ? node26 : 3'b111;
											assign node26 = (inp[1]) ? node28 : 3'b111;
												assign node28 = (inp[2]) ? 3'b011 : 3'b111;
										assign node31 = (inp[1]) ? 3'b011 : node32;
											assign node32 = (inp[0]) ? 3'b011 : 3'b111;
							assign node36 = (inp[3]) ? 3'b011 : node37;
								assign node37 = (inp[4]) ? node39 : 3'b111;
									assign node39 = (inp[0]) ? node47 : node40;
										assign node40 = (inp[5]) ? node42 : 3'b111;
											assign node42 = (inp[1]) ? 3'b011 : node43;
												assign node43 = (inp[2]) ? 3'b011 : 3'b111;
										assign node47 = (inp[2]) ? 3'b011 : node48;
											assign node48 = (inp[5]) ? 3'b011 : node49;
												assign node49 = (inp[1]) ? 3'b011 : 3'b111;
						assign node55 = (inp[8]) ? node81 : node56;
							assign node56 = (inp[4]) ? node64 : node57;
								assign node57 = (inp[3]) ? 3'b011 : node58;
									assign node58 = (inp[0]) ? node60 : 3'b111;
										assign node60 = (inp[5]) ? 3'b011 : 3'b111;
								assign node64 = (inp[3]) ? node66 : 3'b011;
									assign node66 = (inp[0]) ? node74 : node67;
										assign node67 = (inp[5]) ? node69 : 3'b011;
											assign node69 = (inp[2]) ? 3'b101 : node70;
												assign node70 = (inp[1]) ? 3'b101 : 3'b011;
										assign node74 = (inp[1]) ? 3'b101 : node75;
											assign node75 = (inp[5]) ? 3'b101 : node76;
												assign node76 = (inp[2]) ? 3'b101 : 3'b011;
							assign node81 = (inp[3]) ? node89 : node82;
								assign node82 = (inp[4]) ? node84 : 3'b011;
									assign node84 = (inp[0]) ? 3'b101 : node85;
										assign node85 = (inp[5]) ? 3'b101 : 3'b011;
								assign node89 = (inp[4]) ? node91 : 3'b101;
									assign node91 = (inp[0]) ? node93 : 3'b101;
										assign node93 = (inp[1]) ? node95 : 3'b101;
											assign node95 = (inp[5]) ? 3'b001 : 3'b101;
				assign node98 = (inp[7]) ? node162 : node99;
					assign node99 = (inp[11]) ? node141 : node100;
						assign node100 = (inp[8]) ? node122 : node101;
							assign node101 = (inp[3]) ? node111 : node102;
								assign node102 = (inp[1]) ? node104 : 3'b111;
									assign node104 = (inp[0]) ? node106 : 3'b111;
										assign node106 = (inp[5]) ? node108 : 3'b111;
											assign node108 = (inp[4]) ? 3'b011 : 3'b111;
								assign node111 = (inp[1]) ? 3'b011 : node112;
									assign node112 = (inp[2]) ? 3'b011 : node113;
										assign node113 = (inp[0]) ? 3'b011 : node114;
											assign node114 = (inp[5]) ? 3'b011 : node115;
												assign node115 = (inp[4]) ? 3'b011 : 3'b111;
							assign node122 = (inp[3]) ? node124 : 3'b011;
								assign node124 = (inp[4]) ? 3'b101 : node125;
									assign node125 = (inp[5]) ? node133 : node126;
										assign node126 = (inp[2]) ? node128 : 3'b011;
											assign node128 = (inp[0]) ? node130 : 3'b011;
												assign node130 = (inp[1]) ? 3'b101 : 3'b011;
										assign node133 = (inp[0]) ? 3'b101 : node134;
											assign node134 = (inp[1]) ? node136 : 3'b011;
												assign node136 = (inp[2]) ? 3'b101 : 3'b011;
						assign node141 = (inp[3]) ? node151 : node142;
							assign node142 = (inp[8]) ? 3'b101 : node143;
								assign node143 = (inp[5]) ? node145 : 3'b011;
									assign node145 = (inp[4]) ? node147 : 3'b011;
										assign node147 = (inp[0]) ? 3'b101 : 3'b011;
							assign node151 = (inp[8]) ? node153 : 3'b101;
								assign node153 = (inp[4]) ? 3'b001 : node154;
									assign node154 = (inp[0]) ? 3'b001 : node155;
										assign node155 = (inp[5]) ? node157 : 3'b101;
											assign node157 = (inp[1]) ? 3'b001 : 3'b101;
					assign node162 = (inp[11]) ? node212 : node163;
						assign node163 = (inp[8]) ? node187 : node164;
							assign node164 = (inp[4]) ? node180 : node165;
								assign node165 = (inp[3]) ? 3'b101 : node166;
									assign node166 = (inp[1]) ? node172 : node167;
										assign node167 = (inp[5]) ? node169 : 3'b011;
											assign node169 = (inp[0]) ? 3'b101 : 3'b011;
										assign node172 = (inp[5]) ? node176 : node173;
											assign node173 = (inp[0]) ? 3'b111 : 3'b011;
											assign node176 = (inp[0]) ? 3'b101 : 3'b111;
								assign node180 = (inp[3]) ? node182 : 3'b101;
									assign node182 = (inp[0]) ? 3'b001 : node183;
										assign node183 = (inp[5]) ? 3'b001 : 3'b101;
							assign node187 = (inp[3]) ? node203 : node188;
								assign node188 = (inp[4]) ? node196 : node189;
									assign node189 = (inp[5]) ? node191 : 3'b101;
										assign node191 = (inp[2]) ? node193 : 3'b101;
											assign node193 = (inp[0]) ? 3'b001 : 3'b101;
									assign node196 = (inp[2]) ? 3'b001 : node197;
										assign node197 = (inp[0]) ? 3'b001 : node198;
											assign node198 = (inp[5]) ? 3'b001 : 3'b101;
								assign node203 = (inp[5]) ? node205 : 3'b001;
									assign node205 = (inp[0]) ? node207 : 3'b001;
										assign node207 = (inp[1]) ? node209 : 3'b001;
											assign node209 = (inp[4]) ? 3'b110 : 3'b001;
						assign node212 = (inp[8]) ? node240 : node213;
							assign node213 = (inp[3]) ? node221 : node214;
								assign node214 = (inp[0]) ? 3'b001 : node215;
									assign node215 = (inp[4]) ? 3'b001 : node216;
										assign node216 = (inp[5]) ? 3'b001 : 3'b101;
								assign node221 = (inp[4]) ? node231 : node222;
									assign node222 = (inp[1]) ? node224 : 3'b001;
										assign node224 = (inp[0]) ? node226 : 3'b001;
											assign node226 = (inp[5]) ? node228 : 3'b001;
												assign node228 = (inp[2]) ? 3'b110 : 3'b001;
									assign node231 = (inp[5]) ? 3'b110 : node232;
										assign node232 = (inp[0]) ? 3'b110 : node233;
											assign node233 = (inp[1]) ? node235 : 3'b001;
												assign node235 = (inp[2]) ? 3'b110 : 3'b001;
							assign node240 = (inp[3]) ? node254 : node241;
								assign node241 = (inp[4]) ? node249 : node242;
									assign node242 = (inp[5]) ? node244 : 3'b001;
										assign node244 = (inp[2]) ? node246 : 3'b001;
											assign node246 = (inp[0]) ? 3'b110 : 3'b001;
									assign node249 = (inp[2]) ? 3'b110 : node250;
										assign node250 = (inp[1]) ? 3'b110 : 3'b001;
								assign node254 = (inp[0]) ? node256 : 3'b110;
									assign node256 = (inp[4]) ? node258 : 3'b110;
										assign node258 = (inp[5]) ? 3'b010 : 3'b110;
			assign node261 = (inp[10]) ? node431 : node262;
				assign node262 = (inp[7]) ? node332 : node263;
					assign node263 = (inp[11]) ? node301 : node264;
						assign node264 = (inp[3]) ? node284 : node265;
							assign node265 = (inp[8]) ? node277 : node266;
								assign node266 = (inp[2]) ? node268 : 3'b011;
									assign node268 = (inp[1]) ? node270 : 3'b101;
										assign node270 = (inp[4]) ? node272 : 3'b011;
											assign node272 = (inp[0]) ? node274 : 3'b011;
												assign node274 = (inp[5]) ? 3'b101 : 3'b011;
								assign node277 = (inp[5]) ? 3'b101 : node278;
									assign node278 = (inp[4]) ? 3'b101 : node279;
										assign node279 = (inp[0]) ? 3'b101 : 3'b011;
							assign node284 = (inp[8]) ? node294 : node285;
								assign node285 = (inp[5]) ? 3'b101 : node286;
									assign node286 = (inp[0]) ? 3'b101 : node287;
										assign node287 = (inp[4]) ? 3'b101 : node288;
											assign node288 = (inp[1]) ? 3'b101 : 3'b011;
								assign node294 = (inp[4]) ? 3'b001 : node295;
									assign node295 = (inp[5]) ? node297 : 3'b101;
										assign node297 = (inp[0]) ? 3'b001 : 3'b101;
						assign node301 = (inp[8]) ? node319 : node302;
							assign node302 = (inp[3]) ? node310 : node303;
								assign node303 = (inp[5]) ? node305 : 3'b101;
									assign node305 = (inp[0]) ? node307 : 3'b101;
										assign node307 = (inp[4]) ? 3'b001 : 3'b101;
								assign node310 = (inp[2]) ? 3'b001 : node311;
									assign node311 = (inp[1]) ? 3'b001 : node312;
										assign node312 = (inp[5]) ? 3'b001 : node313;
											assign node313 = (inp[4]) ? 3'b001 : 3'b101;
							assign node319 = (inp[3]) ? node321 : 3'b001;
								assign node321 = (inp[4]) ? 3'b110 : node322;
									assign node322 = (inp[0]) ? 3'b110 : node323;
										assign node323 = (inp[5]) ? node325 : 3'b001;
											assign node325 = (inp[1]) ? 3'b110 : node326;
												assign node326 = (inp[2]) ? 3'b110 : 3'b001;
					assign node332 = (inp[11]) ? node382 : node333;
						assign node333 = (inp[8]) ? node363 : node334;
							assign node334 = (inp[4]) ? node348 : node335;
								assign node335 = (inp[3]) ? 3'b001 : node336;
									assign node336 = (inp[1]) ? node342 : node337;
										assign node337 = (inp[0]) ? node339 : 3'b101;
											assign node339 = (inp[5]) ? 3'b001 : 3'b101;
										assign node342 = (inp[0]) ? 3'b001 : node343;
											assign node343 = (inp[5]) ? 3'b001 : 3'b101;
								assign node348 = (inp[3]) ? node350 : 3'b001;
									assign node350 = (inp[0]) ? node358 : node351;
										assign node351 = (inp[5]) ? node353 : 3'b001;
											assign node353 = (inp[1]) ? 3'b110 : node354;
												assign node354 = (inp[2]) ? 3'b110 : 3'b111;
										assign node358 = (inp[2]) ? 3'b110 : node359;
											assign node359 = (inp[1]) ? 3'b110 : 3'b111;
							assign node363 = (inp[3]) ? node371 : node364;
								assign node364 = (inp[4]) ? node366 : 3'b001;
									assign node366 = (inp[5]) ? 3'b110 : node367;
										assign node367 = (inp[0]) ? 3'b110 : 3'b001;
								assign node371 = (inp[5]) ? node373 : 3'b110;
									assign node373 = (inp[0]) ? node375 : 3'b110;
										assign node375 = (inp[4]) ? node377 : 3'b110;
											assign node377 = (inp[2]) ? 3'b010 : node378;
												assign node378 = (inp[1]) ? 3'b010 : 3'b110;
						assign node382 = (inp[3]) ? node414 : node383;
							assign node383 = (inp[4]) ? node401 : node384;
								assign node384 = (inp[8]) ? node396 : node385;
									assign node385 = (inp[0]) ? node391 : node386;
										assign node386 = (inp[1]) ? node388 : 3'b001;
											assign node388 = (inp[5]) ? 3'b110 : 3'b001;
										assign node391 = (inp[1]) ? 3'b110 : node392;
											assign node392 = (inp[5]) ? 3'b110 : 3'b001;
									assign node396 = (inp[2]) ? node398 : 3'b110;
										assign node398 = (inp[1]) ? 3'b010 : 3'b110;
								assign node401 = (inp[8]) ? node403 : 3'b110;
									assign node403 = (inp[1]) ? node409 : node404;
										assign node404 = (inp[2]) ? 3'b110 : node405;
											assign node405 = (inp[5]) ? 3'b010 : 3'b110;
										assign node409 = (inp[2]) ? 3'b010 : node410;
											assign node410 = (inp[5]) ? 3'b010 : 3'b110;
							assign node414 = (inp[8]) ? node422 : node415;
								assign node415 = (inp[4]) ? node417 : 3'b110;
									assign node417 = (inp[5]) ? 3'b010 : node418;
										assign node418 = (inp[0]) ? 3'b010 : 3'b110;
								assign node422 = (inp[5]) ? node424 : 3'b010;
									assign node424 = (inp[0]) ? node426 : 3'b010;
										assign node426 = (inp[1]) ? node428 : 3'b010;
											assign node428 = (inp[2]) ? 3'b010 : 3'b100;
				assign node431 = (inp[7]) ? node473 : node432;
					assign node432 = (inp[11]) ? node456 : node433;
						assign node433 = (inp[8]) ? node443 : node434;
							assign node434 = (inp[3]) ? 3'b110 : node435;
								assign node435 = (inp[4]) ? node437 : 3'b001;
									assign node437 = (inp[0]) ? node439 : 3'b001;
										assign node439 = (inp[5]) ? 3'b110 : 3'b001;
							assign node443 = (inp[3]) ? node445 : 3'b110;
								assign node445 = (inp[4]) ? 3'b010 : node446;
									assign node446 = (inp[5]) ? 3'b010 : node447;
										assign node447 = (inp[0]) ? node449 : 3'b110;
											assign node449 = (inp[1]) ? 3'b010 : node450;
												assign node450 = (inp[2]) ? 3'b010 : 3'b110;
						assign node456 = (inp[8]) ? node464 : node457;
							assign node457 = (inp[3]) ? 3'b010 : node458;
								assign node458 = (inp[2]) ? node460 : 3'b110;
									assign node460 = (inp[4]) ? 3'b010 : 3'b110;
							assign node464 = (inp[3]) ? node466 : 3'b010;
								assign node466 = (inp[4]) ? 3'b100 : node467;
									assign node467 = (inp[0]) ? 3'b100 : node468;
										assign node468 = (inp[5]) ? 3'b100 : 3'b010;
					assign node473 = (inp[11]) ? node521 : node474;
						assign node474 = (inp[3]) ? node498 : node475;
							assign node475 = (inp[8]) ? node483 : node476;
								assign node476 = (inp[5]) ? 3'b010 : node477;
									assign node477 = (inp[4]) ? 3'b010 : node478;
										assign node478 = (inp[0]) ? 3'b010 : 3'b110;
								assign node483 = (inp[4]) ? node491 : node484;
									assign node484 = (inp[0]) ? node486 : 3'b010;
										assign node486 = (inp[5]) ? node488 : 3'b010;
											assign node488 = (inp[2]) ? 3'b100 : 3'b010;
									assign node491 = (inp[1]) ? 3'b100 : node492;
										assign node492 = (inp[2]) ? 3'b100 : node493;
											assign node493 = (inp[5]) ? 3'b100 : 3'b010;
							assign node498 = (inp[8]) ? node514 : node499;
								assign node499 = (inp[4]) ? node507 : node500;
									assign node500 = (inp[5]) ? node502 : 3'b010;
										assign node502 = (inp[2]) ? node504 : 3'b010;
											assign node504 = (inp[0]) ? 3'b100 : 3'b010;
									assign node507 = (inp[0]) ? 3'b100 : node508;
										assign node508 = (inp[5]) ? 3'b100 : node509;
											assign node509 = (inp[2]) ? 3'b100 : 3'b010;
								assign node514 = (inp[5]) ? node516 : 3'b100;
									assign node516 = (inp[0]) ? node518 : 3'b100;
										assign node518 = (inp[4]) ? 3'b000 : 3'b100;
						assign node521 = (inp[8]) ? node545 : node522;
							assign node522 = (inp[3]) ? node530 : node523;
								assign node523 = (inp[5]) ? 3'b100 : node524;
									assign node524 = (inp[4]) ? 3'b100 : node525;
										assign node525 = (inp[0]) ? 3'b100 : 3'b010;
								assign node530 = (inp[4]) ? node538 : node531;
									assign node531 = (inp[5]) ? node533 : 3'b100;
										assign node533 = (inp[2]) ? node535 : 3'b100;
											assign node535 = (inp[0]) ? 3'b000 : 3'b100;
									assign node538 = (inp[1]) ? 3'b000 : node539;
										assign node539 = (inp[2]) ? 3'b000 : node540;
											assign node540 = (inp[5]) ? 3'b000 : 3'b100;
							assign node545 = (inp[4]) ? 3'b000 : node546;
								assign node546 = (inp[3]) ? 3'b000 : node547;
									assign node547 = (inp[0]) ? node549 : 3'b100;
										assign node549 = (inp[5]) ? 3'b000 : 3'b100;
		assign node554 = (inp[6]) ? node776 : node555;
			assign node555 = (inp[10]) ? node675 : node556;
				assign node556 = (inp[7]) ? node594 : node557;
					assign node557 = (inp[11]) ? node575 : node558;
						assign node558 = (inp[8]) ? node566 : node559;
							assign node559 = (inp[3]) ? 3'b001 : node560;
								assign node560 = (inp[4]) ? node562 : 3'b101;
									assign node562 = (inp[5]) ? 3'b001 : 3'b101;
							assign node566 = (inp[3]) ? node568 : 3'b001;
								assign node568 = (inp[5]) ? 3'b110 : node569;
									assign node569 = (inp[4]) ? 3'b110 : node570;
										assign node570 = (inp[0]) ? 3'b110 : 3'b001;
						assign node575 = (inp[3]) ? node585 : node576;
							assign node576 = (inp[8]) ? 3'b110 : node577;
								assign node577 = (inp[4]) ? node579 : 3'b001;
									assign node579 = (inp[5]) ? 3'b110 : node580;
										assign node580 = (inp[0]) ? 3'b110 : 3'b001;
							assign node585 = (inp[8]) ? node587 : 3'b110;
								assign node587 = (inp[0]) ? 3'b010 : node588;
									assign node588 = (inp[4]) ? 3'b010 : node589;
										assign node589 = (inp[5]) ? 3'b010 : 3'b110;
					assign node594 = (inp[11]) ? node640 : node595;
						assign node595 = (inp[8]) ? node619 : node596;
							assign node596 = (inp[3]) ? node604 : node597;
								assign node597 = (inp[5]) ? 3'b110 : node598;
									assign node598 = (inp[0]) ? 3'b110 : node599;
										assign node599 = (inp[4]) ? 3'b110 : 3'b001;
								assign node604 = (inp[4]) ? node612 : node605;
									assign node605 = (inp[1]) ? node607 : 3'b110;
										assign node607 = (inp[0]) ? node609 : 3'b110;
											assign node609 = (inp[5]) ? 3'b010 : 3'b110;
									assign node612 = (inp[0]) ? 3'b010 : node613;
										assign node613 = (inp[1]) ? 3'b010 : node614;
											assign node614 = (inp[5]) ? 3'b010 : 3'b110;
							assign node619 = (inp[3]) ? node627 : node620;
								assign node620 = (inp[4]) ? 3'b010 : node621;
									assign node621 = (inp[5]) ? node623 : 3'b110;
										assign node623 = (inp[0]) ? 3'b010 : 3'b110;
								assign node627 = (inp[4]) ? node629 : 3'b010;
									assign node629 = (inp[0]) ? node635 : node630;
										assign node630 = (inp[2]) ? node632 : 3'b010;
											assign node632 = (inp[5]) ? 3'b100 : 3'b010;
										assign node635 = (inp[5]) ? 3'b100 : node636;
											assign node636 = (inp[2]) ? 3'b100 : 3'b010;
						assign node640 = (inp[8]) ? node654 : node641;
							assign node641 = (inp[3]) ? node645 : node642;
								assign node642 = (inp[4]) ? 3'b010 : 3'b110;
								assign node645 = (inp[4]) ? 3'b100 : node646;
									assign node646 = (inp[2]) ? node648 : 3'b010;
										assign node648 = (inp[0]) ? node650 : 3'b010;
											assign node650 = (inp[5]) ? 3'b100 : 3'b010;
							assign node654 = (inp[4]) ? node662 : node655;
								assign node655 = (inp[3]) ? 3'b100 : node656;
									assign node656 = (inp[0]) ? node658 : 3'b010;
										assign node658 = (inp[5]) ? 3'b100 : 3'b010;
								assign node662 = (inp[3]) ? node664 : 3'b100;
									assign node664 = (inp[1]) ? node670 : node665;
										assign node665 = (inp[5]) ? node667 : 3'b100;
											assign node667 = (inp[0]) ? 3'b000 : 3'b100;
										assign node670 = (inp[0]) ? 3'b000 : node671;
											assign node671 = (inp[2]) ? 3'b100 : 3'b000;
				assign node675 = (inp[7]) ? node751 : node676;
					assign node676 = (inp[11]) ? node706 : node677;
						assign node677 = (inp[8]) ? node685 : node678;
							assign node678 = (inp[3]) ? 3'b010 : node679;
								assign node679 = (inp[4]) ? node681 : 3'b110;
									assign node681 = (inp[1]) ? 3'b010 : 3'b110;
							assign node685 = (inp[3]) ? node697 : node686;
								assign node686 = (inp[2]) ? node688 : 3'b010;
									assign node688 = (inp[1]) ? node690 : 3'b100;
										assign node690 = (inp[5]) ? node692 : 3'b010;
											assign node692 = (inp[0]) ? node694 : 3'b010;
												assign node694 = (inp[4]) ? 3'b100 : 3'b010;
								assign node697 = (inp[4]) ? 3'b100 : node698;
									assign node698 = (inp[0]) ? 3'b100 : node699;
										assign node699 = (inp[5]) ? 3'b100 : node700;
											assign node700 = (inp[2]) ? 3'b100 : 3'b010;
						assign node706 = (inp[8]) ? node730 : node707;
							assign node707 = (inp[3]) ? node723 : node708;
								assign node708 = (inp[4]) ? node716 : node709;
									assign node709 = (inp[5]) ? node711 : 3'b000;
										assign node711 = (inp[0]) ? node713 : 3'b000;
											assign node713 = (inp[2]) ? 3'b100 : 3'b000;
									assign node716 = (inp[2]) ? 3'b100 : node717;
										assign node717 = (inp[5]) ? 3'b100 : node718;
											assign node718 = (inp[1]) ? 3'b100 : 3'b000;
								assign node723 = (inp[0]) ? node725 : 3'b100;
									assign node725 = (inp[4]) ? node727 : 3'b100;
										assign node727 = (inp[5]) ? 3'b000 : 3'b100;
							assign node730 = (inp[3]) ? node742 : node731;
								assign node731 = (inp[2]) ? node733 : 3'b100;
									assign node733 = (inp[1]) ? node735 : 3'b000;
										assign node735 = (inp[0]) ? node737 : 3'b100;
											assign node737 = (inp[4]) ? node739 : 3'b100;
												assign node739 = (inp[5]) ? 3'b000 : 3'b100;
								assign node742 = (inp[5]) ? 3'b000 : node743;
									assign node743 = (inp[2]) ? 3'b000 : node744;
										assign node744 = (inp[4]) ? 3'b000 : node745;
											assign node745 = (inp[0]) ? 3'b000 : 3'b100;
					assign node751 = (inp[11]) ? 3'b000 : node752;
						assign node752 = (inp[8]) ? node768 : node753;
							assign node753 = (inp[3]) ? node761 : node754;
								assign node754 = (inp[5]) ? 3'b100 : node755;
									assign node755 = (inp[4]) ? 3'b100 : node756;
										assign node756 = (inp[0]) ? 3'b100 : 3'b000;
								assign node761 = (inp[4]) ? 3'b000 : node762;
									assign node762 = (inp[5]) ? node764 : 3'b100;
										assign node764 = (inp[0]) ? 3'b000 : 3'b100;
							assign node768 = (inp[0]) ? 3'b000 : node769;
								assign node769 = (inp[4]) ? 3'b000 : node770;
									assign node770 = (inp[5]) ? 3'b000 : 3'b100;
			assign node776 = (inp[10]) ? 3'b000 : node777;
				assign node777 = (inp[7]) ? 3'b000 : node778;
					assign node778 = (inp[11]) ? node802 : node779;
						assign node779 = (inp[8]) ? node787 : node780;
							assign node780 = (inp[3]) ? 3'b100 : node781;
								assign node781 = (inp[4]) ? node783 : 3'b010;
									assign node783 = (inp[1]) ? 3'b100 : 3'b010;
							assign node787 = (inp[3]) ? node793 : node788;
								assign node788 = (inp[2]) ? node790 : 3'b100;
									assign node790 = (inp[1]) ? 3'b100 : 3'b000;
								assign node793 = (inp[0]) ? 3'b000 : node794;
									assign node794 = (inp[4]) ? 3'b000 : node795;
										assign node795 = (inp[5]) ? 3'b000 : node796;
											assign node796 = (inp[2]) ? 3'b000 : 3'b100;
						assign node802 = (inp[3]) ? 3'b000 : node803;
							assign node803 = (inp[8]) ? 3'b000 : node804;
								assign node804 = (inp[2]) ? node806 : 3'b100;
									assign node806 = (inp[4]) ? 3'b000 : 3'b100;

endmodule