module dtc_split75_bm67 (
	input  wire [10-1:0] inp,
	output wire [77-1:0] outp
);

	wire [77-1:0] node1;
	wire [77-1:0] node2;
	wire [77-1:0] node3;
	wire [77-1:0] node6;
	wire [77-1:0] node9;
	wire [77-1:0] node10;
	wire [77-1:0] node13;
	wire [77-1:0] node16;
	wire [77-1:0] node17;
	wire [77-1:0] node18;
	wire [77-1:0] node21;
	wire [77-1:0] node24;
	wire [77-1:0] node25;
	wire [77-1:0] node28;

	assign outp = (inp[8]) ? node16 : node1;
		assign node1 = (inp[1]) ? node9 : node2;
			assign node2 = (inp[6]) ? node6 : node3;
				assign node3 = (inp[7]) ? 77'b00100100000001000101000100010000000000000000100000010000011011000110100000000 : 77'b11100000000101100101000011100000000100000000110000010101000010000100010100100;
				assign node6 = (inp[2]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b10100000100000100000000011010000000000000000001100010000010001000110010000100;
			assign node9 = (inp[0]) ? node13 : node10;
				assign node10 = (inp[6]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000100000100000011000001100100000000010100000100000001000000000001000;
				assign node13 = (inp[4]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;
		assign node16 = (inp[7]) ? node24 : node17;
			assign node17 = (inp[1]) ? node21 : node18;
				assign node18 = (inp[6]) ? 77'b00000000000000000000010000000000000000000000000000000000000000000000000000000 : 77'b00000000100000100000010010000000000000000000001000000000010011000110100000000;
				assign node21 = (inp[0]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000100000000000000000000000000000000000000000000010000010000;
			assign node24 = (inp[9]) ? node28 : node25;
				assign node25 = (inp[1]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000100000000000000000000000000000000000000000000000000000000000000000000;
				assign node28 = (inp[5]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule