module dtc_split75_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node730;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node892;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node912;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node929;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1024;
	wire [3-1:0] node1027;
	wire [3-1:0] node1029;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1117;
	wire [3-1:0] node1120;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1130;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1198;
	wire [3-1:0] node1201;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1231;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1277;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1313;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1328;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1335;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1351;
	wire [3-1:0] node1352;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1366;
	wire [3-1:0] node1367;
	wire [3-1:0] node1370;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1379;
	wire [3-1:0] node1382;
	wire [3-1:0] node1384;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1389;
	wire [3-1:0] node1393;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1401;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1454;
	wire [3-1:0] node1457;
	wire [3-1:0] node1461;
	wire [3-1:0] node1462;
	wire [3-1:0] node1463;
	wire [3-1:0] node1465;
	wire [3-1:0] node1468;
	wire [3-1:0] node1470;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1481;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1485;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1495;
	wire [3-1:0] node1498;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1507;
	wire [3-1:0] node1510;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;

	assign outp = (inp[6]) ? node522 : node1;
		assign node1 = (inp[3]) ? node367 : node2;
			assign node2 = (inp[0]) ? node66 : node3;
				assign node3 = (inp[9]) ? node41 : node4;
					assign node4 = (inp[8]) ? node34 : node5;
						assign node5 = (inp[7]) ? node21 : node6;
							assign node6 = (inp[10]) ? node14 : node7;
								assign node7 = (inp[5]) ? node9 : 3'b000;
									assign node9 = (inp[11]) ? node11 : 3'b010;
										assign node11 = (inp[4]) ? 3'b010 : 3'b000;
								assign node14 = (inp[5]) ? node16 : 3'b010;
									assign node16 = (inp[11]) ? node18 : 3'b100;
										assign node18 = (inp[4]) ? 3'b100 : 3'b110;
							assign node21 = (inp[5]) ? node23 : 3'b000;
								assign node23 = (inp[4]) ? node27 : node24;
									assign node24 = (inp[10]) ? 3'b010 : 3'b000;
									assign node27 = (inp[2]) ? node29 : 3'b000;
										assign node29 = (inp[10]) ? 3'b000 : node30;
											assign node30 = (inp[11]) ? 3'b000 : 3'b010;
						assign node34 = (inp[5]) ? node36 : 3'b000;
							assign node36 = (inp[10]) ? node38 : 3'b000;
								assign node38 = (inp[7]) ? 3'b000 : 3'b010;
					assign node41 = (inp[5]) ? node43 : 3'b000;
						assign node43 = (inp[8]) ? 3'b000 : node44;
							assign node44 = (inp[7]) ? node54 : node45;
								assign node45 = (inp[10]) ? 3'b000 : node46;
									assign node46 = (inp[2]) ? 3'b000 : node47;
										assign node47 = (inp[4]) ? 3'b000 : node48;
											assign node48 = (inp[1]) ? 3'b010 : 3'b000;
								assign node54 = (inp[10]) ? node62 : node55;
									assign node55 = (inp[4]) ? node57 : 3'b000;
										assign node57 = (inp[11]) ? 3'b000 : node58;
											assign node58 = (inp[1]) ? 3'b010 : 3'b000;
									assign node62 = (inp[4]) ? 3'b000 : 3'b010;
				assign node66 = (inp[7]) ? node182 : node67;
					assign node67 = (inp[9]) ? node155 : node68;
						assign node68 = (inp[10]) ? node124 : node69;
							assign node69 = (inp[11]) ? node93 : node70;
								assign node70 = (inp[4]) ? node80 : node71;
									assign node71 = (inp[1]) ? 3'b110 : node72;
										assign node72 = (inp[5]) ? node76 : node73;
											assign node73 = (inp[8]) ? 3'b100 : 3'b110;
											assign node76 = (inp[8]) ? 3'b110 : 3'b000;
									assign node80 = (inp[8]) ? node86 : node81;
										assign node81 = (inp[1]) ? 3'b100 : node82;
											assign node82 = (inp[5]) ? 3'b000 : 3'b110;
										assign node86 = (inp[5]) ? node90 : node87;
											assign node87 = (inp[1]) ? 3'b010 : 3'b000;
											assign node90 = (inp[1]) ? 3'b100 : 3'b110;
								assign node93 = (inp[4]) ? node105 : node94;
									assign node94 = (inp[8]) ? node100 : node95;
										assign node95 = (inp[5]) ? node97 : 3'b010;
											assign node97 = (inp[1]) ? 3'b100 : 3'b000;
										assign node100 = (inp[5]) ? 3'b010 : node101;
											assign node101 = (inp[1]) ? 3'b110 : 3'b100;
									assign node105 = (inp[1]) ? node117 : node106;
										assign node106 = (inp[2]) ? node112 : node107;
											assign node107 = (inp[5]) ? node109 : 3'b000;
												assign node109 = (inp[8]) ? 3'b110 : 3'b000;
											assign node112 = (inp[5]) ? node114 : 3'b110;
												assign node114 = (inp[8]) ? 3'b110 : 3'b000;
										assign node117 = (inp[5]) ? node121 : node118;
											assign node118 = (inp[8]) ? 3'b000 : 3'b100;
											assign node121 = (inp[8]) ? 3'b100 : 3'b000;
							assign node124 = (inp[4]) ? node146 : node125;
								assign node125 = (inp[1]) ? node135 : node126;
									assign node126 = (inp[11]) ? node128 : 3'b000;
										assign node128 = (inp[8]) ? node132 : node129;
											assign node129 = (inp[5]) ? 3'b000 : 3'b100;
											assign node132 = (inp[5]) ? 3'b100 : 3'b000;
									assign node135 = (inp[5]) ? node141 : node136;
										assign node136 = (inp[8]) ? 3'b010 : node137;
											assign node137 = (inp[11]) ? 3'b100 : 3'b010;
										assign node141 = (inp[8]) ? node143 : 3'b100;
											assign node143 = (inp[11]) ? 3'b100 : 3'b010;
								assign node146 = (inp[8]) ? node148 : 3'b000;
									assign node148 = (inp[11]) ? 3'b000 : node149;
										assign node149 = (inp[2]) ? node151 : 3'b000;
											assign node151 = (inp[5]) ? 3'b000 : 3'b100;
						assign node155 = (inp[8]) ? node157 : 3'b000;
							assign node157 = (inp[5]) ? node173 : node158;
								assign node158 = (inp[10]) ? node166 : node159;
									assign node159 = (inp[4]) ? node161 : 3'b100;
										assign node161 = (inp[2]) ? node163 : 3'b000;
											assign node163 = (inp[11]) ? 3'b100 : 3'b000;
									assign node166 = (inp[4]) ? node168 : 3'b000;
										assign node168 = (inp[2]) ? node170 : 3'b000;
											assign node170 = (inp[11]) ? 3'b000 : 3'b100;
								assign node173 = (inp[4]) ? 3'b000 : node174;
									assign node174 = (inp[10]) ? 3'b000 : node175;
										assign node175 = (inp[1]) ? node177 : 3'b000;
											assign node177 = (inp[11]) ? 3'b000 : 3'b100;
					assign node182 = (inp[4]) ? node254 : node183;
						assign node183 = (inp[10]) ? node217 : node184;
							assign node184 = (inp[9]) ? node200 : node185;
								assign node185 = (inp[5]) ? node195 : node186;
									assign node186 = (inp[8]) ? node192 : node187;
										assign node187 = (inp[11]) ? node189 : 3'b001;
											assign node189 = (inp[1]) ? 3'b001 : 3'b000;
										assign node192 = (inp[1]) ? 3'b000 : 3'b010;
									assign node195 = (inp[8]) ? 3'b001 : node196;
										assign node196 = (inp[1]) ? 3'b110 : 3'b100;
								assign node200 = (inp[1]) ? node208 : node201;
									assign node201 = (inp[5]) ? node205 : node202;
										assign node202 = (inp[8]) ? 3'b000 : 3'b010;
										assign node205 = (inp[8]) ? 3'b010 : 3'b100;
									assign node208 = (inp[8]) ? node212 : node209;
										assign node209 = (inp[5]) ? 3'b100 : 3'b010;
										assign node212 = (inp[5]) ? 3'b010 : node213;
											assign node213 = (inp[11]) ? 3'b010 : 3'b110;
							assign node217 = (inp[5]) ? node237 : node218;
								assign node218 = (inp[8]) ? node226 : node219;
									assign node219 = (inp[1]) ? node223 : node220;
										assign node220 = (inp[9]) ? 3'b110 : 3'b100;
										assign node223 = (inp[9]) ? 3'b100 : 3'b110;
									assign node226 = (inp[9]) ? node234 : node227;
										assign node227 = (inp[11]) ? node231 : node228;
											assign node228 = (inp[1]) ? 3'b000 : 3'b100;
											assign node231 = (inp[1]) ? 3'b110 : 3'b100;
										assign node234 = (inp[1]) ? 3'b010 : 3'b110;
								assign node237 = (inp[8]) ? node243 : node238;
									assign node238 = (inp[9]) ? 3'b000 : node239;
										assign node239 = (inp[1]) ? 3'b010 : 3'b000;
									assign node243 = (inp[2]) ? node251 : node244;
										assign node244 = (inp[1]) ? node248 : node245;
											assign node245 = (inp[9]) ? 3'b110 : 3'b100;
											assign node248 = (inp[9]) ? 3'b100 : 3'b110;
										assign node251 = (inp[9]) ? 3'b100 : 3'b110;
						assign node254 = (inp[9]) ? node308 : node255;
							assign node255 = (inp[1]) ? node285 : node256;
								assign node256 = (inp[10]) ? node272 : node257;
									assign node257 = (inp[11]) ? node265 : node258;
										assign node258 = (inp[2]) ? 3'b000 : node259;
											assign node259 = (inp[5]) ? 3'b001 : node260;
												assign node260 = (inp[8]) ? 3'b100 : 3'b001;
										assign node265 = (inp[8]) ? node269 : node266;
											assign node266 = (inp[2]) ? 3'b100 : 3'b000;
											assign node269 = (inp[5]) ? 3'b010 : 3'b000;
									assign node272 = (inp[8]) ? node280 : node273;
										assign node273 = (inp[5]) ? node275 : 3'b010;
											assign node275 = (inp[2]) ? node277 : 3'b000;
												assign node277 = (inp[11]) ? 3'b000 : 3'b100;
										assign node280 = (inp[5]) ? 3'b010 : node281;
											assign node281 = (inp[2]) ? 3'b110 : 3'b000;
								assign node285 = (inp[10]) ? node301 : node286;
									assign node286 = (inp[5]) ? node292 : node287;
										assign node287 = (inp[8]) ? 3'b110 : node288;
											assign node288 = (inp[11]) ? 3'b010 : 3'b110;
										assign node292 = (inp[11]) ? node298 : node293;
											assign node293 = (inp[2]) ? node295 : 3'b010;
												assign node295 = (inp[8]) ? 3'b110 : 3'b010;
											assign node298 = (inp[8]) ? 3'b010 : 3'b100;
									assign node301 = (inp[5]) ? node303 : 3'b010;
										assign node303 = (inp[11]) ? 3'b000 : node304;
											assign node304 = (inp[8]) ? 3'b010 : 3'b100;
							assign node308 = (inp[10]) ? node342 : node309;
								assign node309 = (inp[8]) ? node327 : node310;
									assign node310 = (inp[2]) ? node318 : node311;
										assign node311 = (inp[1]) ? 3'b000 : node312;
											assign node312 = (inp[11]) ? 3'b000 : node313;
												assign node313 = (inp[5]) ? 3'b000 : 3'b010;
										assign node318 = (inp[1]) ? node324 : node319;
											assign node319 = (inp[5]) ? node321 : 3'b000;
												assign node321 = (inp[11]) ? 3'b100 : 3'b000;
											assign node324 = (inp[11]) ? 3'b000 : 3'b100;
									assign node327 = (inp[1]) ? node337 : node328;
										assign node328 = (inp[11]) ? node334 : node329;
											assign node329 = (inp[2]) ? 3'b100 : node330;
												assign node330 = (inp[5]) ? 3'b010 : 3'b110;
											assign node334 = (inp[5]) ? 3'b000 : 3'b010;
										assign node337 = (inp[5]) ? node339 : 3'b100;
											assign node339 = (inp[11]) ? 3'b000 : 3'b100;
								assign node342 = (inp[2]) ? node350 : node343;
									assign node343 = (inp[8]) ? node345 : 3'b000;
										assign node345 = (inp[1]) ? 3'b000 : node346;
											assign node346 = (inp[5]) ? 3'b000 : 3'b010;
									assign node350 = (inp[11]) ? node360 : node351;
										assign node351 = (inp[8]) ? node355 : node352;
											assign node352 = (inp[5]) ? 3'b100 : 3'b000;
											assign node355 = (inp[1]) ? 3'b000 : node356;
												assign node356 = (inp[5]) ? 3'b000 : 3'b010;
										assign node360 = (inp[5]) ? 3'b000 : node361;
											assign node361 = (inp[1]) ? 3'b000 : node362;
												assign node362 = (inp[8]) ? 3'b100 : 3'b000;
			assign node367 = (inp[7]) ? node397 : node368;
				assign node368 = (inp[4]) ? 3'b000 : node369;
					assign node369 = (inp[9]) ? 3'b000 : node370;
						assign node370 = (inp[5]) ? 3'b000 : node371;
							assign node371 = (inp[1]) ? node379 : node372;
								assign node372 = (inp[11]) ? 3'b000 : node373;
									assign node373 = (inp[0]) ? node375 : 3'b000;
										assign node375 = (inp[8]) ? 3'b100 : 3'b000;
								assign node379 = (inp[0]) ? node387 : node380;
									assign node380 = (inp[8]) ? 3'b000 : node381;
										assign node381 = (inp[10]) ? node383 : 3'b100;
											assign node383 = (inp[11]) ? 3'b000 : 3'b100;
									assign node387 = (inp[8]) ? node389 : 3'b000;
										assign node389 = (inp[11]) ? 3'b000 : node390;
											assign node390 = (inp[10]) ? 3'b000 : 3'b100;
				assign node397 = (inp[9]) ? node497 : node398;
					assign node398 = (inp[8]) ? node438 : node399;
						assign node399 = (inp[0]) ? node425 : node400;
							assign node400 = (inp[1]) ? node408 : node401;
								assign node401 = (inp[11]) ? 3'b000 : node402;
									assign node402 = (inp[10]) ? 3'b000 : node403;
										assign node403 = (inp[5]) ? 3'b010 : 3'b000;
								assign node408 = (inp[5]) ? node416 : node409;
									assign node409 = (inp[4]) ? node411 : 3'b010;
										assign node411 = (inp[11]) ? 3'b000 : node412;
											assign node412 = (inp[10]) ? 3'b000 : 3'b010;
									assign node416 = (inp[4]) ? node420 : node417;
										assign node417 = (inp[10]) ? 3'b100 : 3'b110;
										assign node420 = (inp[10]) ? 3'b000 : node421;
											assign node421 = (inp[11]) ? 3'b000 : 3'b100;
							assign node425 = (inp[5]) ? 3'b000 : node426;
								assign node426 = (inp[10]) ? 3'b000 : node427;
									assign node427 = (inp[11]) ? node431 : node428;
										assign node428 = (inp[1]) ? 3'b000 : 3'b100;
										assign node431 = (inp[1]) ? node433 : 3'b000;
											assign node433 = (inp[4]) ? 3'b000 : 3'b100;
						assign node438 = (inp[0]) ? node472 : node439;
							assign node439 = (inp[5]) ? node441 : 3'b100;
								assign node441 = (inp[1]) ? node461 : node442;
									assign node442 = (inp[2]) ? node456 : node443;
										assign node443 = (inp[4]) ? node451 : node444;
											assign node444 = (inp[10]) ? node448 : node445;
												assign node445 = (inp[11]) ? 3'b100 : 3'b000;
												assign node448 = (inp[11]) ? 3'b000 : 3'b100;
											assign node451 = (inp[11]) ? 3'b000 : node452;
												assign node452 = (inp[10]) ? 3'b100 : 3'b000;
										assign node456 = (inp[4]) ? 3'b100 : node457;
											assign node457 = (inp[11]) ? 3'b000 : 3'b100;
									assign node461 = (inp[11]) ? node465 : node462;
										assign node462 = (inp[10]) ? 3'b110 : 3'b010;
										assign node465 = (inp[4]) ? node469 : node466;
											assign node466 = (inp[10]) ? 3'b010 : 3'b110;
											assign node469 = (inp[10]) ? 3'b000 : 3'b100;
							assign node472 = (inp[4]) ? node490 : node473;
								assign node473 = (inp[10]) ? node485 : node474;
									assign node474 = (inp[5]) ? node480 : node475;
										assign node475 = (inp[1]) ? 3'b010 : node476;
											assign node476 = (inp[11]) ? 3'b100 : 3'b110;
										assign node480 = (inp[1]) ? 3'b100 : node481;
											assign node481 = (inp[11]) ? 3'b000 : 3'b100;
									assign node485 = (inp[5]) ? 3'b000 : node486;
										assign node486 = (inp[1]) ? 3'b100 : 3'b000;
								assign node490 = (inp[1]) ? 3'b000 : node491;
									assign node491 = (inp[10]) ? 3'b000 : node492;
										assign node492 = (inp[11]) ? 3'b000 : 3'b100;
					assign node497 = (inp[8]) ? node499 : 3'b000;
						assign node499 = (inp[0]) ? node513 : node500;
							assign node500 = (inp[5]) ? 3'b000 : node501;
								assign node501 = (inp[10]) ? node507 : node502;
									assign node502 = (inp[4]) ? node504 : 3'b100;
										assign node504 = (inp[1]) ? 3'b000 : 3'b100;
									assign node507 = (inp[1]) ? node509 : 3'b000;
										assign node509 = (inp[11]) ? 3'b000 : 3'b100;
							assign node513 = (inp[11]) ? 3'b000 : node514;
								assign node514 = (inp[5]) ? 3'b000 : node515;
									assign node515 = (inp[4]) ? 3'b000 : node516;
										assign node516 = (inp[10]) ? 3'b000 : 3'b010;
		assign node522 = (inp[3]) ? node900 : node523;
			assign node523 = (inp[0]) ? node639 : node524;
				assign node524 = (inp[7]) ? node534 : node525;
					assign node525 = (inp[5]) ? node527 : 3'b001;
						assign node527 = (inp[8]) ? 3'b001 : node528;
							assign node528 = (inp[10]) ? node530 : 3'b000;
								assign node530 = (inp[9]) ? 3'b000 : 3'b001;
					assign node534 = (inp[8]) ? node586 : node535;
						assign node535 = (inp[5]) ? 3'b000 : node536;
							assign node536 = (inp[9]) ? node544 : node537;
								assign node537 = (inp[10]) ? node539 : 3'b111;
									assign node539 = (inp[1]) ? node541 : 3'b111;
										assign node541 = (inp[11]) ? 3'b011 : 3'b111;
								assign node544 = (inp[4]) ? node566 : node545;
									assign node545 = (inp[11]) ? node561 : node546;
										assign node546 = (inp[2]) ? node554 : node547;
											assign node547 = (inp[1]) ? node551 : node548;
												assign node548 = (inp[10]) ? 3'b111 : 3'b011;
												assign node551 = (inp[10]) ? 3'b011 : 3'b111;
											assign node554 = (inp[10]) ? node558 : node555;
												assign node555 = (inp[1]) ? 3'b111 : 3'b011;
												assign node558 = (inp[1]) ? 3'b011 : 3'b111;
										assign node561 = (inp[10]) ? node563 : 3'b111;
											assign node563 = (inp[1]) ? 3'b011 : 3'b111;
									assign node566 = (inp[11]) ? node578 : node567;
										assign node567 = (inp[10]) ? node575 : node568;
											assign node568 = (inp[2]) ? node572 : node569;
												assign node569 = (inp[1]) ? 3'b011 : 3'b111;
												assign node572 = (inp[1]) ? 3'b111 : 3'b011;
											assign node575 = (inp[1]) ? 3'b101 : 3'b111;
										assign node578 = (inp[10]) ? node582 : node579;
											assign node579 = (inp[1]) ? 3'b101 : 3'b011;
											assign node582 = (inp[1]) ? 3'b001 : 3'b101;
						assign node586 = (inp[9]) ? node596 : node587;
							assign node587 = (inp[11]) ? node589 : 3'b111;
								assign node589 = (inp[1]) ? node591 : 3'b111;
									assign node591 = (inp[5]) ? node593 : 3'b111;
										assign node593 = (inp[10]) ? 3'b011 : 3'b111;
							assign node596 = (inp[4]) ? node614 : node597;
								assign node597 = (inp[10]) ? node605 : node598;
									assign node598 = (inp[11]) ? 3'b111 : node599;
										assign node599 = (inp[1]) ? 3'b111 : node600;
											assign node600 = (inp[5]) ? 3'b011 : 3'b111;
									assign node605 = (inp[1]) ? node609 : node606;
										assign node606 = (inp[5]) ? 3'b111 : 3'b011;
										assign node609 = (inp[11]) ? 3'b011 : node610;
											assign node610 = (inp[5]) ? 3'b011 : 3'b111;
								assign node614 = (inp[1]) ? node626 : node615;
									assign node615 = (inp[10]) ? node619 : node616;
										assign node616 = (inp[5]) ? 3'b011 : 3'b111;
										assign node619 = (inp[5]) ? node621 : 3'b011;
											assign node621 = (inp[11]) ? 3'b101 : node622;
												assign node622 = (inp[2]) ? 3'b111 : 3'b011;
									assign node626 = (inp[10]) ? node634 : node627;
										assign node627 = (inp[5]) ? node631 : node628;
											assign node628 = (inp[2]) ? 3'b001 : 3'b011;
											assign node631 = (inp[11]) ? 3'b101 : 3'b111;
										assign node634 = (inp[11]) ? node636 : 3'b101;
											assign node636 = (inp[5]) ? 3'b001 : 3'b101;
				assign node639 = (inp[10]) ? node787 : node640;
					assign node640 = (inp[4]) ? node704 : node641;
						assign node641 = (inp[8]) ? node675 : node642;
							assign node642 = (inp[7]) ? node654 : node643;
								assign node643 = (inp[5]) ? node647 : node644;
									assign node644 = (inp[11]) ? 3'b111 : 3'b011;
									assign node647 = (inp[9]) ? 3'b101 : node648;
										assign node648 = (inp[1]) ? node650 : 3'b001;
											assign node650 = (inp[11]) ? 3'b001 : 3'b101;
								assign node654 = (inp[9]) ? node666 : node655;
									assign node655 = (inp[1]) ? node661 : node656;
										assign node656 = (inp[11]) ? 3'b111 : node657;
											assign node657 = (inp[5]) ? 3'b011 : 3'b111;
										assign node661 = (inp[11]) ? 3'b011 : node662;
											assign node662 = (inp[5]) ? 3'b011 : 3'b111;
									assign node666 = (inp[1]) ? node670 : node667;
										assign node667 = (inp[11]) ? 3'b011 : 3'b111;
										assign node670 = (inp[5]) ? 3'b111 : node671;
											assign node671 = (inp[11]) ? 3'b110 : 3'b101;
							assign node675 = (inp[11]) ? node689 : node676;
								assign node676 = (inp[5]) ? node682 : node677;
									assign node677 = (inp[7]) ? node679 : 3'b111;
										assign node679 = (inp[1]) ? 3'b011 : 3'b111;
									assign node682 = (inp[7]) ? node684 : 3'b011;
										assign node684 = (inp[2]) ? node686 : 3'b011;
											assign node686 = (inp[9]) ? 3'b101 : 3'b111;
								assign node689 = (inp[7]) ? node691 : 3'b111;
									assign node691 = (inp[5]) ? node697 : node692;
										assign node692 = (inp[9]) ? 3'b111 : node693;
											assign node693 = (inp[1]) ? 3'b011 : 3'b111;
										assign node697 = (inp[1]) ? node701 : node698;
											assign node698 = (inp[9]) ? 3'b011 : 3'b111;
											assign node701 = (inp[9]) ? 3'b110 : 3'b011;
						assign node704 = (inp[11]) ? node748 : node705;
							assign node705 = (inp[7]) ? node717 : node706;
								assign node706 = (inp[5]) ? node710 : node707;
									assign node707 = (inp[8]) ? 3'b101 : 3'b001;
									assign node710 = (inp[8]) ? 3'b001 : node711;
										assign node711 = (inp[2]) ? 3'b110 : node712;
											assign node712 = (inp[9]) ? 3'b100 : 3'b000;
								assign node717 = (inp[8]) ? node735 : node718;
									assign node718 = (inp[2]) ? node730 : node719;
										assign node719 = (inp[5]) ? node725 : node720;
											assign node720 = (inp[9]) ? 3'b101 : node721;
												assign node721 = (inp[1]) ? 3'b101 : 3'b111;
											assign node725 = (inp[9]) ? 3'b111 : node726;
												assign node726 = (inp[1]) ? 3'b111 : 3'b011;
										assign node730 = (inp[5]) ? node732 : 3'b111;
											assign node732 = (inp[1]) ? 3'b101 : 3'b001;
									assign node735 = (inp[1]) ? node743 : node736;
										assign node736 = (inp[2]) ? 3'b101 : node737;
											assign node737 = (inp[5]) ? node739 : 3'b011;
												assign node739 = (inp[9]) ? 3'b101 : 3'b111;
										assign node743 = (inp[9]) ? 3'b001 : node744;
											assign node744 = (inp[5]) ? 3'b101 : 3'b011;
							assign node748 = (inp[7]) ? node760 : node749;
								assign node749 = (inp[8]) ? node757 : node750;
									assign node750 = (inp[5]) ? node752 : 3'b011;
										assign node752 = (inp[1]) ? 3'b110 : node753;
											assign node753 = (inp[9]) ? 3'b110 : 3'b010;
									assign node757 = (inp[5]) ? 3'b011 : 3'b111;
								assign node760 = (inp[5]) ? node774 : node761;
									assign node761 = (inp[9]) ? node769 : node762;
										assign node762 = (inp[1]) ? node766 : node763;
											assign node763 = (inp[8]) ? 3'b111 : 3'b011;
											assign node766 = (inp[8]) ? 3'b011 : 3'b101;
										assign node769 = (inp[1]) ? 3'b110 : node770;
											assign node770 = (inp[8]) ? 3'b101 : 3'b001;
									assign node774 = (inp[8]) ? node780 : node775;
										assign node775 = (inp[9]) ? 3'b101 : node776;
											assign node776 = (inp[2]) ? 3'b001 : 3'b101;
										assign node780 = (inp[1]) ? node784 : node781;
											assign node781 = (inp[9]) ? 3'b001 : 3'b011;
											assign node784 = (inp[9]) ? 3'b110 : 3'b101;
					assign node787 = (inp[7]) ? node817 : node788;
						assign node788 = (inp[11]) ? node800 : node789;
							assign node789 = (inp[4]) ? 3'b110 : node790;
								assign node790 = (inp[8]) ? 3'b110 : node791;
									assign node791 = (inp[5]) ? node793 : 3'b110;
										assign node793 = (inp[1]) ? node795 : 3'b100;
											assign node795 = (inp[9]) ? 3'b100 : 3'b000;
							assign node800 = (inp[4]) ? node812 : node801;
								assign node801 = (inp[8]) ? node809 : node802;
									assign node802 = (inp[5]) ? node804 : 3'b010;
										assign node804 = (inp[9]) ? 3'b100 : node805;
											assign node805 = (inp[1]) ? 3'b000 : 3'b100;
									assign node809 = (inp[5]) ? 3'b010 : 3'b110;
								assign node812 = (inp[5]) ? node814 : 3'b100;
									assign node814 = (inp[8]) ? 3'b100 : 3'b110;
						assign node817 = (inp[8]) ? node859 : node818;
							assign node818 = (inp[5]) ? node848 : node819;
								assign node819 = (inp[9]) ? node835 : node820;
									assign node820 = (inp[11]) ? node828 : node821;
										assign node821 = (inp[1]) ? node825 : node822;
											assign node822 = (inp[4]) ? 3'b011 : 3'b111;
											assign node825 = (inp[4]) ? 3'b001 : 3'b011;
										assign node828 = (inp[4]) ? node832 : node829;
											assign node829 = (inp[1]) ? 3'b101 : 3'b111;
											assign node832 = (inp[1]) ? 3'b001 : 3'b101;
									assign node835 = (inp[1]) ? node843 : node836;
										assign node836 = (inp[11]) ? node840 : node837;
											assign node837 = (inp[4]) ? 3'b001 : 3'b101;
											assign node840 = (inp[4]) ? 3'b110 : 3'b101;
										assign node843 = (inp[11]) ? node845 : 3'b110;
											assign node845 = (inp[4]) ? 3'b010 : 3'b110;
								assign node848 = (inp[4]) ? node854 : node849;
									assign node849 = (inp[1]) ? node851 : 3'b110;
										assign node851 = (inp[9]) ? 3'b110 : 3'b010;
									assign node854 = (inp[9]) ? 3'b100 : node855;
										assign node855 = (inp[1]) ? 3'b000 : 3'b100;
							assign node859 = (inp[9]) ? node877 : node860;
								assign node860 = (inp[1]) ? node870 : node861;
									assign node861 = (inp[4]) ? node863 : 3'b111;
										assign node863 = (inp[11]) ? node867 : node864;
											assign node864 = (inp[5]) ? 3'b011 : 3'b111;
											assign node867 = (inp[5]) ? 3'b101 : 3'b011;
									assign node870 = (inp[5]) ? node872 : 3'b101;
										assign node872 = (inp[4]) ? 3'b001 : node873;
											assign node873 = (inp[11]) ? 3'b101 : 3'b011;
								assign node877 = (inp[1]) ? node889 : node878;
									assign node878 = (inp[5]) ? node884 : node879;
										assign node879 = (inp[4]) ? node881 : 3'b011;
											assign node881 = (inp[11]) ? 3'b001 : 3'b101;
										assign node884 = (inp[4]) ? node886 : 3'b101;
											assign node886 = (inp[11]) ? 3'b110 : 3'b001;
									assign node889 = (inp[5]) ? node895 : node890;
										assign node890 = (inp[4]) ? node892 : 3'b001;
											assign node892 = (inp[11]) ? 3'b110 : 3'b100;
										assign node895 = (inp[4]) ? node897 : 3'b110;
											assign node897 = (inp[11]) ? 3'b010 : 3'b110;
			assign node900 = (inp[7]) ? node1152 : node901;
				assign node901 = (inp[9]) ? node1065 : node902;
					assign node902 = (inp[10]) ? node1004 : node903;
						assign node903 = (inp[4]) ? node947 : node904;
							assign node904 = (inp[1]) ? node926 : node905;
								assign node905 = (inp[8]) ? node917 : node906;
									assign node906 = (inp[5]) ? node912 : node907;
										assign node907 = (inp[0]) ? 3'b010 : node908;
											assign node908 = (inp[11]) ? 3'b010 : 3'b110;
										assign node912 = (inp[0]) ? node914 : 3'b000;
											assign node914 = (inp[2]) ? 3'b100 : 3'b110;
									assign node917 = (inp[5]) ? node921 : node918;
										assign node918 = (inp[0]) ? 3'b100 : 3'b000;
										assign node921 = (inp[0]) ? 3'b010 : node922;
											assign node922 = (inp[11]) ? 3'b010 : 3'b110;
								assign node926 = (inp[11]) ? node932 : node927;
									assign node927 = (inp[5]) ? node929 : 3'b110;
										assign node929 = (inp[8]) ? 3'b110 : 3'b010;
									assign node932 = (inp[0]) ? node940 : node933;
										assign node933 = (inp[5]) ? node937 : node934;
											assign node934 = (inp[8]) ? 3'b000 : 3'b010;
											assign node937 = (inp[8]) ? 3'b010 : 3'b000;
										assign node940 = (inp[8]) ? node944 : node941;
											assign node941 = (inp[5]) ? 3'b100 : 3'b010;
											assign node944 = (inp[5]) ? 3'b010 : 3'b110;
							assign node947 = (inp[0]) ? node973 : node948;
								assign node948 = (inp[11]) ? node960 : node949;
									assign node949 = (inp[2]) ? 3'b110 : node950;
										assign node950 = (inp[1]) ? 3'b000 : node951;
											assign node951 = (inp[5]) ? node955 : node952;
												assign node952 = (inp[8]) ? 3'b000 : 3'b110;
												assign node955 = (inp[8]) ? 3'b110 : 3'b000;
									assign node960 = (inp[1]) ? node968 : node961;
										assign node961 = (inp[5]) ? node965 : node962;
											assign node962 = (inp[8]) ? 3'b000 : 3'b010;
											assign node965 = (inp[8]) ? 3'b010 : 3'b000;
										assign node968 = (inp[5]) ? 3'b010 : node969;
											assign node969 = (inp[8]) ? 3'b000 : 3'b010;
								assign node973 = (inp[11]) ? node989 : node974;
									assign node974 = (inp[8]) ? node984 : node975;
										assign node975 = (inp[1]) ? node979 : node976;
											assign node976 = (inp[5]) ? 3'b100 : 3'b010;
											assign node979 = (inp[5]) ? 3'b000 : node980;
												assign node980 = (inp[2]) ? 3'b100 : 3'b000;
										assign node984 = (inp[5]) ? 3'b010 : node985;
											assign node985 = (inp[1]) ? 3'b010 : 3'b000;
									assign node989 = (inp[1]) ? node995 : node990;
										assign node990 = (inp[8]) ? node992 : 3'b100;
											assign node992 = (inp[5]) ? 3'b010 : 3'b000;
										assign node995 = (inp[2]) ? 3'b100 : node996;
											assign node996 = (inp[5]) ? node1000 : node997;
												assign node997 = (inp[8]) ? 3'b000 : 3'b100;
												assign node1000 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1004 = (inp[5]) ? node1034 : node1005;
							assign node1005 = (inp[8]) ? node1021 : node1006;
								assign node1006 = (inp[11]) ? node1016 : node1007;
									assign node1007 = (inp[0]) ? node1009 : 3'b010;
										assign node1009 = (inp[1]) ? node1011 : 3'b100;
											assign node1011 = (inp[4]) ? node1013 : 3'b010;
												assign node1013 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1016 = (inp[1]) ? node1018 : 3'b100;
										assign node1018 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1021 = (inp[4]) ? node1027 : node1022;
									assign node1022 = (inp[0]) ? node1024 : 3'b000;
										assign node1024 = (inp[1]) ? 3'b010 : 3'b000;
									assign node1027 = (inp[2]) ? node1029 : 3'b000;
										assign node1029 = (inp[0]) ? node1031 : 3'b000;
											assign node1031 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1034 = (inp[0]) ? node1048 : node1035;
								assign node1035 = (inp[11]) ? node1043 : node1036;
									assign node1036 = (inp[8]) ? 3'b010 : node1037;
										assign node1037 = (inp[1]) ? node1039 : 3'b110;
											assign node1039 = (inp[2]) ? 3'b100 : 3'b110;
									assign node1043 = (inp[8]) ? 3'b100 : node1044;
										assign node1044 = (inp[1]) ? 3'b100 : 3'b110;
								assign node1048 = (inp[4]) ? node1058 : node1049;
									assign node1049 = (inp[8]) ? node1053 : node1050;
										assign node1050 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1053 = (inp[1]) ? node1055 : 3'b100;
											assign node1055 = (inp[2]) ? 3'b000 : 3'b010;
									assign node1058 = (inp[8]) ? node1060 : 3'b000;
										assign node1060 = (inp[2]) ? 3'b000 : node1061;
											assign node1061 = (inp[11]) ? 3'b000 : 3'b100;
					assign node1065 = (inp[0]) ? node1125 : node1066;
						assign node1066 = (inp[10]) ? node1112 : node1067;
							assign node1067 = (inp[11]) ? node1075 : node1068;
								assign node1068 = (inp[8]) ? node1072 : node1069;
									assign node1069 = (inp[5]) ? 3'b000 : 3'b110;
									assign node1072 = (inp[5]) ? 3'b110 : 3'b000;
								assign node1075 = (inp[2]) ? node1097 : node1076;
									assign node1076 = (inp[4]) ? node1090 : node1077;
										assign node1077 = (inp[1]) ? node1083 : node1078;
											assign node1078 = (inp[8]) ? 3'b000 : node1079;
												assign node1079 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1083 = (inp[8]) ? node1087 : node1084;
												assign node1084 = (inp[5]) ? 3'b000 : 3'b010;
												assign node1087 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1090 = (inp[5]) ? node1094 : node1091;
											assign node1091 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1094 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1097 = (inp[4]) ? node1105 : node1098;
										assign node1098 = (inp[8]) ? node1102 : node1099;
											assign node1099 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1102 = (inp[1]) ? 3'b010 : 3'b000;
										assign node1105 = (inp[5]) ? node1109 : node1106;
											assign node1106 = (inp[8]) ? 3'b000 : 3'b010;
											assign node1109 = (inp[8]) ? 3'b010 : 3'b000;
							assign node1112 = (inp[11]) ? node1120 : node1113;
								assign node1113 = (inp[5]) ? node1117 : node1114;
									assign node1114 = (inp[8]) ? 3'b000 : 3'b010;
									assign node1117 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1120 = (inp[8]) ? node1122 : 3'b100;
									assign node1122 = (inp[5]) ? 3'b100 : 3'b000;
						assign node1125 = (inp[8]) ? node1135 : node1126;
							assign node1126 = (inp[10]) ? 3'b000 : node1127;
								assign node1127 = (inp[4]) ? 3'b000 : node1128;
									assign node1128 = (inp[5]) ? node1130 : 3'b000;
										assign node1130 = (inp[11]) ? 3'b000 : 3'b010;
							assign node1135 = (inp[5]) ? 3'b000 : node1136;
								assign node1136 = (inp[10]) ? node1144 : node1137;
									assign node1137 = (inp[4]) ? node1139 : 3'b100;
										assign node1139 = (inp[2]) ? node1141 : 3'b000;
											assign node1141 = (inp[1]) ? 3'b100 : 3'b000;
									assign node1144 = (inp[11]) ? 3'b000 : node1145;
										assign node1145 = (inp[2]) ? node1147 : 3'b000;
											assign node1147 = (inp[4]) ? 3'b100 : 3'b000;
				assign node1152 = (inp[9]) ? node1338 : node1153;
					assign node1153 = (inp[8]) ? node1239 : node1154;
						assign node1154 = (inp[5]) ? node1204 : node1155;
							assign node1155 = (inp[0]) ? node1179 : node1156;
								assign node1156 = (inp[4]) ? node1164 : node1157;
									assign node1157 = (inp[1]) ? node1161 : node1158;
										assign node1158 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1161 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1164 = (inp[1]) ? node1172 : node1165;
										assign node1165 = (inp[11]) ? node1169 : node1166;
											assign node1166 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1169 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1172 = (inp[10]) ? node1174 : 3'b001;
											assign node1174 = (inp[2]) ? 3'b110 : node1175;
												assign node1175 = (inp[11]) ? 3'b110 : 3'b001;
								assign node1179 = (inp[4]) ? node1187 : node1180;
									assign node1180 = (inp[1]) ? node1184 : node1181;
										assign node1181 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1184 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1187 = (inp[1]) ? node1195 : node1188;
										assign node1188 = (inp[10]) ? 3'b010 : node1189;
											assign node1189 = (inp[11]) ? 3'b110 : node1190;
												assign node1190 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1195 = (inp[10]) ? node1201 : node1196;
											assign node1196 = (inp[2]) ? node1198 : 3'b110;
												assign node1198 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1201 = (inp[11]) ? 3'b100 : 3'b110;
							assign node1204 = (inp[1]) ? node1216 : node1205;
								assign node1205 = (inp[0]) ? node1211 : node1206;
									assign node1206 = (inp[11]) ? 3'b110 : node1207;
										assign node1207 = (inp[10]) ? 3'b110 : 3'b000;
									assign node1211 = (inp[10]) ? 3'b010 : node1212;
										assign node1212 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1216 = (inp[0]) ? node1226 : node1217;
									assign node1217 = (inp[11]) ? node1223 : node1218;
										assign node1218 = (inp[10]) ? node1220 : 3'b001;
											assign node1220 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1223 = (inp[4]) ? 3'b110 : 3'b111;
									assign node1226 = (inp[4]) ? node1228 : 3'b110;
										assign node1228 = (inp[10]) ? node1234 : node1229;
											assign node1229 = (inp[11]) ? node1231 : 3'b010;
												assign node1231 = (inp[2]) ? 3'b100 : 3'b010;
											assign node1234 = (inp[2]) ? node1236 : 3'b100;
												assign node1236 = (inp[11]) ? 3'b000 : 3'b100;
						assign node1239 = (inp[0]) ? node1289 : node1240;
							assign node1240 = (inp[4]) ? node1260 : node1241;
								assign node1241 = (inp[10]) ? node1249 : node1242;
									assign node1242 = (inp[1]) ? node1244 : 3'b111;
										assign node1244 = (inp[5]) ? 3'b011 : node1245;
											assign node1245 = (inp[11]) ? 3'b011 : 3'b111;
									assign node1249 = (inp[1]) ? node1255 : node1250;
										assign node1250 = (inp[5]) ? 3'b011 : node1251;
											assign node1251 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1255 = (inp[5]) ? 3'b101 : node1256;
											assign node1256 = (inp[11]) ? 3'b101 : 3'b011;
								assign node1260 = (inp[10]) ? node1274 : node1261;
									assign node1261 = (inp[5]) ? node1267 : node1262;
										assign node1262 = (inp[11]) ? node1264 : 3'b011;
											assign node1264 = (inp[1]) ? 3'b111 : 3'b001;
										assign node1267 = (inp[1]) ? node1269 : 3'b101;
											assign node1269 = (inp[2]) ? 3'b001 : node1270;
												assign node1270 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1274 = (inp[5]) ? node1280 : node1275;
										assign node1275 = (inp[11]) ? node1277 : 3'b101;
											assign node1277 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1280 = (inp[1]) ? node1284 : node1281;
											assign node1281 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1284 = (inp[11]) ? 3'b110 : node1285;
												assign node1285 = (inp[2]) ? 3'b110 : 3'b001;
							assign node1289 = (inp[4]) ? node1305 : node1290;
								assign node1290 = (inp[10]) ? node1300 : node1291;
									assign node1291 = (inp[1]) ? node1295 : node1292;
										assign node1292 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1295 = (inp[5]) ? 3'b001 : node1296;
											assign node1296 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1300 = (inp[1]) ? 3'b110 : node1301;
										assign node1301 = (inp[5]) ? 3'b001 : 3'b101;
								assign node1305 = (inp[1]) ? node1325 : node1306;
									assign node1306 = (inp[5]) ? node1316 : node1307;
										assign node1307 = (inp[10]) ? node1313 : node1308;
											assign node1308 = (inp[2]) ? 3'b001 : node1309;
												assign node1309 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1313 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1316 = (inp[2]) ? node1322 : node1317;
											assign node1317 = (inp[10]) ? 3'b110 : node1318;
												assign node1318 = (inp[11]) ? 3'b110 : 3'b001;
											assign node1322 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1325 = (inp[10]) ? node1333 : node1326;
										assign node1326 = (inp[11]) ? node1328 : 3'b110;
											assign node1328 = (inp[2]) ? node1330 : 3'b110;
												assign node1330 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1333 = (inp[5]) ? node1335 : 3'b010;
											assign node1335 = (inp[11]) ? 3'b100 : 3'b110;
					assign node1338 = (inp[0]) ? node1450 : node1339;
						assign node1339 = (inp[4]) ? node1373 : node1340;
							assign node1340 = (inp[5]) ? node1360 : node1341;
								assign node1341 = (inp[1]) ? node1351 : node1342;
									assign node1342 = (inp[8]) ? node1346 : node1343;
										assign node1343 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1346 = (inp[11]) ? 3'b101 : node1347;
											assign node1347 = (inp[10]) ? 3'b101 : 3'b011;
									assign node1351 = (inp[10]) ? node1357 : node1352;
										assign node1352 = (inp[8]) ? node1354 : 3'b001;
											assign node1354 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1357 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1360 = (inp[8]) ? node1366 : node1361;
									assign node1361 = (inp[11]) ? 3'b110 : node1362;
										assign node1362 = (inp[10]) ? 3'b110 : 3'b000;
									assign node1366 = (inp[1]) ? node1370 : node1367;
										assign node1367 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1370 = (inp[10]) ? 3'b110 : 3'b001;
							assign node1373 = (inp[10]) ? node1419 : node1374;
								assign node1374 = (inp[11]) ? node1398 : node1375;
									assign node1375 = (inp[2]) ? node1387 : node1376;
										assign node1376 = (inp[1]) ? node1382 : node1377;
											assign node1377 = (inp[5]) ? node1379 : 3'b001;
												assign node1379 = (inp[8]) ? 3'b001 : 3'b000;
											assign node1382 = (inp[8]) ? node1384 : 3'b110;
												assign node1384 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1387 = (inp[8]) ? node1393 : node1388;
											assign node1388 = (inp[5]) ? 3'b000 : node1389;
												assign node1389 = (inp[1]) ? 3'b010 : 3'b110;
											assign node1393 = (inp[5]) ? node1395 : 3'b101;
												assign node1395 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1398 = (inp[1]) ? node1406 : node1399;
										assign node1399 = (inp[2]) ? node1401 : 3'b110;
											assign node1401 = (inp[8]) ? node1403 : 3'b110;
												assign node1403 = (inp[5]) ? 3'b110 : 3'b000;
										assign node1406 = (inp[2]) ? node1412 : node1407;
											assign node1407 = (inp[5]) ? 3'b010 : node1408;
												assign node1408 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1412 = (inp[5]) ? node1416 : node1413;
												assign node1413 = (inp[8]) ? 3'b110 : 3'b010;
												assign node1416 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1419 = (inp[11]) ? node1435 : node1420;
									assign node1420 = (inp[1]) ? node1422 : 3'b110;
										assign node1422 = (inp[8]) ? node1428 : node1423;
											assign node1423 = (inp[2]) ? 3'b110 : node1424;
												assign node1424 = (inp[5]) ? 3'b110 : 3'b010;
											assign node1428 = (inp[5]) ? node1432 : node1429;
												assign node1429 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1432 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1435 = (inp[1]) ? node1443 : node1436;
										assign node1436 = (inp[8]) ? node1440 : node1437;
											assign node1437 = (inp[5]) ? 3'b110 : 3'b010;
											assign node1440 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1443 = (inp[5]) ? node1447 : node1444;
											assign node1444 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1447 = (inp[8]) ? 3'b100 : 3'b110;
						assign node1450 = (inp[4]) ? node1480 : node1451;
							assign node1451 = (inp[8]) ? node1461 : node1452;
								assign node1452 = (inp[5]) ? 3'b000 : node1453;
									assign node1453 = (inp[10]) ? node1457 : node1454;
										assign node1454 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1457 = (inp[1]) ? 3'b100 : 3'b010;
								assign node1461 = (inp[5]) ? node1473 : node1462;
									assign node1462 = (inp[10]) ? node1468 : node1463;
										assign node1463 = (inp[1]) ? node1465 : 3'b001;
											assign node1465 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1468 = (inp[1]) ? node1470 : 3'b110;
											assign node1470 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1473 = (inp[1]) ? node1477 : node1474;
										assign node1474 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1477 = (inp[10]) ? 3'b100 : 3'b010;
							assign node1480 = (inp[1]) ? node1510 : node1481;
								assign node1481 = (inp[8]) ? node1489 : node1482;
									assign node1482 = (inp[5]) ? 3'b000 : node1483;
										assign node1483 = (inp[10]) ? node1485 : 3'b100;
											assign node1485 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1489 = (inp[5]) ? node1501 : node1490;
										assign node1490 = (inp[10]) ? node1498 : node1491;
											assign node1491 = (inp[11]) ? node1495 : node1492;
												assign node1492 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1495 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1498 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1501 = (inp[10]) ? node1507 : node1502;
											assign node1502 = (inp[2]) ? 3'b100 : node1503;
												assign node1503 = (inp[11]) ? 3'b100 : 3'b010;
											assign node1507 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1510 = (inp[10]) ? 3'b000 : node1511;
									assign node1511 = (inp[5]) ? node1517 : node1512;
										assign node1512 = (inp[8]) ? 3'b100 : node1513;
											assign node1513 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1517 = (inp[11]) ? 3'b000 : node1518;
											assign node1518 = (inp[2]) ? node1520 : 3'b000;
												assign node1520 = (inp[8]) ? 3'b100 : 3'b000;

endmodule