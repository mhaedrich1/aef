module dtc_split33_bm72 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node763;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node789;
	wire [3-1:0] node792;
	wire [3-1:0] node793;

	assign outp = (inp[3]) ? node432 : node1;
		assign node1 = (inp[6]) ? node223 : node2;
			assign node2 = (inp[9]) ? node120 : node3;
				assign node3 = (inp[0]) ? node65 : node4;
					assign node4 = (inp[4]) ? node34 : node5;
						assign node5 = (inp[7]) ? node21 : node6;
							assign node6 = (inp[5]) ? node14 : node7;
								assign node7 = (inp[10]) ? node11 : node8;
									assign node8 = (inp[8]) ? 3'b011 : 3'b101;
									assign node11 = (inp[8]) ? 3'b101 : 3'b001;
								assign node14 = (inp[10]) ? node18 : node15;
									assign node15 = (inp[1]) ? 3'b001 : 3'b101;
									assign node18 = (inp[1]) ? 3'b110 : 3'b001;
							assign node21 = (inp[10]) ? node27 : node22;
								assign node22 = (inp[8]) ? node24 : 3'b011;
									assign node24 = (inp[1]) ? 3'b011 : 3'b111;
								assign node27 = (inp[8]) ? node31 : node28;
									assign node28 = (inp[5]) ? 3'b101 : 3'b001;
									assign node31 = (inp[1]) ? 3'b001 : 3'b011;
						assign node34 = (inp[1]) ? node50 : node35;
							assign node35 = (inp[7]) ? node43 : node36;
								assign node36 = (inp[8]) ? node40 : node37;
									assign node37 = (inp[5]) ? 3'b110 : 3'b010;
									assign node40 = (inp[5]) ? 3'b001 : 3'b001;
								assign node43 = (inp[2]) ? node47 : node44;
									assign node44 = (inp[8]) ? 3'b011 : 3'b001;
									assign node47 = (inp[11]) ? 3'b101 : 3'b001;
							assign node50 = (inp[5]) ? node58 : node51;
								assign node51 = (inp[10]) ? node55 : node52;
									assign node52 = (inp[7]) ? 3'b001 : 3'b110;
									assign node55 = (inp[8]) ? 3'b110 : 3'b010;
								assign node58 = (inp[10]) ? node62 : node59;
									assign node59 = (inp[11]) ? 3'b110 : 3'b010;
									assign node62 = (inp[7]) ? 3'b110 : 3'b100;
					assign node65 = (inp[7]) ? node93 : node66;
						assign node66 = (inp[10]) ? node80 : node67;
							assign node67 = (inp[1]) ? node73 : node68;
								assign node68 = (inp[4]) ? node70 : 3'b001;
									assign node70 = (inp[11]) ? 3'b010 : 3'b110;
								assign node73 = (inp[2]) ? node77 : node74;
									assign node74 = (inp[11]) ? 3'b100 : 3'b010;
									assign node77 = (inp[4]) ? 3'b100 : 3'b110;
							assign node80 = (inp[4]) ? node86 : node81;
								assign node81 = (inp[11]) ? node83 : 3'b010;
									assign node83 = (inp[2]) ? 3'b010 : 3'b010;
								assign node86 = (inp[8]) ? node90 : node87;
									assign node87 = (inp[5]) ? 3'b000 : 3'b000;
									assign node90 = (inp[1]) ? 3'b100 : 3'b000;
						assign node93 = (inp[4]) ? node105 : node94;
							assign node94 = (inp[8]) ? node100 : node95;
								assign node95 = (inp[11]) ? node97 : 3'b001;
									assign node97 = (inp[2]) ? 3'b110 : 3'b010;
								assign node100 = (inp[1]) ? node102 : 3'b101;
									assign node102 = (inp[2]) ? 3'b101 : 3'b001;
							assign node105 = (inp[5]) ? node113 : node106;
								assign node106 = (inp[10]) ? node110 : node107;
									assign node107 = (inp[1]) ? 3'b010 : 3'b001;
									assign node110 = (inp[8]) ? 3'b000 : 3'b110;
								assign node113 = (inp[11]) ? node117 : node114;
									assign node114 = (inp[10]) ? 3'b010 : 3'b110;
									assign node117 = (inp[8]) ? 3'b110 : 3'b100;
				assign node120 = (inp[7]) ? node168 : node121;
					assign node121 = (inp[1]) ? node145 : node122;
						assign node122 = (inp[0]) ? node136 : node123;
							assign node123 = (inp[5]) ? node131 : node124;
								assign node124 = (inp[4]) ? node128 : node125;
									assign node125 = (inp[2]) ? 3'b010 : 3'b001;
									assign node128 = (inp[2]) ? 3'b000 : 3'b010;
								assign node131 = (inp[8]) ? node133 : 3'b100;
									assign node133 = (inp[2]) ? 3'b010 : 3'b010;
							assign node136 = (inp[8]) ? node140 : node137;
								assign node137 = (inp[11]) ? 3'b000 : 3'b010;
								assign node140 = (inp[2]) ? node142 : 3'b100;
									assign node142 = (inp[11]) ? 3'b000 : 3'b100;
						assign node145 = (inp[0]) ? node161 : node146;
							assign node146 = (inp[8]) ? node154 : node147;
								assign node147 = (inp[5]) ? node151 : node148;
									assign node148 = (inp[11]) ? 3'b100 : 3'b100;
									assign node151 = (inp[4]) ? 3'b000 : 3'b100;
								assign node154 = (inp[5]) ? node158 : node155;
									assign node155 = (inp[2]) ? 3'b010 : 3'b000;
									assign node158 = (inp[4]) ? 3'b100 : 3'b000;
							assign node161 = (inp[10]) ? 3'b000 : node162;
								assign node162 = (inp[4]) ? 3'b000 : node163;
									assign node163 = (inp[2]) ? 3'b000 : 3'b100;
					assign node168 = (inp[4]) ? node194 : node169;
						assign node169 = (inp[0]) ? node183 : node170;
							assign node170 = (inp[1]) ? node176 : node171;
								assign node171 = (inp[10]) ? 3'b001 : node172;
									assign node172 = (inp[8]) ? 3'b101 : 3'b001;
								assign node176 = (inp[2]) ? node180 : node177;
									assign node177 = (inp[8]) ? 3'b001 : 3'b110;
									assign node180 = (inp[8]) ? 3'b110 : 3'b010;
							assign node183 = (inp[1]) ? node189 : node184;
								assign node184 = (inp[5]) ? node186 : 3'b110;
									assign node186 = (inp[11]) ? 3'b010 : 3'b010;
								assign node189 = (inp[5]) ? node191 : 3'b010;
									assign node191 = (inp[11]) ? 3'b100 : 3'b010;
						assign node194 = (inp[0]) ? node210 : node195;
							assign node195 = (inp[10]) ? node203 : node196;
								assign node196 = (inp[1]) ? node200 : node197;
									assign node197 = (inp[2]) ? 3'b110 : 3'b001;
									assign node200 = (inp[2]) ? 3'b010 : 3'b110;
								assign node203 = (inp[5]) ? node207 : node204;
									assign node204 = (inp[2]) ? 3'b010 : 3'b010;
									assign node207 = (inp[1]) ? 3'b100 : 3'b010;
							assign node210 = (inp[2]) ? node218 : node211;
								assign node211 = (inp[10]) ? node215 : node212;
									assign node212 = (inp[1]) ? 3'b100 : 3'b010;
									assign node215 = (inp[5]) ? 3'b000 : 3'b100;
								assign node218 = (inp[1]) ? 3'b000 : node219;
									assign node219 = (inp[8]) ? 3'b010 : 3'b000;
			assign node223 = (inp[9]) ? node319 : node224;
				assign node224 = (inp[0]) ? node258 : node225;
					assign node225 = (inp[7]) ? node247 : node226;
						assign node226 = (inp[4]) ? node234 : node227;
							assign node227 = (inp[10]) ? node229 : 3'b111;
								assign node229 = (inp[1]) ? node231 : 3'b111;
									assign node231 = (inp[5]) ? 3'b011 : 3'b011;
							assign node234 = (inp[10]) ? node242 : node235;
								assign node235 = (inp[2]) ? node239 : node236;
									assign node236 = (inp[1]) ? 3'b011 : 3'b111;
									assign node239 = (inp[8]) ? 3'b111 : 3'b101;
								assign node242 = (inp[5]) ? 3'b101 : node243;
									assign node243 = (inp[11]) ? 3'b001 : 3'b011;
						assign node247 = (inp[4]) ? node249 : 3'b111;
							assign node249 = (inp[10]) ? node251 : 3'b111;
								assign node251 = (inp[1]) ? node255 : node252;
									assign node252 = (inp[11]) ? 3'b111 : 3'b111;
									assign node255 = (inp[2]) ? 3'b011 : 3'b111;
					assign node258 = (inp[7]) ? node290 : node259;
						assign node259 = (inp[11]) ? node275 : node260;
							assign node260 = (inp[4]) ? node268 : node261;
								assign node261 = (inp[10]) ? node265 : node262;
									assign node262 = (inp[2]) ? 3'b011 : 3'b011;
									assign node265 = (inp[2]) ? 3'b101 : 3'b011;
								assign node268 = (inp[10]) ? node272 : node269;
									assign node269 = (inp[8]) ? 3'b101 : 3'b001;
									assign node272 = (inp[1]) ? 3'b000 : 3'b001;
							assign node275 = (inp[4]) ? node283 : node276;
								assign node276 = (inp[5]) ? node280 : node277;
									assign node277 = (inp[8]) ? 3'b011 : 3'b101;
									assign node280 = (inp[10]) ? 3'b101 : 3'b101;
								assign node283 = (inp[10]) ? node287 : node284;
									assign node284 = (inp[2]) ? 3'b001 : 3'b001;
									assign node287 = (inp[2]) ? 3'b110 : 3'b001;
						assign node290 = (inp[4]) ? node304 : node291;
							assign node291 = (inp[8]) ? node299 : node292;
								assign node292 = (inp[10]) ? node296 : node293;
									assign node293 = (inp[11]) ? 3'b011 : 3'b111;
									assign node296 = (inp[5]) ? 3'b011 : 3'b011;
								assign node299 = (inp[5]) ? node301 : 3'b111;
									assign node301 = (inp[11]) ? 3'b001 : 3'b111;
							assign node304 = (inp[1]) ? node312 : node305;
								assign node305 = (inp[10]) ? node309 : node306;
									assign node306 = (inp[8]) ? 3'b111 : 3'b011;
									assign node309 = (inp[5]) ? 3'b101 : 3'b011;
								assign node312 = (inp[5]) ? node316 : node313;
									assign node313 = (inp[8]) ? 3'b001 : 3'b101;
									assign node316 = (inp[10]) ? 3'b001 : 3'b101;
				assign node319 = (inp[0]) ? node375 : node320;
					assign node320 = (inp[4]) ? node344 : node321;
						assign node321 = (inp[7]) ? node333 : node322;
							assign node322 = (inp[2]) ? node328 : node323;
								assign node323 = (inp[5]) ? 3'b101 : node324;
									assign node324 = (inp[1]) ? 3'b001 : 3'b011;
								assign node328 = (inp[10]) ? node330 : 3'b101;
									assign node330 = (inp[1]) ? 3'b110 : 3'b101;
							assign node333 = (inp[10]) ? node339 : node334;
								assign node334 = (inp[5]) ? node336 : 3'b111;
									assign node336 = (inp[8]) ? 3'b111 : 3'b011;
								assign node339 = (inp[5]) ? 3'b101 : node340;
									assign node340 = (inp[11]) ? 3'b011 : 3'b111;
						assign node344 = (inp[10]) ? node360 : node345;
							assign node345 = (inp[7]) ? node353 : node346;
								assign node346 = (inp[8]) ? node350 : node347;
									assign node347 = (inp[2]) ? 3'b000 : 3'b001;
									assign node350 = (inp[5]) ? 3'b001 : 3'b101;
								assign node353 = (inp[2]) ? node357 : node354;
									assign node354 = (inp[11]) ? 3'b101 : 3'b111;
									assign node357 = (inp[8]) ? 3'b011 : 3'b101;
							assign node360 = (inp[7]) ? node368 : node361;
								assign node361 = (inp[1]) ? node365 : node362;
									assign node362 = (inp[8]) ? 3'b001 : 3'b110;
									assign node365 = (inp[5]) ? 3'b010 : 3'b110;
								assign node368 = (inp[8]) ? node372 : node369;
									assign node369 = (inp[1]) ? 3'b001 : 3'b101;
									assign node372 = (inp[1]) ? 3'b001 : 3'b011;
					assign node375 = (inp[4]) ? node405 : node376;
						assign node376 = (inp[7]) ? node392 : node377;
							assign node377 = (inp[10]) ? node385 : node378;
								assign node378 = (inp[11]) ? node382 : node379;
									assign node379 = (inp[2]) ? 3'b001 : 3'b001;
									assign node382 = (inp[1]) ? 3'b010 : 3'b001;
								assign node385 = (inp[8]) ? node389 : node386;
									assign node386 = (inp[1]) ? 3'b010 : 3'b110;
									assign node389 = (inp[2]) ? 3'b110 : 3'b001;
							assign node392 = (inp[5]) ? node398 : node393;
								assign node393 = (inp[11]) ? node395 : 3'b011;
									assign node395 = (inp[10]) ? 3'b001 : 3'b011;
								assign node398 = (inp[2]) ? node402 : node399;
									assign node399 = (inp[1]) ? 3'b001 : 3'b101;
									assign node402 = (inp[10]) ? 3'b001 : 3'b001;
						assign node405 = (inp[10]) ? node421 : node406;
							assign node406 = (inp[7]) ? node414 : node407;
								assign node407 = (inp[2]) ? node411 : node408;
									assign node408 = (inp[5]) ? 3'b100 : 3'b110;
									assign node411 = (inp[8]) ? 3'b110 : 3'b010;
								assign node414 = (inp[11]) ? node418 : node415;
									assign node415 = (inp[1]) ? 3'b001 : 3'b001;
									assign node418 = (inp[2]) ? 3'b010 : 3'b001;
							assign node421 = (inp[7]) ? node425 : node422;
								assign node422 = (inp[1]) ? 3'b100 : 3'b010;
								assign node425 = (inp[1]) ? node429 : node426;
									assign node426 = (inp[5]) ? 3'b110 : 3'b101;
									assign node429 = (inp[2]) ? 3'b110 : 3'b010;
		assign node432 = (inp[6]) ? node574 : node433;
			assign node433 = (inp[4]) ? node525 : node434;
				assign node434 = (inp[0]) ? node494 : node435;
					assign node435 = (inp[9]) ? node467 : node436;
						assign node436 = (inp[10]) ? node452 : node437;
							assign node437 = (inp[7]) ? node445 : node438;
								assign node438 = (inp[2]) ? node442 : node439;
									assign node439 = (inp[1]) ? 3'b000 : 3'b010;
									assign node442 = (inp[11]) ? 3'b100 : 3'b010;
								assign node445 = (inp[11]) ? node449 : node446;
									assign node446 = (inp[1]) ? 3'b001 : 3'b001;
									assign node449 = (inp[1]) ? 3'b000 : 3'b001;
							assign node452 = (inp[1]) ? node460 : node453;
								assign node453 = (inp[2]) ? node457 : node454;
									assign node454 = (inp[8]) ? 3'b010 : 3'b100;
									assign node457 = (inp[7]) ? 3'b010 : 3'b010;
								assign node460 = (inp[7]) ? node464 : node461;
									assign node461 = (inp[11]) ? 3'b000 : 3'b100;
									assign node464 = (inp[8]) ? 3'b010 : 3'b100;
						assign node467 = (inp[7]) ? node479 : node468;
							assign node468 = (inp[11]) ? node474 : node469;
								assign node469 = (inp[8]) ? node471 : 3'b000;
									assign node471 = (inp[1]) ? 3'b000 : 3'b100;
								assign node474 = (inp[5]) ? 3'b000 : node475;
									assign node475 = (inp[2]) ? 3'b000 : 3'b100;
							assign node479 = (inp[1]) ? node487 : node480;
								assign node480 = (inp[8]) ? node484 : node481;
									assign node481 = (inp[11]) ? 3'b100 : 3'b000;
									assign node484 = (inp[5]) ? 3'b010 : 3'b010;
								assign node487 = (inp[10]) ? node491 : node488;
									assign node488 = (inp[2]) ? 3'b100 : 3'b000;
									assign node491 = (inp[5]) ? 3'b000 : 3'b100;
					assign node494 = (inp[10]) ? node514 : node495;
						assign node495 = (inp[1]) ? node507 : node496;
							assign node496 = (inp[7]) ? node502 : node497;
								assign node497 = (inp[9]) ? 3'b000 : node498;
									assign node498 = (inp[11]) ? 3'b100 : 3'b100;
								assign node502 = (inp[9]) ? 3'b100 : node503;
									assign node503 = (inp[11]) ? 3'b000 : 3'b010;
							assign node507 = (inp[9]) ? 3'b000 : node508;
								assign node508 = (inp[8]) ? 3'b100 : node509;
									assign node509 = (inp[11]) ? 3'b000 : 3'b000;
						assign node514 = (inp[7]) ? node516 : 3'b000;
							assign node516 = (inp[9]) ? 3'b000 : node517;
								assign node517 = (inp[11]) ? node521 : node518;
									assign node518 = (inp[5]) ? 3'b000 : 3'b100;
									assign node521 = (inp[1]) ? 3'b000 : 3'b000;
				assign node525 = (inp[9]) ? node563 : node526;
					assign node526 = (inp[0]) ? node554 : node527;
						assign node527 = (inp[7]) ? node539 : node528;
							assign node528 = (inp[1]) ? node534 : node529;
								assign node529 = (inp[11]) ? node531 : 3'b100;
									assign node531 = (inp[10]) ? 3'b000 : 3'b100;
								assign node534 = (inp[2]) ? 3'b000 : node535;
									assign node535 = (inp[8]) ? 3'b100 : 3'b000;
							assign node539 = (inp[5]) ? node547 : node540;
								assign node540 = (inp[10]) ? node544 : node541;
									assign node541 = (inp[8]) ? 3'b001 : 3'b010;
									assign node544 = (inp[8]) ? 3'b010 : 3'b100;
								assign node547 = (inp[10]) ? node551 : node548;
									assign node548 = (inp[1]) ? 3'b100 : 3'b110;
									assign node551 = (inp[1]) ? 3'b000 : 3'b100;
						assign node554 = (inp[10]) ? 3'b000 : node555;
							assign node555 = (inp[7]) ? node557 : 3'b000;
								assign node557 = (inp[2]) ? 3'b000 : node558;
									assign node558 = (inp[8]) ? 3'b100 : 3'b000;
					assign node563 = (inp[0]) ? 3'b000 : node564;
						assign node564 = (inp[7]) ? node566 : 3'b000;
							assign node566 = (inp[1]) ? 3'b000 : node567;
								assign node567 = (inp[5]) ? 3'b000 : node568;
									assign node568 = (inp[11]) ? 3'b000 : 3'b100;
			assign node574 = (inp[9]) ? node688 : node575;
				assign node575 = (inp[0]) ? node631 : node576;
					assign node576 = (inp[10]) ? node604 : node577;
						assign node577 = (inp[8]) ? node591 : node578;
							assign node578 = (inp[2]) ? node586 : node579;
								assign node579 = (inp[4]) ? node583 : node580;
									assign node580 = (inp[7]) ? 3'b011 : 3'b101;
									assign node583 = (inp[1]) ? 3'b001 : 3'b101;
								assign node586 = (inp[1]) ? node588 : 3'b001;
									assign node588 = (inp[4]) ? 3'b010 : 3'b001;
							assign node591 = (inp[2]) ? node599 : node592;
								assign node592 = (inp[11]) ? node596 : node593;
									assign node593 = (inp[4]) ? 3'b001 : 3'b011;
									assign node596 = (inp[7]) ? 3'b001 : 3'b001;
								assign node599 = (inp[7]) ? node601 : 3'b001;
									assign node601 = (inp[5]) ? 3'b001 : 3'b101;
						assign node604 = (inp[7]) ? node618 : node605;
							assign node605 = (inp[4]) ? node613 : node606;
								assign node606 = (inp[1]) ? node610 : node607;
									assign node607 = (inp[5]) ? 3'b001 : 3'b101;
									assign node610 = (inp[8]) ? 3'b110 : 3'b110;
								assign node613 = (inp[8]) ? node615 : 3'b010;
									assign node615 = (inp[11]) ? 3'b010 : 3'b110;
							assign node618 = (inp[1]) ? node626 : node619;
								assign node619 = (inp[8]) ? node623 : node620;
									assign node620 = (inp[5]) ? 3'b001 : 3'b101;
									assign node623 = (inp[4]) ? 3'b101 : 3'b011;
								assign node626 = (inp[4]) ? 3'b110 : node627;
									assign node627 = (inp[11]) ? 3'b001 : 3'b101;
					assign node631 = (inp[4]) ? node663 : node632;
						assign node632 = (inp[7]) ? node648 : node633;
							assign node633 = (inp[10]) ? node641 : node634;
								assign node634 = (inp[5]) ? node638 : node635;
									assign node635 = (inp[1]) ? 3'b110 : 3'b001;
									assign node638 = (inp[2]) ? 3'b010 : 3'b110;
								assign node641 = (inp[1]) ? node645 : node642;
									assign node642 = (inp[11]) ? 3'b010 : 3'b110;
									assign node645 = (inp[5]) ? 3'b000 : 3'b010;
							assign node648 = (inp[10]) ? node656 : node649;
								assign node649 = (inp[11]) ? node653 : node650;
									assign node650 = (inp[8]) ? 3'b101 : 3'b001;
									assign node653 = (inp[2]) ? 3'b001 : 3'b001;
								assign node656 = (inp[5]) ? node660 : node657;
									assign node657 = (inp[8]) ? 3'b001 : 3'b000;
									assign node660 = (inp[2]) ? 3'b110 : 3'b000;
						assign node663 = (inp[7]) ? node679 : node664;
							assign node664 = (inp[8]) ? node672 : node665;
								assign node665 = (inp[10]) ? node669 : node666;
									assign node666 = (inp[5]) ? 3'b100 : 3'b100;
									assign node669 = (inp[1]) ? 3'b000 : 3'b100;
								assign node672 = (inp[1]) ? node676 : node673;
									assign node673 = (inp[5]) ? 3'b010 : 3'b010;
									assign node676 = (inp[10]) ? 3'b100 : 3'b010;
							assign node679 = (inp[10]) ? node681 : 3'b110;
								assign node681 = (inp[5]) ? node685 : node682;
									assign node682 = (inp[8]) ? 3'b110 : 3'b010;
									assign node685 = (inp[8]) ? 3'b010 : 3'b100;
				assign node688 = (inp[0]) ? node748 : node689;
					assign node689 = (inp[7]) ? node719 : node690;
						assign node690 = (inp[4]) ? node704 : node691;
							assign node691 = (inp[1]) ? node697 : node692;
								assign node692 = (inp[2]) ? 3'b110 : node693;
									assign node693 = (inp[8]) ? 3'b001 : 3'b010;
								assign node697 = (inp[10]) ? node701 : node698;
									assign node698 = (inp[11]) ? 3'b110 : 3'b010;
									assign node701 = (inp[2]) ? 3'b100 : 3'b100;
							assign node704 = (inp[10]) ? node712 : node705;
								assign node705 = (inp[1]) ? node709 : node706;
									assign node706 = (inp[8]) ? 3'b010 : 3'b100;
									assign node709 = (inp[8]) ? 3'b100 : 3'b000;
								assign node712 = (inp[1]) ? node716 : node713;
									assign node713 = (inp[2]) ? 3'b000 : 3'b100;
									assign node716 = (inp[5]) ? 3'b000 : 3'b000;
						assign node719 = (inp[11]) ? node733 : node720;
							assign node720 = (inp[1]) ? node726 : node721;
								assign node721 = (inp[4]) ? node723 : 3'b001;
									assign node723 = (inp[2]) ? 3'b010 : 3'b001;
								assign node726 = (inp[10]) ? node730 : node727;
									assign node727 = (inp[2]) ? 3'b010 : 3'b001;
									assign node730 = (inp[2]) ? 3'b100 : 3'b010;
							assign node733 = (inp[2]) ? node741 : node734;
								assign node734 = (inp[8]) ? node738 : node735;
									assign node735 = (inp[4]) ? 3'b010 : 3'b000;
									assign node738 = (inp[4]) ? 3'b100 : 3'b001;
								assign node741 = (inp[10]) ? node745 : node742;
									assign node742 = (inp[5]) ? 3'b010 : 3'b110;
									assign node745 = (inp[5]) ? 3'b110 : 3'b010;
					assign node748 = (inp[7]) ? node770 : node749;
						assign node749 = (inp[11]) ? node763 : node750;
							assign node750 = (inp[4]) ? node758 : node751;
								assign node751 = (inp[1]) ? node755 : node752;
									assign node752 = (inp[8]) ? 3'b010 : 3'b100;
									assign node755 = (inp[2]) ? 3'b100 : 3'b000;
								assign node758 = (inp[1]) ? 3'b000 : node759;
									assign node759 = (inp[2]) ? 3'b000 : 3'b100;
							assign node763 = (inp[8]) ? node765 : 3'b000;
								assign node765 = (inp[1]) ? node767 : 3'b010;
									assign node767 = (inp[10]) ? 3'b000 : 3'b000;
						assign node770 = (inp[4]) ? node784 : node771;
							assign node771 = (inp[10]) ? node777 : node772;
								assign node772 = (inp[2]) ? node774 : 3'b110;
									assign node774 = (inp[1]) ? 3'b010 : 3'b010;
								assign node777 = (inp[11]) ? node781 : node778;
									assign node778 = (inp[5]) ? 3'b010 : 3'b010;
									assign node781 = (inp[1]) ? 3'b100 : 3'b100;
							assign node784 = (inp[1]) ? node792 : node785;
								assign node785 = (inp[5]) ? node789 : node786;
									assign node786 = (inp[8]) ? 3'b010 : 3'b000;
									assign node789 = (inp[2]) ? 3'b000 : 3'b100;
								assign node792 = (inp[10]) ? 3'b000 : node793;
									assign node793 = (inp[5]) ? 3'b000 : 3'b100;

endmodule