module dtc_split05_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node145;

	assign outp = (inp[9]) ? node90 : node1;
		assign node1 = (inp[6]) ? node45 : node2;
			assign node2 = (inp[10]) ? node14 : node3;
				assign node3 = (inp[7]) ? node5 : 3'b111;
					assign node5 = (inp[11]) ? 3'b011 : node6;
						assign node6 = (inp[4]) ? 3'b011 : node7;
							assign node7 = (inp[1]) ? 3'b111 : node8;
								assign node8 = (inp[3]) ? 3'b011 : 3'b111;
				assign node14 = (inp[11]) ? node32 : node15;
					assign node15 = (inp[7]) ? node25 : node16;
						assign node16 = (inp[3]) ? node20 : node17;
							assign node17 = (inp[8]) ? 3'b011 : 3'b111;
							assign node20 = (inp[8]) ? node22 : 3'b011;
								assign node22 = (inp[1]) ? 3'b101 : 3'b011;
						assign node25 = (inp[8]) ? 3'b001 : node26;
							assign node26 = (inp[2]) ? node28 : 3'b101;
								assign node28 = (inp[5]) ? 3'b001 : 3'b011;
					assign node32 = (inp[3]) ? node38 : node33;
						assign node33 = (inp[5]) ? 3'b011 : node34;
							assign node34 = (inp[7]) ? 3'b001 : 3'b101;
						assign node38 = (inp[7]) ? node40 : 3'b101;
							assign node40 = (inp[0]) ? node42 : 3'b110;
								assign node42 = (inp[5]) ? 3'b010 : 3'b110;
			assign node45 = (inp[10]) ? node73 : node46;
				assign node46 = (inp[11]) ? node60 : node47;
					assign node47 = (inp[5]) ? node53 : node48;
						assign node48 = (inp[3]) ? node50 : 3'b101;
							assign node50 = (inp[8]) ? 3'b001 : 3'b101;
						assign node53 = (inp[4]) ? 3'b011 : node54;
							assign node54 = (inp[1]) ? 3'b001 : node55;
								assign node55 = (inp[7]) ? 3'b001 : 3'b101;
					assign node60 = (inp[7]) ? node66 : node61;
						assign node61 = (inp[3]) ? 3'b110 : node62;
							assign node62 = (inp[8]) ? 3'b001 : 3'b101;
						assign node66 = (inp[2]) ? node68 : 3'b010;
							assign node68 = (inp[8]) ? 3'b100 : node69;
								assign node69 = (inp[3]) ? 3'b010 : 3'b110;
				assign node73 = (inp[2]) ? node83 : node74;
					assign node74 = (inp[7]) ? node78 : node75;
						assign node75 = (inp[8]) ? 3'b010 : 3'b001;
						assign node78 = (inp[11]) ? node80 : 3'b010;
							assign node80 = (inp[8]) ? 3'b000 : 3'b100;
					assign node83 = (inp[4]) ? node85 : 3'b100;
						assign node85 = (inp[11]) ? 3'b100 : node86;
							assign node86 = (inp[7]) ? 3'b010 : 3'b110;
		assign node90 = (inp[6]) ? node138 : node91;
			assign node91 = (inp[10]) ? node113 : node92;
				assign node92 = (inp[7]) ? node102 : node93;
					assign node93 = (inp[8]) ? node97 : node94;
						assign node94 = (inp[1]) ? 3'b101 : 3'b001;
						assign node97 = (inp[11]) ? node99 : 3'b001;
							assign node99 = (inp[3]) ? 3'b010 : 3'b110;
					assign node102 = (inp[1]) ? node108 : node103;
						assign node103 = (inp[11]) ? node105 : 3'b110;
							assign node105 = (inp[4]) ? 3'b100 : 3'b010;
						assign node108 = (inp[8]) ? node110 : 3'b010;
							assign node110 = (inp[5]) ? 3'b010 : 3'b110;
				assign node113 = (inp[7]) ? node131 : node114;
					assign node114 = (inp[11]) ? node122 : node115;
						assign node115 = (inp[8]) ? node117 : 3'b010;
							assign node117 = (inp[3]) ? 3'b100 : node118;
								assign node118 = (inp[2]) ? 3'b010 : 3'b000;
						assign node122 = (inp[1]) ? node128 : node123;
							assign node123 = (inp[0]) ? node125 : 3'b010;
								assign node125 = (inp[5]) ? 3'b010 : 3'b100;
							assign node128 = (inp[3]) ? 3'b000 : 3'b100;
					assign node131 = (inp[11]) ? 3'b000 : node132;
						assign node132 = (inp[8]) ? 3'b000 : node133;
							assign node133 = (inp[3]) ? 3'b000 : 3'b100;
			assign node138 = (inp[7]) ? 3'b000 : node139;
				assign node139 = (inp[10]) ? 3'b000 : node140;
					assign node140 = (inp[11]) ? 3'b000 : node141;
						assign node141 = (inp[5]) ? node143 : 3'b010;
							assign node143 = (inp[1]) ? node145 : 3'b100;
								assign node145 = (inp[2]) ? 3'b000 : 3'b100;

endmodule