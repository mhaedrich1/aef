module dtc_split66_bm67 (
	input  wire [10-1:0] inp,
	output wire [77-1:0] outp
);

	wire [77-1:0] node1;
	wire [77-1:0] node4;

	assign outp = (inp[8]) ? node4 : node1;
		assign node1 = (inp[1]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000100000000000;
		assign node4 = (inp[7]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule