module dtc_split5_bm82 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;

	assign outp = (inp[0]) ? node60 : node1;
		assign node1 = (inp[3]) ? node31 : node2;
			assign node2 = (inp[6]) ? node16 : node3;
				assign node3 = (inp[4]) ? node9 : node4;
					assign node4 = (inp[7]) ? node6 : 3'b001;
						assign node6 = (inp[1]) ? 3'b011 : 3'b111;
					assign node9 = (inp[1]) ? node13 : node10;
						assign node10 = (inp[7]) ? 3'b111 : 3'b111;
						assign node13 = (inp[8]) ? 3'b101 : 3'b011;
				assign node16 = (inp[1]) ? node24 : node17;
					assign node17 = (inp[7]) ? node21 : node18;
						assign node18 = (inp[9]) ? 3'b111 : 3'b001;
						assign node21 = (inp[9]) ? 3'b101 : 3'b110;
					assign node24 = (inp[9]) ? node28 : node25;
						assign node25 = (inp[4]) ? 3'b000 : 3'b000;
						assign node28 = (inp[10]) ? 3'b101 : 3'b010;
			assign node31 = (inp[6]) ? node45 : node32;
				assign node32 = (inp[4]) ? node40 : node33;
					assign node33 = (inp[9]) ? node37 : node34;
						assign node34 = (inp[1]) ? 3'b111 : 3'b111;
						assign node37 = (inp[8]) ? 3'b111 : 3'b111;
					assign node40 = (inp[7]) ? node42 : 3'b111;
						assign node42 = (inp[2]) ? 3'b111 : 3'b111;
				assign node45 = (inp[1]) ? node53 : node46;
					assign node46 = (inp[9]) ? node50 : node47;
						assign node47 = (inp[7]) ? 3'b011 : 3'b111;
						assign node50 = (inp[4]) ? 3'b111 : 3'b111;
					assign node53 = (inp[9]) ? node57 : node54;
						assign node54 = (inp[7]) ? 3'b010 : 3'b001;
						assign node57 = (inp[7]) ? 3'b101 : 3'b111;
		assign node60 = (inp[6]) ? node92 : node61;
			assign node61 = (inp[3]) ? node77 : node62;
				assign node62 = (inp[1]) ? node70 : node63;
					assign node63 = (inp[7]) ? node67 : node64;
						assign node64 = (inp[4]) ? 3'b001 : 3'b100;
						assign node67 = (inp[9]) ? 3'b111 : 3'b100;
					assign node70 = (inp[7]) ? node74 : node71;
						assign node71 = (inp[4]) ? 3'b000 : 3'b010;
						assign node74 = (inp[9]) ? 3'b000 : 3'b000;
				assign node77 = (inp[1]) ? node85 : node78;
					assign node78 = (inp[9]) ? node82 : node79;
						assign node79 = (inp[7]) ? 3'b011 : 3'b111;
						assign node82 = (inp[7]) ? 3'b111 : 3'b111;
					assign node85 = (inp[9]) ? node89 : node86;
						assign node86 = (inp[7]) ? 3'b110 : 3'b101;
						assign node89 = (inp[7]) ? 3'b101 : 3'b111;
			assign node92 = (inp[3]) ? node106 : node93;
				assign node93 = (inp[9]) ? node99 : node94;
					assign node94 = (inp[4]) ? node96 : 3'b000;
						assign node96 = (inp[7]) ? 3'b000 : 3'b000;
					assign node99 = (inp[1]) ? node103 : node100;
						assign node100 = (inp[7]) ? 3'b000 : 3'b010;
						assign node103 = (inp[7]) ? 3'b000 : 3'b000;
				assign node106 = (inp[1]) ? node114 : node107;
					assign node107 = (inp[9]) ? node111 : node108;
						assign node108 = (inp[7]) ? 3'b000 : 3'b010;
						assign node111 = (inp[4]) ? 3'b101 : 3'b100;
					assign node114 = (inp[7]) ? node118 : node115;
						assign node115 = (inp[9]) ? 3'b000 : 3'b000;
						assign node118 = (inp[4]) ? 3'b000 : 3'b000;

endmodule