module dtc_split75_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node10;
	wire [14-1:0] node13;
	wire [14-1:0] node14;
	wire [14-1:0] node17;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node25;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node32;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node41;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node48;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node56;
	wire [14-1:0] node59;
	wire [14-1:0] node60;
	wire [14-1:0] node63;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node73;
	wire [14-1:0] node76;
	wire [14-1:0] node77;
	wire [14-1:0] node80;
	wire [14-1:0] node83;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node88;
	wire [14-1:0] node91;
	wire [14-1:0] node92;
	wire [14-1:0] node95;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node101;
	wire [14-1:0] node104;
	wire [14-1:0] node107;
	wire [14-1:0] node108;
	wire [14-1:0] node111;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node116;
	wire [14-1:0] node119;
	wire [14-1:0] node122;
	wire [14-1:0] node123;
	wire [14-1:0] node126;
	wire [14-1:0] node129;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node132;
	wire [14-1:0] node133;
	wire [14-1:0] node134;
	wire [14-1:0] node137;
	wire [14-1:0] node140;
	wire [14-1:0] node141;
	wire [14-1:0] node144;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node149;
	wire [14-1:0] node152;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node159;
	wire [14-1:0] node162;
	wire [14-1:0] node163;
	wire [14-1:0] node164;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node175;
	wire [14-1:0] node178;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node183;
	wire [14-1:0] node186;
	wire [14-1:0] node187;
	wire [14-1:0] node190;
	wire [14-1:0] node193;
	wire [14-1:0] node194;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node200;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node207;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node222;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node231;
	wire [14-1:0] node234;
	wire [14-1:0] node235;
	wire [14-1:0] node238;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node243;
	wire [14-1:0] node246;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node253;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node258;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node262;
	wire [14-1:0] node265;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node272;
	wire [14-1:0] node275;
	wire [14-1:0] node276;
	wire [14-1:0] node277;
	wire [14-1:0] node280;
	wire [14-1:0] node283;
	wire [14-1:0] node284;
	wire [14-1:0] node287;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node293;
	wire [14-1:0] node296;
	wire [14-1:0] node299;
	wire [14-1:0] node300;
	wire [14-1:0] node303;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node311;
	wire [14-1:0] node314;
	wire [14-1:0] node315;
	wire [14-1:0] node318;
	wire [14-1:0] node321;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node328;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node340;
	wire [14-1:0] node343;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node350;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node359;
	wire [14-1:0] node362;
	wire [14-1:0] node363;
	wire [14-1:0] node366;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node374;
	wire [14-1:0] node377;
	wire [14-1:0] node378;
	wire [14-1:0] node381;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node392;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node399;
	wire [14-1:0] node402;
	wire [14-1:0] node403;
	wire [14-1:0] node404;
	wire [14-1:0] node407;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node414;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node423;
	wire [14-1:0] node426;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node433;
	wire [14-1:0] node434;
	wire [14-1:0] node435;
	wire [14-1:0] node438;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node445;
	wire [14-1:0] node448;
	wire [14-1:0] node449;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node452;
	wire [14-1:0] node455;
	wire [14-1:0] node458;
	wire [14-1:0] node459;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node470;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node482;
	wire [14-1:0] node483;
	wire [14-1:0] node486;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node493;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node501;
	wire [14-1:0] node504;
	wire [14-1:0] node505;
	wire [14-1:0] node508;

	assign outp = (inp[4]) ? node256 : node1;
		assign node1 = (inp[11]) ? node129 : node2;
			assign node2 = (inp[12]) ? node66 : node3;
				assign node3 = (inp[6]) ? node35 : node4;
					assign node4 = (inp[8]) ? node20 : node5;
						assign node5 = (inp[13]) ? node13 : node6;
							assign node6 = (inp[3]) ? node10 : node7;
								assign node7 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
								assign node10 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
							assign node13 = (inp[1]) ? node17 : node14;
								assign node14 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node17 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node20 = (inp[0]) ? node28 : node21;
							assign node21 = (inp[2]) ? node25 : node22;
								assign node22 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node25 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node28 = (inp[10]) ? node32 : node29;
								assign node29 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node32 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
					assign node35 = (inp[13]) ? node51 : node36;
						assign node36 = (inp[5]) ? node44 : node37;
							assign node37 = (inp[0]) ? node41 : node38;
								assign node38 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node41 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node44 = (inp[1]) ? node48 : node45;
								assign node45 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node48 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node51 = (inp[0]) ? node59 : node52;
							assign node52 = (inp[5]) ? node56 : node53;
								assign node53 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node56 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node59 = (inp[9]) ? node63 : node60;
								assign node60 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node63 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
				assign node66 = (inp[5]) ? node98 : node67;
					assign node67 = (inp[7]) ? node83 : node68;
						assign node68 = (inp[10]) ? node76 : node69;
							assign node69 = (inp[2]) ? node73 : node70;
								assign node70 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node73 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node76 = (inp[8]) ? node80 : node77;
								assign node77 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node80 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node83 = (inp[13]) ? node91 : node84;
							assign node84 = (inp[0]) ? node88 : node85;
								assign node85 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node88 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node91 = (inp[6]) ? node95 : node92;
								assign node92 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node95 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node98 = (inp[9]) ? node114 : node99;
						assign node99 = (inp[1]) ? node107 : node100;
							assign node100 = (inp[6]) ? node104 : node101;
								assign node101 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node104 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node107 = (inp[13]) ? node111 : node108;
								assign node108 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node111 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node114 = (inp[2]) ? node122 : node115;
							assign node115 = (inp[0]) ? node119 : node116;
								assign node116 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node119 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node122 = (inp[13]) ? node126 : node123;
								assign node123 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node126 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
			assign node129 = (inp[9]) ? node193 : node130;
				assign node130 = (inp[1]) ? node162 : node131;
					assign node131 = (inp[2]) ? node147 : node132;
						assign node132 = (inp[12]) ? node140 : node133;
							assign node133 = (inp[6]) ? node137 : node134;
								assign node134 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node137 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node140 = (inp[6]) ? node144 : node141;
								assign node141 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node144 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node147 = (inp[5]) ? node155 : node148;
							assign node148 = (inp[7]) ? node152 : node149;
								assign node149 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node152 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node155 = (inp[8]) ? node159 : node156;
								assign node156 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node159 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node162 = (inp[3]) ? node178 : node163;
						assign node163 = (inp[7]) ? node171 : node164;
							assign node164 = (inp[12]) ? node168 : node165;
								assign node165 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node168 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node171 = (inp[6]) ? node175 : node172;
								assign node172 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node175 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node178 = (inp[6]) ? node186 : node179;
							assign node179 = (inp[2]) ? node183 : node180;
								assign node180 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node183 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node186 = (inp[7]) ? node190 : node187;
								assign node187 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node190 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
				assign node193 = (inp[13]) ? node225 : node194;
					assign node194 = (inp[2]) ? node210 : node195;
						assign node195 = (inp[6]) ? node203 : node196;
							assign node196 = (inp[7]) ? node200 : node197;
								assign node197 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node200 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node203 = (inp[8]) ? node207 : node204;
								assign node204 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node207 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node210 = (inp[7]) ? node218 : node211;
							assign node211 = (inp[8]) ? node215 : node212;
								assign node212 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node215 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node218 = (inp[3]) ? node222 : node219;
								assign node219 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node222 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node225 = (inp[10]) ? node241 : node226;
						assign node226 = (inp[3]) ? node234 : node227;
							assign node227 = (inp[5]) ? node231 : node228;
								assign node228 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node231 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node234 = (inp[7]) ? node238 : node235;
								assign node235 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node238 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node241 = (inp[3]) ? node249 : node242;
							assign node242 = (inp[7]) ? node246 : node243;
								assign node243 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node246 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node249 = (inp[8]) ? node253 : node250;
								assign node250 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node253 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
		assign node256 = (inp[7]) ? node384 : node257;
			assign node257 = (inp[10]) ? node321 : node258;
				assign node258 = (inp[0]) ? node290 : node259;
					assign node259 = (inp[6]) ? node275 : node260;
						assign node260 = (inp[1]) ? node268 : node261;
							assign node261 = (inp[2]) ? node265 : node262;
								assign node262 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node265 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node268 = (inp[9]) ? node272 : node269;
								assign node269 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node272 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node275 = (inp[13]) ? node283 : node276;
							assign node276 = (inp[5]) ? node280 : node277;
								assign node277 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node280 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node283 = (inp[8]) ? node287 : node284;
								assign node284 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node287 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
					assign node290 = (inp[2]) ? node306 : node291;
						assign node291 = (inp[8]) ? node299 : node292;
							assign node292 = (inp[3]) ? node296 : node293;
								assign node293 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node296 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node299 = (inp[1]) ? node303 : node300;
								assign node300 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node303 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node306 = (inp[8]) ? node314 : node307;
							assign node307 = (inp[13]) ? node311 : node308;
								assign node308 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node311 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node314 = (inp[6]) ? node318 : node315;
								assign node315 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node318 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
				assign node321 = (inp[3]) ? node353 : node322;
					assign node322 = (inp[11]) ? node338 : node323;
						assign node323 = (inp[8]) ? node331 : node324;
							assign node324 = (inp[13]) ? node328 : node325;
								assign node325 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node328 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node331 = (inp[12]) ? node335 : node332;
								assign node332 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node335 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node338 = (inp[9]) ? node346 : node339;
							assign node339 = (inp[0]) ? node343 : node340;
								assign node340 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node343 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node346 = (inp[5]) ? node350 : node347;
								assign node347 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node350 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node353 = (inp[6]) ? node369 : node354;
						assign node354 = (inp[2]) ? node362 : node355;
							assign node355 = (inp[5]) ? node359 : node356;
								assign node356 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node359 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node362 = (inp[0]) ? node366 : node363;
								assign node363 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node366 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node369 = (inp[1]) ? node377 : node370;
							assign node370 = (inp[8]) ? node374 : node371;
								assign node371 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node374 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node377 = (inp[13]) ? node381 : node378;
								assign node378 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node381 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
			assign node384 = (inp[13]) ? node448 : node385;
				assign node385 = (inp[5]) ? node417 : node386;
					assign node386 = (inp[10]) ? node402 : node387;
						assign node387 = (inp[8]) ? node395 : node388;
							assign node388 = (inp[0]) ? node392 : node389;
								assign node389 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node392 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node395 = (inp[1]) ? node399 : node396;
								assign node396 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node399 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node402 = (inp[1]) ? node410 : node403;
							assign node403 = (inp[12]) ? node407 : node404;
								assign node404 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node407 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node410 = (inp[3]) ? node414 : node411;
								assign node411 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node414 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node417 = (inp[6]) ? node433 : node418;
						assign node418 = (inp[9]) ? node426 : node419;
							assign node419 = (inp[12]) ? node423 : node420;
								assign node420 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node423 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node426 = (inp[3]) ? node430 : node427;
								assign node427 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node430 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node433 = (inp[11]) ? node441 : node434;
							assign node434 = (inp[2]) ? node438 : node435;
								assign node435 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node438 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node441 = (inp[8]) ? node445 : node442;
								assign node442 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node445 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node448 = (inp[10]) ? node480 : node449;
					assign node449 = (inp[1]) ? node465 : node450;
						assign node450 = (inp[6]) ? node458 : node451;
							assign node451 = (inp[3]) ? node455 : node452;
								assign node452 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node455 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node458 = (inp[5]) ? node462 : node459;
								assign node459 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node462 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node465 = (inp[8]) ? node473 : node466;
							assign node466 = (inp[2]) ? node470 : node467;
								assign node467 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node470 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node473 = (inp[5]) ? node477 : node474;
								assign node474 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node477 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node480 = (inp[8]) ? node496 : node481;
						assign node481 = (inp[11]) ? node489 : node482;
							assign node482 = (inp[1]) ? node486 : node483;
								assign node483 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node486 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node489 = (inp[0]) ? node493 : node490;
								assign node490 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node493 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node496 = (inp[2]) ? node504 : node497;
							assign node497 = (inp[12]) ? node501 : node498;
								assign node498 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node501 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node504 = (inp[3]) ? node508 : node505;
								assign node505 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node508 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;

endmodule