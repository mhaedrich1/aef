module dtc_split125_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node21;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node42;
	wire [4-1:0] node44;
	wire [4-1:0] node46;
	wire [4-1:0] node48;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node59;
	wire [4-1:0] node61;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node85;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node91;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node105;
	wire [4-1:0] node106;
	wire [4-1:0] node108;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node113;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node122;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node143;
	wire [4-1:0] node146;
	wire [4-1:0] node148;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node153;
	wire [4-1:0] node155;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node167;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node181;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node189;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node205;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node210;
	wire [4-1:0] node212;
	wire [4-1:0] node214;
	wire [4-1:0] node217;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node225;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node232;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node240;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node250;
	wire [4-1:0] node255;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node283;
	wire [4-1:0] node285;
	wire [4-1:0] node287;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node295;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node302;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node322;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node341;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node346;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node356;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node363;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node370;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node394;
	wire [4-1:0] node396;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node402;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node411;
	wire [4-1:0] node413;
	wire [4-1:0] node418;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node448;
	wire [4-1:0] node453;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node459;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node468;
	wire [4-1:0] node470;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node483;
	wire [4-1:0] node489;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node506;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node555;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node586;
	wire [4-1:0] node588;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node595;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node610;
	wire [4-1:0] node614;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node641;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node650;
	wire [4-1:0] node652;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node661;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node704;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node709;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node746;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node767;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node778;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node796;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node814;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node822;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node840;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node847;
	wire [4-1:0] node849;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node860;
	wire [4-1:0] node862;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node880;
	wire [4-1:0] node882;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node897;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node902;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node915;
	wire [4-1:0] node917;
	wire [4-1:0] node919;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node935;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node949;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node955;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node967;
	wire [4-1:0] node971;
	wire [4-1:0] node973;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node984;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node998;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1005;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1011;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1015;
	wire [4-1:0] node1020;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1034;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1052;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1061;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1089;
	wire [4-1:0] node1093;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1098;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1106;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1113;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1120;
	wire [4-1:0] node1122;
	wire [4-1:0] node1125;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1131;
	wire [4-1:0] node1134;

	assign outp = (inp[10]) ? node434 : node1;
		assign node1 = (inp[5]) ? node159 : node2;
			assign node2 = (inp[4]) ? node78 : node3;
				assign node3 = (inp[14]) ? node39 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node24 : node7;
							assign node7 = (inp[6]) ? node9 : 4'b1111;
								assign node9 = (inp[9]) ? node11 : 4'b1111;
									assign node11 = (inp[8]) ? node13 : 4'b1111;
										assign node13 = (inp[7]) ? node21 : node14;
											assign node14 = (inp[1]) ? node16 : 4'b1111;
												assign node16 = (inp[15]) ? node18 : 4'b1111;
													assign node18 = (inp[11]) ? 4'b1101 : 4'b1111;
											assign node21 = (inp[2]) ? 4'b1101 : 4'b1111;
							assign node24 = (inp[2]) ? 4'b1101 : node25;
								assign node25 = (inp[6]) ? node31 : node26;
									assign node26 = (inp[9]) ? node28 : 4'b1111;
										assign node28 = (inp[8]) ? 4'b1101 : 4'b1111;
									assign node31 = (inp[7]) ? 4'b1101 : node32;
										assign node32 = (inp[9]) ? 4'b1101 : node33;
											assign node33 = (inp[8]) ? 4'b1101 : 4'b1111;
					assign node39 = (inp[13]) ? node51 : node40;
						assign node40 = (inp[12]) ? node42 : 4'b1101;
							assign node42 = (inp[6]) ? node44 : 4'b1101;
								assign node44 = (inp[9]) ? node46 : 4'b1101;
									assign node46 = (inp[2]) ? node48 : 4'b1101;
										assign node48 = (inp[8]) ? 4'b1011 : 4'b1101;
						assign node51 = (inp[12]) ? node65 : node52;
							assign node52 = (inp[8]) ? node54 : 4'b1101;
								assign node54 = (inp[9]) ? node56 : 4'b1101;
									assign node56 = (inp[2]) ? node58 : 4'b1101;
										assign node58 = (inp[6]) ? 4'b1011 : node59;
											assign node59 = (inp[7]) ? node61 : 4'b1101;
												assign node61 = (inp[15]) ? 4'b1111 : 4'b1101;
							assign node65 = (inp[6]) ? 4'b1011 : node66;
								assign node66 = (inp[9]) ? 4'b1111 : node67;
									assign node67 = (inp[2]) ? 4'b1111 : node68;
										assign node68 = (inp[8]) ? node70 : 4'b1101;
											assign node70 = (inp[15]) ? node72 : 4'b1101;
												assign node72 = (inp[7]) ? 4'b1111 : 4'b1101;
				assign node78 = (inp[6]) ? node122 : node79;
					assign node79 = (inp[14]) ? node105 : node80;
						assign node80 = (inp[12]) ? node96 : node81;
							assign node81 = (inp[13]) ? node83 : 4'b1011;
								assign node83 = (inp[9]) ? node85 : 4'b1011;
									assign node85 = (inp[2]) ? node87 : 4'b1011;
										assign node87 = (inp[8]) ? 4'b1001 : node88;
											assign node88 = (inp[7]) ? 4'b1001 : node89;
												assign node89 = (inp[11]) ? node91 : 4'b1011;
													assign node91 = (inp[0]) ? 4'b1001 : 4'b1011;
							assign node96 = (inp[13]) ? 4'b1001 : node97;
								assign node97 = (inp[2]) ? node99 : 4'b1011;
									assign node99 = (inp[8]) ? 4'b1001 : node100;
										assign node100 = (inp[9]) ? 4'b1001 : 4'b1011;
						assign node105 = (inp[12]) ? node117 : node106;
							assign node106 = (inp[13]) ? node108 : 4'b1001;
								assign node108 = (inp[2]) ? node110 : 4'b1001;
									assign node110 = (inp[9]) ? 4'b1011 : node111;
										assign node111 = (inp[7]) ? node113 : 4'b1001;
											assign node113 = (inp[0]) ? 4'b1001 : 4'b1011;
							assign node117 = (inp[13]) ? 4'b1011 : node118;
								assign node118 = (inp[2]) ? 4'b1011 : 4'b1001;
					assign node122 = (inp[14]) ? node140 : node123;
						assign node123 = (inp[12]) ? node133 : node124;
							assign node124 = (inp[13]) ? node126 : 4'b1011;
								assign node126 = (inp[2]) ? node128 : 4'b1011;
									assign node128 = (inp[9]) ? 4'b1001 : node129;
										assign node129 = (inp[8]) ? 4'b1001 : 4'b1011;
							assign node133 = (inp[13]) ? 4'b1001 : node134;
								assign node134 = (inp[9]) ? 4'b1001 : node135;
									assign node135 = (inp[2]) ? 4'b1001 : 4'b1011;
						assign node140 = (inp[12]) ? node146 : node141;
							assign node141 = (inp[13]) ? node143 : 4'b1001;
								assign node143 = (inp[2]) ? 4'b1111 : 4'b1001;
							assign node146 = (inp[2]) ? node148 : 4'b1110;
								assign node148 = (inp[13]) ? node150 : 4'b1110;
									assign node150 = (inp[9]) ? 4'b1100 : node151;
										assign node151 = (inp[8]) ? node153 : 4'b1110;
											assign node153 = (inp[11]) ? node155 : 4'b1110;
												assign node155 = (inp[15]) ? 4'b1100 : 4'b1110;
			assign node159 = (inp[12]) ? node273 : node160;
				assign node160 = (inp[6]) ? node220 : node161;
					assign node161 = (inp[13]) ? node205 : node162;
						assign node162 = (inp[4]) ? node186 : node163;
							assign node163 = (inp[8]) ? node175 : node164;
								assign node164 = (inp[14]) ? node170 : node165;
									assign node165 = (inp[2]) ? node167 : 4'b1001;
										assign node167 = (inp[9]) ? 4'b1011 : 4'b1001;
									assign node170 = (inp[9]) ? 4'b1001 : node171;
										assign node171 = (inp[2]) ? 4'b1001 : 4'b1011;
								assign node175 = (inp[2]) ? node177 : 4'b1001;
									assign node177 = (inp[14]) ? 4'b1001 : node178;
										assign node178 = (inp[9]) ? 4'b1011 : node179;
											assign node179 = (inp[3]) ? node181 : 4'b1001;
												assign node181 = (inp[1]) ? 4'b1001 : 4'b1011;
							assign node186 = (inp[14]) ? node194 : node187;
								assign node187 = (inp[9]) ? node189 : 4'b1101;
									assign node189 = (inp[2]) ? node191 : 4'b1101;
										assign node191 = (inp[8]) ? 4'b1011 : 4'b1101;
								assign node194 = (inp[9]) ? 4'b1001 : node195;
									assign node195 = (inp[2]) ? 4'b1001 : node196;
										assign node196 = (inp[8]) ? node198 : 4'b1011;
											assign node198 = (inp[7]) ? 4'b1001 : node199;
												assign node199 = (inp[0]) ? 4'b1011 : 4'b1001;
						assign node205 = (inp[14]) ? node207 : 4'b1011;
							assign node207 = (inp[2]) ? node217 : node208;
								assign node208 = (inp[8]) ? node210 : 4'b1001;
									assign node210 = (inp[15]) ? node212 : 4'b1001;
										assign node212 = (inp[7]) ? node214 : 4'b1001;
											assign node214 = (inp[4]) ? 4'b1011 : 4'b1001;
								assign node217 = (inp[4]) ? 4'b1011 : 4'b1111;
					assign node220 = (inp[14]) ? node244 : node221;
						assign node221 = (inp[4]) ? node237 : node222;
							assign node222 = (inp[13]) ? 4'b1101 : node223;
								assign node223 = (inp[9]) ? node225 : 4'b1111;
									assign node225 = (inp[2]) ? node227 : 4'b1111;
										assign node227 = (inp[8]) ? 4'b1101 : node228;
											assign node228 = (inp[3]) ? node230 : 4'b1111;
												assign node230 = (inp[1]) ? node232 : 4'b1111;
													assign node232 = (inp[7]) ? 4'b1101 : 4'b1111;
							assign node237 = (inp[13]) ? 4'b1001 : node238;
								assign node238 = (inp[2]) ? node240 : 4'b1011;
									assign node240 = (inp[9]) ? 4'b1001 : 4'b1011;
						assign node244 = (inp[4]) ? node266 : node245;
							assign node245 = (inp[2]) ? node255 : node246;
								assign node246 = (inp[13]) ? 4'b1111 : node247;
									assign node247 = (inp[9]) ? 4'b1111 : node248;
										assign node248 = (inp[8]) ? node250 : 4'b1101;
											assign node250 = (inp[15]) ? 4'b1111 : 4'b1101;
								assign node255 = (inp[13]) ? node257 : 4'b1111;
									assign node257 = (inp[9]) ? 4'b1101 : node258;
										assign node258 = (inp[8]) ? 4'b1101 : node259;
											assign node259 = (inp[7]) ? 4'b1101 : node260;
												assign node260 = (inp[11]) ? 4'b1101 : 4'b1111;
							assign node266 = (inp[13]) ? node268 : 4'b1110;
								assign node268 = (inp[2]) ? 4'b1100 : node269;
									assign node269 = (inp[9]) ? 4'b1100 : 4'b1110;
				assign node273 = (inp[6]) ? node377 : node274;
					assign node274 = (inp[14]) ? node350 : node275;
						assign node275 = (inp[4]) ? node333 : node276;
							assign node276 = (inp[9]) ? node290 : node277;
								assign node277 = (inp[2]) ? node281 : node278;
									assign node278 = (inp[13]) ? 4'b1110 : 4'b1100;
									assign node281 = (inp[3]) ? node283 : 4'b1110;
										assign node283 = (inp[13]) ? node285 : 4'b1110;
											assign node285 = (inp[8]) ? node287 : 4'b1110;
												assign node287 = (inp[7]) ? 4'b1100 : 4'b1110;
								assign node290 = (inp[15]) ? node298 : node291;
									assign node291 = (inp[2]) ? node295 : node292;
										assign node292 = (inp[13]) ? 4'b1110 : 4'b1100;
										assign node295 = (inp[13]) ? 4'b1100 : 4'b1110;
									assign node298 = (inp[7]) ? node318 : node299;
										assign node299 = (inp[11]) ? node305 : node300;
											assign node300 = (inp[2]) ? node302 : 4'b1100;
												assign node302 = (inp[13]) ? 4'b1100 : 4'b1110;
											assign node305 = (inp[0]) ? node311 : node306;
												assign node306 = (inp[13]) ? node308 : 4'b1110;
													assign node308 = (inp[2]) ? 4'b1100 : 4'b1110;
												assign node311 = (inp[1]) ? 4'b1110 : node312;
													assign node312 = (inp[13]) ? 4'b1100 : node313;
														assign node313 = (inp[2]) ? 4'b1110 : 4'b1100;
										assign node318 = (inp[0]) ? node326 : node319;
											assign node319 = (inp[1]) ? 4'b1110 : node320;
												assign node320 = (inp[8]) ? node322 : 4'b1100;
													assign node322 = (inp[13]) ? 4'b1100 : 4'b1110;
											assign node326 = (inp[2]) ? 4'b1110 : node327;
												assign node327 = (inp[13]) ? 4'b1110 : node328;
													assign node328 = (inp[8]) ? 4'b1110 : 4'b1100;
							assign node333 = (inp[13]) ? node341 : node334;
								assign node334 = (inp[2]) ? node336 : 4'b1110;
									assign node336 = (inp[9]) ? 4'b1100 : node337;
										assign node337 = (inp[8]) ? 4'b1100 : 4'b1110;
								assign node341 = (inp[2]) ? node343 : 4'b1100;
									assign node343 = (inp[9]) ? 4'b1110 : node344;
										assign node344 = (inp[7]) ? node346 : 4'b1100;
											assign node346 = (inp[15]) ? 4'b1110 : 4'b1100;
						assign node350 = (inp[4]) ? node360 : node351;
							assign node351 = (inp[13]) ? 4'b1010 : node352;
								assign node352 = (inp[9]) ? node354 : 4'b1100;
									assign node354 = (inp[2]) ? node356 : 4'b1100;
										assign node356 = (inp[8]) ? 4'b1010 : 4'b1100;
							assign node360 = (inp[13]) ? node370 : node361;
								assign node361 = (inp[9]) ? node363 : 4'b1110;
									assign node363 = (inp[2]) ? node365 : 4'b1110;
										assign node365 = (inp[7]) ? 4'b1100 : node366;
											assign node366 = (inp[8]) ? 4'b1100 : 4'b1110;
								assign node370 = (inp[8]) ? node372 : 4'b1100;
									assign node372 = (inp[9]) ? node374 : 4'b1100;
										assign node374 = (inp[2]) ? 4'b1010 : 4'b1100;
					assign node377 = (inp[13]) ? node405 : node378;
						assign node378 = (inp[4]) ? node394 : node379;
							assign node379 = (inp[2]) ? 4'b1000 : node380;
								assign node380 = (inp[14]) ? node388 : node381;
									assign node381 = (inp[8]) ? 4'b1000 : node382;
										assign node382 = (inp[9]) ? 4'b1000 : node383;
											assign node383 = (inp[7]) ? 4'b1000 : 4'b1010;
									assign node388 = (inp[9]) ? node390 : 4'b1010;
										assign node390 = (inp[8]) ? 4'b1000 : 4'b1010;
							assign node394 = (inp[7]) ? node396 : 4'b1010;
								assign node396 = (inp[1]) ? node398 : 4'b1010;
									assign node398 = (inp[8]) ? node400 : 4'b1010;
										assign node400 = (inp[2]) ? node402 : 4'b1010;
											assign node402 = (inp[9]) ? 4'b1000 : 4'b1010;
						assign node405 = (inp[4]) ? node421 : node406;
							assign node406 = (inp[2]) ? node418 : node407;
								assign node407 = (inp[14]) ? 4'b1000 : node408;
									assign node408 = (inp[9]) ? 4'b1010 : node409;
										assign node409 = (inp[7]) ? node411 : 4'b1000;
											assign node411 = (inp[15]) ? node413 : 4'b1000;
												assign node413 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node418 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node421 = (inp[14]) ? 4'b1000 : node422;
								assign node422 = (inp[9]) ? node424 : 4'b1000;
									assign node424 = (inp[7]) ? node426 : 4'b1000;
										assign node426 = (inp[8]) ? node428 : 4'b1000;
											assign node428 = (inp[2]) ? node430 : 4'b1000;
												assign node430 = (inp[15]) ? 4'b1010 : 4'b1000;
		assign node434 = (inp[5]) ? node632 : node435;
			assign node435 = (inp[4]) ? node539 : node436;
				assign node436 = (inp[6]) ? node506 : node437;
					assign node437 = (inp[14]) ? node473 : node438;
						assign node438 = (inp[2]) ? node464 : node439;
							assign node439 = (inp[13]) ? node453 : node440;
								assign node440 = (inp[12]) ? node442 : 4'b1100;
									assign node442 = (inp[9]) ? node444 : 4'b1110;
										assign node444 = (inp[7]) ? 4'b1100 : node445;
											assign node445 = (inp[8]) ? 4'b1100 : node446;
												assign node446 = (inp[1]) ? node448 : 4'b1110;
													assign node448 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node453 = (inp[0]) ? node455 : 4'b1100;
									assign node455 = (inp[11]) ? 4'b1100 : node456;
										assign node456 = (inp[12]) ? 4'b1100 : node457;
											assign node457 = (inp[15]) ? node459 : 4'b1100;
												assign node459 = (inp[9]) ? 4'b1110 : 4'b1100;
							assign node464 = (inp[13]) ? node466 : 4'b1100;
								assign node466 = (inp[12]) ? node468 : 4'b1110;
									assign node468 = (inp[9]) ? node470 : 4'b1100;
										assign node470 = (inp[8]) ? 4'b1010 : 4'b1100;
						assign node473 = (inp[12]) ? node489 : node474;
							assign node474 = (inp[13]) ? node476 : 4'b1110;
								assign node476 = (inp[2]) ? 4'b1100 : node477;
									assign node477 = (inp[9]) ? 4'b1100 : node478;
										assign node478 = (inp[8]) ? node480 : 4'b1110;
											assign node480 = (inp[0]) ? 4'b1100 : node481;
												assign node481 = (inp[1]) ? node483 : 4'b1110;
													assign node483 = (inp[3]) ? 4'b1100 : 4'b1110;
							assign node489 = (inp[13]) ? node491 : 4'b1010;
								assign node491 = (inp[2]) ? 4'b1000 : node492;
									assign node492 = (inp[1]) ? node498 : node493;
										assign node493 = (inp[9]) ? node495 : 4'b1010;
											assign node495 = (inp[7]) ? 4'b1000 : 4'b1010;
										assign node498 = (inp[7]) ? node500 : 4'b1010;
											assign node500 = (inp[9]) ? node502 : 4'b1010;
												assign node502 = (inp[0]) ? 4'b1010 : 4'b1000;
					assign node506 = (inp[14]) ? node518 : node507;
						assign node507 = (inp[13]) ? 4'b1010 : node508;
							assign node508 = (inp[12]) ? 4'b1000 : node509;
								assign node509 = (inp[8]) ? node511 : 4'b1100;
									assign node511 = (inp[9]) ? node513 : 4'b1100;
										assign node513 = (inp[2]) ? 4'b1010 : 4'b1100;
						assign node518 = (inp[2]) ? node528 : node519;
							assign node519 = (inp[13]) ? 4'b1000 : node520;
								assign node520 = (inp[15]) ? node522 : 4'b1010;
									assign node522 = (inp[11]) ? node524 : 4'b1010;
										assign node524 = (inp[12]) ? 4'b1000 : 4'b1010;
							assign node528 = (inp[9]) ? 4'b1000 : node529;
								assign node529 = (inp[12]) ? 4'b1000 : node530;
									assign node530 = (inp[15]) ? 4'b1000 : node531;
										assign node531 = (inp[1]) ? 4'b1000 : node532;
											assign node532 = (inp[7]) ? 4'b1000 : 4'b1010;
				assign node539 = (inp[12]) ? node593 : node540;
					assign node540 = (inp[6]) ? node570 : node541;
						assign node541 = (inp[14]) ? node565 : node542;
							assign node542 = (inp[8]) ? node550 : node543;
								assign node543 = (inp[13]) ? 4'b1010 : node544;
									assign node544 = (inp[9]) ? 4'b1010 : node545;
										assign node545 = (inp[2]) ? 4'b1010 : 4'b1000;
								assign node550 = (inp[13]) ? node560 : node551;
									assign node551 = (inp[2]) ? 4'b1010 : node552;
										assign node552 = (inp[9]) ? 4'b1010 : node553;
											assign node553 = (inp[3]) ? node555 : 4'b1000;
												assign node555 = (inp[7]) ? 4'b1010 : 4'b1000;
									assign node560 = (inp[2]) ? node562 : 4'b1010;
										assign node562 = (inp[9]) ? 4'b1000 : 4'b1010;
							assign node565 = (inp[2]) ? node567 : 4'b1000;
								assign node567 = (inp[13]) ? 4'b1110 : 4'b1000;
						assign node570 = (inp[14]) ? node580 : node571;
							assign node571 = (inp[13]) ? node573 : 4'b1110;
								assign node573 = (inp[9]) ? 4'b1100 : node574;
									assign node574 = (inp[2]) ? 4'b1100 : node575;
										assign node575 = (inp[8]) ? 4'b1100 : 4'b1110;
							assign node580 = (inp[13]) ? 4'b1110 : node581;
								assign node581 = (inp[2]) ? node583 : 4'b1100;
									assign node583 = (inp[9]) ? 4'b1110 : node584;
										assign node584 = (inp[15]) ? node586 : 4'b1100;
											assign node586 = (inp[8]) ? node588 : 4'b1100;
												assign node588 = (inp[11]) ? 4'b1100 : 4'b1110;
					assign node593 = (inp[6]) ? node603 : node594;
						assign node594 = (inp[14]) ? node600 : node595;
							assign node595 = (inp[2]) ? node597 : 4'b1111;
								assign node597 = (inp[13]) ? 4'b1101 : 4'b1111;
							assign node600 = (inp[13]) ? 4'b1111 : 4'b1101;
						assign node603 = (inp[14]) ? node621 : node604;
							assign node604 = (inp[13]) ? node614 : node605;
								assign node605 = (inp[2]) ? 4'b1101 : node606;
									assign node606 = (inp[7]) ? node608 : 4'b1111;
										assign node608 = (inp[8]) ? node610 : 4'b1111;
											assign node610 = (inp[9]) ? 4'b1101 : 4'b1111;
								assign node614 = (inp[9]) ? node616 : 4'b1101;
									assign node616 = (inp[2]) ? node618 : 4'b1101;
										assign node618 = (inp[8]) ? 4'b1011 : 4'b1101;
							assign node621 = (inp[13]) ? node623 : 4'b1011;
								assign node623 = (inp[2]) ? 4'b1001 : node624;
									assign node624 = (inp[9]) ? node626 : 4'b1011;
										assign node626 = (inp[8]) ? 4'b1001 : node627;
											assign node627 = (inp[7]) ? 4'b1001 : 4'b1011;
			assign node632 = (inp[12]) ? node866 : node633;
				assign node633 = (inp[6]) ? node717 : node634;
					assign node634 = (inp[14]) ? node666 : node635;
						assign node635 = (inp[13]) ? node645 : node636;
							assign node636 = (inp[4]) ? node638 : 4'b0111;
								assign node638 = (inp[2]) ? 4'b0101 : node639;
									assign node639 = (inp[9]) ? node641 : 4'b0111;
										assign node641 = (inp[8]) ? 4'b0101 : 4'b0111;
							assign node645 = (inp[4]) ? node655 : node646;
								assign node646 = (inp[15]) ? node648 : 4'b0101;
									assign node648 = (inp[9]) ? node650 : 4'b0101;
										assign node650 = (inp[2]) ? node652 : 4'b0101;
											assign node652 = (inp[7]) ? 4'b0111 : 4'b0101;
								assign node655 = (inp[9]) ? 4'b0111 : node656;
									assign node656 = (inp[2]) ? 4'b0111 : node657;
										assign node657 = (inp[7]) ? node659 : 4'b0101;
											assign node659 = (inp[15]) ? node661 : 4'b0101;
												assign node661 = (inp[3]) ? 4'b0111 : 4'b0101;
						assign node666 = (inp[13]) ? node696 : node667;
							assign node667 = (inp[4]) ? node681 : node668;
								assign node668 = (inp[8]) ? node670 : 4'b0111;
									assign node670 = (inp[2]) ? node672 : 4'b0111;
										assign node672 = (inp[1]) ? node674 : 4'b0111;
											assign node674 = (inp[0]) ? 4'b0111 : node675;
												assign node675 = (inp[15]) ? 4'b0101 : node676;
													assign node676 = (inp[3]) ? 4'b0101 : 4'b0111;
								assign node681 = (inp[2]) ? node691 : node682;
									assign node682 = (inp[9]) ? 4'b0101 : node683;
										assign node683 = (inp[3]) ? 4'b0101 : node684;
											assign node684 = (inp[0]) ? 4'b0101 : node685;
												assign node685 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node691 = (inp[9]) ? node693 : 4'b0101;
										assign node693 = (inp[8]) ? 4'b0011 : 4'b0101;
							assign node696 = (inp[4]) ? node704 : node697;
								assign node697 = (inp[9]) ? node699 : 4'b0101;
									assign node699 = (inp[2]) ? node701 : 4'b0101;
										assign node701 = (inp[8]) ? 4'b0011 : 4'b0101;
								assign node704 = (inp[2]) ? node706 : 4'b0011;
									assign node706 = (inp[9]) ? 4'b0001 : node707;
										assign node707 = (inp[8]) ? node709 : 4'b0011;
											assign node709 = (inp[15]) ? node711 : 4'b0011;
												assign node711 = (inp[7]) ? 4'b0001 : node712;
													assign node712 = (inp[3]) ? 4'b0011 : 4'b0001;
					assign node717 = (inp[14]) ? node827 : node718;
						assign node718 = (inp[13]) ? node740 : node719;
							assign node719 = (inp[2]) ? node731 : node720;
								assign node720 = (inp[4]) ? node722 : 4'b0011;
									assign node722 = (inp[7]) ? node724 : 4'b0001;
										assign node724 = (inp[8]) ? node726 : 4'b0001;
											assign node726 = (inp[0]) ? 4'b0011 : node727;
												assign node727 = (inp[3]) ? 4'b0011 : 4'b0001;
								assign node731 = (inp[4]) ? 4'b0011 : node732;
									assign node732 = (inp[9]) ? node734 : 4'b0011;
										assign node734 = (inp[7]) ? 4'b0001 : node735;
											assign node735 = (inp[8]) ? 4'b0001 : 4'b0011;
							assign node740 = (inp[1]) ? node796 : node741;
								assign node741 = (inp[8]) ? node765 : node742;
									assign node742 = (inp[0]) ? node754 : node743;
										assign node743 = (inp[2]) ? node749 : node744;
											assign node744 = (inp[4]) ? node746 : 4'b0001;
												assign node746 = (inp[9]) ? 4'b0001 : 4'b0011;
											assign node749 = (inp[4]) ? 4'b0001 : node750;
												assign node750 = (inp[9]) ? 4'b0011 : 4'b0001;
										assign node754 = (inp[2]) ? node760 : node755;
											assign node755 = (inp[9]) ? 4'b0001 : node756;
												assign node756 = (inp[4]) ? 4'b0011 : 4'b0001;
											assign node760 = (inp[9]) ? node762 : 4'b0001;
												assign node762 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node765 = (inp[0]) ? node787 : node766;
										assign node766 = (inp[15]) ? node778 : node767;
											assign node767 = (inp[7]) ? node769 : 4'b0001;
												assign node769 = (inp[2]) ? node773 : node770;
													assign node770 = (inp[11]) ? 4'b0011 : 4'b0001;
													assign node773 = (inp[11]) ? 4'b0001 : node774;
														assign node774 = (inp[4]) ? 4'b0001 : 4'b0011;
											assign node778 = (inp[9]) ? 4'b0011 : node779;
												assign node779 = (inp[7]) ? node783 : node780;
													assign node780 = (inp[4]) ? 4'b0011 : 4'b0001;
													assign node783 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node787 = (inp[2]) ? node791 : node788;
											assign node788 = (inp[9]) ? 4'b0001 : 4'b0011;
											assign node791 = (inp[11]) ? 4'b0001 : node792;
												assign node792 = (inp[4]) ? 4'b0001 : 4'b0011;
								assign node796 = (inp[7]) ? node808 : node797;
									assign node797 = (inp[0]) ? 4'b0001 : node798;
										assign node798 = (inp[8]) ? 4'b0001 : node799;
											assign node799 = (inp[15]) ? 4'b0011 : node800;
												assign node800 = (inp[9]) ? 4'b0001 : node801;
													assign node801 = (inp[2]) ? 4'b0001 : 4'b0011;
									assign node808 = (inp[2]) ? node818 : node809;
										assign node809 = (inp[4]) ? node811 : 4'b0001;
											assign node811 = (inp[9]) ? 4'b0001 : node812;
												assign node812 = (inp[3]) ? node814 : 4'b0011;
													assign node814 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node818 = (inp[4]) ? 4'b0001 : node819;
											assign node819 = (inp[9]) ? 4'b0011 : node820;
												assign node820 = (inp[8]) ? node822 : 4'b0001;
													assign node822 = (inp[15]) ? 4'b0011 : 4'b0001;
						assign node827 = (inp[4]) ? node843 : node828;
							assign node828 = (inp[13]) ? node840 : node829;
								assign node829 = (inp[2]) ? node831 : 4'b0011;
									assign node831 = (inp[8]) ? 4'b0001 : node832;
										assign node832 = (inp[9]) ? 4'b0001 : node833;
											assign node833 = (inp[11]) ? node835 : 4'b0011;
												assign node835 = (inp[1]) ? 4'b0001 : 4'b0011;
								assign node840 = (inp[2]) ? 4'b0111 : 4'b0001;
							assign node843 = (inp[13]) ? node853 : node844;
								assign node844 = (inp[2]) ? node846 : 4'b0110;
									assign node846 = (inp[9]) ? 4'b0100 : node847;
										assign node847 = (inp[15]) ? node849 : 4'b0110;
											assign node849 = (inp[7]) ? 4'b0100 : 4'b0110;
								assign node853 = (inp[2]) ? 4'b0110 : node854;
									assign node854 = (inp[15]) ? node856 : 4'b0100;
										assign node856 = (inp[1]) ? node858 : 4'b0100;
											assign node858 = (inp[9]) ? node860 : 4'b0100;
												assign node860 = (inp[7]) ? node862 : 4'b0100;
													assign node862 = (inp[8]) ? 4'b0110 : 4'b0100;
				assign node866 = (inp[4]) ? node984 : node867;
					assign node867 = (inp[14]) ? node935 : node868;
						assign node868 = (inp[13]) ? node906 : node869;
							assign node869 = (inp[6]) ? node885 : node870;
								assign node870 = (inp[9]) ? node880 : node871;
									assign node871 = (inp[2]) ? 4'b0100 : node872;
										assign node872 = (inp[8]) ? node874 : 4'b0110;
											assign node874 = (inp[7]) ? 4'b0100 : node875;
												assign node875 = (inp[3]) ? 4'b0110 : 4'b0100;
									assign node880 = (inp[2]) ? node882 : 4'b0100;
										assign node882 = (inp[8]) ? 4'b0010 : 4'b0100;
								assign node885 = (inp[8]) ? node897 : node886;
									assign node886 = (inp[15]) ? node892 : node887;
										assign node887 = (inp[9]) ? 4'b0100 : node888;
											assign node888 = (inp[2]) ? 4'b0100 : 4'b0110;
										assign node892 = (inp[9]) ? 4'b0110 : node893;
											assign node893 = (inp[2]) ? 4'b0100 : 4'b0110;
									assign node897 = (inp[2]) ? node899 : 4'b0100;
										assign node899 = (inp[9]) ? 4'b0110 : node900;
											assign node900 = (inp[7]) ? node902 : 4'b0100;
												assign node902 = (inp[15]) ? 4'b0110 : 4'b0100;
							assign node906 = (inp[6]) ? node922 : node907;
								assign node907 = (inp[2]) ? node909 : 4'b0010;
									assign node909 = (inp[0]) ? node915 : node910;
										assign node910 = (inp[8]) ? 4'b0000 : node911;
											assign node911 = (inp[7]) ? 4'b0000 : 4'b0010;
										assign node915 = (inp[3]) ? node917 : 4'b0000;
											assign node917 = (inp[11]) ? node919 : 4'b0000;
												assign node919 = (inp[1]) ? 4'b0000 : 4'b0010;
								assign node922 = (inp[2]) ? node930 : node923;
									assign node923 = (inp[9]) ? node925 : 4'b0110;
										assign node925 = (inp[7]) ? 4'b0100 : node926;
											assign node926 = (inp[8]) ? 4'b0100 : 4'b0110;
									assign node930 = (inp[9]) ? node932 : 4'b0100;
										assign node932 = (inp[8]) ? 4'b0010 : 4'b0100;
						assign node935 = (inp[6]) ? node959 : node936;
							assign node936 = (inp[2]) ? node952 : node937;
								assign node937 = (inp[9]) ? node949 : node938;
									assign node938 = (inp[8]) ? node940 : 4'b0000;
										assign node940 = (inp[3]) ? 4'b0000 : node941;
											assign node941 = (inp[7]) ? node943 : 4'b0000;
												assign node943 = (inp[0]) ? 4'b0000 : node944;
													assign node944 = (inp[11]) ? 4'b0000 : 4'b0010;
									assign node949 = (inp[13]) ? 4'b0000 : 4'b0010;
								assign node952 = (inp[13]) ? 4'b0110 : node953;
									assign node953 = (inp[9]) ? node955 : 4'b0010;
										assign node955 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node959 = (inp[2]) ? node971 : node960;
								assign node960 = (inp[8]) ? node962 : 4'b0010;
									assign node962 = (inp[9]) ? node964 : 4'b0010;
										assign node964 = (inp[7]) ? 4'b0000 : node965;
											assign node965 = (inp[1]) ? node967 : 4'b0010;
												assign node967 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node971 = (inp[0]) ? node973 : 4'b0000;
									assign node973 = (inp[15]) ? node975 : 4'b0000;
										assign node975 = (inp[13]) ? 4'b0000 : node976;
											assign node976 = (inp[8]) ? node978 : 4'b0000;
												assign node978 = (inp[7]) ? node980 : 4'b0000;
													assign node980 = (inp[9]) ? 4'b0010 : 4'b0000;
					assign node984 = (inp[14]) ? node1056 : node985;
						assign node985 = (inp[13]) ? node1023 : node986;
							assign node986 = (inp[2]) ? node1002 : node987;
								assign node987 = (inp[6]) ? node995 : node988;
									assign node988 = (inp[11]) ? node990 : 4'b0111;
										assign node990 = (inp[3]) ? 4'b0111 : node991;
											assign node991 = (inp[9]) ? 4'b0101 : 4'b0111;
									assign node995 = (inp[9]) ? 4'b0111 : node996;
										assign node996 = (inp[7]) ? node998 : 4'b0101;
											assign node998 = (inp[15]) ? 4'b0111 : 4'b0101;
								assign node1002 = (inp[6]) ? node1010 : node1003;
									assign node1003 = (inp[1]) ? node1005 : 4'b0101;
										assign node1005 = (inp[15]) ? node1007 : 4'b0101;
											assign node1007 = (inp[3]) ? 4'b0111 : 4'b0101;
									assign node1010 = (inp[9]) ? node1020 : node1011;
										assign node1011 = (inp[7]) ? 4'b0101 : node1012;
											assign node1012 = (inp[8]) ? 4'b0101 : node1013;
												assign node1013 = (inp[11]) ? node1015 : 4'b0111;
													assign node1015 = (inp[1]) ? 4'b0101 : 4'b0111;
										assign node1020 = (inp[8]) ? 4'b0011 : 4'b0101;
							assign node1023 = (inp[6]) ? node1039 : node1024;
								assign node1024 = (inp[2]) ? node1034 : node1025;
									assign node1025 = (inp[8]) ? node1027 : 4'b0111;
										assign node1027 = (inp[9]) ? node1029 : 4'b0111;
											assign node1029 = (inp[7]) ? 4'b0101 : node1030;
												assign node1030 = (inp[11]) ? 4'b0101 : 4'b0111;
									assign node1034 = (inp[8]) ? node1036 : 4'b0101;
										assign node1036 = (inp[9]) ? 4'b0011 : 4'b0101;
								assign node1039 = (inp[9]) ? node1047 : node1040;
									assign node1040 = (inp[8]) ? node1042 : 4'b0011;
										assign node1042 = (inp[2]) ? 4'b0011 : node1043;
											assign node1043 = (inp[7]) ? 4'b0001 : 4'b0011;
									assign node1047 = (inp[15]) ? node1049 : 4'b0001;
										assign node1049 = (inp[2]) ? 4'b0001 : node1050;
											assign node1050 = (inp[7]) ? node1052 : 4'b0001;
												assign node1052 = (inp[8]) ? 4'b0011 : 4'b0001;
						assign node1056 = (inp[6]) ? node1080 : node1057;
							assign node1057 = (inp[2]) ? node1071 : node1058;
								assign node1058 = (inp[9]) ? node1064 : node1059;
									assign node1059 = (inp[8]) ? node1061 : 4'b0011;
										assign node1061 = (inp[13]) ? 4'b0001 : 4'b0011;
									assign node1064 = (inp[13]) ? 4'b0001 : node1065;
										assign node1065 = (inp[7]) ? 4'b0001 : node1066;
											assign node1066 = (inp[8]) ? 4'b0001 : 4'b0011;
								assign node1071 = (inp[13]) ? node1075 : node1072;
									assign node1072 = (inp[9]) ? 4'b0011 : 4'b0001;
									assign node1075 = (inp[8]) ? node1077 : 4'b0111;
										assign node1077 = (inp[9]) ? 4'b0101 : 4'b0111;
							assign node1080 = (inp[13]) ? node1102 : node1081;
								assign node1081 = (inp[9]) ? node1093 : node1082;
									assign node1082 = (inp[8]) ? node1084 : 4'b0110;
										assign node1084 = (inp[2]) ? node1086 : 4'b0110;
											assign node1086 = (inp[7]) ? 4'b0100 : node1087;
												assign node1087 = (inp[11]) ? node1089 : 4'b0110;
													assign node1089 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node1093 = (inp[8]) ? node1095 : 4'b0100;
										assign node1095 = (inp[2]) ? 4'b0010 : node1096;
											assign node1096 = (inp[7]) ? node1098 : 4'b0100;
												assign node1098 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node1102 = (inp[2]) ? node1116 : node1103;
									assign node1103 = (inp[8]) ? node1109 : node1104;
										assign node1104 = (inp[7]) ? node1106 : 4'b0010;
											assign node1106 = (inp[9]) ? 4'b0010 : 4'b0000;
										assign node1109 = (inp[7]) ? node1111 : 4'b0000;
											assign node1111 = (inp[15]) ? node1113 : 4'b0000;
												assign node1113 = (inp[9]) ? 4'b0000 : 4'b0010;
									assign node1116 = (inp[7]) ? node1128 : node1117;
										assign node1117 = (inp[8]) ? node1125 : node1118;
											assign node1118 = (inp[9]) ? node1120 : 4'b0110;
												assign node1120 = (inp[11]) ? node1122 : 4'b0110;
													assign node1122 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node1125 = (inp[15]) ? 4'b0100 : 4'b0010;
										assign node1128 = (inp[15]) ? node1134 : node1129;
											assign node1129 = (inp[8]) ? node1131 : 4'b0100;
												assign node1131 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node1134 = (inp[8]) ? 4'b0110 : 4'b0100;

endmodule