module dtc_split125_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node92 : node3;
			assign node3 = (inp[4]) ? node37 : node4;
				assign node4 = (inp[9]) ? node16 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[8]) ? 3'b100 : node7;
							assign node7 = (inp[11]) ? 3'b000 : node8;
								assign node8 = (inp[10]) ? 3'b100 : node9;
									assign node9 = (inp[7]) ? 3'b000 : 3'b100;
					assign node16 = (inp[8]) ? node26 : node17;
						assign node17 = (inp[1]) ? 3'b100 : node18;
							assign node18 = (inp[11]) ? node20 : 3'b000;
								assign node20 = (inp[3]) ? node22 : 3'b100;
									assign node22 = (inp[5]) ? 3'b100 : 3'b000;
						assign node26 = (inp[5]) ? node32 : node27;
							assign node27 = (inp[1]) ? 3'b000 : node28;
								assign node28 = (inp[10]) ? 3'b100 : 3'b000;
							assign node32 = (inp[1]) ? node34 : 3'b000;
								assign node34 = (inp[11]) ? 3'b100 : 3'b000;
				assign node37 = (inp[9]) ? node49 : node38;
					assign node38 = (inp[1]) ? node40 : 3'b100;
						assign node40 = (inp[8]) ? node44 : node41;
							assign node41 = (inp[11]) ? 3'b000 : 3'b100;
							assign node44 = (inp[10]) ? 3'b100 : node45;
								assign node45 = (inp[11]) ? 3'b000 : 3'b100;
					assign node49 = (inp[11]) ? node73 : node50;
						assign node50 = (inp[7]) ? node62 : node51;
							assign node51 = (inp[3]) ? node55 : node52;
								assign node52 = (inp[10]) ? 3'b111 : 3'b101;
								assign node55 = (inp[10]) ? node59 : node56;
									assign node56 = (inp[2]) ? 3'b000 : 3'b100;
									assign node59 = (inp[8]) ? 3'b000 : 3'b101;
							assign node62 = (inp[2]) ? node68 : node63;
								assign node63 = (inp[8]) ? node65 : 3'b001;
									assign node65 = (inp[10]) ? 3'b011 : 3'b001;
								assign node68 = (inp[8]) ? 3'b000 : node69;
									assign node69 = (inp[10]) ? 3'b101 : 3'b001;
						assign node73 = (inp[8]) ? node81 : node74;
							assign node74 = (inp[1]) ? node76 : 3'b101;
								assign node76 = (inp[10]) ? 3'b100 : node77;
									assign node77 = (inp[2]) ? 3'b000 : 3'b000;
							assign node81 = (inp[1]) ? node89 : node82;
								assign node82 = (inp[7]) ? node86 : node83;
									assign node83 = (inp[5]) ? 3'b100 : 3'b000;
									assign node86 = (inp[10]) ? 3'b010 : 3'b000;
								assign node89 = (inp[2]) ? 3'b000 : 3'b001;
			assign node92 = (inp[9]) ? node94 : 3'b000;
				assign node94 = (inp[1]) ? node122 : node95;
					assign node95 = (inp[4]) ? node101 : node96;
						assign node96 = (inp[11]) ? node98 : 3'b100;
							assign node98 = (inp[2]) ? 3'b100 : 3'b000;
						assign node101 = (inp[8]) ? node113 : node102;
							assign node102 = (inp[5]) ? node108 : node103;
								assign node103 = (inp[11]) ? 3'b100 : node104;
									assign node104 = (inp[10]) ? 3'b100 : 3'b000;
								assign node108 = (inp[2]) ? 3'b000 : node109;
									assign node109 = (inp[10]) ? 3'b000 : 3'b100;
							assign node113 = (inp[7]) ? node117 : node114;
								assign node114 = (inp[2]) ? 3'b001 : 3'b101;
								assign node117 = (inp[11]) ? node119 : 3'b001;
									assign node119 = (inp[10]) ? 3'b000 : 3'b101;
					assign node122 = (inp[4]) ? node124 : 3'b000;
						assign node124 = (inp[3]) ? node134 : node125;
							assign node125 = (inp[5]) ? node131 : node126;
								assign node126 = (inp[2]) ? node128 : 3'b100;
									assign node128 = (inp[8]) ? 3'b000 : 3'b100;
								assign node131 = (inp[8]) ? 3'b100 : 3'b000;
							assign node134 = (inp[11]) ? 3'b000 : node135;
								assign node135 = (inp[7]) ? node137 : 3'b100;
									assign node137 = (inp[10]) ? 3'b000 : 3'b000;

endmodule