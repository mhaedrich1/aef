module dtc_split33_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node230;

	assign outp = (inp[3]) ? node162 : node1;
		assign node1 = (inp[4]) ? node95 : node2;
			assign node2 = (inp[0]) ? node64 : node3;
				assign node3 = (inp[6]) ? node35 : node4;
					assign node4 = (inp[9]) ? node20 : node5;
						assign node5 = (inp[5]) ? node13 : node6;
							assign node6 = (inp[1]) ? node10 : node7;
								assign node7 = (inp[8]) ? 3'b100 : 3'b000;
								assign node10 = (inp[7]) ? 3'b110 : 3'b010;
							assign node13 = (inp[2]) ? node17 : node14;
								assign node14 = (inp[10]) ? 3'b000 : 3'b000;
								assign node17 = (inp[7]) ? 3'b100 : 3'b000;
						assign node20 = (inp[1]) ? node28 : node21;
							assign node21 = (inp[5]) ? node25 : node22;
								assign node22 = (inp[2]) ? 3'b110 : 3'b010;
								assign node25 = (inp[2]) ? 3'b000 : 3'b100;
							assign node28 = (inp[5]) ? node32 : node29;
								assign node29 = (inp[2]) ? 3'b101 : 3'b101;
								assign node32 = (inp[2]) ? 3'b111 : 3'b110;
					assign node35 = (inp[9]) ? node49 : node36;
						assign node36 = (inp[5]) ? node42 : node37;
							assign node37 = (inp[2]) ? 3'b011 : node38;
								assign node38 = (inp[1]) ? 3'b011 : 3'b011;
							assign node42 = (inp[1]) ? node46 : node43;
								assign node43 = (inp[7]) ? 3'b010 : 3'b011;
								assign node46 = (inp[7]) ? 3'b011 : 3'b011;
						assign node49 = (inp[5]) ? node57 : node50;
							assign node50 = (inp[10]) ? node54 : node51;
								assign node51 = (inp[11]) ? 3'b111 : 3'b011;
								assign node54 = (inp[1]) ? 3'b111 : 3'b111;
							assign node57 = (inp[7]) ? node61 : node58;
								assign node58 = (inp[11]) ? 3'b011 : 3'b101;
								assign node61 = (inp[2]) ? 3'b111 : 3'b011;
				assign node64 = (inp[6]) ? 3'b111 : node65;
					assign node65 = (inp[1]) ? node81 : node66;
						assign node66 = (inp[2]) ? node74 : node67;
							assign node67 = (inp[7]) ? node71 : node68;
								assign node68 = (inp[5]) ? 3'b110 : 3'b111;
								assign node71 = (inp[9]) ? 3'b011 : 3'b001;
							assign node74 = (inp[11]) ? node78 : node75;
								assign node75 = (inp[9]) ? 3'b011 : 3'b101;
								assign node78 = (inp[9]) ? 3'b111 : 3'b011;
						assign node81 = (inp[9]) ? node89 : node82;
							assign node82 = (inp[7]) ? node86 : node83;
								assign node83 = (inp[5]) ? 3'b101 : 3'b111;
								assign node86 = (inp[10]) ? 3'b111 : 3'b011;
							assign node89 = (inp[5]) ? node91 : 3'b111;
								assign node91 = (inp[7]) ? 3'b111 : 3'b111;
			assign node95 = (inp[0]) ? node125 : node96;
				assign node96 = (inp[6]) ? node112 : node97;
					assign node97 = (inp[9]) ? node99 : 3'b000;
						assign node99 = (inp[7]) ? node105 : node100;
							assign node100 = (inp[8]) ? node102 : 3'b000;
								assign node102 = (inp[11]) ? 3'b000 : 3'b000;
							assign node105 = (inp[10]) ? node109 : node106;
								assign node106 = (inp[1]) ? 3'b100 : 3'b000;
								assign node109 = (inp[2]) ? 3'b010 : 3'b100;
					assign node112 = (inp[1]) ? node114 : 3'b000;
						assign node114 = (inp[7]) ? node120 : node115;
							assign node115 = (inp[10]) ? node117 : 3'b000;
								assign node117 = (inp[8]) ? 3'b000 : 3'b000;
							assign node120 = (inp[9]) ? node122 : 3'b000;
								assign node122 = (inp[11]) ? 3'b001 : 3'b001;
				assign node125 = (inp[9]) ? node141 : node126;
					assign node126 = (inp[6]) ? 3'b000 : node127;
						assign node127 = (inp[7]) ? node135 : node128;
							assign node128 = (inp[8]) ? node132 : node129;
								assign node129 = (inp[2]) ? 3'b110 : 3'b100;
								assign node132 = (inp[10]) ? 3'b010 : 3'b000;
							assign node135 = (inp[2]) ? node137 : 3'b110;
								assign node137 = (inp[5]) ? 3'b110 : 3'b111;
					assign node141 = (inp[6]) ? node157 : node142;
						assign node142 = (inp[5]) ? node150 : node143;
							assign node143 = (inp[1]) ? node147 : node144;
								assign node144 = (inp[7]) ? 3'b101 : 3'b010;
								assign node147 = (inp[10]) ? 3'b111 : 3'b101;
							assign node150 = (inp[1]) ? node154 : node151;
								assign node151 = (inp[7]) ? 3'b110 : 3'b010;
								assign node154 = (inp[8]) ? 3'b100 : 3'b001;
						assign node157 = (inp[7]) ? 3'b111 : node158;
							assign node158 = (inp[10]) ? 3'b111 : 3'b011;
		assign node162 = (inp[0]) ? node176 : node163;
			assign node163 = (inp[9]) ? node165 : 3'b000;
				assign node165 = (inp[8]) ? node167 : 3'b000;
					assign node167 = (inp[7]) ? node169 : 3'b000;
						assign node169 = (inp[6]) ? 3'b000 : node170;
							assign node170 = (inp[11]) ? node172 : 3'b000;
								assign node172 = (inp[5]) ? 3'b000 : 3'b100;
			assign node176 = (inp[9]) ? node188 : node177;
				assign node177 = (inp[4]) ? 3'b000 : node178;
					assign node178 = (inp[6]) ? 3'b000 : node179;
						assign node179 = (inp[7]) ? 3'b100 : node180;
							assign node180 = (inp[5]) ? 3'b000 : node181;
								assign node181 = (inp[1]) ? 3'b100 : 3'b000;
				assign node188 = (inp[4]) ? node218 : node189;
					assign node189 = (inp[6]) ? node205 : node190;
						assign node190 = (inp[1]) ? node198 : node191;
							assign node191 = (inp[5]) ? node195 : node192;
								assign node192 = (inp[11]) ? 3'b000 : 3'b000;
								assign node195 = (inp[2]) ? 3'b000 : 3'b000;
							assign node198 = (inp[8]) ? node202 : node199;
								assign node199 = (inp[7]) ? 3'b110 : 3'b000;
								assign node202 = (inp[10]) ? 3'b010 : 3'b000;
						assign node205 = (inp[7]) ? node213 : node206;
							assign node206 = (inp[1]) ? node210 : node207;
								assign node207 = (inp[8]) ? 3'b011 : 3'b011;
								assign node210 = (inp[11]) ? 3'b001 : 3'b011;
							assign node213 = (inp[1]) ? 3'b101 : node214;
								assign node214 = (inp[8]) ? 3'b101 : 3'b100;
					assign node218 = (inp[1]) ? node220 : 3'b000;
						assign node220 = (inp[6]) ? node226 : node221;
							assign node221 = (inp[2]) ? node223 : 3'b000;
								assign node223 = (inp[5]) ? 3'b000 : 3'b100;
							assign node226 = (inp[5]) ? node230 : node227;
								assign node227 = (inp[7]) ? 3'b110 : 3'b100;
								assign node230 = (inp[11]) ? 3'b000 : 3'b000;

endmodule