module dtc_split25_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node17;
	wire [4-1:0] node18;
	wire [4-1:0] node22;
	wire [4-1:0] node24;
	wire [4-1:0] node27;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node56;
	wire [4-1:0] node59;
	wire [4-1:0] node60;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node66;
	wire [4-1:0] node69;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node76;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node88;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node102;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node117;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node129;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node144;
	wire [4-1:0] node147;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node165;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node176;
	wire [4-1:0] node177;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node191;
	wire [4-1:0] node193;
	wire [4-1:0] node196;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node207;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node215;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node222;
	wire [4-1:0] node225;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node234;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node241;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node255;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node285;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node305;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node316;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node329;
	wire [4-1:0] node333;
	wire [4-1:0] node335;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node347;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node364;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node372;
	wire [4-1:0] node373;
	wire [4-1:0] node376;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node395;
	wire [4-1:0] node399;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node428;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node437;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node457;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node464;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node473;
	wire [4-1:0] node475;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node493;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node506;
	wire [4-1:0] node509;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node530;
	wire [4-1:0] node533;
	wire [4-1:0] node535;
	wire [4-1:0] node537;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node547;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node563;
	wire [4-1:0] node564;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node571;
	wire [4-1:0] node574;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node587;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node611;
	wire [4-1:0] node613;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node623;
	wire [4-1:0] node626;
	wire [4-1:0] node629;
	wire [4-1:0] node631;
	wire [4-1:0] node633;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node648;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node664;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node685;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node698;
	wire [4-1:0] node700;
	wire [4-1:0] node702;
	wire [4-1:0] node704;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node712;
	wire [4-1:0] node715;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node738;
	wire [4-1:0] node740;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node750;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node775;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node789;
	wire [4-1:0] node791;
	wire [4-1:0] node794;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node806;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node812;
	wire [4-1:0] node814;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node822;
	wire [4-1:0] node825;
	wire [4-1:0] node826;
	wire [4-1:0] node830;
	wire [4-1:0] node832;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node868;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node880;
	wire [4-1:0] node881;
	wire [4-1:0] node883;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node896;
	wire [4-1:0] node897;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node916;
	wire [4-1:0] node919;
	wire [4-1:0] node922;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node939;
	wire [4-1:0] node941;
	wire [4-1:0] node943;
	wire [4-1:0] node945;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node957;
	wire [4-1:0] node959;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node966;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node984;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node994;
	wire [4-1:0] node996;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1003;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1011;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1018;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1062;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1075;
	wire [4-1:0] node1079;
	wire [4-1:0] node1081;
	wire [4-1:0] node1083;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1110;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1137;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1157;
	wire [4-1:0] node1162;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1169;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1179;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1205;
	wire [4-1:0] node1207;
	wire [4-1:0] node1209;
	wire [4-1:0] node1212;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1246;
	wire [4-1:0] node1248;
	wire [4-1:0] node1251;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1262;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1298;
	wire [4-1:0] node1299;
	wire [4-1:0] node1302;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1314;
	wire [4-1:0] node1318;
	wire [4-1:0] node1320;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1327;
	wire [4-1:0] node1329;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1336;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1352;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1358;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1378;
	wire [4-1:0] node1380;
	wire [4-1:0] node1382;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1388;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1395;
	wire [4-1:0] node1398;
	wire [4-1:0] node1399;
	wire [4-1:0] node1402;
	wire [4-1:0] node1405;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1446;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1454;
	wire [4-1:0] node1457;
	wire [4-1:0] node1458;
	wire [4-1:0] node1459;
	wire [4-1:0] node1463;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1470;
	wire [4-1:0] node1471;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1509;
	wire [4-1:0] node1513;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1518;
	wire [4-1:0] node1523;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1543;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1554;
	wire [4-1:0] node1555;
	wire [4-1:0] node1557;
	wire [4-1:0] node1560;
	wire [4-1:0] node1563;
	wire [4-1:0] node1565;
	wire [4-1:0] node1567;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1574;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1585;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1597;
	wire [4-1:0] node1599;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1613;
	wire [4-1:0] node1616;
	wire [4-1:0] node1618;
	wire [4-1:0] node1621;
	wire [4-1:0] node1623;
	wire [4-1:0] node1624;
	wire [4-1:0] node1627;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1635;
	wire [4-1:0] node1637;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1643;
	wire [4-1:0] node1646;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1653;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1662;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1674;
	wire [4-1:0] node1676;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1683;
	wire [4-1:0] node1685;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1703;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1713;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1719;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1729;
	wire [4-1:0] node1730;
	wire [4-1:0] node1734;
	wire [4-1:0] node1735;
	wire [4-1:0] node1737;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1746;
	wire [4-1:0] node1749;
	wire [4-1:0] node1750;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1759;
	wire [4-1:0] node1760;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1771;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1783;
	wire [4-1:0] node1786;
	wire [4-1:0] node1788;
	wire [4-1:0] node1789;
	wire [4-1:0] node1790;
	wire [4-1:0] node1792;
	wire [4-1:0] node1795;
	wire [4-1:0] node1797;
	wire [4-1:0] node1801;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1804;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1822;
	wire [4-1:0] node1823;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1839;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1851;
	wire [4-1:0] node1854;
	wire [4-1:0] node1855;
	wire [4-1:0] node1859;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1867;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1882;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1888;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1896;
	wire [4-1:0] node1897;
	wire [4-1:0] node1900;
	wire [4-1:0] node1903;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1909;
	wire [4-1:0] node1911;
	wire [4-1:0] node1913;
	wire [4-1:0] node1916;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1937;
	wire [4-1:0] node1938;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1946;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1957;
	wire [4-1:0] node1960;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1968;
	wire [4-1:0] node1971;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1995;
	wire [4-1:0] node1997;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2006;
	wire [4-1:0] node2008;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2026;
	wire [4-1:0] node2030;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2037;
	wire [4-1:0] node2040;
	wire [4-1:0] node2042;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2047;
	wire [4-1:0] node2049;
	wire [4-1:0] node2053;
	wire [4-1:0] node2054;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2062;
	wire [4-1:0] node2063;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2070;
	wire [4-1:0] node2072;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2080;
	wire [4-1:0] node2083;
	wire [4-1:0] node2085;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2095;
	wire [4-1:0] node2098;
	wire [4-1:0] node2100;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2119;
	wire [4-1:0] node2121;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2140;
	wire [4-1:0] node2142;
	wire [4-1:0] node2146;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2150;
	wire [4-1:0] node2153;
	wire [4-1:0] node2154;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2167;
	wire [4-1:0] node2170;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2180;
	wire [4-1:0] node2182;
	wire [4-1:0] node2184;
	wire [4-1:0] node2187;
	wire [4-1:0] node2188;
	wire [4-1:0] node2191;
	wire [4-1:0] node2194;
	wire [4-1:0] node2195;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2207;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2216;
	wire [4-1:0] node2219;
	wire [4-1:0] node2221;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2234;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2253;
	wire [4-1:0] node2256;
	wire [4-1:0] node2258;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2266;
	wire [4-1:0] node2268;
	wire [4-1:0] node2271;
	wire [4-1:0] node2272;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2280;
	wire [4-1:0] node2281;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2291;
	wire [4-1:0] node2293;
	wire [4-1:0] node2296;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;
	wire [4-1:0] node2314;
	wire [4-1:0] node2316;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2325;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2331;
	wire [4-1:0] node2333;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2343;
	wire [4-1:0] node2344;
	wire [4-1:0] node2345;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2350;
	wire [4-1:0] node2353;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2360;
	wire [4-1:0] node2362;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2376;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2383;
	wire [4-1:0] node2386;
	wire [4-1:0] node2387;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2390;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2399;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2410;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2421;
	wire [4-1:0] node2422;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2430;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2436;
	wire [4-1:0] node2438;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2446;
	wire [4-1:0] node2447;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2452;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2459;
	wire [4-1:0] node2462;
	wire [4-1:0] node2465;
	wire [4-1:0] node2466;
	wire [4-1:0] node2467;
	wire [4-1:0] node2468;
	wire [4-1:0] node2472;
	wire [4-1:0] node2475;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2481;
	wire [4-1:0] node2482;
	wire [4-1:0] node2486;
	wire [4-1:0] node2487;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2499;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2507;
	wire [4-1:0] node2510;
	wire [4-1:0] node2513;
	wire [4-1:0] node2515;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2533;
	wire [4-1:0] node2537;
	wire [4-1:0] node2539;
	wire [4-1:0] node2541;
	wire [4-1:0] node2544;
	wire [4-1:0] node2545;
	wire [4-1:0] node2546;
	wire [4-1:0] node2548;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2561;
	wire [4-1:0] node2564;
	wire [4-1:0] node2565;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2570;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2585;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2592;
	wire [4-1:0] node2593;
	wire [4-1:0] node2596;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2602;
	wire [4-1:0] node2605;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2616;
	wire [4-1:0] node2617;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2628;
	wire [4-1:0] node2629;
	wire [4-1:0] node2632;
	wire [4-1:0] node2635;
	wire [4-1:0] node2638;
	wire [4-1:0] node2639;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2649;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2657;
	wire [4-1:0] node2658;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2669;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2674;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2683;
	wire [4-1:0] node2686;
	wire [4-1:0] node2688;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2695;
	wire [4-1:0] node2697;
	wire [4-1:0] node2700;
	wire [4-1:0] node2703;
	wire [4-1:0] node2705;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2710;
	wire [4-1:0] node2711;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2716;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2725;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2738;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2743;
	wire [4-1:0] node2747;
	wire [4-1:0] node2748;
	wire [4-1:0] node2749;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2758;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2762;
	wire [4-1:0] node2766;
	wire [4-1:0] node2768;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2790;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2802;
	wire [4-1:0] node2804;
	wire [4-1:0] node2805;
	wire [4-1:0] node2809;
	wire [4-1:0] node2810;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2818;
	wire [4-1:0] node2819;
	wire [4-1:0] node2820;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2832;
	wire [4-1:0] node2833;
	wire [4-1:0] node2834;
	wire [4-1:0] node2837;
	wire [4-1:0] node2840;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2851;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2864;
	wire [4-1:0] node2867;
	wire [4-1:0] node2869;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2874;
	wire [4-1:0] node2875;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2889;
	wire [4-1:0] node2890;
	wire [4-1:0] node2891;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2897;
	wire [4-1:0] node2899;
	wire [4-1:0] node2902;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2915;
	wire [4-1:0] node2919;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2937;
	wire [4-1:0] node2940;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2946;
	wire [4-1:0] node2949;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2954;
	wire [4-1:0] node2957;
	wire [4-1:0] node2959;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2967;
	wire [4-1:0] node2971;
	wire [4-1:0] node2974;
	wire [4-1:0] node2975;
	wire [4-1:0] node2977;
	wire [4-1:0] node2980;
	wire [4-1:0] node2982;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2995;
	wire [4-1:0] node2996;
	wire [4-1:0] node2999;
	wire [4-1:0] node3001;
	wire [4-1:0] node3004;
	wire [4-1:0] node3006;
	wire [4-1:0] node3007;
	wire [4-1:0] node3008;
	wire [4-1:0] node3009;
	wire [4-1:0] node3014;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3020;
	wire [4-1:0] node3022;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3028;
	wire [4-1:0] node3030;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3055;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3061;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3076;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3087;
	wire [4-1:0] node3091;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3096;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3102;
	wire [4-1:0] node3104;
	wire [4-1:0] node3107;
	wire [4-1:0] node3110;
	wire [4-1:0] node3111;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3118;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3125;
	wire [4-1:0] node3127;
	wire [4-1:0] node3129;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3136;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3141;
	wire [4-1:0] node3144;
	wire [4-1:0] node3146;
	wire [4-1:0] node3148;
	wire [4-1:0] node3151;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3171;
	wire [4-1:0] node3174;
	wire [4-1:0] node3175;
	wire [4-1:0] node3179;
	wire [4-1:0] node3180;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3186;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3197;
	wire [4-1:0] node3201;
	wire [4-1:0] node3202;
	wire [4-1:0] node3206;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3218;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3225;
	wire [4-1:0] node3226;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3232;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3238;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3249;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3254;
	wire [4-1:0] node3255;
	wire [4-1:0] node3260;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3272;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3282;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3291;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3298;
	wire [4-1:0] node3299;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3307;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3313;
	wire [4-1:0] node3315;
	wire [4-1:0] node3317;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3331;
	wire [4-1:0] node3332;
	wire [4-1:0] node3333;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3343;
	wire [4-1:0] node3344;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3352;
	wire [4-1:0] node3356;
	wire [4-1:0] node3357;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3360;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3372;
	wire [4-1:0] node3373;
	wire [4-1:0] node3377;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3383;
	wire [4-1:0] node3384;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3402;
	wire [4-1:0] node3403;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3406;
	wire [4-1:0] node3410;
	wire [4-1:0] node3411;
	wire [4-1:0] node3415;
	wire [4-1:0] node3416;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3424;
	wire [4-1:0] node3425;
	wire [4-1:0] node3426;
	wire [4-1:0] node3427;
	wire [4-1:0] node3430;
	wire [4-1:0] node3433;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3440;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3448;
	wire [4-1:0] node3450;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3457;
	wire [4-1:0] node3458;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3470;
	wire [4-1:0] node3473;
	wire [4-1:0] node3476;
	wire [4-1:0] node3477;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3484;
	wire [4-1:0] node3488;
	wire [4-1:0] node3489;
	wire [4-1:0] node3490;
	wire [4-1:0] node3494;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3505;
	wire [4-1:0] node3507;
	wire [4-1:0] node3510;
	wire [4-1:0] node3513;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3516;
	wire [4-1:0] node3519;
	wire [4-1:0] node3521;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3527;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3535;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3544;
	wire [4-1:0] node3545;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3550;
	wire [4-1:0] node3553;
	wire [4-1:0] node3556;
	wire [4-1:0] node3557;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3563;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3570;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3578;
	wire [4-1:0] node3579;
	wire [4-1:0] node3580;
	wire [4-1:0] node3581;
	wire [4-1:0] node3582;
	wire [4-1:0] node3585;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3595;
	wire [4-1:0] node3596;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3607;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3612;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3618;
	wire [4-1:0] node3622;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3625;
	wire [4-1:0] node3629;
	wire [4-1:0] node3632;
	wire [4-1:0] node3635;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3640;
	wire [4-1:0] node3641;
	wire [4-1:0] node3645;
	wire [4-1:0] node3646;
	wire [4-1:0] node3648;
	wire [4-1:0] node3651;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3660;
	wire [4-1:0] node3663;
	wire [4-1:0] node3666;
	wire [4-1:0] node3668;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3675;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3684;
	wire [4-1:0] node3685;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3707;
	wire [4-1:0] node3708;
	wire [4-1:0] node3709;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3719;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3725;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3733;
	wire [4-1:0] node3736;
	wire [4-1:0] node3737;
	wire [4-1:0] node3738;
	wire [4-1:0] node3741;
	wire [4-1:0] node3745;
	wire [4-1:0] node3746;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3752;
	wire [4-1:0] node3753;
	wire [4-1:0] node3756;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3763;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3780;
	wire [4-1:0] node3783;
	wire [4-1:0] node3785;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3796;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3806;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3811;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3818;
	wire [4-1:0] node3819;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3832;
	wire [4-1:0] node3833;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3847;
	wire [4-1:0] node3848;
	wire [4-1:0] node3852;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3860;
	wire [4-1:0] node3861;
	wire [4-1:0] node3865;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3872;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3882;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3891;
	wire [4-1:0] node3894;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3900;
	wire [4-1:0] node3903;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3913;
	wire [4-1:0] node3916;
	wire [4-1:0] node3917;
	wire [4-1:0] node3919;
	wire [4-1:0] node3922;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3932;
	wire [4-1:0] node3934;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3942;
	wire [4-1:0] node3945;
	wire [4-1:0] node3948;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3951;
	wire [4-1:0] node3952;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3969;
	wire [4-1:0] node3970;
	wire [4-1:0] node3973;
	wire [4-1:0] node3975;
	wire [4-1:0] node3978;
	wire [4-1:0] node3979;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3985;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3997;
	wire [4-1:0] node4000;
	wire [4-1:0] node4003;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4006;
	wire [4-1:0] node4008;
	wire [4-1:0] node4011;
	wire [4-1:0] node4014;
	wire [4-1:0] node4015;
	wire [4-1:0] node4016;
	wire [4-1:0] node4020;
	wire [4-1:0] node4021;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4034;
	wire [4-1:0] node4036;
	wire [4-1:0] node4039;
	wire [4-1:0] node4041;
	wire [4-1:0] node4042;
	wire [4-1:0] node4045;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4059;
	wire [4-1:0] node4062;
	wire [4-1:0] node4063;
	wire [4-1:0] node4066;
	wire [4-1:0] node4068;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4075;
	wire [4-1:0] node4076;
	wire [4-1:0] node4080;
	wire [4-1:0] node4081;
	wire [4-1:0] node4082;
	wire [4-1:0] node4085;
	wire [4-1:0] node4089;
	wire [4-1:0] node4090;
	wire [4-1:0] node4091;
	wire [4-1:0] node4094;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4103;
	wire [4-1:0] node4105;
	wire [4-1:0] node4108;
	wire [4-1:0] node4109;
	wire [4-1:0] node4110;
	wire [4-1:0] node4115;
	wire [4-1:0] node4116;
	wire [4-1:0] node4120;
	wire [4-1:0] node4121;
	wire [4-1:0] node4122;
	wire [4-1:0] node4123;
	wire [4-1:0] node4126;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4138;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4147;
	wire [4-1:0] node4150;
	wire [4-1:0] node4151;
	wire [4-1:0] node4153;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4161;
	wire [4-1:0] node4162;
	wire [4-1:0] node4163;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4170;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4177;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4182;
	wire [4-1:0] node4184;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4190;
	wire [4-1:0] node4194;
	wire [4-1:0] node4195;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4210;
	wire [4-1:0] node4213;
	wire [4-1:0] node4215;
	wire [4-1:0] node4218;
	wire [4-1:0] node4219;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4227;
	wire [4-1:0] node4230;
	wire [4-1:0] node4233;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4243;
	wire [4-1:0] node4244;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4253;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4260;
	wire [4-1:0] node4264;
	wire [4-1:0] node4267;
	wire [4-1:0] node4268;
	wire [4-1:0] node4269;
	wire [4-1:0] node4272;
	wire [4-1:0] node4275;
	wire [4-1:0] node4276;
	wire [4-1:0] node4278;
	wire [4-1:0] node4281;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4295;
	wire [4-1:0] node4299;
	wire [4-1:0] node4302;
	wire [4-1:0] node4305;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4310;
	wire [4-1:0] node4311;
	wire [4-1:0] node4315;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4331;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4338;
	wire [4-1:0] node4341;
	wire [4-1:0] node4342;
	wire [4-1:0] node4346;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4353;
	wire [4-1:0] node4355;
	wire [4-1:0] node4358;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4362;
	wire [4-1:0] node4365;
	wire [4-1:0] node4368;
	wire [4-1:0] node4371;
	wire [4-1:0] node4372;
	wire [4-1:0] node4373;
	wire [4-1:0] node4374;
	wire [4-1:0] node4375;
	wire [4-1:0] node4377;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4384;
	wire [4-1:0] node4385;
	wire [4-1:0] node4387;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4397;
	wire [4-1:0] node4398;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4402;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4419;
	wire [4-1:0] node4420;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4429;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4437;
	wire [4-1:0] node4438;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4446;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4450;
	wire [4-1:0] node4453;
	wire [4-1:0] node4454;
	wire [4-1:0] node4457;
	wire [4-1:0] node4460;
	wire [4-1:0] node4461;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4478;
	wire [4-1:0] node4481;
	wire [4-1:0] node4484;
	wire [4-1:0] node4485;
	wire [4-1:0] node4486;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4494;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4500;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4507;
	wire [4-1:0] node4509;
	wire [4-1:0] node4513;
	wire [4-1:0] node4514;
	wire [4-1:0] node4518;
	wire [4-1:0] node4521;
	wire [4-1:0] node4522;
	wire [4-1:0] node4523;
	wire [4-1:0] node4526;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4533;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4539;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4550;
	wire [4-1:0] node4551;
	wire [4-1:0] node4556;
	wire [4-1:0] node4557;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4565;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4569;
	wire [4-1:0] node4572;
	wire [4-1:0] node4574;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4581;
	wire [4-1:0] node4583;
	wire [4-1:0] node4584;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4593;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4600;
	wire [4-1:0] node4601;
	wire [4-1:0] node4604;
	wire [4-1:0] node4607;
	wire [4-1:0] node4608;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4612;
	wire [4-1:0] node4616;
	wire [4-1:0] node4617;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4624;
	wire [4-1:0] node4626;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4633;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4649;
	wire [4-1:0] node4653;
	wire [4-1:0] node4654;
	wire [4-1:0] node4655;
	wire [4-1:0] node4656;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4662;
	wire [4-1:0] node4663;
	wire [4-1:0] node4664;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4672;
	wire [4-1:0] node4675;
	wire [4-1:0] node4676;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4682;
	wire [4-1:0] node4684;
	wire [4-1:0] node4685;
	wire [4-1:0] node4690;
	wire [4-1:0] node4691;
	wire [4-1:0] node4692;
	wire [4-1:0] node4694;
	wire [4-1:0] node4698;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4713;
	wire [4-1:0] node4716;
	wire [4-1:0] node4717;
	wire [4-1:0] node4718;
	wire [4-1:0] node4719;
	wire [4-1:0] node4724;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4746;
	wire [4-1:0] node4748;
	wire [4-1:0] node4751;
	wire [4-1:0] node4753;
	wire [4-1:0] node4755;
	wire [4-1:0] node4758;
	wire [4-1:0] node4759;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4765;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4772;
	wire [4-1:0] node4775;
	wire [4-1:0] node4776;
	wire [4-1:0] node4778;
	wire [4-1:0] node4781;
	wire [4-1:0] node4784;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4789;
	wire [4-1:0] node4790;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4802;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4810;
	wire [4-1:0] node4813;
	wire [4-1:0] node4815;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4821;
	wire [4-1:0] node4824;
	wire [4-1:0] node4825;
	wire [4-1:0] node4827;
	wire [4-1:0] node4830;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4835;
	wire [4-1:0] node4838;
	wire [4-1:0] node4839;
	wire [4-1:0] node4843;
	wire [4-1:0] node4844;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4849;
	wire [4-1:0] node4852;
	wire [4-1:0] node4855;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4862;
	wire [4-1:0] node4863;
	wire [4-1:0] node4864;
	wire [4-1:0] node4865;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4871;
	wire [4-1:0] node4874;
	wire [4-1:0] node4876;
	wire [4-1:0] node4878;
	wire [4-1:0] node4879;
	wire [4-1:0] node4881;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4895;
	wire [4-1:0] node4896;
	wire [4-1:0] node4899;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4919;
	wire [4-1:0] node4920;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4927;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4936;
	wire [4-1:0] node4939;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4944;
	wire [4-1:0] node4945;
	wire [4-1:0] node4948;
	wire [4-1:0] node4951;
	wire [4-1:0] node4952;
	wire [4-1:0] node4955;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4962;
	wire [4-1:0] node4964;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4977;
	wire [4-1:0] node4980;
	wire [4-1:0] node4983;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4989;
	wire [4-1:0] node4991;
	wire [4-1:0] node4994;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node4997;
	wire [4-1:0] node5000;
	wire [4-1:0] node5003;
	wire [4-1:0] node5005;
	wire [4-1:0] node5007;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5017;
	wire [4-1:0] node5019;
	wire [4-1:0] node5022;
	wire [4-1:0] node5024;
	wire [4-1:0] node5026;
	wire [4-1:0] node5029;
	wire [4-1:0] node5030;
	wire [4-1:0] node5031;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5038;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5042;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5050;
	wire [4-1:0] node5052;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5059;
	wire [4-1:0] node5062;
	wire [4-1:0] node5063;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5070;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5079;
	wire [4-1:0] node5082;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5089;
	wire [4-1:0] node5092;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5097;
	wire [4-1:0] node5100;
	wire [4-1:0] node5101;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5109;
	wire [4-1:0] node5110;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5115;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5124;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5130;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5138;
	wire [4-1:0] node5139;
	wire [4-1:0] node5140;
	wire [4-1:0] node5141;
	wire [4-1:0] node5142;
	wire [4-1:0] node5147;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5156;
	wire [4-1:0] node5158;
	wire [4-1:0] node5161;
	wire [4-1:0] node5164;
	wire [4-1:0] node5165;
	wire [4-1:0] node5166;
	wire [4-1:0] node5171;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5175;
	wire [4-1:0] node5176;
	wire [4-1:0] node5177;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5189;
	wire [4-1:0] node5192;
	wire [4-1:0] node5194;
	wire [4-1:0] node5197;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5214;
	wire [4-1:0] node5217;
	wire [4-1:0] node5221;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5228;
	wire [4-1:0] node5231;
	wire [4-1:0] node5233;
	wire [4-1:0] node5236;
	wire [4-1:0] node5237;
	wire [4-1:0] node5240;
	wire [4-1:0] node5243;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5257;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5265;
	wire [4-1:0] node5266;
	wire [4-1:0] node5269;
	wire [4-1:0] node5272;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5279;
	wire [4-1:0] node5282;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5288;
	wire [4-1:0] node5291;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5294;
	wire [4-1:0] node5297;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5308;
	wire [4-1:0] node5310;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5317;
	wire [4-1:0] node5318;
	wire [4-1:0] node5319;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5324;
	wire [4-1:0] node5326;
	wire [4-1:0] node5329;
	wire [4-1:0] node5330;
	wire [4-1:0] node5333;
	wire [4-1:0] node5334;
	wire [4-1:0] node5335;
	wire [4-1:0] node5338;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5345;
	wire [4-1:0] node5346;
	wire [4-1:0] node5348;
	wire [4-1:0] node5352;
	wire [4-1:0] node5353;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5358;
	wire [4-1:0] node5362;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5367;
	wire [4-1:0] node5368;
	wire [4-1:0] node5371;
	wire [4-1:0] node5372;
	wire [4-1:0] node5375;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5382;
	wire [4-1:0] node5383;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5399;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5406;
	wire [4-1:0] node5409;
	wire [4-1:0] node5410;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5415;
	wire [4-1:0] node5419;
	wire [4-1:0] node5421;
	wire [4-1:0] node5424;
	wire [4-1:0] node5425;
	wire [4-1:0] node5426;
	wire [4-1:0] node5427;
	wire [4-1:0] node5429;
	wire [4-1:0] node5430;
	wire [4-1:0] node5433;
	wire [4-1:0] node5434;
	wire [4-1:0] node5438;
	wire [4-1:0] node5439;
	wire [4-1:0] node5441;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5452;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5469;
	wire [4-1:0] node5470;
	wire [4-1:0] node5474;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5481;
	wire [4-1:0] node5484;
	wire [4-1:0] node5486;
	wire [4-1:0] node5487;
	wire [4-1:0] node5491;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5497;
	wire [4-1:0] node5500;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5507;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5516;
	wire [4-1:0] node5519;
	wire [4-1:0] node5521;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5528;
	wire [4-1:0] node5532;
	wire [4-1:0] node5535;
	wire [4-1:0] node5536;
	wire [4-1:0] node5537;
	wire [4-1:0] node5538;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5547;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5555;
	wire [4-1:0] node5558;
	wire [4-1:0] node5560;
	wire [4-1:0] node5563;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5568;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5577;
	wire [4-1:0] node5579;
	wire [4-1:0] node5582;
	wire [4-1:0] node5583;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5590;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5596;
	wire [4-1:0] node5597;
	wire [4-1:0] node5601;
	wire [4-1:0] node5602;
	wire [4-1:0] node5604;
	wire [4-1:0] node5607;
	wire [4-1:0] node5609;
	wire [4-1:0] node5612;
	wire [4-1:0] node5613;
	wire [4-1:0] node5614;
	wire [4-1:0] node5616;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5628;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5644;
	wire [4-1:0] node5645;
	wire [4-1:0] node5646;
	wire [4-1:0] node5649;
	wire [4-1:0] node5651;
	wire [4-1:0] node5654;
	wire [4-1:0] node5657;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5664;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5669;
	wire [4-1:0] node5670;
	wire [4-1:0] node5673;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5680;
	wire [4-1:0] node5682;
	wire [4-1:0] node5683;
	wire [4-1:0] node5684;
	wire [4-1:0] node5688;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5700;
	wire [4-1:0] node5703;
	wire [4-1:0] node5705;
	wire [4-1:0] node5706;
	wire [4-1:0] node5710;
	wire [4-1:0] node5712;
	wire [4-1:0] node5714;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5719;
	wire [4-1:0] node5720;
	wire [4-1:0] node5724;
	wire [4-1:0] node5725;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5735;
	wire [4-1:0] node5737;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5743;
	wire [4-1:0] node5744;
	wire [4-1:0] node5745;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5749;
	wire [4-1:0] node5753;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5762;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5769;
	wire [4-1:0] node5773;
	wire [4-1:0] node5774;
	wire [4-1:0] node5777;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5781;
	wire [4-1:0] node5785;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5790;
	wire [4-1:0] node5792;
	wire [4-1:0] node5793;
	wire [4-1:0] node5797;
	wire [4-1:0] node5799;
	wire [4-1:0] node5801;
	wire [4-1:0] node5804;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5807;
	wire [4-1:0] node5809;
	wire [4-1:0] node5813;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5820;
	wire [4-1:0] node5821;
	wire [4-1:0] node5822;
	wire [4-1:0] node5824;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5832;
	wire [4-1:0] node5833;
	wire [4-1:0] node5835;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5842;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5847;
	wire [4-1:0] node5851;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5856;
	wire [4-1:0] node5859;
	wire [4-1:0] node5861;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5867;
	wire [4-1:0] node5870;
	wire [4-1:0] node5871;
	wire [4-1:0] node5875;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5878;
	wire [4-1:0] node5879;
	wire [4-1:0] node5882;
	wire [4-1:0] node5885;
	wire [4-1:0] node5887;
	wire [4-1:0] node5888;
	wire [4-1:0] node5892;
	wire [4-1:0] node5893;
	wire [4-1:0] node5894;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5905;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5912;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5919;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5926;
	wire [4-1:0] node5927;
	wire [4-1:0] node5928;
	wire [4-1:0] node5932;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5939;
	wire [4-1:0] node5941;
	wire [4-1:0] node5944;
	wire [4-1:0] node5945;
	wire [4-1:0] node5946;
	wire [4-1:0] node5947;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5955;
	wire [4-1:0] node5958;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5961;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5971;
	wire [4-1:0] node5972;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5982;
	wire [4-1:0] node5983;
	wire [4-1:0] node5984;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5995;
	wire [4-1:0] node5996;
	wire [4-1:0] node5998;
	wire [4-1:0] node6001;
	wire [4-1:0] node6003;
	wire [4-1:0] node6004;
	wire [4-1:0] node6008;
	wire [4-1:0] node6009;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6016;
	wire [4-1:0] node6019;
	wire [4-1:0] node6020;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6028;
	wire [4-1:0] node6031;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6038;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6043;
	wire [4-1:0] node6047;
	wire [4-1:0] node6048;
	wire [4-1:0] node6050;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6059;
	wire [4-1:0] node6060;
	wire [4-1:0] node6064;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6068;
	wire [4-1:0] node6071;
	wire [4-1:0] node6074;
	wire [4-1:0] node6076;
	wire [4-1:0] node6077;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6085;
	wire [4-1:0] node6087;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6092;
	wire [4-1:0] node6095;
	wire [4-1:0] node6098;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6107;
	wire [4-1:0] node6108;
	wire [4-1:0] node6109;
	wire [4-1:0] node6111;
	wire [4-1:0] node6114;
	wire [4-1:0] node6115;
	wire [4-1:0] node6116;
	wire [4-1:0] node6120;
	wire [4-1:0] node6123;
	wire [4-1:0] node6124;
	wire [4-1:0] node6125;
	wire [4-1:0] node6127;
	wire [4-1:0] node6129;
	wire [4-1:0] node6132;
	wire [4-1:0] node6134;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6140;
	wire [4-1:0] node6143;
	wire [4-1:0] node6146;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6157;
	wire [4-1:0] node6158;
	wire [4-1:0] node6159;
	wire [4-1:0] node6162;
	wire [4-1:0] node6166;
	wire [4-1:0] node6167;
	wire [4-1:0] node6169;
	wire [4-1:0] node6172;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6179;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6185;
	wire [4-1:0] node6187;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6192;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6208;
	wire [4-1:0] node6210;
	wire [4-1:0] node6211;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6218;
	wire [4-1:0] node6220;
	wire [4-1:0] node6224;
	wire [4-1:0] node6225;
	wire [4-1:0] node6226;
	wire [4-1:0] node6227;
	wire [4-1:0] node6229;
	wire [4-1:0] node6231;
	wire [4-1:0] node6236;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6241;
	wire [4-1:0] node6247;
	wire [4-1:0] node6248;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6267;
	wire [4-1:0] node6268;
	wire [4-1:0] node6272;
	wire [4-1:0] node6274;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6280;
	wire [4-1:0] node6281;
	wire [4-1:0] node6283;
	wire [4-1:0] node6286;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6293;
	wire [4-1:0] node6297;
	wire [4-1:0] node6298;
	wire [4-1:0] node6300;
	wire [4-1:0] node6303;
	wire [4-1:0] node6306;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6309;
	wire [4-1:0] node6311;
	wire [4-1:0] node6314;
	wire [4-1:0] node6316;
	wire [4-1:0] node6319;
	wire [4-1:0] node6320;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6336;
	wire [4-1:0] node6337;
	wire [4-1:0] node6339;
	wire [4-1:0] node6342;
	wire [4-1:0] node6343;
	wire [4-1:0] node6347;
	wire [4-1:0] node6348;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6367;
	wire [4-1:0] node6369;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6380;
	wire [4-1:0] node6381;
	wire [4-1:0] node6382;
	wire [4-1:0] node6384;
	wire [4-1:0] node6388;
	wire [4-1:0] node6390;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6395;
	wire [4-1:0] node6396;
	wire [4-1:0] node6397;
	wire [4-1:0] node6400;
	wire [4-1:0] node6404;
	wire [4-1:0] node6405;
	wire [4-1:0] node6407;
	wire [4-1:0] node6408;
	wire [4-1:0] node6411;
	wire [4-1:0] node6414;
	wire [4-1:0] node6415;
	wire [4-1:0] node6419;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6423;
	wire [4-1:0] node6427;
	wire [4-1:0] node6429;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6434;
	wire [4-1:0] node6435;
	wire [4-1:0] node6436;
	wire [4-1:0] node6437;
	wire [4-1:0] node6438;
	wire [4-1:0] node6440;
	wire [4-1:0] node6443;
	wire [4-1:0] node6445;
	wire [4-1:0] node6447;
	wire [4-1:0] node6450;
	wire [4-1:0] node6451;
	wire [4-1:0] node6453;
	wire [4-1:0] node6457;
	wire [4-1:0] node6458;
	wire [4-1:0] node6461;
	wire [4-1:0] node6463;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6469;
	wire [4-1:0] node6471;
	wire [4-1:0] node6472;
	wire [4-1:0] node6478;
	wire [4-1:0] node6479;
	wire [4-1:0] node6480;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6486;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6493;
	wire [4-1:0] node6494;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6503;
	wire [4-1:0] node6504;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6512;
	wire [4-1:0] node6514;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6520;
	wire [4-1:0] node6523;
	wire [4-1:0] node6525;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6530;
	wire [4-1:0] node6532;
	wire [4-1:0] node6533;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6540;
	wire [4-1:0] node6544;
	wire [4-1:0] node6545;
	wire [4-1:0] node6547;
	wire [4-1:0] node6551;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6554;
	wire [4-1:0] node6555;
	wire [4-1:0] node6556;
	wire [4-1:0] node6561;
	wire [4-1:0] node6563;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6573;
	wire [4-1:0] node6574;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6583;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6596;
	wire [4-1:0] node6597;
	wire [4-1:0] node6598;
	wire [4-1:0] node6599;
	wire [4-1:0] node6602;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6607;
	wire [4-1:0] node6608;
	wire [4-1:0] node6613;
	wire [4-1:0] node6615;
	wire [4-1:0] node6616;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6623;
	wire [4-1:0] node6624;
	wire [4-1:0] node6627;
	wire [4-1:0] node6630;
	wire [4-1:0] node6631;
	wire [4-1:0] node6633;
	wire [4-1:0] node6636;
	wire [4-1:0] node6638;
	wire [4-1:0] node6639;
	wire [4-1:0] node6643;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6648;
	wire [4-1:0] node6650;
	wire [4-1:0] node6652;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6666;
	wire [4-1:0] node6669;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6675;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6684;
	wire [4-1:0] node6685;
	wire [4-1:0] node6686;
	wire [4-1:0] node6687;
	wire [4-1:0] node6689;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6698;
	wire [4-1:0] node6699;
	wire [4-1:0] node6702;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6710;
	wire [4-1:0] node6711;
	wire [4-1:0] node6712;
	wire [4-1:0] node6715;
	wire [4-1:0] node6719;
	wire [4-1:0] node6720;
	wire [4-1:0] node6722;
	wire [4-1:0] node6725;
	wire [4-1:0] node6727;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6735;
	wire [4-1:0] node6738;
	wire [4-1:0] node6741;
	wire [4-1:0] node6743;
	wire [4-1:0] node6745;
	wire [4-1:0] node6748;
	wire [4-1:0] node6749;
	wire [4-1:0] node6751;
	wire [4-1:0] node6753;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6769;
	wire [4-1:0] node6770;
	wire [4-1:0] node6774;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6785;
	wire [4-1:0] node6787;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6800;
	wire [4-1:0] node6803;
	wire [4-1:0] node6804;
	wire [4-1:0] node6808;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6817;
	wire [4-1:0] node6818;
	wire [4-1:0] node6823;
	wire [4-1:0] node6824;
	wire [4-1:0] node6825;
	wire [4-1:0] node6826;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6833;
	wire [4-1:0] node6835;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6841;
	wire [4-1:0] node6844;
	wire [4-1:0] node6845;
	wire [4-1:0] node6847;
	wire [4-1:0] node6850;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6856;
	wire [4-1:0] node6857;
	wire [4-1:0] node6858;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6879;
	wire [4-1:0] node6881;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6887;
	wire [4-1:0] node6888;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6895;
	wire [4-1:0] node6896;
	wire [4-1:0] node6899;
	wire [4-1:0] node6900;
	wire [4-1:0] node6901;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6922;
	wire [4-1:0] node6924;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6934;
	wire [4-1:0] node6935;
	wire [4-1:0] node6938;
	wire [4-1:0] node6941;
	wire [4-1:0] node6944;
	wire [4-1:0] node6945;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6951;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6959;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6969;
	wire [4-1:0] node6970;
	wire [4-1:0] node6973;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6980;
	wire [4-1:0] node6984;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6991;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6994;
	wire [4-1:0] node6998;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7005;
	wire [4-1:0] node7006;
	wire [4-1:0] node7007;
	wire [4-1:0] node7011;
	wire [4-1:0] node7014;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7023;
	wire [4-1:0] node7024;
	wire [4-1:0] node7026;
	wire [4-1:0] node7027;
	wire [4-1:0] node7029;
	wire [4-1:0] node7034;
	wire [4-1:0] node7035;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7041;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7050;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7055;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7065;
	wire [4-1:0] node7067;
	wire [4-1:0] node7070;
	wire [4-1:0] node7072;
	wire [4-1:0] node7073;
	wire [4-1:0] node7076;
	wire [4-1:0] node7079;
	wire [4-1:0] node7081;
	wire [4-1:0] node7084;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7094;
	wire [4-1:0] node7096;
	wire [4-1:0] node7099;
	wire [4-1:0] node7100;
	wire [4-1:0] node7101;
	wire [4-1:0] node7102;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7109;
	wire [4-1:0] node7110;
	wire [4-1:0] node7114;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7122;
	wire [4-1:0] node7125;
	wire [4-1:0] node7126;
	wire [4-1:0] node7127;
	wire [4-1:0] node7129;
	wire [4-1:0] node7130;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7137;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7145;
	wire [4-1:0] node7146;
	wire [4-1:0] node7150;
	wire [4-1:0] node7151;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7154;
	wire [4-1:0] node7155;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7160;
	wire [4-1:0] node7164;
	wire [4-1:0] node7165;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7178;
	wire [4-1:0] node7179;
	wire [4-1:0] node7183;
	wire [4-1:0] node7184;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7196;
	wire [4-1:0] node7198;
	wire [4-1:0] node7201;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7208;
	wire [4-1:0] node7209;
	wire [4-1:0] node7212;
	wire [4-1:0] node7215;
	wire [4-1:0] node7217;
	wire [4-1:0] node7218;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7228;
	wire [4-1:0] node7229;
	wire [4-1:0] node7230;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7236;
	wire [4-1:0] node7239;
	wire [4-1:0] node7242;
	wire [4-1:0] node7244;
	wire [4-1:0] node7247;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7255;
	wire [4-1:0] node7258;
	wire [4-1:0] node7260;
	wire [4-1:0] node7262;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7270;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7279;
	wire [4-1:0] node7281;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7286;
	wire [4-1:0] node7287;
	wire [4-1:0] node7291;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7299;
	wire [4-1:0] node7302;
	wire [4-1:0] node7303;
	wire [4-1:0] node7305;
	wire [4-1:0] node7308;
	wire [4-1:0] node7309;
	wire [4-1:0] node7311;
	wire [4-1:0] node7314;
	wire [4-1:0] node7317;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7320;
	wire [4-1:0] node7323;
	wire [4-1:0] node7326;
	wire [4-1:0] node7327;
	wire [4-1:0] node7328;
	wire [4-1:0] node7329;
	wire [4-1:0] node7330;
	wire [4-1:0] node7331;
	wire [4-1:0] node7337;
	wire [4-1:0] node7338;
	wire [4-1:0] node7339;
	wire [4-1:0] node7342;
	wire [4-1:0] node7346;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7351;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7366;
	wire [4-1:0] node7370;
	wire [4-1:0] node7373;
	wire [4-1:0] node7374;
	wire [4-1:0] node7376;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7383;
	wire [4-1:0] node7384;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7390;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7396;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7404;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7408;
	wire [4-1:0] node7409;
	wire [4-1:0] node7410;
	wire [4-1:0] node7411;
	wire [4-1:0] node7412;
	wire [4-1:0] node7415;
	wire [4-1:0] node7418;
	wire [4-1:0] node7420;
	wire [4-1:0] node7423;
	wire [4-1:0] node7424;
	wire [4-1:0] node7425;
	wire [4-1:0] node7426;
	wire [4-1:0] node7427;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7437;
	wire [4-1:0] node7439;
	wire [4-1:0] node7441;
	wire [4-1:0] node7444;
	wire [4-1:0] node7445;
	wire [4-1:0] node7446;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7457;
	wire [4-1:0] node7458;
	wire [4-1:0] node7461;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7467;
	wire [4-1:0] node7471;
	wire [4-1:0] node7473;
	wire [4-1:0] node7476;
	wire [4-1:0] node7477;
	wire [4-1:0] node7480;
	wire [4-1:0] node7483;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7489;
	wire [4-1:0] node7491;
	wire [4-1:0] node7495;
	wire [4-1:0] node7496;
	wire [4-1:0] node7498;
	wire [4-1:0] node7501;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7506;
	wire [4-1:0] node7509;
	wire [4-1:0] node7512;
	wire [4-1:0] node7513;
	wire [4-1:0] node7514;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7524;
	wire [4-1:0] node7528;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7531;
	wire [4-1:0] node7535;
	wire [4-1:0] node7538;
	wire [4-1:0] node7539;
	wire [4-1:0] node7541;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7547;
	wire [4-1:0] node7550;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7559;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7568;
	wire [4-1:0] node7569;
	wire [4-1:0] node7573;
	wire [4-1:0] node7574;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7581;
	wire [4-1:0] node7583;
	wire [4-1:0] node7586;
	wire [4-1:0] node7587;
	wire [4-1:0] node7588;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7596;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7603;
	wire [4-1:0] node7605;
	wire [4-1:0] node7607;
	wire [4-1:0] node7610;
	wire [4-1:0] node7612;
	wire [4-1:0] node7613;
	wire [4-1:0] node7615;
	wire [4-1:0] node7619;
	wire [4-1:0] node7620;
	wire [4-1:0] node7621;
	wire [4-1:0] node7622;
	wire [4-1:0] node7626;
	wire [4-1:0] node7627;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7646;
	wire [4-1:0] node7647;
	wire [4-1:0] node7648;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7652;
	wire [4-1:0] node7655;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7662;
	wire [4-1:0] node7665;
	wire [4-1:0] node7666;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7674;
	wire [4-1:0] node7677;
	wire [4-1:0] node7678;
	wire [4-1:0] node7679;
	wire [4-1:0] node7681;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7688;
	wire [4-1:0] node7691;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7701;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7711;
	wire [4-1:0] node7713;
	wire [4-1:0] node7716;
	wire [4-1:0] node7717;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7723;
	wire [4-1:0] node7726;
	wire [4-1:0] node7727;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7743;
	wire [4-1:0] node7744;
	wire [4-1:0] node7745;
	wire [4-1:0] node7748;
	wire [4-1:0] node7749;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7756;
	wire [4-1:0] node7758;
	wire [4-1:0] node7761;
	wire [4-1:0] node7763;
	wire [4-1:0] node7766;
	wire [4-1:0] node7769;
	wire [4-1:0] node7770;
	wire [4-1:0] node7771;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7777;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7784;
	wire [4-1:0] node7787;
	wire [4-1:0] node7789;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7797;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7802;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7810;
	wire [4-1:0] node7811;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7815;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7822;
	wire [4-1:0] node7824;
	wire [4-1:0] node7825;
	wire [4-1:0] node7829;
	wire [4-1:0] node7831;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7836;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7842;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7849;
	wire [4-1:0] node7851;
	wire [4-1:0] node7853;
	wire [4-1:0] node7856;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7859;
	wire [4-1:0] node7862;
	wire [4-1:0] node7866;
	wire [4-1:0] node7868;
	wire [4-1:0] node7871;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7876;
	wire [4-1:0] node7878;
	wire [4-1:0] node7882;
	wire [4-1:0] node7883;
	wire [4-1:0] node7885;
	wire [4-1:0] node7888;
	wire [4-1:0] node7891;
	wire [4-1:0] node7892;
	wire [4-1:0] node7894;
	wire [4-1:0] node7897;
	wire [4-1:0] node7899;
	wire [4-1:0] node7902;
	wire [4-1:0] node7903;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7917;
	wire [4-1:0] node7919;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7927;
	wire [4-1:0] node7930;
	wire [4-1:0] node7933;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7936;
	wire [4-1:0] node7938;
	wire [4-1:0] node7939;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7955;
	wire [4-1:0] node7957;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7962;
	wire [4-1:0] node7965;
	wire [4-1:0] node7968;
	wire [4-1:0] node7971;
	wire [4-1:0] node7972;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7978;
	wire [4-1:0] node7982;
	wire [4-1:0] node7983;
	wire [4-1:0] node7986;
	wire [4-1:0] node7988;
	wire [4-1:0] node7991;
	wire [4-1:0] node7992;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7998;
	wire [4-1:0] node8000;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8006;
	wire [4-1:0] node8007;
	wire [4-1:0] node8011;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8017;
	wire [4-1:0] node8018;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8033;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8048;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8058;
	wire [4-1:0] node8061;
	wire [4-1:0] node8062;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8068;
	wire [4-1:0] node8071;
	wire [4-1:0] node8073;
	wire [4-1:0] node8075;
	wire [4-1:0] node8077;
	wire [4-1:0] node8080;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8087;
	wire [4-1:0] node8090;
	wire [4-1:0] node8093;
	wire [4-1:0] node8094;
	wire [4-1:0] node8098;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8103;
	wire [4-1:0] node8107;
	wire [4-1:0] node8108;
	wire [4-1:0] node8109;
	wire [4-1:0] node8110;
	wire [4-1:0] node8114;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8127;
	wire [4-1:0] node8128;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8138;
	wire [4-1:0] node8139;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8153;
	wire [4-1:0] node8156;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8162;
	wire [4-1:0] node8163;
	wire [4-1:0] node8165;
	wire [4-1:0] node8169;
	wire [4-1:0] node8171;
	wire [4-1:0] node8173;
	wire [4-1:0] node8176;
	wire [4-1:0] node8178;
	wire [4-1:0] node8181;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8184;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8191;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8195;
	wire [4-1:0] node8198;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8211;
	wire [4-1:0] node8212;
	wire [4-1:0] node8213;
	wire [4-1:0] node8215;
	wire [4-1:0] node8216;
	wire [4-1:0] node8218;
	wire [4-1:0] node8222;
	wire [4-1:0] node8225;
	wire [4-1:0] node8226;
	wire [4-1:0] node8227;
	wire [4-1:0] node8231;
	wire [4-1:0] node8233;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8242;
	wire [4-1:0] node8245;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8256;
	wire [4-1:0] node8257;
	wire [4-1:0] node8258;
	wire [4-1:0] node8261;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8275;
	wire [4-1:0] node8276;
	wire [4-1:0] node8279;
	wire [4-1:0] node8282;
	wire [4-1:0] node8283;
	wire [4-1:0] node8285;
	wire [4-1:0] node8287;
	wire [4-1:0] node8291;
	wire [4-1:0] node8293;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8308;
	wire [4-1:0] node8313;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8318;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8325;
	wire [4-1:0] node8327;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8335;
	wire [4-1:0] node8337;
	wire [4-1:0] node8340;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8345;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8352;
	wire [4-1:0] node8353;
	wire [4-1:0] node8355;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8361;
	wire [4-1:0] node8364;
	wire [4-1:0] node8366;
	wire [4-1:0] node8369;
	wire [4-1:0] node8372;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8375;
	wire [4-1:0] node8377;
	wire [4-1:0] node8380;
	wire [4-1:0] node8383;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8387;
	wire [4-1:0] node8391;
	wire [4-1:0] node8393;
	wire [4-1:0] node8394;
	wire [4-1:0] node8398;
	wire [4-1:0] node8399;
	wire [4-1:0] node8400;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8406;
	wire [4-1:0] node8411;
	wire [4-1:0] node8412;
	wire [4-1:0] node8413;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8418;
	wire [4-1:0] node8421;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8428;
	wire [4-1:0] node8429;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8437;
	wire [4-1:0] node8438;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8448;
	wire [4-1:0] node8449;
	wire [4-1:0] node8453;
	wire [4-1:0] node8454;
	wire [4-1:0] node8458;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8468;
	wire [4-1:0] node8471;
	wire [4-1:0] node8472;
	wire [4-1:0] node8476;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8484;
	wire [4-1:0] node8485;
	wire [4-1:0] node8486;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8495;
	wire [4-1:0] node8496;
	wire [4-1:0] node8499;
	wire [4-1:0] node8500;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8510;
	wire [4-1:0] node8514;
	wire [4-1:0] node8515;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8529;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8540;
	wire [4-1:0] node8543;
	wire [4-1:0] node8546;
	wire [4-1:0] node8547;
	wire [4-1:0] node8550;
	wire [4-1:0] node8551;
	wire [4-1:0] node8553;
	wire [4-1:0] node8556;
	wire [4-1:0] node8559;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8564;
	wire [4-1:0] node8565;
	wire [4-1:0] node8569;
	wire [4-1:0] node8570;
	wire [4-1:0] node8571;
	wire [4-1:0] node8573;
	wire [4-1:0] node8576;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8588;
	wire [4-1:0] node8590;
	wire [4-1:0] node8593;
	wire [4-1:0] node8594;
	wire [4-1:0] node8597;
	wire [4-1:0] node8600;
	wire [4-1:0] node8601;
	wire [4-1:0] node8602;
	wire [4-1:0] node8606;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8611;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8614;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8622;
	wire [4-1:0] node8623;
	wire [4-1:0] node8624;
	wire [4-1:0] node8628;
	wire [4-1:0] node8629;
	wire [4-1:0] node8630;
	wire [4-1:0] node8633;
	wire [4-1:0] node8636;
	wire [4-1:0] node8638;
	wire [4-1:0] node8641;
	wire [4-1:0] node8642;
	wire [4-1:0] node8644;
	wire [4-1:0] node8647;
	wire [4-1:0] node8648;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8659;
	wire [4-1:0] node8660;
	wire [4-1:0] node8661;
	wire [4-1:0] node8666;
	wire [4-1:0] node8667;
	wire [4-1:0] node8669;
	wire [4-1:0] node8671;
	wire [4-1:0] node8674;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8690;
	wire [4-1:0] node8692;
	wire [4-1:0] node8693;
	wire [4-1:0] node8694;
	wire [4-1:0] node8698;
	wire [4-1:0] node8701;
	wire [4-1:0] node8702;
	wire [4-1:0] node8704;
	wire [4-1:0] node8707;
	wire [4-1:0] node8709;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8715;
	wire [4-1:0] node8718;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8726;
	wire [4-1:0] node8728;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8737;
	wire [4-1:0] node8738;
	wire [4-1:0] node8739;
	wire [4-1:0] node8741;
	wire [4-1:0] node8743;
	wire [4-1:0] node8744;
	wire [4-1:0] node8747;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8753;
	wire [4-1:0] node8754;
	wire [4-1:0] node8759;
	wire [4-1:0] node8760;
	wire [4-1:0] node8761;
	wire [4-1:0] node8762;
	wire [4-1:0] node8765;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8772;
	wire [4-1:0] node8773;
	wire [4-1:0] node8774;
	wire [4-1:0] node8775;
	wire [4-1:0] node8778;
	wire [4-1:0] node8780;
	wire [4-1:0] node8783;
	wire [4-1:0] node8784;
	wire [4-1:0] node8786;
	wire [4-1:0] node8789;
	wire [4-1:0] node8791;
	wire [4-1:0] node8794;
	wire [4-1:0] node8795;
	wire [4-1:0] node8796;
	wire [4-1:0] node8799;
	wire [4-1:0] node8802;
	wire [4-1:0] node8804;
	wire [4-1:0] node8805;
	wire [4-1:0] node8806;
	wire [4-1:0] node8811;
	wire [4-1:0] node8812;
	wire [4-1:0] node8813;
	wire [4-1:0] node8814;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8821;
	wire [4-1:0] node8823;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8832;
	wire [4-1:0] node8835;
	wire [4-1:0] node8836;
	wire [4-1:0] node8837;
	wire [4-1:0] node8840;
	wire [4-1:0] node8842;
	wire [4-1:0] node8844;
	wire [4-1:0] node8845;
	wire [4-1:0] node8848;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8858;
	wire [4-1:0] node8861;
	wire [4-1:0] node8863;
	wire [4-1:0] node8866;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8875;
	wire [4-1:0] node8877;
	wire [4-1:0] node8879;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8892;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8899;
	wire [4-1:0] node8901;
	wire [4-1:0] node8905;
	wire [4-1:0] node8906;
	wire [4-1:0] node8907;
	wire [4-1:0] node8910;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8916;
	wire [4-1:0] node8917;
	wire [4-1:0] node8918;
	wire [4-1:0] node8922;
	wire [4-1:0] node8924;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8932;
	wire [4-1:0] node8935;
	wire [4-1:0] node8937;
	wire [4-1:0] node8940;
	wire [4-1:0] node8941;
	wire [4-1:0] node8942;
	wire [4-1:0] node8945;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8951;
	wire [4-1:0] node8954;
	wire [4-1:0] node8956;
	wire [4-1:0] node8959;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8967;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8988;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8993;
	wire [4-1:0] node8994;
	wire [4-1:0] node8995;
	wire [4-1:0] node8996;
	wire [4-1:0] node8998;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9008;
	wire [4-1:0] node9010;
	wire [4-1:0] node9013;
	wire [4-1:0] node9014;
	wire [4-1:0] node9015;
	wire [4-1:0] node9017;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9023;
	wire [4-1:0] node9026;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9033;
	wire [4-1:0] node9036;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9045;
	wire [4-1:0] node9049;
	wire [4-1:0] node9050;
	wire [4-1:0] node9051;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9058;
	wire [4-1:0] node9059;
	wire [4-1:0] node9063;
	wire [4-1:0] node9064;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9070;
	wire [4-1:0] node9073;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9079;
	wire [4-1:0] node9082;
	wire [4-1:0] node9083;
	wire [4-1:0] node9085;
	wire [4-1:0] node9086;
	wire [4-1:0] node9088;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9095;
	wire [4-1:0] node9098;
	wire [4-1:0] node9099;
	wire [4-1:0] node9100;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9107;
	wire [4-1:0] node9109;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9119;
	wire [4-1:0] node9123;
	wire [4-1:0] node9124;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9134;
	wire [4-1:0] node9137;
	wire [4-1:0] node9138;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9147;
	wire [4-1:0] node9151;
	wire [4-1:0] node9154;
	wire [4-1:0] node9155;
	wire [4-1:0] node9156;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9167;
	wire [4-1:0] node9169;
	wire [4-1:0] node9171;
	wire [4-1:0] node9174;
	wire [4-1:0] node9175;
	wire [4-1:0] node9176;
	wire [4-1:0] node9179;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9187;
	wire [4-1:0] node9188;
	wire [4-1:0] node9189;
	wire [4-1:0] node9191;
	wire [4-1:0] node9193;
	wire [4-1:0] node9196;
	wire [4-1:0] node9197;
	wire [4-1:0] node9199;
	wire [4-1:0] node9201;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9209;
	wire [4-1:0] node9211;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9222;
	wire [4-1:0] node9223;
	wire [4-1:0] node9227;
	wire [4-1:0] node9228;
	wire [4-1:0] node9229;
	wire [4-1:0] node9231;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9242;
	wire [4-1:0] node9243;
	wire [4-1:0] node9246;
	wire [4-1:0] node9248;
	wire [4-1:0] node9249;
	wire [4-1:0] node9253;
	wire [4-1:0] node9255;
	wire [4-1:0] node9256;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9263;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9272;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9278;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9287;
	wire [4-1:0] node9290;
	wire [4-1:0] node9291;
	wire [4-1:0] node9294;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9300;
	wire [4-1:0] node9302;
	wire [4-1:0] node9305;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9311;
	wire [4-1:0] node9315;
	wire [4-1:0] node9317;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9324;
	wire [4-1:0] node9325;
	wire [4-1:0] node9326;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9337;
	wire [4-1:0] node9339;
	wire [4-1:0] node9342;
	wire [4-1:0] node9343;
	wire [4-1:0] node9345;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9357;
	wire [4-1:0] node9360;
	wire [4-1:0] node9363;
	wire [4-1:0] node9364;
	wire [4-1:0] node9366;
	wire [4-1:0] node9370;
	wire [4-1:0] node9371;
	wire [4-1:0] node9372;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9383;
	wire [4-1:0] node9385;
	wire [4-1:0] node9388;
	wire [4-1:0] node9390;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9400;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9407;
	wire [4-1:0] node9408;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9413;
	wire [4-1:0] node9415;
	wire [4-1:0] node9416;
	wire [4-1:0] node9419;
	wire [4-1:0] node9422;
	wire [4-1:0] node9423;
	wire [4-1:0] node9425;
	wire [4-1:0] node9426;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9433;
	wire [4-1:0] node9434;
	wire [4-1:0] node9437;
	wire [4-1:0] node9438;
	wire [4-1:0] node9439;
	wire [4-1:0] node9442;
	wire [4-1:0] node9447;
	wire [4-1:0] node9449;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9456;
	wire [4-1:0] node9457;
	wire [4-1:0] node9458;
	wire [4-1:0] node9461;
	wire [4-1:0] node9463;
	wire [4-1:0] node9464;
	wire [4-1:0] node9466;
	wire [4-1:0] node9469;
	wire [4-1:0] node9471;
	wire [4-1:0] node9474;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9481;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9484;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9489;
	wire [4-1:0] node9492;
	wire [4-1:0] node9494;
	wire [4-1:0] node9497;
	wire [4-1:0] node9499;
	wire [4-1:0] node9502;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9511;
	wire [4-1:0] node9512;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9527;
	wire [4-1:0] node9528;
	wire [4-1:0] node9529;
	wire [4-1:0] node9532;
	wire [4-1:0] node9535;
	wire [4-1:0] node9536;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9544;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9550;
	wire [4-1:0] node9553;
	wire [4-1:0] node9554;
	wire [4-1:0] node9556;
	wire [4-1:0] node9560;
	wire [4-1:0] node9561;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9566;
	wire [4-1:0] node9567;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9581;
	wire [4-1:0] node9583;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9591;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9600;
	wire [4-1:0] node9601;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9616;
	wire [4-1:0] node9617;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9625;
	wire [4-1:0] node9627;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9633;
	wire [4-1:0] node9636;
	wire [4-1:0] node9637;
	wire [4-1:0] node9642;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9648;
	wire [4-1:0] node9649;
	wire [4-1:0] node9650;
	wire [4-1:0] node9654;
	wire [4-1:0] node9656;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9662;
	wire [4-1:0] node9663;
	wire [4-1:0] node9667;
	wire [4-1:0] node9671;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9675;
	wire [4-1:0] node9678;
	wire [4-1:0] node9681;
	wire [4-1:0] node9684;
	wire [4-1:0] node9685;
	wire [4-1:0] node9686;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9691;
	wire [4-1:0] node9695;
	wire [4-1:0] node9696;
	wire [4-1:0] node9697;
	wire [4-1:0] node9700;
	wire [4-1:0] node9702;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9708;
	wire [4-1:0] node9710;
	wire [4-1:0] node9713;
	wire [4-1:0] node9715;
	wire [4-1:0] node9718;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9722;
	wire [4-1:0] node9725;
	wire [4-1:0] node9726;
	wire [4-1:0] node9728;
	wire [4-1:0] node9732;
	wire [4-1:0] node9733;
	wire [4-1:0] node9734;
	wire [4-1:0] node9738;
	wire [4-1:0] node9739;
	wire [4-1:0] node9741;
	wire [4-1:0] node9742;
	wire [4-1:0] node9745;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9753;
	wire [4-1:0] node9756;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9765;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9774;
	wire [4-1:0] node9776;
	wire [4-1:0] node9778;
	wire [4-1:0] node9781;
	wire [4-1:0] node9783;
	wire [4-1:0] node9786;
	wire [4-1:0] node9787;
	wire [4-1:0] node9789;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9796;
	wire [4-1:0] node9798;
	wire [4-1:0] node9801;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9805;
	wire [4-1:0] node9807;
	wire [4-1:0] node9808;
	wire [4-1:0] node9811;
	wire [4-1:0] node9814;
	wire [4-1:0] node9815;
	wire [4-1:0] node9816;
	wire [4-1:0] node9818;
	wire [4-1:0] node9823;
	wire [4-1:0] node9824;
	wire [4-1:0] node9825;
	wire [4-1:0] node9827;
	wire [4-1:0] node9830;
	wire [4-1:0] node9831;
	wire [4-1:0] node9833;
	wire [4-1:0] node9837;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9844;
	wire [4-1:0] node9845;
	wire [4-1:0] node9846;
	wire [4-1:0] node9847;
	wire [4-1:0] node9848;
	wire [4-1:0] node9851;
	wire [4-1:0] node9854;
	wire [4-1:0] node9856;
	wire [4-1:0] node9858;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9866;
	wire [4-1:0] node9869;
	wire [4-1:0] node9870;
	wire [4-1:0] node9871;
	wire [4-1:0] node9875;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9881;
	wire [4-1:0] node9882;
	wire [4-1:0] node9888;
	wire [4-1:0] node9889;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9894;
	wire [4-1:0] node9897;
	wire [4-1:0] node9900;
	wire [4-1:0] node9901;
	wire [4-1:0] node9902;
	wire [4-1:0] node9903;
	wire [4-1:0] node9909;
	wire [4-1:0] node9910;
	wire [4-1:0] node9911;
	wire [4-1:0] node9912;
	wire [4-1:0] node9913;
	wire [4-1:0] node9914;
	wire [4-1:0] node9915;
	wire [4-1:0] node9918;
	wire [4-1:0] node9923;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9928;
	wire [4-1:0] node9929;
	wire [4-1:0] node9930;
	wire [4-1:0] node9933;
	wire [4-1:0] node9937;
	wire [4-1:0] node9938;
	wire [4-1:0] node9940;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9948;
	wire [4-1:0] node9951;
	wire [4-1:0] node9955;
	wire [4-1:0] node9956;
	wire [4-1:0] node9957;
	wire [4-1:0] node9961;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9968;
	wire [4-1:0] node9970;
	wire [4-1:0] node9971;
	wire [4-1:0] node9972;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9981;
	wire [4-1:0] node9982;
	wire [4-1:0] node9983;
	wire [4-1:0] node9985;
	wire [4-1:0] node9988;
	wire [4-1:0] node9989;
	wire [4-1:0] node9991;
	wire [4-1:0] node9992;
	wire [4-1:0] node9993;
	wire [4-1:0] node9999;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10002;
	wire [4-1:0] node10005;
	wire [4-1:0] node10009;
	wire [4-1:0] node10010;
	wire [4-1:0] node10011;
	wire [4-1:0] node10012;
	wire [4-1:0] node10013;
	wire [4-1:0] node10017;
	wire [4-1:0] node10019;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10025;
	wire [4-1:0] node10028;
	wire [4-1:0] node10030;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10040;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10044;
	wire [4-1:0] node10046;
	wire [4-1:0] node10048;
	wire [4-1:0] node10050;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10056;
	wire [4-1:0] node10058;
	wire [4-1:0] node10059;
	wire [4-1:0] node10063;
	wire [4-1:0] node10064;
	wire [4-1:0] node10067;
	wire [4-1:0] node10070;
	wire [4-1:0] node10071;
	wire [4-1:0] node10073;
	wire [4-1:0] node10075;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10082;
	wire [4-1:0] node10085;
	wire [4-1:0] node10086;
	wire [4-1:0] node10087;
	wire [4-1:0] node10088;
	wire [4-1:0] node10090;
	wire [4-1:0] node10091;
	wire [4-1:0] node10092;
	wire [4-1:0] node10095;
	wire [4-1:0] node10098;
	wire [4-1:0] node10100;
	wire [4-1:0] node10103;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10109;
	wire [4-1:0] node10112;
	wire [4-1:0] node10113;
	wire [4-1:0] node10114;
	wire [4-1:0] node10118;
	wire [4-1:0] node10119;
	wire [4-1:0] node10120;
	wire [4-1:0] node10123;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10129;
	wire [4-1:0] node10130;
	wire [4-1:0] node10133;
	wire [4-1:0] node10134;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10142;
	wire [4-1:0] node10145;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10149;
	wire [4-1:0] node10152;
	wire [4-1:0] node10153;
	wire [4-1:0] node10155;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10170;
	wire [4-1:0] node10173;
	wire [4-1:0] node10175;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10182;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10191;
	wire [4-1:0] node10192;
	wire [4-1:0] node10195;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10203;
	wire [4-1:0] node10205;
	wire [4-1:0] node10208;
	wire [4-1:0] node10211;
	wire [4-1:0] node10212;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10222;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10238;
	wire [4-1:0] node10242;
	wire [4-1:0] node10245;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10253;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10256;
	wire [4-1:0] node10257;
	wire [4-1:0] node10258;
	wire [4-1:0] node10260;
	wire [4-1:0] node10263;
	wire [4-1:0] node10265;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10270;
	wire [4-1:0] node10274;
	wire [4-1:0] node10276;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10284;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10296;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10307;
	wire [4-1:0] node10310;
	wire [4-1:0] node10311;
	wire [4-1:0] node10312;
	wire [4-1:0] node10313;
	wire [4-1:0] node10315;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10323;
	wire [4-1:0] node10324;
	wire [4-1:0] node10325;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10334;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10337;
	wire [4-1:0] node10341;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10354;
	wire [4-1:0] node10355;
	wire [4-1:0] node10359;
	wire [4-1:0] node10362;
	wire [4-1:0] node10363;
	wire [4-1:0] node10364;
	wire [4-1:0] node10365;
	wire [4-1:0] node10368;
	wire [4-1:0] node10371;
	wire [4-1:0] node10374;
	wire [4-1:0] node10375;
	wire [4-1:0] node10376;
	wire [4-1:0] node10381;
	wire [4-1:0] node10382;
	wire [4-1:0] node10383;
	wire [4-1:0] node10384;
	wire [4-1:0] node10385;
	wire [4-1:0] node10386;
	wire [4-1:0] node10390;
	wire [4-1:0] node10392;
	wire [4-1:0] node10395;
	wire [4-1:0] node10396;
	wire [4-1:0] node10397;
	wire [4-1:0] node10401;
	wire [4-1:0] node10403;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10412;
	wire [4-1:0] node10415;
	wire [4-1:0] node10416;
	wire [4-1:0] node10417;
	wire [4-1:0] node10419;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10427;
	wire [4-1:0] node10429;
	wire [4-1:0] node10432;
	wire [4-1:0] node10433;
	wire [4-1:0] node10434;
	wire [4-1:0] node10436;
	wire [4-1:0] node10437;
	wire [4-1:0] node10440;
	wire [4-1:0] node10442;
	wire [4-1:0] node10445;
	wire [4-1:0] node10446;
	wire [4-1:0] node10449;
	wire [4-1:0] node10451;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10459;
	wire [4-1:0] node10460;
	wire [4-1:0] node10461;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10473;
	wire [4-1:0] node10474;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10480;
	wire [4-1:0] node10481;
	wire [4-1:0] node10486;
	wire [4-1:0] node10487;
	wire [4-1:0] node10488;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10497;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10505;
	wire [4-1:0] node10506;
	wire [4-1:0] node10507;
	wire [4-1:0] node10510;
	wire [4-1:0] node10513;
	wire [4-1:0] node10514;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10542;
	wire [4-1:0] node10545;
	wire [4-1:0] node10546;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10550;
	wire [4-1:0] node10553;
	wire [4-1:0] node10556;
	wire [4-1:0] node10558;
	wire [4-1:0] node10561;
	wire [4-1:0] node10562;
	wire [4-1:0] node10563;
	wire [4-1:0] node10567;
	wire [4-1:0] node10570;
	wire [4-1:0] node10571;
	wire [4-1:0] node10572;
	wire [4-1:0] node10573;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10579;
	wire [4-1:0] node10581;
	wire [4-1:0] node10582;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10592;
	wire [4-1:0] node10596;
	wire [4-1:0] node10597;
	wire [4-1:0] node10600;
	wire [4-1:0] node10603;
	wire [4-1:0] node10604;
	wire [4-1:0] node10605;
	wire [4-1:0] node10606;
	wire [4-1:0] node10609;
	wire [4-1:0] node10612;
	wire [4-1:0] node10613;
	wire [4-1:0] node10614;
	wire [4-1:0] node10618;
	wire [4-1:0] node10621;
	wire [4-1:0] node10622;
	wire [4-1:0] node10623;
	wire [4-1:0] node10625;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10638;
	wire [4-1:0] node10639;
	wire [4-1:0] node10640;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10646;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10651;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10658;
	wire [4-1:0] node10659;
	wire [4-1:0] node10660;
	wire [4-1:0] node10664;
	wire [4-1:0] node10665;
	wire [4-1:0] node10669;
	wire [4-1:0] node10670;
	wire [4-1:0] node10671;
	wire [4-1:0] node10675;
	wire [4-1:0] node10678;
	wire [4-1:0] node10679;
	wire [4-1:0] node10681;
	wire [4-1:0] node10684;
	wire [4-1:0] node10687;
	wire [4-1:0] node10688;
	wire [4-1:0] node10689;
	wire [4-1:0] node10690;
	wire [4-1:0] node10692;
	wire [4-1:0] node10695;
	wire [4-1:0] node10696;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10705;
	wire [4-1:0] node10706;
	wire [4-1:0] node10708;
	wire [4-1:0] node10709;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10717;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10724;
	wire [4-1:0] node10727;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10736;
	wire [4-1:0] node10739;
	wire [4-1:0] node10740;
	wire [4-1:0] node10741;
	wire [4-1:0] node10743;
	wire [4-1:0] node10746;
	wire [4-1:0] node10749;
	wire [4-1:0] node10752;
	wire [4-1:0] node10753;
	wire [4-1:0] node10754;
	wire [4-1:0] node10755;
	wire [4-1:0] node10756;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10764;
	wire [4-1:0] node10767;
	wire [4-1:0] node10770;
	wire [4-1:0] node10771;
	wire [4-1:0] node10773;
	wire [4-1:0] node10774;
	wire [4-1:0] node10778;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10783;
	wire [4-1:0] node10784;
	wire [4-1:0] node10785;
	wire [4-1:0] node10786;
	wire [4-1:0] node10788;
	wire [4-1:0] node10791;
	wire [4-1:0] node10793;
	wire [4-1:0] node10796;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10803;
	wire [4-1:0] node10804;
	wire [4-1:0] node10805;
	wire [4-1:0] node10808;
	wire [4-1:0] node10812;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10824;
	wire [4-1:0] node10825;
	wire [4-1:0] node10828;
	wire [4-1:0] node10830;
	wire [4-1:0] node10833;
	wire [4-1:0] node10834;
	wire [4-1:0] node10835;
	wire [4-1:0] node10836;
	wire [4-1:0] node10837;
	wire [4-1:0] node10838;
	wire [4-1:0] node10839;
	wire [4-1:0] node10844;
	wire [4-1:0] node10847;
	wire [4-1:0] node10849;
	wire [4-1:0] node10850;
	wire [4-1:0] node10854;
	wire [4-1:0] node10856;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10867;
	wire [4-1:0] node10869;
	wire [4-1:0] node10873;
	wire [4-1:0] node10874;
	wire [4-1:0] node10878;
	wire [4-1:0] node10879;
	wire [4-1:0] node10880;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10883;
	wire [4-1:0] node10884;
	wire [4-1:0] node10885;
	wire [4-1:0] node10888;
	wire [4-1:0] node10891;
	wire [4-1:0] node10893;
	wire [4-1:0] node10894;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10901;
	wire [4-1:0] node10902;
	wire [4-1:0] node10903;
	wire [4-1:0] node10906;
	wire [4-1:0] node10911;
	wire [4-1:0] node10912;
	wire [4-1:0] node10914;
	wire [4-1:0] node10916;
	wire [4-1:0] node10919;
	wire [4-1:0] node10920;
	wire [4-1:0] node10922;
	wire [4-1:0] node10924;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10930;
	wire [4-1:0] node10932;
	wire [4-1:0] node10935;
	wire [4-1:0] node10936;
	wire [4-1:0] node10937;
	wire [4-1:0] node10938;
	wire [4-1:0] node10939;
	wire [4-1:0] node10943;
	wire [4-1:0] node10945;
	wire [4-1:0] node10949;
	wire [4-1:0] node10950;
	wire [4-1:0] node10954;
	wire [4-1:0] node10955;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10959;
	wire [4-1:0] node10962;
	wire [4-1:0] node10966;
	wire [4-1:0] node10967;
	wire [4-1:0] node10970;
	wire [4-1:0] node10973;
	wire [4-1:0] node10974;
	wire [4-1:0] node10975;
	wire [4-1:0] node10976;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10982;
	wire [4-1:0] node10986;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10991;
	wire [4-1:0] node10994;
	wire [4-1:0] node10996;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11004;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11011;
	wire [4-1:0] node11015;
	wire [4-1:0] node11016;
	wire [4-1:0] node11017;
	wire [4-1:0] node11021;
	wire [4-1:0] node11022;
	wire [4-1:0] node11023;
	wire [4-1:0] node11028;
	wire [4-1:0] node11029;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11032;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11036;
	wire [4-1:0] node11040;
	wire [4-1:0] node11041;
	wire [4-1:0] node11045;
	wire [4-1:0] node11047;
	wire [4-1:0] node11049;
	wire [4-1:0] node11052;
	wire [4-1:0] node11053;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11057;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11066;
	wire [4-1:0] node11068;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11073;
	wire [4-1:0] node11075;
	wire [4-1:0] node11077;
	wire [4-1:0] node11080;
	wire [4-1:0] node11081;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11087;
	wire [4-1:0] node11090;
	wire [4-1:0] node11093;
	wire [4-1:0] node11094;
	wire [4-1:0] node11095;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11114;
	wire [4-1:0] node11118;
	wire [4-1:0] node11119;
	wire [4-1:0] node11121;
	wire [4-1:0] node11125;
	wire [4-1:0] node11126;
	wire [4-1:0] node11128;
	wire [4-1:0] node11131;
	wire [4-1:0] node11132;
	wire [4-1:0] node11135;
	wire [4-1:0] node11137;
	wire [4-1:0] node11139;
	wire [4-1:0] node11141;
	wire [4-1:0] node11144;
	wire [4-1:0] node11145;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11149;
	wire [4-1:0] node11152;
	wire [4-1:0] node11154;
	wire [4-1:0] node11157;
	wire [4-1:0] node11158;
	wire [4-1:0] node11162;
	wire [4-1:0] node11163;
	wire [4-1:0] node11164;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11171;
	wire [4-1:0] node11173;
	wire [4-1:0] node11177;
	wire [4-1:0] node11178;
	wire [4-1:0] node11179;
	wire [4-1:0] node11180;
	wire [4-1:0] node11181;
	wire [4-1:0] node11182;
	wire [4-1:0] node11183;
	wire [4-1:0] node11185;
	wire [4-1:0] node11188;
	wire [4-1:0] node11189;
	wire [4-1:0] node11191;
	wire [4-1:0] node11194;
	wire [4-1:0] node11196;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11201;
	wire [4-1:0] node11202;
	wire [4-1:0] node11205;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11213;
	wire [4-1:0] node11216;
	wire [4-1:0] node11221;
	wire [4-1:0] node11222;
	wire [4-1:0] node11224;
	wire [4-1:0] node11227;
	wire [4-1:0] node11228;
	wire [4-1:0] node11231;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11238;
	wire [4-1:0] node11239;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11246;
	wire [4-1:0] node11248;
	wire [4-1:0] node11251;
	wire [4-1:0] node11252;
	wire [4-1:0] node11253;
	wire [4-1:0] node11255;
	wire [4-1:0] node11259;
	wire [4-1:0] node11262;
	wire [4-1:0] node11263;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11266;
	wire [4-1:0] node11271;
	wire [4-1:0] node11272;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11280;
	wire [4-1:0] node11284;
	wire [4-1:0] node11287;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11292;
	wire [4-1:0] node11293;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11308;
	wire [4-1:0] node11309;
	wire [4-1:0] node11314;
	wire [4-1:0] node11315;
	wire [4-1:0] node11316;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11322;
	wire [4-1:0] node11325;
	wire [4-1:0] node11329;
	wire [4-1:0] node11330;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11333;
	wire [4-1:0] node11334;
	wire [4-1:0] node11338;
	wire [4-1:0] node11341;
	wire [4-1:0] node11344;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11350;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11354;
	wire [4-1:0] node11359;
	wire [4-1:0] node11360;
	wire [4-1:0] node11361;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11367;
	wire [4-1:0] node11372;
	wire [4-1:0] node11373;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11376;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11383;
	wire [4-1:0] node11385;
	wire [4-1:0] node11388;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11395;
	wire [4-1:0] node11397;
	wire [4-1:0] node11399;
	wire [4-1:0] node11402;
	wire [4-1:0] node11403;
	wire [4-1:0] node11406;
	wire [4-1:0] node11407;
	wire [4-1:0] node11410;
	wire [4-1:0] node11413;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11417;
	wire [4-1:0] node11419;
	wire [4-1:0] node11421;
	wire [4-1:0] node11424;
	wire [4-1:0] node11425;
	wire [4-1:0] node11427;
	wire [4-1:0] node11428;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11435;
	wire [4-1:0] node11438;
	wire [4-1:0] node11439;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11452;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11457;
	wire [4-1:0] node11458;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11466;
	wire [4-1:0] node11469;
	wire [4-1:0] node11470;
	wire [4-1:0] node11471;
	wire [4-1:0] node11473;
	wire [4-1:0] node11476;
	wire [4-1:0] node11479;
	wire [4-1:0] node11481;
	wire [4-1:0] node11484;
	wire [4-1:0] node11485;
	wire [4-1:0] node11486;
	wire [4-1:0] node11488;
	wire [4-1:0] node11489;
	wire [4-1:0] node11493;
	wire [4-1:0] node11495;
	wire [4-1:0] node11497;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11507;
	wire [4-1:0] node11510;
	wire [4-1:0] node11511;
	wire [4-1:0] node11513;
	wire [4-1:0] node11516;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11523;
	wire [4-1:0] node11524;
	wire [4-1:0] node11525;
	wire [4-1:0] node11526;
	wire [4-1:0] node11529;
	wire [4-1:0] node11532;
	wire [4-1:0] node11533;
	wire [4-1:0] node11536;
	wire [4-1:0] node11539;
	wire [4-1:0] node11541;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11548;
	wire [4-1:0] node11549;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11553;
	wire [4-1:0] node11557;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11564;
	wire [4-1:0] node11566;
	wire [4-1:0] node11569;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11574;
	wire [4-1:0] node11578;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11583;
	wire [4-1:0] node11587;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11598;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11609;
	wire [4-1:0] node11610;
	wire [4-1:0] node11614;
	wire [4-1:0] node11615;
	wire [4-1:0] node11616;
	wire [4-1:0] node11617;
	wire [4-1:0] node11621;
	wire [4-1:0] node11622;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11630;
	wire [4-1:0] node11631;
	wire [4-1:0] node11637;
	wire [4-1:0] node11638;
	wire [4-1:0] node11642;
	wire [4-1:0] node11643;
	wire [4-1:0] node11644;
	wire [4-1:0] node11645;
	wire [4-1:0] node11647;
	wire [4-1:0] node11650;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11656;
	wire [4-1:0] node11660;
	wire [4-1:0] node11661;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11678;
	wire [4-1:0] node11680;
	wire [4-1:0] node11682;
	wire [4-1:0] node11685;
	wire [4-1:0] node11686;
	wire [4-1:0] node11688;
	wire [4-1:0] node11692;
	wire [4-1:0] node11693;
	wire [4-1:0] node11694;
	wire [4-1:0] node11697;
	wire [4-1:0] node11700;
	wire [4-1:0] node11703;
	wire [4-1:0] node11704;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11710;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11717;
	wire [4-1:0] node11718;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11724;
	wire [4-1:0] node11725;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11738;
	wire [4-1:0] node11741;
	wire [4-1:0] node11742;
	wire [4-1:0] node11746;
	wire [4-1:0] node11747;
	wire [4-1:0] node11750;
	wire [4-1:0] node11751;
	wire [4-1:0] node11752;
	wire [4-1:0] node11756;
	wire [4-1:0] node11759;
	wire [4-1:0] node11760;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11768;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11774;
	wire [4-1:0] node11777;
	wire [4-1:0] node11779;
	wire [4-1:0] node11782;
	wire [4-1:0] node11783;
	wire [4-1:0] node11784;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11792;
	wire [4-1:0] node11795;
	wire [4-1:0] node11796;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11806;
	wire [4-1:0] node11808;
	wire [4-1:0] node11811;
	wire [4-1:0] node11812;
	wire [4-1:0] node11813;
	wire [4-1:0] node11815;
	wire [4-1:0] node11818;
	wire [4-1:0] node11821;
	wire [4-1:0] node11822;
	wire [4-1:0] node11825;
	wire [4-1:0] node11828;
	wire [4-1:0] node11829;
	wire [4-1:0] node11830;
	wire [4-1:0] node11831;
	wire [4-1:0] node11832;
	wire [4-1:0] node11833;
	wire [4-1:0] node11834;
	wire [4-1:0] node11835;
	wire [4-1:0] node11838;
	wire [4-1:0] node11839;
	wire [4-1:0] node11843;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11846;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11853;
	wire [4-1:0] node11857;
	wire [4-1:0] node11860;
	wire [4-1:0] node11861;
	wire [4-1:0] node11862;
	wire [4-1:0] node11863;
	wire [4-1:0] node11864;
	wire [4-1:0] node11867;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11875;
	wire [4-1:0] node11876;
	wire [4-1:0] node11878;
	wire [4-1:0] node11881;
	wire [4-1:0] node11884;
	wire [4-1:0] node11885;
	wire [4-1:0] node11886;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11892;
	wire [4-1:0] node11895;
	wire [4-1:0] node11896;
	wire [4-1:0] node11897;
	wire [4-1:0] node11902;
	wire [4-1:0] node11904;
	wire [4-1:0] node11907;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11912;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11925;
	wire [4-1:0] node11926;
	wire [4-1:0] node11931;
	wire [4-1:0] node11933;
	wire [4-1:0] node11936;
	wire [4-1:0] node11937;
	wire [4-1:0] node11938;
	wire [4-1:0] node11939;
	wire [4-1:0] node11943;
	wire [4-1:0] node11944;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11950;
	wire [4-1:0] node11952;
	wire [4-1:0] node11955;
	wire [4-1:0] node11958;
	wire [4-1:0] node11960;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11966;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11977;
	wire [4-1:0] node11980;
	wire [4-1:0] node11981;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11987;
	wire [4-1:0] node11989;
	wire [4-1:0] node11992;
	wire [4-1:0] node11995;
	wire [4-1:0] node11996;
	wire [4-1:0] node11998;
	wire [4-1:0] node12000;
	wire [4-1:0] node12003;
	wire [4-1:0] node12004;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12012;
	wire [4-1:0] node12013;
	wire [4-1:0] node12014;
	wire [4-1:0] node12017;
	wire [4-1:0] node12020;
	wire [4-1:0] node12021;
	wire [4-1:0] node12023;
	wire [4-1:0] node12026;
	wire [4-1:0] node12029;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12033;
	wire [4-1:0] node12034;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12043;
	wire [4-1:0] node12045;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12058;
	wire [4-1:0] node12059;
	wire [4-1:0] node12064;
	wire [4-1:0] node12065;
	wire [4-1:0] node12066;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12076;
	wire [4-1:0] node12081;
	wire [4-1:0] node12082;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12089;
	wire [4-1:0] node12092;
	wire [4-1:0] node12093;
	wire [4-1:0] node12094;
	wire [4-1:0] node12095;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12105;
	wire [4-1:0] node12106;
	wire [4-1:0] node12108;
	wire [4-1:0] node12110;
	wire [4-1:0] node12113;
	wire [4-1:0] node12115;
	wire [4-1:0] node12117;
	wire [4-1:0] node12120;
	wire [4-1:0] node12121;
	wire [4-1:0] node12122;
	wire [4-1:0] node12123;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12127;
	wire [4-1:0] node12131;
	wire [4-1:0] node12132;
	wire [4-1:0] node12134;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12142;
	wire [4-1:0] node12144;
	wire [4-1:0] node12147;
	wire [4-1:0] node12149;
	wire [4-1:0] node12153;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12158;
	wire [4-1:0] node12159;
	wire [4-1:0] node12163;
	wire [4-1:0] node12165;
	wire [4-1:0] node12167;
	wire [4-1:0] node12168;
	wire [4-1:0] node12170;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12178;
	wire [4-1:0] node12182;
	wire [4-1:0] node12184;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12190;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12208;
	wire [4-1:0] node12209;
	wire [4-1:0] node12210;
	wire [4-1:0] node12214;
	wire [4-1:0] node12216;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12224;
	wire [4-1:0] node12225;
	wire [4-1:0] node12227;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12233;
	wire [4-1:0] node12237;
	wire [4-1:0] node12239;
	wire [4-1:0] node12242;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12246;
	wire [4-1:0] node12247;
	wire [4-1:0] node12250;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12255;
	wire [4-1:0] node12259;
	wire [4-1:0] node12262;
	wire [4-1:0] node12263;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12271;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12279;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12284;
	wire [4-1:0] node12288;
	wire [4-1:0] node12291;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12297;
	wire [4-1:0] node12300;
	wire [4-1:0] node12301;
	wire [4-1:0] node12302;
	wire [4-1:0] node12303;
	wire [4-1:0] node12305;
	wire [4-1:0] node12306;
	wire [4-1:0] node12310;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12315;
	wire [4-1:0] node12319;
	wire [4-1:0] node12320;
	wire [4-1:0] node12322;
	wire [4-1:0] node12324;
	wire [4-1:0] node12325;
	wire [4-1:0] node12329;
	wire [4-1:0] node12330;
	wire [4-1:0] node12333;
	wire [4-1:0] node12335;
	wire [4-1:0] node12337;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12342;
	wire [4-1:0] node12344;
	wire [4-1:0] node12346;
	wire [4-1:0] node12349;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12360;
	wire [4-1:0] node12361;
	wire [4-1:0] node12363;
	wire [4-1:0] node12366;
	wire [4-1:0] node12370;
	wire [4-1:0] node12371;
	wire [4-1:0] node12373;
	wire [4-1:0] node12377;
	wire [4-1:0] node12378;
	wire [4-1:0] node12379;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12386;
	wire [4-1:0] node12389;
	wire [4-1:0] node12391;
	wire [4-1:0] node12394;
	wire [4-1:0] node12395;
	wire [4-1:0] node12396;
	wire [4-1:0] node12397;
	wire [4-1:0] node12402;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12412;
	wire [4-1:0] node12413;
	wire [4-1:0] node12417;
	wire [4-1:0] node12419;
	wire [4-1:0] node12420;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12427;
	wire [4-1:0] node12428;
	wire [4-1:0] node12429;
	wire [4-1:0] node12434;
	wire [4-1:0] node12436;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12445;
	wire [4-1:0] node12448;
	wire [4-1:0] node12449;
	wire [4-1:0] node12453;
	wire [4-1:0] node12455;
	wire [4-1:0] node12457;
	wire [4-1:0] node12460;
	wire [4-1:0] node12461;
	wire [4-1:0] node12464;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12468;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12479;
	wire [4-1:0] node12481;
	wire [4-1:0] node12483;
	wire [4-1:0] node12485;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12492;
	wire [4-1:0] node12493;
	wire [4-1:0] node12497;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12503;
	wire [4-1:0] node12504;
	wire [4-1:0] node12505;
	wire [4-1:0] node12508;
	wire [4-1:0] node12512;
	wire [4-1:0] node12513;
	wire [4-1:0] node12514;
	wire [4-1:0] node12515;
	wire [4-1:0] node12516;
	wire [4-1:0] node12517;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12520;
	wire [4-1:0] node12521;
	wire [4-1:0] node12525;
	wire [4-1:0] node12527;
	wire [4-1:0] node12531;
	wire [4-1:0] node12532;
	wire [4-1:0] node12535;
	wire [4-1:0] node12537;
	wire [4-1:0] node12540;
	wire [4-1:0] node12541;
	wire [4-1:0] node12542;
	wire [4-1:0] node12543;
	wire [4-1:0] node12547;
	wire [4-1:0] node12549;
	wire [4-1:0] node12552;
	wire [4-1:0] node12553;
	wire [4-1:0] node12556;
	wire [4-1:0] node12558;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12563;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12569;
	wire [4-1:0] node12570;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12579;
	wire [4-1:0] node12584;
	wire [4-1:0] node12586;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12594;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12601;
	wire [4-1:0] node12602;
	wire [4-1:0] node12607;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12614;
	wire [4-1:0] node12615;
	wire [4-1:0] node12619;
	wire [4-1:0] node12622;
	wire [4-1:0] node12623;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12630;
	wire [4-1:0] node12632;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12637;
	wire [4-1:0] node12638;
	wire [4-1:0] node12642;
	wire [4-1:0] node12645;
	wire [4-1:0] node12647;
	wire [4-1:0] node12650;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12655;
	wire [4-1:0] node12657;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12668;
	wire [4-1:0] node12669;
	wire [4-1:0] node12671;
	wire [4-1:0] node12672;
	wire [4-1:0] node12674;
	wire [4-1:0] node12675;
	wire [4-1:0] node12680;
	wire [4-1:0] node12682;
	wire [4-1:0] node12683;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12689;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12692;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12702;
	wire [4-1:0] node12703;
	wire [4-1:0] node12705;
	wire [4-1:0] node12708;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12725;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12732;
	wire [4-1:0] node12733;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12739;
	wire [4-1:0] node12740;
	wire [4-1:0] node12743;
	wire [4-1:0] node12746;
	wire [4-1:0] node12747;
	wire [4-1:0] node12750;
	wire [4-1:0] node12751;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12757;
	wire [4-1:0] node12758;
	wire [4-1:0] node12759;
	wire [4-1:0] node12762;
	wire [4-1:0] node12763;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12770;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12780;
	wire [4-1:0] node12781;
	wire [4-1:0] node12782;
	wire [4-1:0] node12784;
	wire [4-1:0] node12788;
	wire [4-1:0] node12789;
	wire [4-1:0] node12790;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12799;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12803;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12812;
	wire [4-1:0] node12814;
	wire [4-1:0] node12816;
	wire [4-1:0] node12819;
	wire [4-1:0] node12820;
	wire [4-1:0] node12822;
	wire [4-1:0] node12823;
	wire [4-1:0] node12826;
	wire [4-1:0] node12829;
	wire [4-1:0] node12831;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12836;
	wire [4-1:0] node12837;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12845;
	wire [4-1:0] node12848;
	wire [4-1:0] node12850;
	wire [4-1:0] node12852;
	wire [4-1:0] node12855;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12859;
	wire [4-1:0] node12861;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12872;
	wire [4-1:0] node12873;
	wire [4-1:0] node12875;
	wire [4-1:0] node12877;
	wire [4-1:0] node12880;
	wire [4-1:0] node12882;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12887;
	wire [4-1:0] node12888;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12897;
	wire [4-1:0] node12902;
	wire [4-1:0] node12903;
	wire [4-1:0] node12904;
	wire [4-1:0] node12905;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12912;
	wire [4-1:0] node12915;
	wire [4-1:0] node12916;
	wire [4-1:0] node12919;
	wire [4-1:0] node12921;
	wire [4-1:0] node12924;
	wire [4-1:0] node12925;
	wire [4-1:0] node12926;
	wire [4-1:0] node12928;
	wire [4-1:0] node12931;
	wire [4-1:0] node12932;
	wire [4-1:0] node12936;
	wire [4-1:0] node12937;
	wire [4-1:0] node12940;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12954;
	wire [4-1:0] node12955;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12963;
	wire [4-1:0] node12966;
	wire [4-1:0] node12967;
	wire [4-1:0] node12969;
	wire [4-1:0] node12972;
	wire [4-1:0] node12973;
	wire [4-1:0] node12974;
	wire [4-1:0] node12977;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12984;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12995;
	wire [4-1:0] node12996;
	wire [4-1:0] node13000;
	wire [4-1:0] node13003;
	wire [4-1:0] node13004;
	wire [4-1:0] node13006;
	wire [4-1:0] node13008;
	wire [4-1:0] node13011;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13018;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13024;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13034;
	wire [4-1:0] node13035;
	wire [4-1:0] node13036;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13043;
	wire [4-1:0] node13046;
	wire [4-1:0] node13047;
	wire [4-1:0] node13048;
	wire [4-1:0] node13049;
	wire [4-1:0] node13052;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13060;
	wire [4-1:0] node13063;
	wire [4-1:0] node13064;
	wire [4-1:0] node13065;
	wire [4-1:0] node13066;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13072;
	wire [4-1:0] node13073;
	wire [4-1:0] node13079;
	wire [4-1:0] node13080;
	wire [4-1:0] node13081;
	wire [4-1:0] node13084;
	wire [4-1:0] node13085;
	wire [4-1:0] node13087;
	wire [4-1:0] node13091;
	wire [4-1:0] node13092;
	wire [4-1:0] node13095;
	wire [4-1:0] node13097;
	wire [4-1:0] node13099;
	wire [4-1:0] node13102;
	wire [4-1:0] node13103;
	wire [4-1:0] node13104;
	wire [4-1:0] node13105;
	wire [4-1:0] node13106;
	wire [4-1:0] node13109;
	wire [4-1:0] node13110;
	wire [4-1:0] node13114;
	wire [4-1:0] node13115;
	wire [4-1:0] node13116;
	wire [4-1:0] node13120;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13127;
	wire [4-1:0] node13128;
	wire [4-1:0] node13130;
	wire [4-1:0] node13131;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13149;
	wire [4-1:0] node13150;
	wire [4-1:0] node13154;
	wire [4-1:0] node13155;
	wire [4-1:0] node13156;
	wire [4-1:0] node13157;
	wire [4-1:0] node13160;
	wire [4-1:0] node13163;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13169;
	wire [4-1:0] node13172;
	wire [4-1:0] node13173;
	wire [4-1:0] node13174;
	wire [4-1:0] node13175;
	wire [4-1:0] node13179;
	wire [4-1:0] node13180;
	wire [4-1:0] node13181;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13190;
	wire [4-1:0] node13191;
	wire [4-1:0] node13195;
	wire [4-1:0] node13196;
	wire [4-1:0] node13197;
	wire [4-1:0] node13198;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13201;
	wire [4-1:0] node13202;
	wire [4-1:0] node13203;
	wire [4-1:0] node13204;
	wire [4-1:0] node13207;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13213;
	wire [4-1:0] node13214;
	wire [4-1:0] node13216;
	wire [4-1:0] node13220;
	wire [4-1:0] node13221;
	wire [4-1:0] node13225;
	wire [4-1:0] node13226;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13232;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13238;
	wire [4-1:0] node13239;
	wire [4-1:0] node13240;
	wire [4-1:0] node13241;
	wire [4-1:0] node13246;
	wire [4-1:0] node13248;
	wire [4-1:0] node13251;
	wire [4-1:0] node13252;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13265;
	wire [4-1:0] node13267;
	wire [4-1:0] node13270;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13281;
	wire [4-1:0] node13284;
	wire [4-1:0] node13285;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13293;
	wire [4-1:0] node13294;
	wire [4-1:0] node13297;
	wire [4-1:0] node13299;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13309;
	wire [4-1:0] node13312;
	wire [4-1:0] node13314;
	wire [4-1:0] node13317;
	wire [4-1:0] node13318;
	wire [4-1:0] node13319;
	wire [4-1:0] node13321;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13327;
	wire [4-1:0] node13329;
	wire [4-1:0] node13332;
	wire [4-1:0] node13334;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13341;
	wire [4-1:0] node13343;
	wire [4-1:0] node13346;
	wire [4-1:0] node13348;
	wire [4-1:0] node13351;
	wire [4-1:0] node13352;
	wire [4-1:0] node13353;
	wire [4-1:0] node13356;
	wire [4-1:0] node13358;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13364;
	wire [4-1:0] node13365;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13374;
	wire [4-1:0] node13376;
	wire [4-1:0] node13379;
	wire [4-1:0] node13380;
	wire [4-1:0] node13383;
	wire [4-1:0] node13385;
	wire [4-1:0] node13388;
	wire [4-1:0] node13389;
	wire [4-1:0] node13391;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13402;
	wire [4-1:0] node13405;
	wire [4-1:0] node13406;
	wire [4-1:0] node13407;
	wire [4-1:0] node13408;
	wire [4-1:0] node13410;
	wire [4-1:0] node13413;
	wire [4-1:0] node13415;
	wire [4-1:0] node13417;
	wire [4-1:0] node13420;
	wire [4-1:0] node13421;
	wire [4-1:0] node13424;
	wire [4-1:0] node13427;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13432;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13441;
	wire [4-1:0] node13442;
	wire [4-1:0] node13445;
	wire [4-1:0] node13447;
	wire [4-1:0] node13450;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13453;
	wire [4-1:0] node13455;
	wire [4-1:0] node13456;
	wire [4-1:0] node13459;
	wire [4-1:0] node13462;
	wire [4-1:0] node13463;
	wire [4-1:0] node13464;
	wire [4-1:0] node13468;
	wire [4-1:0] node13471;
	wire [4-1:0] node13472;
	wire [4-1:0] node13475;
	wire [4-1:0] node13478;
	wire [4-1:0] node13479;
	wire [4-1:0] node13480;
	wire [4-1:0] node13482;
	wire [4-1:0] node13484;
	wire [4-1:0] node13487;
	wire [4-1:0] node13489;
	wire [4-1:0] node13490;
	wire [4-1:0] node13494;
	wire [4-1:0] node13495;
	wire [4-1:0] node13496;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13500;
	wire [4-1:0] node13505;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13512;
	wire [4-1:0] node13513;
	wire [4-1:0] node13515;
	wire [4-1:0] node13519;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13524;
	wire [4-1:0] node13526;
	wire [4-1:0] node13528;
	wire [4-1:0] node13530;
	wire [4-1:0] node13533;
	wire [4-1:0] node13534;
	wire [4-1:0] node13535;
	wire [4-1:0] node13536;
	wire [4-1:0] node13539;
	wire [4-1:0] node13543;
	wire [4-1:0] node13546;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13551;
	wire [4-1:0] node13553;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13566;
	wire [4-1:0] node13569;
	wire [4-1:0] node13570;
	wire [4-1:0] node13571;
	wire [4-1:0] node13572;
	wire [4-1:0] node13575;
	wire [4-1:0] node13577;
	wire [4-1:0] node13580;
	wire [4-1:0] node13581;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13587;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13599;
	wire [4-1:0] node13602;
	wire [4-1:0] node13605;
	wire [4-1:0] node13608;
	wire [4-1:0] node13609;
	wire [4-1:0] node13610;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13613;
	wire [4-1:0] node13614;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13623;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13628;
	wire [4-1:0] node13631;
	wire [4-1:0] node13634;
	wire [4-1:0] node13636;
	wire [4-1:0] node13639;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13645;
	wire [4-1:0] node13648;
	wire [4-1:0] node13650;
	wire [4-1:0] node13651;
	wire [4-1:0] node13655;
	wire [4-1:0] node13656;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13662;
	wire [4-1:0] node13665;
	wire [4-1:0] node13666;
	wire [4-1:0] node13670;
	wire [4-1:0] node13671;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13675;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13680;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13693;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13704;
	wire [4-1:0] node13705;
	wire [4-1:0] node13709;
	wire [4-1:0] node13712;
	wire [4-1:0] node13713;
	wire [4-1:0] node13714;
	wire [4-1:0] node13718;
	wire [4-1:0] node13720;
	wire [4-1:0] node13722;
	wire [4-1:0] node13725;
	wire [4-1:0] node13727;
	wire [4-1:0] node13729;
	wire [4-1:0] node13731;
	wire [4-1:0] node13732;
	wire [4-1:0] node13735;
	wire [4-1:0] node13738;
	wire [4-1:0] node13739;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13744;
	wire [4-1:0] node13746;
	wire [4-1:0] node13749;
	wire [4-1:0] node13751;
	wire [4-1:0] node13753;
	wire [4-1:0] node13755;
	wire [4-1:0] node13758;
	wire [4-1:0] node13759;
	wire [4-1:0] node13760;
	wire [4-1:0] node13763;
	wire [4-1:0] node13766;
	wire [4-1:0] node13768;
	wire [4-1:0] node13769;
	wire [4-1:0] node13773;
	wire [4-1:0] node13774;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13780;
	wire [4-1:0] node13781;
	wire [4-1:0] node13786;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13799;
	wire [4-1:0] node13800;
	wire [4-1:0] node13804;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13808;
	wire [4-1:0] node13809;
	wire [4-1:0] node13813;
	wire [4-1:0] node13816;
	wire [4-1:0] node13818;
	wire [4-1:0] node13821;
	wire [4-1:0] node13822;
	wire [4-1:0] node13823;
	wire [4-1:0] node13824;
	wire [4-1:0] node13825;
	wire [4-1:0] node13827;
	wire [4-1:0] node13830;
	wire [4-1:0] node13833;
	wire [4-1:0] node13834;
	wire [4-1:0] node13838;
	wire [4-1:0] node13839;
	wire [4-1:0] node13841;
	wire [4-1:0] node13844;
	wire [4-1:0] node13846;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13860;
	wire [4-1:0] node13865;
	wire [4-1:0] node13866;
	wire [4-1:0] node13867;
	wire [4-1:0] node13868;
	wire [4-1:0] node13873;
	wire [4-1:0] node13874;
	wire [4-1:0] node13878;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13881;
	wire [4-1:0] node13882;
	wire [4-1:0] node13883;
	wire [4-1:0] node13884;
	wire [4-1:0] node13885;
	wire [4-1:0] node13887;
	wire [4-1:0] node13888;
	wire [4-1:0] node13889;
	wire [4-1:0] node13894;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13903;
	wire [4-1:0] node13907;
	wire [4-1:0] node13910;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13915;
	wire [4-1:0] node13919;
	wire [4-1:0] node13922;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13928;
	wire [4-1:0] node13929;
	wire [4-1:0] node13933;
	wire [4-1:0] node13935;
	wire [4-1:0] node13938;
	wire [4-1:0] node13939;
	wire [4-1:0] node13941;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13950;
	wire [4-1:0] node13954;
	wire [4-1:0] node13957;
	wire [4-1:0] node13958;
	wire [4-1:0] node13959;
	wire [4-1:0] node13962;
	wire [4-1:0] node13964;
	wire [4-1:0] node13967;
	wire [4-1:0] node13969;
	wire [4-1:0] node13972;
	wire [4-1:0] node13973;
	wire [4-1:0] node13974;
	wire [4-1:0] node13976;
	wire [4-1:0] node13977;
	wire [4-1:0] node13981;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13987;
	wire [4-1:0] node13988;
	wire [4-1:0] node13989;
	wire [4-1:0] node13993;
	wire [4-1:0] node13995;
	wire [4-1:0] node13998;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14002;
	wire [4-1:0] node14005;
	wire [4-1:0] node14006;
	wire [4-1:0] node14010;
	wire [4-1:0] node14013;
	wire [4-1:0] node14014;
	wire [4-1:0] node14015;
	wire [4-1:0] node14016;
	wire [4-1:0] node14017;
	wire [4-1:0] node14019;
	wire [4-1:0] node14020;
	wire [4-1:0] node14022;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14031;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14036;
	wire [4-1:0] node14037;
	wire [4-1:0] node14040;
	wire [4-1:0] node14043;
	wire [4-1:0] node14044;
	wire [4-1:0] node14047;
	wire [4-1:0] node14050;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14053;
	wire [4-1:0] node14055;
	wire [4-1:0] node14059;
	wire [4-1:0] node14060;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14068;
	wire [4-1:0] node14070;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14078;
	wire [4-1:0] node14079;
	wire [4-1:0] node14080;
	wire [4-1:0] node14081;
	wire [4-1:0] node14085;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14092;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14098;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14103;
	wire [4-1:0] node14107;
	wire [4-1:0] node14109;
	wire [4-1:0] node14111;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14117;
	wire [4-1:0] node14120;
	wire [4-1:0] node14122;
	wire [4-1:0] node14125;
	wire [4-1:0] node14126;
	wire [4-1:0] node14127;
	wire [4-1:0] node14129;
	wire [4-1:0] node14132;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14140;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14144;
	wire [4-1:0] node14145;
	wire [4-1:0] node14149;
	wire [4-1:0] node14150;
	wire [4-1:0] node14151;
	wire [4-1:0] node14155;
	wire [4-1:0] node14156;
	wire [4-1:0] node14160;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14167;
	wire [4-1:0] node14168;
	wire [4-1:0] node14171;
	wire [4-1:0] node14173;
	wire [4-1:0] node14176;
	wire [4-1:0] node14177;
	wire [4-1:0] node14181;
	wire [4-1:0] node14182;
	wire [4-1:0] node14184;
	wire [4-1:0] node14187;
	wire [4-1:0] node14188;
	wire [4-1:0] node14189;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14200;
	wire [4-1:0] node14201;
	wire [4-1:0] node14205;
	wire [4-1:0] node14207;
	wire [4-1:0] node14210;
	wire [4-1:0] node14211;
	wire [4-1:0] node14213;
	wire [4-1:0] node14214;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14222;
	wire [4-1:0] node14223;
	wire [4-1:0] node14225;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14231;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14237;
	wire [4-1:0] node14238;
	wire [4-1:0] node14242;
	wire [4-1:0] node14243;
	wire [4-1:0] node14244;
	wire [4-1:0] node14247;
	wire [4-1:0] node14249;
	wire [4-1:0] node14252;
	wire [4-1:0] node14255;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14259;
	wire [4-1:0] node14262;
	wire [4-1:0] node14263;
	wire [4-1:0] node14267;
	wire [4-1:0] node14270;
	wire [4-1:0] node14271;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14274;
	wire [4-1:0] node14275;
	wire [4-1:0] node14278;
	wire [4-1:0] node14281;
	wire [4-1:0] node14282;
	wire [4-1:0] node14286;
	wire [4-1:0] node14287;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14299;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14306;
	wire [4-1:0] node14307;
	wire [4-1:0] node14308;
	wire [4-1:0] node14312;
	wire [4-1:0] node14315;
	wire [4-1:0] node14316;
	wire [4-1:0] node14317;
	wire [4-1:0] node14320;
	wire [4-1:0] node14322;
	wire [4-1:0] node14325;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14331;
	wire [4-1:0] node14332;
	wire [4-1:0] node14333;
	wire [4-1:0] node14338;
	wire [4-1:0] node14339;
	wire [4-1:0] node14342;
	wire [4-1:0] node14344;
	wire [4-1:0] node14347;
	wire [4-1:0] node14348;
	wire [4-1:0] node14349;
	wire [4-1:0] node14350;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14357;
	wire [4-1:0] node14358;
	wire [4-1:0] node14362;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14367;
	wire [4-1:0] node14368;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14384;
	wire [4-1:0] node14388;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14395;
	wire [4-1:0] node14396;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14399;
	wire [4-1:0] node14400;
	wire [4-1:0] node14403;
	wire [4-1:0] node14406;
	wire [4-1:0] node14407;
	wire [4-1:0] node14410;
	wire [4-1:0] node14412;
	wire [4-1:0] node14415;
	wire [4-1:0] node14416;
	wire [4-1:0] node14417;
	wire [4-1:0] node14421;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14426;
	wire [4-1:0] node14428;
	wire [4-1:0] node14431;
	wire [4-1:0] node14433;
	wire [4-1:0] node14434;
	wire [4-1:0] node14435;
	wire [4-1:0] node14439;
	wire [4-1:0] node14442;
	wire [4-1:0] node14443;
	wire [4-1:0] node14446;
	wire [4-1:0] node14447;
	wire [4-1:0] node14449;
	wire [4-1:0] node14452;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14458;
	wire [4-1:0] node14459;
	wire [4-1:0] node14460;
	wire [4-1:0] node14466;
	wire [4-1:0] node14467;
	wire [4-1:0] node14469;
	wire [4-1:0] node14472;
	wire [4-1:0] node14473;
	wire [4-1:0] node14477;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14485;
	wire [4-1:0] node14486;
	wire [4-1:0] node14490;
	wire [4-1:0] node14491;
	wire [4-1:0] node14494;
	wire [4-1:0] node14497;
	wire [4-1:0] node14498;
	wire [4-1:0] node14499;
	wire [4-1:0] node14500;
	wire [4-1:0] node14503;
	wire [4-1:0] node14506;
	wire [4-1:0] node14508;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14518;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14524;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14531;
	wire [4-1:0] node14535;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14538;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14554;
	wire [4-1:0] node14555;
	wire [4-1:0] node14556;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14573;
	wire [4-1:0] node14576;
	wire [4-1:0] node14577;
	wire [4-1:0] node14578;
	wire [4-1:0] node14579;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14592;
	wire [4-1:0] node14595;
	wire [4-1:0] node14596;
	wire [4-1:0] node14597;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14603;
	wire [4-1:0] node14605;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14613;
	wire [4-1:0] node14616;
	wire [4-1:0] node14619;
	wire [4-1:0] node14622;
	wire [4-1:0] node14624;
	wire [4-1:0] node14626;
	wire [4-1:0] node14629;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14634;
	wire [4-1:0] node14637;
	wire [4-1:0] node14639;
	wire [4-1:0] node14641;
	wire [4-1:0] node14643;
	wire [4-1:0] node14644;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14651;
	wire [4-1:0] node14652;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14660;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14666;
	wire [4-1:0] node14668;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14674;
	wire [4-1:0] node14677;
	wire [4-1:0] node14680;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14683;
	wire [4-1:0] node14684;
	wire [4-1:0] node14688;
	wire [4-1:0] node14690;
	wire [4-1:0] node14694;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14701;
	wire [4-1:0] node14705;
	wire [4-1:0] node14706;
	wire [4-1:0] node14707;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14712;
	wire [4-1:0] node14714;
	wire [4-1:0] node14715;
	wire [4-1:0] node14718;
	wire [4-1:0] node14721;
	wire [4-1:0] node14722;
	wire [4-1:0] node14723;
	wire [4-1:0] node14725;
	wire [4-1:0] node14730;
	wire [4-1:0] node14731;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14737;
	wire [4-1:0] node14738;
	wire [4-1:0] node14739;
	wire [4-1:0] node14741;
	wire [4-1:0] node14745;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14750;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14756;
	wire [4-1:0] node14757;
	wire [4-1:0] node14760;
	wire [4-1:0] node14763;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14769;
	wire [4-1:0] node14771;
	wire [4-1:0] node14772;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14786;
	wire [4-1:0] node14788;
	wire [4-1:0] node14790;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14800;
	wire [4-1:0] node14801;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14814;
	wire [4-1:0] node14815;
	wire [4-1:0] node14817;
	wire [4-1:0] node14819;
	wire [4-1:0] node14822;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14829;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14833;
	wire [4-1:0] node14837;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14845;
	wire [4-1:0] node14848;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14853;
	wire [4-1:0] node14856;
	wire [4-1:0] node14857;
	wire [4-1:0] node14861;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14864;
	wire [4-1:0] node14869;
	wire [4-1:0] node14870;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14877;
	wire [4-1:0] node14879;
	wire [4-1:0] node14881;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14887;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14894;
	wire [4-1:0] node14897;
	wire [4-1:0] node14899;
	wire [4-1:0] node14900;
	wire [4-1:0] node14902;
	wire [4-1:0] node14905;
	wire [4-1:0] node14908;
	wire [4-1:0] node14909;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14915;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14921;
	wire [4-1:0] node14924;
	wire [4-1:0] node14925;
	wire [4-1:0] node14929;
	wire [4-1:0] node14930;
	wire [4-1:0] node14931;
	wire [4-1:0] node14933;
	wire [4-1:0] node14935;
	wire [4-1:0] node14938;
	wire [4-1:0] node14939;
	wire [4-1:0] node14941;
	wire [4-1:0] node14944;
	wire [4-1:0] node14947;
	wire [4-1:0] node14948;
	wire [4-1:0] node14950;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14957;
	wire [4-1:0] node14958;
	wire [4-1:0] node14962;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14965;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14970;
	wire [4-1:0] node14973;
	wire [4-1:0] node14976;
	wire [4-1:0] node14977;
	wire [4-1:0] node14980;
	wire [4-1:0] node14982;
	wire [4-1:0] node14985;
	wire [4-1:0] node14986;
	wire [4-1:0] node14987;
	wire [4-1:0] node14989;
	wire [4-1:0] node14992;
	wire [4-1:0] node14995;
	wire [4-1:0] node14996;
	wire [4-1:0] node14999;
	wire [4-1:0] node15000;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15006;
	wire [4-1:0] node15008;
	wire [4-1:0] node15009;
	wire [4-1:0] node15013;
	wire [4-1:0] node15015;
	wire [4-1:0] node15018;
	wire [4-1:0] node15019;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15025;
	wire [4-1:0] node15026;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15033;
	wire [4-1:0] node15034;
	wire [4-1:0] node15037;
	wire [4-1:0] node15038;
	wire [4-1:0] node15043;
	wire [4-1:0] node15044;
	wire [4-1:0] node15048;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15058;
	wire [4-1:0] node15059;
	wire [4-1:0] node15062;
	wire [4-1:0] node15065;
	wire [4-1:0] node15066;
	wire [4-1:0] node15067;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15074;
	wire [4-1:0] node15075;
	wire [4-1:0] node15076;
	wire [4-1:0] node15081;
	wire [4-1:0] node15082;
	wire [4-1:0] node15084;
	wire [4-1:0] node15086;
	wire [4-1:0] node15089;
	wire [4-1:0] node15090;
	wire [4-1:0] node15092;
	wire [4-1:0] node15096;
	wire [4-1:0] node15097;
	wire [4-1:0] node15098;
	wire [4-1:0] node15099;
	wire [4-1:0] node15101;
	wire [4-1:0] node15104;
	wire [4-1:0] node15105;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15112;
	wire [4-1:0] node15115;
	wire [4-1:0] node15117;
	wire [4-1:0] node15120;
	wire [4-1:0] node15121;
	wire [4-1:0] node15122;
	wire [4-1:0] node15124;
	wire [4-1:0] node15127;
	wire [4-1:0] node15128;
	wire [4-1:0] node15130;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15137;
	wire [4-1:0] node15140;
	wire [4-1:0] node15141;
	wire [4-1:0] node15142;
	wire [4-1:0] node15147;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15151;
	wire [4-1:0] node15152;
	wire [4-1:0] node15153;
	wire [4-1:0] node15154;
	wire [4-1:0] node15158;
	wire [4-1:0] node15159;
	wire [4-1:0] node15160;
	wire [4-1:0] node15164;
	wire [4-1:0] node15165;
	wire [4-1:0] node15169;
	wire [4-1:0] node15170;
	wire [4-1:0] node15171;
	wire [4-1:0] node15173;
	wire [4-1:0] node15175;
	wire [4-1:0] node15178;
	wire [4-1:0] node15179;
	wire [4-1:0] node15183;
	wire [4-1:0] node15185;
	wire [4-1:0] node15186;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15195;
	wire [4-1:0] node15197;
	wire [4-1:0] node15200;
	wire [4-1:0] node15201;
	wire [4-1:0] node15203;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15210;
	wire [4-1:0] node15212;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15220;
	wire [4-1:0] node15221;
	wire [4-1:0] node15223;
	wire [4-1:0] node15225;
	wire [4-1:0] node15228;
	wire [4-1:0] node15231;
	wire [4-1:0] node15232;
	wire [4-1:0] node15233;
	wire [4-1:0] node15234;
	wire [4-1:0] node15236;
	wire [4-1:0] node15239;
	wire [4-1:0] node15240;
	wire [4-1:0] node15242;
	wire [4-1:0] node15243;
	wire [4-1:0] node15247;
	wire [4-1:0] node15250;
	wire [4-1:0] node15251;
	wire [4-1:0] node15252;
	wire [4-1:0] node15253;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15262;
	wire [4-1:0] node15263;
	wire [4-1:0] node15267;
	wire [4-1:0] node15268;
	wire [4-1:0] node15269;
	wire [4-1:0] node15271;
	wire [4-1:0] node15272;
	wire [4-1:0] node15274;
	wire [4-1:0] node15276;
	wire [4-1:0] node15279;
	wire [4-1:0] node15281;
	wire [4-1:0] node15284;
	wire [4-1:0] node15286;
	wire [4-1:0] node15287;
	wire [4-1:0] node15289;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15295;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15299;
	wire [4-1:0] node15304;
	wire [4-1:0] node15306;
	wire [4-1:0] node15309;
	wire [4-1:0] node15310;
	wire [4-1:0] node15312;
	wire [4-1:0] node15316;
	wire [4-1:0] node15317;
	wire [4-1:0] node15318;
	wire [4-1:0] node15319;
	wire [4-1:0] node15320;
	wire [4-1:0] node15322;
	wire [4-1:0] node15325;
	wire [4-1:0] node15327;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15334;
	wire [4-1:0] node15335;
	wire [4-1:0] node15339;
	wire [4-1:0] node15341;
	wire [4-1:0] node15342;
	wire [4-1:0] node15344;
	wire [4-1:0] node15347;
	wire [4-1:0] node15349;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15354;
	wire [4-1:0] node15357;
	wire [4-1:0] node15360;
	wire [4-1:0] node15361;
	wire [4-1:0] node15363;
	wire [4-1:0] node15364;
	wire [4-1:0] node15368;
	wire [4-1:0] node15369;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15375;
	wire [4-1:0] node15376;
	wire [4-1:0] node15377;
	wire [4-1:0] node15378;
	wire [4-1:0] node15379;
	wire [4-1:0] node15380;
	wire [4-1:0] node15381;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15408;
	wire [4-1:0] node15409;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15417;
	wire [4-1:0] node15419;
	wire [4-1:0] node15420;
	wire [4-1:0] node15423;
	wire [4-1:0] node15426;
	wire [4-1:0] node15427;
	wire [4-1:0] node15428;
	wire [4-1:0] node15432;
	wire [4-1:0] node15434;
	wire [4-1:0] node15437;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15443;
	wire [4-1:0] node15447;
	wire [4-1:0] node15448;
	wire [4-1:0] node15452;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15455;
	wire [4-1:0] node15456;
	wire [4-1:0] node15458;
	wire [4-1:0] node15459;
	wire [4-1:0] node15464;
	wire [4-1:0] node15466;
	wire [4-1:0] node15467;
	wire [4-1:0] node15469;
	wire [4-1:0] node15473;
	wire [4-1:0] node15474;
	wire [4-1:0] node15476;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15483;
	wire [4-1:0] node15484;
	wire [4-1:0] node15486;
	wire [4-1:0] node15490;
	wire [4-1:0] node15491;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15495;
	wire [4-1:0] node15498;
	wire [4-1:0] node15502;
	wire [4-1:0] node15503;
	wire [4-1:0] node15504;
	wire [4-1:0] node15507;
	wire [4-1:0] node15510;
	wire [4-1:0] node15511;
	wire [4-1:0] node15515;
	wire [4-1:0] node15516;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15523;
	wire [4-1:0] node15524;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15532;
	wire [4-1:0] node15536;
	wire [4-1:0] node15537;
	wire [4-1:0] node15542;
	wire [4-1:0] node15543;
	wire [4-1:0] node15544;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15549;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15554;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15560;
	wire [4-1:0] node15563;
	wire [4-1:0] node15565;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15571;
	wire [4-1:0] node15576;
	wire [4-1:0] node15577;
	wire [4-1:0] node15579;
	wire [4-1:0] node15580;
	wire [4-1:0] node15583;
	wire [4-1:0] node15586;
	wire [4-1:0] node15587;
	wire [4-1:0] node15589;
	wire [4-1:0] node15592;
	wire [4-1:0] node15594;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15604;
	wire [4-1:0] node15608;
	wire [4-1:0] node15609;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15618;
	wire [4-1:0] node15619;
	wire [4-1:0] node15621;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15628;
	wire [4-1:0] node15631;
	wire [4-1:0] node15632;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15638;
	wire [4-1:0] node15642;
	wire [4-1:0] node15644;
	wire [4-1:0] node15646;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15651;
	wire [4-1:0] node15654;
	wire [4-1:0] node15657;
	wire [4-1:0] node15658;
	wire [4-1:0] node15661;
	wire [4-1:0] node15664;
	wire [4-1:0] node15665;
	wire [4-1:0] node15666;
	wire [4-1:0] node15667;
	wire [4-1:0] node15668;
	wire [4-1:0] node15669;
	wire [4-1:0] node15670;
	wire [4-1:0] node15671;
	wire [4-1:0] node15674;
	wire [4-1:0] node15677;
	wire [4-1:0] node15680;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15687;
	wire [4-1:0] node15689;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15696;
	wire [4-1:0] node15699;
	wire [4-1:0] node15700;
	wire [4-1:0] node15703;
	wire [4-1:0] node15706;
	wire [4-1:0] node15707;
	wire [4-1:0] node15709;
	wire [4-1:0] node15712;
	wire [4-1:0] node15714;
	wire [4-1:0] node15717;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15721;
	wire [4-1:0] node15722;
	wire [4-1:0] node15723;
	wire [4-1:0] node15728;
	wire [4-1:0] node15730;
	wire [4-1:0] node15732;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15739;
	wire [4-1:0] node15740;
	wire [4-1:0] node15743;
	wire [4-1:0] node15745;
	wire [4-1:0] node15746;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15752;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15755;
	wire [4-1:0] node15759;
	wire [4-1:0] node15760;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15766;
	wire [4-1:0] node15768;
	wire [4-1:0] node15772;
	wire [4-1:0] node15773;
	wire [4-1:0] node15777;
	wire [4-1:0] node15778;
	wire [4-1:0] node15779;
	wire [4-1:0] node15781;
	wire [4-1:0] node15784;
	wire [4-1:0] node15787;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15794;
	wire [4-1:0] node15796;
	wire [4-1:0] node15799;
	wire [4-1:0] node15801;
	wire [4-1:0] node15803;
	wire [4-1:0] node15806;
	wire [4-1:0] node15807;
	wire [4-1:0] node15808;
	wire [4-1:0] node15809;
	wire [4-1:0] node15810;
	wire [4-1:0] node15813;
	wire [4-1:0] node15816;
	wire [4-1:0] node15818;
	wire [4-1:0] node15821;
	wire [4-1:0] node15822;
	wire [4-1:0] node15825;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15830;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15841;
	wire [4-1:0] node15843;
	wire [4-1:0] node15844;
	wire [4-1:0] node15848;
	wire [4-1:0] node15849;
	wire [4-1:0] node15853;
	wire [4-1:0] node15854;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15860;
	wire [4-1:0] node15863;
	wire [4-1:0] node15864;
	wire [4-1:0] node15865;
	wire [4-1:0] node15867;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15877;
	wire [4-1:0] node15878;
	wire [4-1:0] node15879;
	wire [4-1:0] node15880;
	wire [4-1:0] node15883;
	wire [4-1:0] node15887;
	wire [4-1:0] node15889;
	wire [4-1:0] node15891;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15896;
	wire [4-1:0] node15897;
	wire [4-1:0] node15898;
	wire [4-1:0] node15901;
	wire [4-1:0] node15903;
	wire [4-1:0] node15904;
	wire [4-1:0] node15908;
	wire [4-1:0] node15910;
	wire [4-1:0] node15913;
	wire [4-1:0] node15914;
	wire [4-1:0] node15916;
	wire [4-1:0] node15917;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15928;
	wire [4-1:0] node15929;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15935;
	wire [4-1:0] node15936;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15942;
	wire [4-1:0] node15946;
	wire [4-1:0] node15947;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15953;
	wire [4-1:0] node15954;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15958;
	wire [4-1:0] node15962;
	wire [4-1:0] node15963;
	wire [4-1:0] node15967;
	wire [4-1:0] node15968;
	wire [4-1:0] node15969;
	wire [4-1:0] node15972;
	wire [4-1:0] node15975;
	wire [4-1:0] node15976;
	wire [4-1:0] node15978;
	wire [4-1:0] node15982;
	wire [4-1:0] node15983;
	wire [4-1:0] node15984;
	wire [4-1:0] node15986;
	wire [4-1:0] node15989;
	wire [4-1:0] node15991;
	wire [4-1:0] node15992;
	wire [4-1:0] node15994;
	wire [4-1:0] node15998;
	wire [4-1:0] node15999;
	wire [4-1:0] node16001;
	wire [4-1:0] node16002;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16014;
	wire [4-1:0] node16017;
	wire [4-1:0] node16018;
	wire [4-1:0] node16019;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16022;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16029;
	wire [4-1:0] node16030;
	wire [4-1:0] node16034;
	wire [4-1:0] node16037;
	wire [4-1:0] node16038;
	wire [4-1:0] node16041;
	wire [4-1:0] node16044;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16050;
	wire [4-1:0] node16051;
	wire [4-1:0] node16052;
	wire [4-1:0] node16055;
	wire [4-1:0] node16058;
	wire [4-1:0] node16060;
	wire [4-1:0] node16061;
	wire [4-1:0] node16065;
	wire [4-1:0] node16066;
	wire [4-1:0] node16067;
	wire [4-1:0] node16068;
	wire [4-1:0] node16072;
	wire [4-1:0] node16074;
	wire [4-1:0] node16076;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16082;
	wire [4-1:0] node16083;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16090;
	wire [4-1:0] node16091;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16094;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16100;
	wire [4-1:0] node16103;
	wire [4-1:0] node16104;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16111;
	wire [4-1:0] node16113;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16118;
	wire [4-1:0] node16119;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16128;
	wire [4-1:0] node16130;
	wire [4-1:0] node16132;
	wire [4-1:0] node16133;
	wire [4-1:0] node16135;
	wire [4-1:0] node16139;
	wire [4-1:0] node16140;
	wire [4-1:0] node16141;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16149;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16156;
	wire [4-1:0] node16157;
	wire [4-1:0] node16161;
	wire [4-1:0] node16163;
	wire [4-1:0] node16165;
	wire [4-1:0] node16167;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16174;
	wire [4-1:0] node16177;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16184;
	wire [4-1:0] node16187;
	wire [4-1:0] node16188;
	wire [4-1:0] node16190;
	wire [4-1:0] node16193;
	wire [4-1:0] node16194;
	wire [4-1:0] node16197;
	wire [4-1:0] node16200;
	wire [4-1:0] node16201;
	wire [4-1:0] node16202;
	wire [4-1:0] node16203;
	wire [4-1:0] node16206;
	wire [4-1:0] node16209;
	wire [4-1:0] node16210;
	wire [4-1:0] node16213;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16221;
	wire [4-1:0] node16222;
	wire [4-1:0] node16225;
	wire [4-1:0] node16226;
	wire [4-1:0] node16230;
	wire [4-1:0] node16231;
	wire [4-1:0] node16234;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16239;
	wire [4-1:0] node16240;
	wire [4-1:0] node16241;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16247;
	wire [4-1:0] node16249;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16265;
	wire [4-1:0] node16266;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16274;
	wire [4-1:0] node16277;
	wire [4-1:0] node16280;
	wire [4-1:0] node16282;
	wire [4-1:0] node16285;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16295;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16300;
	wire [4-1:0] node16301;
	wire [4-1:0] node16305;
	wire [4-1:0] node16308;
	wire [4-1:0] node16309;
	wire [4-1:0] node16313;
	wire [4-1:0] node16314;
	wire [4-1:0] node16315;
	wire [4-1:0] node16316;
	wire [4-1:0] node16318;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16329;
	wire [4-1:0] node16332;
	wire [4-1:0] node16333;
	wire [4-1:0] node16334;
	wire [4-1:0] node16336;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16344;
	wire [4-1:0] node16345;
	wire [4-1:0] node16349;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16352;
	wire [4-1:0] node16355;
	wire [4-1:0] node16358;
	wire [4-1:0] node16360;
	wire [4-1:0] node16362;
	wire [4-1:0] node16365;
	wire [4-1:0] node16366;
	wire [4-1:0] node16367;
	wire [4-1:0] node16368;
	wire [4-1:0] node16371;
	wire [4-1:0] node16373;
	wire [4-1:0] node16376;
	wire [4-1:0] node16377;
	wire [4-1:0] node16379;
	wire [4-1:0] node16383;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16387;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16395;
	wire [4-1:0] node16396;
	wire [4-1:0] node16397;
	wire [4-1:0] node16398;
	wire [4-1:0] node16399;
	wire [4-1:0] node16403;
	wire [4-1:0] node16406;
	wire [4-1:0] node16407;
	wire [4-1:0] node16408;
	wire [4-1:0] node16412;
	wire [4-1:0] node16413;
	wire [4-1:0] node16416;
	wire [4-1:0] node16419;
	wire [4-1:0] node16421;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16427;
	wire [4-1:0] node16429;
	wire [4-1:0] node16431;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16436;
	wire [4-1:0] node16437;
	wire [4-1:0] node16440;
	wire [4-1:0] node16443;
	wire [4-1:0] node16445;
	wire [4-1:0] node16448;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16453;
	wire [4-1:0] node16456;
	wire [4-1:0] node16457;
	wire [4-1:0] node16459;
	wire [4-1:0] node16462;
	wire [4-1:0] node16463;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16471;
	wire [4-1:0] node16472;
	wire [4-1:0] node16473;
	wire [4-1:0] node16475;
	wire [4-1:0] node16480;
	wire [4-1:0] node16481;
	wire [4-1:0] node16482;
	wire [4-1:0] node16484;
	wire [4-1:0] node16487;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16494;
	wire [4-1:0] node16496;
	wire [4-1:0] node16498;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16503;
	wire [4-1:0] node16505;
	wire [4-1:0] node16507;
	wire [4-1:0] node16508;
	wire [4-1:0] node16512;
	wire [4-1:0] node16513;
	wire [4-1:0] node16517;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16528;
	wire [4-1:0] node16533;
	wire [4-1:0] node16535;
	wire [4-1:0] node16536;
	wire [4-1:0] node16538;
	wire [4-1:0] node16542;
	wire [4-1:0] node16543;
	wire [4-1:0] node16544;
	wire [4-1:0] node16545;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16549;
	wire [4-1:0] node16550;
	wire [4-1:0] node16553;
	wire [4-1:0] node16555;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16562;
	wire [4-1:0] node16565;
	wire [4-1:0] node16568;
	wire [4-1:0] node16569;
	wire [4-1:0] node16571;
	wire [4-1:0] node16573;
	wire [4-1:0] node16574;
	wire [4-1:0] node16575;
	wire [4-1:0] node16578;
	wire [4-1:0] node16582;
	wire [4-1:0] node16583;
	wire [4-1:0] node16584;
	wire [4-1:0] node16589;
	wire [4-1:0] node16590;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16593;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16600;
	wire [4-1:0] node16602;
	wire [4-1:0] node16605;
	wire [4-1:0] node16606;
	wire [4-1:0] node16610;
	wire [4-1:0] node16612;
	wire [4-1:0] node16615;
	wire [4-1:0] node16616;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16629;
	wire [4-1:0] node16633;
	wire [4-1:0] node16634;
	wire [4-1:0] node16638;
	wire [4-1:0] node16639;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16644;
	wire [4-1:0] node16647;
	wire [4-1:0] node16648;
	wire [4-1:0] node16652;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16657;
	wire [4-1:0] node16660;
	wire [4-1:0] node16661;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16669;
	wire [4-1:0] node16672;
	wire [4-1:0] node16673;
	wire [4-1:0] node16674;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16680;
	wire [4-1:0] node16682;
	wire [4-1:0] node16685;
	wire [4-1:0] node16687;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16692;
	wire [4-1:0] node16696;
	wire [4-1:0] node16699;
	wire [4-1:0] node16700;
	wire [4-1:0] node16701;
	wire [4-1:0] node16702;
	wire [4-1:0] node16703;
	wire [4-1:0] node16704;
	wire [4-1:0] node16705;
	wire [4-1:0] node16708;
	wire [4-1:0] node16709;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16717;
	wire [4-1:0] node16718;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16721;
	wire [4-1:0] node16725;
	wire [4-1:0] node16726;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16732;
	wire [4-1:0] node16736;
	wire [4-1:0] node16737;
	wire [4-1:0] node16740;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16745;
	wire [4-1:0] node16748;
	wire [4-1:0] node16751;
	wire [4-1:0] node16753;
	wire [4-1:0] node16755;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16761;
	wire [4-1:0] node16763;
	wire [4-1:0] node16767;
	wire [4-1:0] node16768;
	wire [4-1:0] node16770;
	wire [4-1:0] node16773;
	wire [4-1:0] node16774;
	wire [4-1:0] node16776;
	wire [4-1:0] node16777;
	wire [4-1:0] node16780;
	wire [4-1:0] node16783;
	wire [4-1:0] node16784;
	wire [4-1:0] node16788;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16793;
	wire [4-1:0] node16796;
	wire [4-1:0] node16797;
	wire [4-1:0] node16798;
	wire [4-1:0] node16801;
	wire [4-1:0] node16804;
	wire [4-1:0] node16805;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16813;
	wire [4-1:0] node16814;
	wire [4-1:0] node16815;
	wire [4-1:0] node16816;
	wire [4-1:0] node16817;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16823;
	wire [4-1:0] node16825;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16830;
	wire [4-1:0] node16834;
	wire [4-1:0] node16836;
	wire [4-1:0] node16839;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16842;
	wire [4-1:0] node16847;
	wire [4-1:0] node16849;
	wire [4-1:0] node16851;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16857;
	wire [4-1:0] node16859;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16865;
	wire [4-1:0] node16867;
	wire [4-1:0] node16870;
	wire [4-1:0] node16871;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16878;
	wire [4-1:0] node16879;
	wire [4-1:0] node16883;
	wire [4-1:0] node16884;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16892;
	wire [4-1:0] node16893;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16899;
	wire [4-1:0] node16902;
	wire [4-1:0] node16905;
	wire [4-1:0] node16908;
	wire [4-1:0] node16909;
	wire [4-1:0] node16910;
	wire [4-1:0] node16911;
	wire [4-1:0] node16915;
	wire [4-1:0] node16916;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16923;
	wire [4-1:0] node16925;
	wire [4-1:0] node16929;
	wire [4-1:0] node16930;
	wire [4-1:0] node16931;
	wire [4-1:0] node16933;
	wire [4-1:0] node16936;
	wire [4-1:0] node16939;
	wire [4-1:0] node16940;
	wire [4-1:0] node16941;
	wire [4-1:0] node16944;
	wire [4-1:0] node16946;
	wire [4-1:0] node16949;
	wire [4-1:0] node16950;
	wire [4-1:0] node16952;
	wire [4-1:0] node16955;
	wire [4-1:0] node16957;
	wire [4-1:0] node16958;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16965;
	wire [4-1:0] node16966;
	wire [4-1:0] node16968;
	wire [4-1:0] node16971;
	wire [4-1:0] node16972;
	wire [4-1:0] node16973;
	wire [4-1:0] node16977;
	wire [4-1:0] node16978;
	wire [4-1:0] node16979;
	wire [4-1:0] node16984;
	wire [4-1:0] node16985;
	wire [4-1:0] node16986;
	wire [4-1:0] node16987;
	wire [4-1:0] node16989;
	wire [4-1:0] node16992;
	wire [4-1:0] node16993;
	wire [4-1:0] node16997;
	wire [4-1:0] node16998;
	wire [4-1:0] node17001;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17008;
	wire [4-1:0] node17011;
	wire [4-1:0] node17012;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17017;
	wire [4-1:0] node17020;
	wire [4-1:0] node17021;
	wire [4-1:0] node17022;
	wire [4-1:0] node17024;
	wire [4-1:0] node17027;
	wire [4-1:0] node17031;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17037;
	wire [4-1:0] node17040;
	wire [4-1:0] node17043;
	wire [4-1:0] node17044;
	wire [4-1:0] node17048;
	wire [4-1:0] node17049;
	wire [4-1:0] node17050;
	wire [4-1:0] node17051;
	wire [4-1:0] node17052;
	wire [4-1:0] node17055;
	wire [4-1:0] node17056;
	wire [4-1:0] node17057;
	wire [4-1:0] node17060;
	wire [4-1:0] node17064;
	wire [4-1:0] node17066;
	wire [4-1:0] node17067;
	wire [4-1:0] node17070;
	wire [4-1:0] node17073;
	wire [4-1:0] node17074;
	wire [4-1:0] node17075;
	wire [4-1:0] node17076;
	wire [4-1:0] node17080;
	wire [4-1:0] node17081;
	wire [4-1:0] node17082;
	wire [4-1:0] node17085;
	wire [4-1:0] node17088;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17096;
	wire [4-1:0] node17099;
	wire [4-1:0] node17100;
	wire [4-1:0] node17104;
	wire [4-1:0] node17105;
	wire [4-1:0] node17106;
	wire [4-1:0] node17109;
	wire [4-1:0] node17112;
	wire [4-1:0] node17113;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17119;
	wire [4-1:0] node17120;
	wire [4-1:0] node17122;
	wire [4-1:0] node17125;
	wire [4-1:0] node17127;
	wire [4-1:0] node17129;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17136;
	wire [4-1:0] node17139;
	wire [4-1:0] node17140;
	wire [4-1:0] node17141;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17148;
	wire [4-1:0] node17151;
	wire [4-1:0] node17152;
	wire [4-1:0] node17153;
	wire [4-1:0] node17156;
	wire [4-1:0] node17159;
	wire [4-1:0] node17160;
	wire [4-1:0] node17163;
	wire [4-1:0] node17166;
	wire [4-1:0] node17167;
	wire [4-1:0] node17168;
	wire [4-1:0] node17169;
	wire [4-1:0] node17171;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17176;
	wire [4-1:0] node17182;
	wire [4-1:0] node17183;
	wire [4-1:0] node17184;
	wire [4-1:0] node17185;
	wire [4-1:0] node17186;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17194;
	wire [4-1:0] node17197;
	wire [4-1:0] node17201;
	wire [4-1:0] node17202;
	wire [4-1:0] node17203;
	wire [4-1:0] node17206;
	wire [4-1:0] node17209;
	wire [4-1:0] node17210;
	wire [4-1:0] node17211;
	wire [4-1:0] node17213;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17220;
	wire [4-1:0] node17223;
	wire [4-1:0] node17224;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17230;
	wire [4-1:0] node17231;
	wire [4-1:0] node17232;
	wire [4-1:0] node17235;
	wire [4-1:0] node17239;
	wire [4-1:0] node17240;
	wire [4-1:0] node17241;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17248;
	wire [4-1:0] node17252;
	wire [4-1:0] node17253;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17263;
	wire [4-1:0] node17264;
	wire [4-1:0] node17268;
	wire [4-1:0] node17269;
	wire [4-1:0] node17270;
	wire [4-1:0] node17272;
	wire [4-1:0] node17276;
	wire [4-1:0] node17277;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17288;
	wire [4-1:0] node17289;
	wire [4-1:0] node17290;
	wire [4-1:0] node17293;
	wire [4-1:0] node17294;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17303;
	wire [4-1:0] node17305;
	wire [4-1:0] node17308;
	wire [4-1:0] node17309;
	wire [4-1:0] node17310;
	wire [4-1:0] node17311;
	wire [4-1:0] node17314;
	wire [4-1:0] node17317;
	wire [4-1:0] node17318;
	wire [4-1:0] node17320;
	wire [4-1:0] node17323;
	wire [4-1:0] node17324;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17332;
	wire [4-1:0] node17333;
	wire [4-1:0] node17337;
	wire [4-1:0] node17340;
	wire [4-1:0] node17341;
	wire [4-1:0] node17346;
	wire [4-1:0] node17347;
	wire [4-1:0] node17348;
	wire [4-1:0] node17350;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17357;
	wire [4-1:0] node17360;
	wire [4-1:0] node17362;
	wire [4-1:0] node17365;
	wire [4-1:0] node17366;
	wire [4-1:0] node17367;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17379;
	wire [4-1:0] node17380;
	wire [4-1:0] node17381;
	wire [4-1:0] node17382;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17392;
	wire [4-1:0] node17393;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17396;
	wire [4-1:0] node17397;
	wire [4-1:0] node17398;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17404;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17410;
	wire [4-1:0] node17413;
	wire [4-1:0] node17416;
	wire [4-1:0] node17417;
	wire [4-1:0] node17418;
	wire [4-1:0] node17419;
	wire [4-1:0] node17422;
	wire [4-1:0] node17425;
	wire [4-1:0] node17428;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17433;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17443;
	wire [4-1:0] node17444;
	wire [4-1:0] node17445;
	wire [4-1:0] node17446;
	wire [4-1:0] node17447;
	wire [4-1:0] node17449;
	wire [4-1:0] node17453;
	wire [4-1:0] node17456;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17460;
	wire [4-1:0] node17463;
	wire [4-1:0] node17464;
	wire [4-1:0] node17468;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17475;
	wire [4-1:0] node17476;
	wire [4-1:0] node17477;
	wire [4-1:0] node17480;
	wire [4-1:0] node17482;
	wire [4-1:0] node17485;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17488;
	wire [4-1:0] node17490;
	wire [4-1:0] node17493;
	wire [4-1:0] node17497;
	wire [4-1:0] node17498;
	wire [4-1:0] node17501;
	wire [4-1:0] node17504;
	wire [4-1:0] node17505;
	wire [4-1:0] node17506;
	wire [4-1:0] node17507;
	wire [4-1:0] node17509;
	wire [4-1:0] node17512;
	wire [4-1:0] node17513;
	wire [4-1:0] node17514;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17520;
	wire [4-1:0] node17524;
	wire [4-1:0] node17525;
	wire [4-1:0] node17527;
	wire [4-1:0] node17528;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17535;
	wire [4-1:0] node17537;
	wire [4-1:0] node17540;
	wire [4-1:0] node17541;
	wire [4-1:0] node17544;
	wire [4-1:0] node17547;
	wire [4-1:0] node17549;
	wire [4-1:0] node17552;
	wire [4-1:0] node17553;
	wire [4-1:0] node17554;
	wire [4-1:0] node17556;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17564;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17567;
	wire [4-1:0] node17570;
	wire [4-1:0] node17574;
	wire [4-1:0] node17577;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17580;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17584;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17589;
	wire [4-1:0] node17592;
	wire [4-1:0] node17596;
	wire [4-1:0] node17598;
	wire [4-1:0] node17599;
	wire [4-1:0] node17602;
	wire [4-1:0] node17604;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17612;
	wire [4-1:0] node17616;
	wire [4-1:0] node17617;
	wire [4-1:0] node17619;
	wire [4-1:0] node17620;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17628;
	wire [4-1:0] node17629;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17637;
	wire [4-1:0] node17638;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17648;
	wire [4-1:0] node17650;
	wire [4-1:0] node17653;
	wire [4-1:0] node17654;
	wire [4-1:0] node17656;
	wire [4-1:0] node17659;
	wire [4-1:0] node17660;
	wire [4-1:0] node17663;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17670;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17679;
	wire [4-1:0] node17680;
	wire [4-1:0] node17681;
	wire [4-1:0] node17682;
	wire [4-1:0] node17683;
	wire [4-1:0] node17684;
	wire [4-1:0] node17687;
	wire [4-1:0] node17690;
	wire [4-1:0] node17691;
	wire [4-1:0] node17696;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17705;
	wire [4-1:0] node17708;
	wire [4-1:0] node17709;
	wire [4-1:0] node17710;
	wire [4-1:0] node17713;
	wire [4-1:0] node17717;
	wire [4-1:0] node17718;
	wire [4-1:0] node17719;
	wire [4-1:0] node17720;
	wire [4-1:0] node17721;
	wire [4-1:0] node17723;
	wire [4-1:0] node17726;
	wire [4-1:0] node17728;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17734;
	wire [4-1:0] node17737;
	wire [4-1:0] node17740;
	wire [4-1:0] node17742;
	wire [4-1:0] node17743;
	wire [4-1:0] node17747;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17754;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17759;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17766;
	wire [4-1:0] node17768;
	wire [4-1:0] node17771;
	wire [4-1:0] node17772;
	wire [4-1:0] node17773;
	wire [4-1:0] node17774;
	wire [4-1:0] node17776;
	wire [4-1:0] node17780;
	wire [4-1:0] node17784;
	wire [4-1:0] node17785;
	wire [4-1:0] node17786;
	wire [4-1:0] node17788;
	wire [4-1:0] node17791;
	wire [4-1:0] node17793;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17798;
	wire [4-1:0] node17800;
	wire [4-1:0] node17803;
	wire [4-1:0] node17805;
	wire [4-1:0] node17808;
	wire [4-1:0] node17809;
	wire [4-1:0] node17813;
	wire [4-1:0] node17814;
	wire [4-1:0] node17815;
	wire [4-1:0] node17816;
	wire [4-1:0] node17818;
	wire [4-1:0] node17821;
	wire [4-1:0] node17822;
	wire [4-1:0] node17823;
	wire [4-1:0] node17828;
	wire [4-1:0] node17830;
	wire [4-1:0] node17832;
	wire [4-1:0] node17833;
	wire [4-1:0] node17835;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17841;
	wire [4-1:0] node17842;
	wire [4-1:0] node17845;
	wire [4-1:0] node17848;
	wire [4-1:0] node17849;
	wire [4-1:0] node17850;
	wire [4-1:0] node17855;
	wire [4-1:0] node17856;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17860;
	wire [4-1:0] node17861;
	wire [4-1:0] node17866;
	wire [4-1:0] node17868;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17875;
	wire [4-1:0] node17878;
	wire [4-1:0] node17879;
	wire [4-1:0] node17880;
	wire [4-1:0] node17881;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17887;
	wire [4-1:0] node17888;
	wire [4-1:0] node17891;
	wire [4-1:0] node17892;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17903;
	wire [4-1:0] node17905;
	wire [4-1:0] node17908;
	wire [4-1:0] node17909;
	wire [4-1:0] node17910;
	wire [4-1:0] node17911;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17919;
	wire [4-1:0] node17920;
	wire [4-1:0] node17921;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17930;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17936;
	wire [4-1:0] node17938;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17943;
	wire [4-1:0] node17946;
	wire [4-1:0] node17947;
	wire [4-1:0] node17951;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17957;
	wire [4-1:0] node17958;
	wire [4-1:0] node17962;
	wire [4-1:0] node17964;
	wire [4-1:0] node17966;
	wire [4-1:0] node17967;
	wire [4-1:0] node17968;
	wire [4-1:0] node17972;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17979;
	wire [4-1:0] node17982;
	wire [4-1:0] node17985;
	wire [4-1:0] node17986;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17998;
	wire [4-1:0] node17999;
	wire [4-1:0] node18000;
	wire [4-1:0] node18001;
	wire [4-1:0] node18003;
	wire [4-1:0] node18004;
	wire [4-1:0] node18009;
	wire [4-1:0] node18011;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18020;
	wire [4-1:0] node18022;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18028;
	wire [4-1:0] node18032;
	wire [4-1:0] node18034;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18042;
	wire [4-1:0] node18044;
	wire [4-1:0] node18047;
	wire [4-1:0] node18049;
	wire [4-1:0] node18052;
	wire [4-1:0] node18053;
	wire [4-1:0] node18054;
	wire [4-1:0] node18058;
	wire [4-1:0] node18060;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18068;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18073;
	wire [4-1:0] node18076;
	wire [4-1:0] node18079;
	wire [4-1:0] node18080;
	wire [4-1:0] node18083;
	wire [4-1:0] node18086;
	wire [4-1:0] node18087;
	wire [4-1:0] node18088;
	wire [4-1:0] node18089;
	wire [4-1:0] node18090;
	wire [4-1:0] node18091;
	wire [4-1:0] node18095;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18101;
	wire [4-1:0] node18105;
	wire [4-1:0] node18106;
	wire [4-1:0] node18107;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18114;
	wire [4-1:0] node18115;
	wire [4-1:0] node18117;
	wire [4-1:0] node18119;
	wire [4-1:0] node18120;
	wire [4-1:0] node18123;
	wire [4-1:0] node18126;
	wire [4-1:0] node18128;
	wire [4-1:0] node18129;
	wire [4-1:0] node18130;
	wire [4-1:0] node18133;
	wire [4-1:0] node18138;
	wire [4-1:0] node18139;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18147;
	wire [4-1:0] node18150;
	wire [4-1:0] node18153;
	wire [4-1:0] node18154;
	wire [4-1:0] node18157;
	wire [4-1:0] node18160;
	wire [4-1:0] node18161;
	wire [4-1:0] node18162;
	wire [4-1:0] node18163;
	wire [4-1:0] node18165;
	wire [4-1:0] node18168;
	wire [4-1:0] node18169;
	wire [4-1:0] node18171;
	wire [4-1:0] node18173;
	wire [4-1:0] node18174;
	wire [4-1:0] node18178;
	wire [4-1:0] node18179;
	wire [4-1:0] node18180;
	wire [4-1:0] node18185;
	wire [4-1:0] node18186;
	wire [4-1:0] node18189;
	wire [4-1:0] node18192;
	wire [4-1:0] node18193;
	wire [4-1:0] node18194;
	wire [4-1:0] node18196;
	wire [4-1:0] node18199;
	wire [4-1:0] node18200;
	wire [4-1:0] node18202;
	wire [4-1:0] node18205;
	wire [4-1:0] node18207;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18212;
	wire [4-1:0] node18216;
	wire [4-1:0] node18217;
	wire [4-1:0] node18220;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18225;
	wire [4-1:0] node18229;
	wire [4-1:0] node18230;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18236;
	wire [4-1:0] node18237;
	wire [4-1:0] node18238;
	wire [4-1:0] node18239;
	wire [4-1:0] node18240;
	wire [4-1:0] node18241;
	wire [4-1:0] node18244;
	wire [4-1:0] node18245;
	wire [4-1:0] node18249;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18255;
	wire [4-1:0] node18256;
	wire [4-1:0] node18258;
	wire [4-1:0] node18259;
	wire [4-1:0] node18260;
	wire [4-1:0] node18263;
	wire [4-1:0] node18267;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18272;
	wire [4-1:0] node18273;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18280;
	wire [4-1:0] node18283;
	wire [4-1:0] node18286;
	wire [4-1:0] node18287;
	wire [4-1:0] node18288;
	wire [4-1:0] node18289;
	wire [4-1:0] node18291;
	wire [4-1:0] node18296;
	wire [4-1:0] node18298;
	wire [4-1:0] node18299;
	wire [4-1:0] node18302;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18307;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18319;
	wire [4-1:0] node18320;
	wire [4-1:0] node18322;
	wire [4-1:0] node18325;
	wire [4-1:0] node18327;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18333;
	wire [4-1:0] node18338;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18342;
	wire [4-1:0] node18343;
	wire [4-1:0] node18347;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18353;
	wire [4-1:0] node18354;
	wire [4-1:0] node18358;
	wire [4-1:0] node18361;
	wire [4-1:0] node18362;
	wire [4-1:0] node18363;
	wire [4-1:0] node18364;
	wire [4-1:0] node18369;
	wire [4-1:0] node18370;
	wire [4-1:0] node18371;
	wire [4-1:0] node18376;
	wire [4-1:0] node18377;
	wire [4-1:0] node18378;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18384;
	wire [4-1:0] node18387;
	wire [4-1:0] node18388;
	wire [4-1:0] node18390;
	wire [4-1:0] node18393;
	wire [4-1:0] node18394;
	wire [4-1:0] node18397;
	wire [4-1:0] node18400;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18403;
	wire [4-1:0] node18408;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18419;
	wire [4-1:0] node18421;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18424;
	wire [4-1:0] node18426;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18435;
	wire [4-1:0] node18438;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18448;
	wire [4-1:0] node18451;
	wire [4-1:0] node18454;
	wire [4-1:0] node18455;
	wire [4-1:0] node18456;
	wire [4-1:0] node18457;
	wire [4-1:0] node18462;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18475;
	wire [4-1:0] node18476;
	wire [4-1:0] node18480;
	wire [4-1:0] node18481;
	wire [4-1:0] node18482;
	wire [4-1:0] node18483;
	wire [4-1:0] node18484;
	wire [4-1:0] node18485;
	wire [4-1:0] node18486;
	wire [4-1:0] node18487;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18499;
	wire [4-1:0] node18501;
	wire [4-1:0] node18504;
	wire [4-1:0] node18505;
	wire [4-1:0] node18508;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18513;
	wire [4-1:0] node18514;
	wire [4-1:0] node18515;
	wire [4-1:0] node18521;
	wire [4-1:0] node18522;
	wire [4-1:0] node18523;
	wire [4-1:0] node18525;
	wire [4-1:0] node18526;
	wire [4-1:0] node18532;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18536;
	wire [4-1:0] node18537;
	wire [4-1:0] node18538;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18548;
	wire [4-1:0] node18551;
	wire [4-1:0] node18552;
	wire [4-1:0] node18553;
	wire [4-1:0] node18554;
	wire [4-1:0] node18555;
	wire [4-1:0] node18561;
	wire [4-1:0] node18564;
	wire [4-1:0] node18565;
	wire [4-1:0] node18566;
	wire [4-1:0] node18569;
	wire [4-1:0] node18572;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18577;
	wire [4-1:0] node18580;
	wire [4-1:0] node18581;
	wire [4-1:0] node18584;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18589;
	wire [4-1:0] node18590;
	wire [4-1:0] node18591;
	wire [4-1:0] node18592;
	wire [4-1:0] node18594;
	wire [4-1:0] node18596;
	wire [4-1:0] node18599;
	wire [4-1:0] node18601;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18608;
	wire [4-1:0] node18611;
	wire [4-1:0] node18612;
	wire [4-1:0] node18614;
	wire [4-1:0] node18617;
	wire [4-1:0] node18618;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18629;
	wire [4-1:0] node18630;
	wire [4-1:0] node18631;
	wire [4-1:0] node18632;
	wire [4-1:0] node18633;
	wire [4-1:0] node18636;
	wire [4-1:0] node18638;
	wire [4-1:0] node18641;
	wire [4-1:0] node18642;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18657;
	wire [4-1:0] node18658;
	wire [4-1:0] node18659;
	wire [4-1:0] node18664;
	wire [4-1:0] node18665;
	wire [4-1:0] node18666;
	wire [4-1:0] node18667;
	wire [4-1:0] node18668;
	wire [4-1:0] node18669;
	wire [4-1:0] node18673;
	wire [4-1:0] node18674;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18684;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18689;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;

	assign outp = (inp[3]) ? node10486 : node1;
		assign node1 = (inp[6]) ? node6101 : node2;
			assign node2 = (inp[14]) ? node2922 : node3;
				assign node3 = (inp[8]) ? node1547 : node4;
					assign node4 = (inp[12]) ? node754 : node5;
						assign node5 = (inp[7]) ? node379 : node6;
							assign node6 = (inp[4]) ? node196 : node7;
								assign node7 = (inp[0]) ? node91 : node8;
									assign node8 = (inp[13]) ? node46 : node9;
										assign node9 = (inp[2]) ? node27 : node10;
											assign node10 = (inp[9]) ? node22 : node11;
												assign node11 = (inp[5]) ? node17 : node12;
													assign node12 = (inp[15]) ? 4'b0000 : node13;
														assign node13 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node17 = (inp[10]) ? 4'b0101 : node18;
														assign node18 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node22 = (inp[10]) ? node24 : 4'b0001;
													assign node24 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node27 = (inp[1]) ? node35 : node28;
												assign node28 = (inp[9]) ? node32 : node29;
													assign node29 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node32 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node35 = (inp[5]) ? node39 : node36;
													assign node36 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node39 = (inp[15]) ? node41 : 4'b0000;
														assign node41 = (inp[10]) ? 4'b0000 : node42;
															assign node42 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node46 = (inp[2]) ? node64 : node47;
											assign node47 = (inp[1]) ? node59 : node48;
												assign node48 = (inp[5]) ? node50 : 4'b0101;
													assign node50 = (inp[15]) ? node52 : 4'b0100;
														assign node52 = (inp[10]) ? node56 : node53;
															assign node53 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node56 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node59 = (inp[5]) ? 4'b0001 : node60;
													assign node60 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node64 = (inp[5]) ? node80 : node65;
												assign node65 = (inp[11]) ? node69 : node66;
													assign node66 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node69 = (inp[1]) ? node71 : 4'b0000;
														assign node71 = (inp[10]) ? 4'b0001 : node72;
															assign node72 = (inp[15]) ? node76 : node73;
																assign node73 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node76 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node80 = (inp[1]) ? node88 : node81;
													assign node81 = (inp[9]) ? node83 : 4'b0000;
														assign node83 = (inp[10]) ? 4'b0001 : node84;
															assign node84 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node88 = (inp[15]) ? 4'b0101 : 4'b0100;
									assign node91 = (inp[9]) ? node147 : node92;
										assign node92 = (inp[15]) ? node110 : node93;
											assign node93 = (inp[10]) ? node99 : node94;
												assign node94 = (inp[5]) ? 4'b0001 : node95;
													assign node95 = (inp[11]) ? 4'b0101 : 4'b0001;
												assign node99 = (inp[1]) ? node105 : node100;
													assign node100 = (inp[13]) ? node102 : 4'b0000;
														assign node102 = (inp[2]) ? 4'b0000 : 4'b0101;
													assign node105 = (inp[2]) ? node107 : 4'b0000;
														assign node107 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node110 = (inp[1]) ? node124 : node111;
												assign node111 = (inp[10]) ? node117 : node112;
													assign node112 = (inp[13]) ? 4'b0000 : node113;
														assign node113 = (inp[11]) ? 4'b0101 : 4'b0000;
													assign node117 = (inp[11]) ? node119 : 4'b0101;
														assign node119 = (inp[5]) ? 4'b0000 : node120;
															assign node120 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node124 = (inp[5]) ? node132 : node125;
													assign node125 = (inp[2]) ? node129 : node126;
														assign node126 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node129 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node132 = (inp[13]) ? node138 : node133;
														assign node133 = (inp[11]) ? 4'b0000 : node134;
															assign node134 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node138 = (inp[2]) ? node140 : 4'b0000;
															assign node140 = (inp[11]) ? node144 : node141;
																assign node141 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node144 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node147 = (inp[2]) ? node175 : node148;
											assign node148 = (inp[15]) ? node160 : node149;
												assign node149 = (inp[13]) ? node151 : 4'b0001;
													assign node151 = (inp[1]) ? node157 : node152;
														assign node152 = (inp[5]) ? node154 : 4'b0101;
															assign node154 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node157 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node160 = (inp[11]) ? node172 : node161;
													assign node161 = (inp[1]) ? node165 : node162;
														assign node162 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node165 = (inp[5]) ? node167 : 4'b0001;
															assign node167 = (inp[13]) ? 4'b0001 : node168;
																assign node168 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node172 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node175 = (inp[13]) ? node191 : node176;
												assign node176 = (inp[1]) ? 4'b0100 : node177;
													assign node177 = (inp[5]) ? node179 : 4'b0101;
														assign node179 = (inp[15]) ? node185 : node180;
															assign node180 = (inp[10]) ? 4'b0100 : node181;
																assign node181 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node185 = (inp[10]) ? node187 : 4'b0100;
																assign node187 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node191 = (inp[1]) ? node193 : 4'b0000;
													assign node193 = (inp[11]) ? 4'b0101 : 4'b0100;
								assign node196 = (inp[15]) ? node300 : node197;
									assign node197 = (inp[13]) ? node255 : node198;
										assign node198 = (inp[1]) ? node210 : node199;
											assign node199 = (inp[2]) ? node205 : node200;
												assign node200 = (inp[5]) ? node202 : 4'b0001;
													assign node202 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node205 = (inp[9]) ? node207 : 4'b0101;
													assign node207 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node210 = (inp[11]) ? node228 : node211;
												assign node211 = (inp[2]) ? node225 : node212;
													assign node212 = (inp[10]) ? node218 : node213;
														assign node213 = (inp[9]) ? node215 : 4'b0100;
															assign node215 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node218 = (inp[9]) ? node222 : node219;
															assign node219 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node222 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node225 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node228 = (inp[10]) ? node238 : node229;
													assign node229 = (inp[0]) ? node231 : 4'b0100;
														assign node231 = (inp[9]) ? 4'b0101 : node232;
															assign node232 = (inp[5]) ? node234 : 4'b0001;
																assign node234 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node238 = (inp[9]) ? node244 : node239;
														assign node239 = (inp[5]) ? node241 : 4'b0000;
															assign node241 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node244 = (inp[2]) ? node250 : node245;
															assign node245 = (inp[5]) ? 4'b0101 : node246;
																assign node246 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node250 = (inp[5]) ? 4'b0000 : node251;
																assign node251 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node255 = (inp[2]) ? node273 : node256;
											assign node256 = (inp[5]) ? node266 : node257;
												assign node257 = (inp[1]) ? 4'b0100 : node258;
													assign node258 = (inp[10]) ? 4'b0101 : node259;
														assign node259 = (inp[0]) ? node261 : 4'b0100;
															assign node261 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node266 = (inp[11]) ? 4'b0000 : node267;
													assign node267 = (inp[9]) ? 4'b0001 : node268;
														assign node268 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node273 = (inp[5]) ? node293 : node274;
												assign node274 = (inp[1]) ? node288 : node275;
													assign node275 = (inp[11]) ? node281 : node276;
														assign node276 = (inp[9]) ? node278 : 4'b0001;
															assign node278 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node281 = (inp[0]) ? node285 : node282;
															assign node282 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node285 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node288 = (inp[11]) ? 4'b0000 : node289;
														assign node289 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node293 = (inp[1]) ? 4'b0101 : node294;
													assign node294 = (inp[10]) ? node296 : 4'b0001;
														assign node296 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node300 = (inp[9]) ? node340 : node301;
										assign node301 = (inp[13]) ? node319 : node302;
											assign node302 = (inp[5]) ? node308 : node303;
												assign node303 = (inp[2]) ? node305 : 4'b0010;
													assign node305 = (inp[0]) ? 4'b0010 : 4'b0110;
												assign node308 = (inp[2]) ? node316 : node309;
													assign node309 = (inp[11]) ? 4'b0110 : node310;
														assign node310 = (inp[1]) ? 4'b0110 : node311;
															assign node311 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node316 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node319 = (inp[2]) ? node333 : node320;
												assign node320 = (inp[11]) ? node326 : node321;
													assign node321 = (inp[10]) ? node323 : 4'b0010;
														assign node323 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node326 = (inp[1]) ? 4'b0011 : node327;
														assign node327 = (inp[5]) ? node329 : 4'b0110;
															assign node329 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node333 = (inp[10]) ? node335 : 4'b0111;
													assign node335 = (inp[1]) ? node337 : 4'b0010;
														assign node337 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node340 = (inp[5]) ? node358 : node341;
											assign node341 = (inp[2]) ? node353 : node342;
												assign node342 = (inp[11]) ? node350 : node343;
													assign node343 = (inp[0]) ? node347 : node344;
														assign node344 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node347 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node350 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node353 = (inp[0]) ? 4'b0011 : node354;
													assign node354 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node358 = (inp[1]) ? node372 : node359;
												assign node359 = (inp[11]) ? node367 : node360;
													assign node360 = (inp[0]) ? node364 : node361;
														assign node361 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node364 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node367 = (inp[2]) ? 4'b0111 : node368;
														assign node368 = (inp[10]) ? 4'b0111 : 4'b0010;
												assign node372 = (inp[10]) ? node376 : node373;
													assign node373 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node376 = (inp[11]) ? 4'b0110 : 4'b0111;
							assign node379 = (inp[4]) ? node559 : node380;
								assign node380 = (inp[0]) ? node482 : node381;
									assign node381 = (inp[1]) ? node431 : node382;
										assign node382 = (inp[10]) ? node406 : node383;
											assign node383 = (inp[11]) ? node391 : node384;
												assign node384 = (inp[15]) ? 4'b0110 : node385;
													assign node385 = (inp[2]) ? 4'b0010 : node386;
														assign node386 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node391 = (inp[5]) ? node399 : node392;
													assign node392 = (inp[9]) ? 4'b0010 : node393;
														assign node393 = (inp[13]) ? node395 : 4'b0110;
															assign node395 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node399 = (inp[13]) ? node401 : 4'b0011;
														assign node401 = (inp[2]) ? 4'b0010 : node402;
															assign node402 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node406 = (inp[9]) ? node424 : node407;
												assign node407 = (inp[5]) ? node415 : node408;
													assign node408 = (inp[2]) ? node410 : 4'b0011;
														assign node410 = (inp[15]) ? 4'b0011 : node411;
															assign node411 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node415 = (inp[13]) ? node419 : node416;
														assign node416 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node419 = (inp[15]) ? node421 : 4'b0010;
															assign node421 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node424 = (inp[5]) ? node428 : node425;
													assign node425 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node428 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node431 = (inp[10]) ? node449 : node432;
											assign node432 = (inp[9]) ? node440 : node433;
												assign node433 = (inp[13]) ? node437 : node434;
													assign node434 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node437 = (inp[11]) ? 4'b0111 : 4'b0011;
												assign node440 = (inp[13]) ? node444 : node441;
													assign node441 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node444 = (inp[11]) ? 4'b0110 : node445;
														assign node445 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node449 = (inp[15]) ? node467 : node450;
												assign node450 = (inp[11]) ? node460 : node451;
													assign node451 = (inp[5]) ? node457 : node452;
														assign node452 = (inp[2]) ? node454 : 4'b0111;
															assign node454 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node457 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node460 = (inp[2]) ? node462 : 4'b0011;
														assign node462 = (inp[13]) ? node464 : 4'b0010;
															assign node464 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node467 = (inp[11]) ? node473 : node468;
													assign node468 = (inp[2]) ? 4'b0010 : node469;
														assign node469 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node473 = (inp[5]) ? node475 : 4'b0110;
														assign node475 = (inp[9]) ? 4'b0110 : node476;
															assign node476 = (inp[13]) ? 4'b0110 : node477;
																assign node477 = (inp[2]) ? 4'b0111 : 4'b0011;
									assign node482 = (inp[9]) ? node516 : node483;
										assign node483 = (inp[5]) ? node497 : node484;
											assign node484 = (inp[1]) ? 4'b0011 : node485;
												assign node485 = (inp[15]) ? node489 : node486;
													assign node486 = (inp[13]) ? 4'b0011 : 4'b0110;
													assign node489 = (inp[2]) ? node493 : node490;
														assign node490 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node493 = (inp[13]) ? 4'b0111 : 4'b0011;
											assign node497 = (inp[1]) ? node509 : node498;
												assign node498 = (inp[15]) ? node500 : 4'b0111;
													assign node500 = (inp[2]) ? node506 : node501;
														assign node501 = (inp[10]) ? 4'b0111 : node502;
															assign node502 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node506 = (inp[13]) ? 4'b0111 : 4'b0010;
												assign node509 = (inp[15]) ? node511 : 4'b0110;
													assign node511 = (inp[11]) ? node513 : 4'b0010;
														assign node513 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node516 = (inp[10]) ? node540 : node517;
											assign node517 = (inp[1]) ? node527 : node518;
												assign node518 = (inp[5]) ? node522 : node519;
													assign node519 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node522 = (inp[15]) ? node524 : 4'b0011;
														assign node524 = (inp[11]) ? 4'b0010 : 4'b0110;
												assign node527 = (inp[13]) ? node533 : node528;
													assign node528 = (inp[2]) ? node530 : 4'b0110;
														assign node530 = (inp[11]) ? 4'b0011 : 4'b0111;
													assign node533 = (inp[15]) ? node535 : 4'b0010;
														assign node535 = (inp[5]) ? node537 : 4'b0011;
															assign node537 = (inp[2]) ? 4'b0011 : 4'b0111;
											assign node540 = (inp[2]) ? node550 : node541;
												assign node541 = (inp[5]) ? node547 : node542;
													assign node542 = (inp[15]) ? 4'b0011 : node543;
														assign node543 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node547 = (inp[11]) ? 4'b0110 : 4'b0011;
												assign node550 = (inp[15]) ? node554 : node551;
													assign node551 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node554 = (inp[1]) ? 4'b0111 : node555;
														assign node555 = (inp[5]) ? 4'b0111 : 4'b0110;
								assign node559 = (inp[15]) ? node657 : node560;
									assign node560 = (inp[9]) ? node616 : node561;
										assign node561 = (inp[11]) ? node579 : node562;
											assign node562 = (inp[0]) ? node568 : node563;
												assign node563 = (inp[10]) ? 4'b0110 : node564;
													assign node564 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node568 = (inp[13]) ? node574 : node569;
													assign node569 = (inp[10]) ? node571 : 4'b0010;
														assign node571 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node574 = (inp[1]) ? node576 : 4'b0011;
														assign node576 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node579 = (inp[0]) ? node595 : node580;
												assign node580 = (inp[10]) ? node590 : node581;
													assign node581 = (inp[2]) ? node583 : 4'b0110;
														assign node583 = (inp[1]) ? node585 : 4'b0111;
															assign node585 = (inp[5]) ? node587 : 4'b0010;
																assign node587 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node590 = (inp[5]) ? node592 : 4'b0011;
														assign node592 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node595 = (inp[1]) ? node611 : node596;
													assign node596 = (inp[13]) ? node604 : node597;
														assign node597 = (inp[2]) ? node599 : 4'b0010;
															assign node599 = (inp[10]) ? 4'b0110 : node600;
																assign node600 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node604 = (inp[2]) ? 4'b0011 : node605;
															assign node605 = (inp[5]) ? node607 : 4'b0111;
																assign node607 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node611 = (inp[10]) ? node613 : 4'b0011;
														assign node613 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node616 = (inp[11]) ? node636 : node617;
											assign node617 = (inp[5]) ? node629 : node618;
												assign node618 = (inp[13]) ? node626 : node619;
													assign node619 = (inp[2]) ? node623 : node620;
														assign node620 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node623 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node626 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node629 = (inp[13]) ? node631 : 4'b0110;
													assign node631 = (inp[2]) ? node633 : 4'b0111;
														assign node633 = (inp[1]) ? 4'b0111 : 4'b0011;
											assign node636 = (inp[2]) ? node648 : node637;
												assign node637 = (inp[5]) ? node639 : 4'b0010;
													assign node639 = (inp[1]) ? node641 : 4'b0011;
														assign node641 = (inp[10]) ? node645 : node642;
															assign node642 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node645 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node648 = (inp[13]) ? node650 : 4'b0110;
													assign node650 = (inp[0]) ? node654 : node651;
														assign node651 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node654 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node657 = (inp[13]) ? node707 : node658;
										assign node658 = (inp[2]) ? node672 : node659;
											assign node659 = (inp[5]) ? node669 : node660;
												assign node660 = (inp[0]) ? 4'b0001 : node661;
													assign node661 = (inp[9]) ? 4'b0000 : node662;
														assign node662 = (inp[10]) ? node664 : 4'b0000;
															assign node664 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node669 = (inp[1]) ? 4'b0100 : 4'b0000;
											assign node672 = (inp[1]) ? node688 : node673;
												assign node673 = (inp[5]) ? node675 : 4'b0101;
													assign node675 = (inp[9]) ? node681 : node676;
														assign node676 = (inp[0]) ? 4'b0100 : node677;
															assign node677 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node681 = (inp[10]) ? node685 : node682;
															assign node682 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node685 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node688 = (inp[5]) ? node698 : node689;
													assign node689 = (inp[11]) ? node691 : 4'b0100;
														assign node691 = (inp[10]) ? node693 : 4'b0101;
															assign node693 = (inp[0]) ? 4'b0100 : node694;
																assign node694 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node698 = (inp[10]) ? node700 : 4'b0000;
														assign node700 = (inp[11]) ? node702 : 4'b0000;
															assign node702 = (inp[9]) ? node704 : 4'b0001;
																assign node704 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node707 = (inp[2]) ? node729 : node708;
											assign node708 = (inp[5]) ? node718 : node709;
												assign node709 = (inp[0]) ? node715 : node710;
													assign node710 = (inp[10]) ? node712 : 4'b0100;
														assign node712 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node715 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node718 = (inp[1]) ? node722 : node719;
													assign node719 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node722 = (inp[10]) ? node724 : 4'b0000;
														assign node724 = (inp[9]) ? node726 : 4'b0001;
															assign node726 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node729 = (inp[1]) ? node743 : node730;
												assign node730 = (inp[11]) ? node738 : node731;
													assign node731 = (inp[10]) ? node735 : node732;
														assign node732 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node735 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node738 = (inp[0]) ? node740 : 4'b0000;
														assign node740 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node743 = (inp[5]) ? node747 : node744;
													assign node744 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node747 = (inp[0]) ? 4'b0101 : node748;
														assign node748 = (inp[11]) ? node750 : 4'b0100;
															assign node750 = (inp[9]) ? 4'b0101 : 4'b0100;
						assign node754 = (inp[7]) ? node1140 : node755;
							assign node755 = (inp[15]) ? node977 : node756;
								assign node756 = (inp[11]) ? node852 : node757;
									assign node757 = (inp[9]) ? node809 : node758;
										assign node758 = (inp[10]) ? node784 : node759;
											assign node759 = (inp[4]) ? node773 : node760;
												assign node760 = (inp[1]) ? node762 : 4'b0010;
													assign node762 = (inp[0]) ? node770 : node763;
														assign node763 = (inp[2]) ? node765 : 4'b0011;
															assign node765 = (inp[5]) ? 4'b0111 : node766;
																assign node766 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node770 = (inp[2]) ? 4'b0010 : 4'b0111;
												assign node773 = (inp[13]) ? node775 : 4'b0010;
													assign node775 = (inp[1]) ? node777 : 4'b0110;
														assign node777 = (inp[2]) ? node781 : node778;
															assign node778 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node781 = (inp[5]) ? 4'b0010 : 4'b0111;
											assign node784 = (inp[2]) ? node794 : node785;
												assign node785 = (inp[4]) ? node789 : node786;
													assign node786 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node789 = (inp[13]) ? node791 : 4'b0111;
														assign node791 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node794 = (inp[4]) ? node804 : node795;
													assign node795 = (inp[13]) ? node799 : node796;
														assign node796 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node799 = (inp[0]) ? node801 : 4'b0010;
															assign node801 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node804 = (inp[13]) ? node806 : 4'b0011;
														assign node806 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node809 = (inp[10]) ? node817 : node810;
											assign node810 = (inp[1]) ? node812 : 4'b0111;
												assign node812 = (inp[0]) ? node814 : 4'b0110;
													assign node814 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node817 = (inp[4]) ? node839 : node818;
												assign node818 = (inp[1]) ? node830 : node819;
													assign node819 = (inp[0]) ? node821 : 4'b0110;
														assign node821 = (inp[5]) ? node825 : node822;
															assign node822 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node825 = (inp[13]) ? 4'b0110 : node826;
																assign node826 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node830 = (inp[13]) ? node832 : 4'b0111;
														assign node832 = (inp[0]) ? 4'b0010 : node833;
															assign node833 = (inp[5]) ? node835 : 4'b0011;
																assign node835 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node839 = (inp[2]) ? node849 : node840;
													assign node840 = (inp[1]) ? node844 : node841;
														assign node841 = (inp[5]) ? 4'b0011 : 4'b0110;
														assign node844 = (inp[13]) ? node846 : 4'b0010;
															assign node846 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node849 = (inp[13]) ? 4'b0011 : 4'b0010;
									assign node852 = (inp[0]) ? node910 : node853;
										assign node853 = (inp[9]) ? node887 : node854;
											assign node854 = (inp[10]) ? node876 : node855;
												assign node855 = (inp[5]) ? node871 : node856;
													assign node856 = (inp[13]) ? node864 : node857;
														assign node857 = (inp[1]) ? 4'b0111 : node858;
															assign node858 = (inp[4]) ? 4'b0010 : node859;
																assign node859 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node864 = (inp[4]) ? node868 : node865;
															assign node865 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node868 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node871 = (inp[13]) ? node873 : 4'b0010;
														assign node873 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node876 = (inp[5]) ? node880 : node877;
													assign node877 = (inp[1]) ? 4'b0110 : 4'b0011;
													assign node880 = (inp[1]) ? 4'b0011 : node881;
														assign node881 = (inp[13]) ? node883 : 4'b0111;
															assign node883 = (inp[2]) ? 4'b0010 : 4'b0111;
											assign node887 = (inp[10]) ? node893 : node888;
												assign node888 = (inp[5]) ? 4'b0011 : node889;
													assign node889 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node893 = (inp[5]) ? node901 : node894;
													assign node894 = (inp[1]) ? node896 : 4'b0110;
														assign node896 = (inp[2]) ? 4'b0111 : node897;
															assign node897 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node901 = (inp[4]) ? node905 : node902;
														assign node902 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node905 = (inp[1]) ? 4'b0010 : node906;
															assign node906 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node910 = (inp[2]) ? node948 : node911;
											assign node911 = (inp[10]) ? node933 : node912;
												assign node912 = (inp[13]) ? node922 : node913;
													assign node913 = (inp[4]) ? node919 : node914;
														assign node914 = (inp[5]) ? node916 : 4'b0011;
															assign node916 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node919 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node922 = (inp[1]) ? node924 : 4'b0010;
														assign node924 = (inp[4]) ? node928 : node925;
															assign node925 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node928 = (inp[5]) ? node930 : 4'b0011;
																assign node930 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node933 = (inp[1]) ? node939 : node934;
													assign node934 = (inp[9]) ? 4'b0111 : node935;
														assign node935 = (inp[13]) ? 4'b0011 : 4'b0110;
													assign node939 = (inp[5]) ? node941 : 4'b0010;
														assign node941 = (inp[13]) ? node943 : 4'b0111;
															assign node943 = (inp[4]) ? node945 : 4'b0010;
																assign node945 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node948 = (inp[10]) ? node962 : node949;
												assign node949 = (inp[4]) ? node957 : node950;
													assign node950 = (inp[1]) ? node952 : 4'b0010;
														assign node952 = (inp[13]) ? 4'b0110 : node953;
															assign node953 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node957 = (inp[1]) ? node959 : 4'b0110;
														assign node959 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node962 = (inp[5]) ? node970 : node963;
													assign node963 = (inp[9]) ? 4'b0010 : node964;
														assign node964 = (inp[1]) ? node966 : 4'b0011;
															assign node966 = (inp[4]) ? 4'b0110 : 4'b0011;
													assign node970 = (inp[9]) ? 4'b0010 : node971;
														assign node971 = (inp[13]) ? 4'b0010 : node972;
															assign node972 = (inp[4]) ? 4'b0010 : 4'b0110;
								assign node977 = (inp[4]) ? node1049 : node978;
									assign node978 = (inp[13]) ? node1014 : node979;
										assign node979 = (inp[2]) ? node999 : node980;
											assign node980 = (inp[1]) ? node988 : node981;
												assign node981 = (inp[5]) ? 4'b0011 : node982;
													assign node982 = (inp[11]) ? node984 : 4'b0011;
														assign node984 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node988 = (inp[5]) ? node994 : node989;
													assign node989 = (inp[9]) ? node991 : 4'b0011;
														assign node991 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node994 = (inp[0]) ? node996 : 4'b0110;
														assign node996 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node999 = (inp[5]) ? node1007 : node1000;
												assign node1000 = (inp[1]) ? 4'b0111 : node1001;
													assign node1001 = (inp[10]) ? node1003 : 4'b0111;
														assign node1003 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node1007 = (inp[1]) ? node1011 : node1008;
													assign node1008 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node1011 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node1014 = (inp[2]) ? node1034 : node1015;
											assign node1015 = (inp[5]) ? node1025 : node1016;
												assign node1016 = (inp[11]) ? node1018 : 4'b0110;
													assign node1018 = (inp[1]) ? node1020 : 4'b0110;
														assign node1020 = (inp[9]) ? 4'b0111 : node1021;
															assign node1021 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node1025 = (inp[1]) ? node1027 : 4'b0111;
													assign node1027 = (inp[10]) ? node1029 : 4'b0010;
														assign node1029 = (inp[11]) ? 4'b0010 : node1030;
															assign node1030 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node1034 = (inp[11]) ? node1046 : node1035;
												assign node1035 = (inp[0]) ? 4'b0110 : node1036;
													assign node1036 = (inp[10]) ? node1040 : node1037;
														assign node1037 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node1040 = (inp[5]) ? node1042 : 4'b0011;
															assign node1042 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node1046 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node1049 = (inp[13]) ? node1107 : node1050;
										assign node1050 = (inp[2]) ? node1086 : node1051;
											assign node1051 = (inp[1]) ? node1069 : node1052;
												assign node1052 = (inp[5]) ? node1058 : node1053;
													assign node1053 = (inp[9]) ? 4'b0000 : node1054;
														assign node1054 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node1058 = (inp[0]) ? node1062 : node1059;
														assign node1059 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1062 = (inp[9]) ? node1064 : 4'b0001;
															assign node1064 = (inp[10]) ? 4'b0001 : node1065;
																assign node1065 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node1069 = (inp[5]) ? node1079 : node1070;
													assign node1070 = (inp[10]) ? node1072 : 4'b0001;
														assign node1072 = (inp[9]) ? 4'b0000 : node1073;
															assign node1073 = (inp[11]) ? node1075 : 4'b0001;
																assign node1075 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node1079 = (inp[0]) ? node1081 : 4'b0101;
														assign node1081 = (inp[10]) ? node1083 : 4'b0100;
															assign node1083 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node1086 = (inp[1]) ? node1094 : node1087;
												assign node1087 = (inp[9]) ? 4'b0101 : node1088;
													assign node1088 = (inp[5]) ? 4'b0100 : node1089;
														assign node1089 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node1094 = (inp[5]) ? node1098 : node1095;
													assign node1095 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1098 = (inp[10]) ? node1102 : node1099;
														assign node1099 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1102 = (inp[0]) ? 4'b0000 : node1103;
															assign node1103 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node1107 = (inp[2]) ? node1129 : node1108;
											assign node1108 = (inp[1]) ? node1122 : node1109;
												assign node1109 = (inp[11]) ? node1117 : node1110;
													assign node1110 = (inp[9]) ? node1112 : 4'b0101;
														assign node1112 = (inp[0]) ? 4'b0101 : node1113;
															assign node1113 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node1117 = (inp[0]) ? 4'b0100 : node1118;
														assign node1118 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node1122 = (inp[5]) ? node1126 : node1123;
													assign node1123 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node1126 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1129 = (inp[1]) ? node1137 : node1130;
												assign node1130 = (inp[11]) ? 4'b0000 : node1131;
													assign node1131 = (inp[0]) ? 4'b0001 : node1132;
														assign node1132 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node1137 = (inp[10]) ? 4'b0100 : 4'b0101;
							assign node1140 = (inp[4]) ? node1340 : node1141;
								assign node1141 = (inp[9]) ? node1219 : node1142;
									assign node1142 = (inp[10]) ? node1182 : node1143;
										assign node1143 = (inp[13]) ? node1165 : node1144;
											assign node1144 = (inp[5]) ? node1150 : node1145;
												assign node1145 = (inp[11]) ? node1147 : 4'b0000;
													assign node1147 = (inp[15]) ? 4'b0001 : 4'b0100;
												assign node1150 = (inp[15]) ? node1162 : node1151;
													assign node1151 = (inp[2]) ? 4'b0000 : node1152;
														assign node1152 = (inp[11]) ? 4'b0100 : node1153;
															assign node1153 = (inp[0]) ? node1157 : node1154;
																assign node1154 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node1157 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node1162 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node1165 = (inp[5]) ? node1179 : node1166;
												assign node1166 = (inp[15]) ? node1172 : node1167;
													assign node1167 = (inp[1]) ? node1169 : 4'b0001;
														assign node1169 = (inp[11]) ? 4'b0001 : 4'b0100;
													assign node1172 = (inp[11]) ? node1176 : node1173;
														assign node1173 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node1176 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node1179 = (inp[15]) ? 4'b0001 : 4'b0000;
										assign node1182 = (inp[11]) ? node1202 : node1183;
											assign node1183 = (inp[2]) ? node1195 : node1184;
												assign node1184 = (inp[5]) ? 4'b0100 : node1185;
													assign node1185 = (inp[13]) ? node1191 : node1186;
														assign node1186 = (inp[15]) ? node1188 : 4'b0101;
															assign node1188 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node1191 = (inp[1]) ? 4'b0100 : 4'b0001;
												assign node1195 = (inp[13]) ? node1199 : node1196;
													assign node1196 = (inp[15]) ? 4'b0101 : 4'b0001;
													assign node1199 = (inp[15]) ? 4'b0001 : 4'b0101;
											assign node1202 = (inp[5]) ? node1212 : node1203;
												assign node1203 = (inp[15]) ? node1205 : 4'b0001;
													assign node1205 = (inp[1]) ? node1207 : 4'b0100;
														assign node1207 = (inp[2]) ? node1209 : 4'b0000;
															assign node1209 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node1212 = (inp[1]) ? node1214 : 4'b0001;
													assign node1214 = (inp[15]) ? 4'b0101 : node1215;
														assign node1215 = (inp[13]) ? 4'b0100 : 4'b0000;
									assign node1219 = (inp[13]) ? node1277 : node1220;
										assign node1220 = (inp[1]) ? node1256 : node1221;
											assign node1221 = (inp[11]) ? node1233 : node1222;
												assign node1222 = (inp[15]) ? node1228 : node1223;
													assign node1223 = (inp[10]) ? 4'b0000 : node1224;
														assign node1224 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node1228 = (inp[0]) ? 4'b0100 : node1229;
														assign node1229 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node1233 = (inp[5]) ? node1251 : node1234;
													assign node1234 = (inp[0]) ? node1240 : node1235;
														assign node1235 = (inp[2]) ? 4'b0001 : node1236;
															assign node1236 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node1240 = (inp[15]) ? node1246 : node1241;
															assign node1241 = (inp[10]) ? 4'b0101 : node1242;
																assign node1242 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node1246 = (inp[2]) ? node1248 : 4'b0101;
																assign node1248 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1251 = (inp[10]) ? node1253 : 4'b0101;
														assign node1253 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node1256 = (inp[0]) ? node1266 : node1257;
												assign node1257 = (inp[15]) ? 4'b0001 : node1258;
													assign node1258 = (inp[2]) ? node1260 : 4'b0100;
														assign node1260 = (inp[5]) ? node1262 : 4'b0001;
															assign node1262 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node1266 = (inp[11]) ? 4'b0001 : node1267;
													assign node1267 = (inp[15]) ? node1271 : node1268;
														assign node1268 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node1271 = (inp[2]) ? 4'b0100 : node1272;
															assign node1272 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node1277 = (inp[0]) ? node1309 : node1278;
											assign node1278 = (inp[10]) ? node1298 : node1279;
												assign node1279 = (inp[15]) ? node1285 : node1280;
													assign node1280 = (inp[2]) ? node1282 : 4'b0100;
														assign node1282 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node1285 = (inp[2]) ? node1293 : node1286;
														assign node1286 = (inp[1]) ? node1288 : 4'b0001;
															assign node1288 = (inp[11]) ? node1290 : 4'b0101;
																assign node1290 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node1293 = (inp[5]) ? 4'b0001 : node1294;
															assign node1294 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node1298 = (inp[15]) ? node1302 : node1299;
													assign node1299 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node1302 = (inp[2]) ? node1304 : 4'b0101;
														assign node1304 = (inp[11]) ? 4'b0000 : node1305;
															assign node1305 = (inp[5]) ? 4'b0001 : 4'b0100;
											assign node1309 = (inp[11]) ? node1323 : node1310;
												assign node1310 = (inp[2]) ? node1318 : node1311;
													assign node1311 = (inp[5]) ? 4'b0101 : node1312;
														assign node1312 = (inp[15]) ? node1314 : 4'b0100;
															assign node1314 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1318 = (inp[15]) ? node1320 : 4'b0101;
														assign node1320 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node1323 = (inp[10]) ? node1333 : node1324;
													assign node1324 = (inp[5]) ? 4'b0001 : node1325;
														assign node1325 = (inp[1]) ? node1327 : 4'b0001;
															assign node1327 = (inp[15]) ? node1329 : 4'b0000;
																assign node1329 = (inp[2]) ? 4'b0000 : 4'b0101;
													assign node1333 = (inp[1]) ? 4'b0001 : node1334;
														assign node1334 = (inp[15]) ? node1336 : 4'b0101;
															assign node1336 = (inp[2]) ? 4'b0101 : 4'b0001;
								assign node1340 = (inp[15]) ? node1428 : node1341;
									assign node1341 = (inp[5]) ? node1385 : node1342;
										assign node1342 = (inp[13]) ? node1362 : node1343;
											assign node1343 = (inp[11]) ? node1355 : node1344;
												assign node1344 = (inp[2]) ? node1348 : node1345;
													assign node1345 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node1348 = (inp[1]) ? node1352 : node1349;
														assign node1349 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node1352 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node1355 = (inp[9]) ? 4'b0100 : node1356;
													assign node1356 = (inp[10]) ? node1358 : 4'b0001;
														assign node1358 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node1362 = (inp[2]) ? node1372 : node1363;
												assign node1363 = (inp[1]) ? 4'b0100 : node1364;
													assign node1364 = (inp[9]) ? node1366 : 4'b0000;
														assign node1366 = (inp[0]) ? 4'b0001 : node1367;
															assign node1367 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node1372 = (inp[1]) ? node1378 : node1373;
													assign node1373 = (inp[11]) ? 4'b0100 : node1374;
														assign node1374 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node1378 = (inp[10]) ? node1380 : 4'b0001;
														assign node1380 = (inp[11]) ? node1382 : 4'b0000;
															assign node1382 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node1385 = (inp[1]) ? node1405 : node1386;
											assign node1386 = (inp[2]) ? node1398 : node1387;
												assign node1387 = (inp[13]) ? node1391 : node1388;
													assign node1388 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node1391 = (inp[11]) ? node1393 : 4'b0100;
														assign node1393 = (inp[10]) ? node1395 : 4'b0101;
															assign node1395 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node1398 = (inp[13]) ? node1402 : node1399;
													assign node1399 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1402 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1405 = (inp[11]) ? node1419 : node1406;
												assign node1406 = (inp[10]) ? node1410 : node1407;
													assign node1407 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node1410 = (inp[9]) ? 4'b0001 : node1411;
														assign node1411 = (inp[2]) ? 4'b0000 : node1412;
															assign node1412 = (inp[13]) ? 4'b0101 : node1413;
																assign node1413 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node1419 = (inp[0]) ? node1421 : 4'b0101;
													assign node1421 = (inp[9]) ? node1423 : 4'b0100;
														assign node1423 = (inp[2]) ? 4'b0001 : node1424;
															assign node1424 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node1428 = (inp[11]) ? node1494 : node1429;
										assign node1429 = (inp[5]) ? node1449 : node1430;
											assign node1430 = (inp[9]) ? node1442 : node1431;
												assign node1431 = (inp[13]) ? node1435 : node1432;
													assign node1432 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node1435 = (inp[1]) ? 4'b0010 : node1436;
														assign node1436 = (inp[10]) ? node1438 : 4'b0011;
															assign node1438 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node1442 = (inp[0]) ? node1444 : 4'b0110;
													assign node1444 = (inp[13]) ? node1446 : 4'b0110;
														assign node1446 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node1449 = (inp[1]) ? node1467 : node1450;
												assign node1450 = (inp[10]) ? 4'b0011 : node1451;
													assign node1451 = (inp[9]) ? node1457 : node1452;
														assign node1452 = (inp[13]) ? node1454 : 4'b0010;
															assign node1454 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node1457 = (inp[13]) ? node1463 : node1458;
															assign node1458 = (inp[0]) ? 4'b0110 : node1459;
																assign node1459 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node1463 = (inp[2]) ? 4'b0110 : 4'b0011;
												assign node1467 = (inp[10]) ? node1483 : node1468;
													assign node1468 = (inp[13]) ? node1476 : node1469;
														assign node1469 = (inp[2]) ? 4'b0110 : node1470;
															assign node1470 = (inp[0]) ? 4'b0011 : node1471;
																assign node1471 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node1476 = (inp[2]) ? 4'b0011 : node1477;
															assign node1477 = (inp[9]) ? node1479 : 4'b0111;
																assign node1479 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node1483 = (inp[9]) ? node1491 : node1484;
														assign node1484 = (inp[13]) ? node1488 : node1485;
															assign node1485 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1488 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node1491 = (inp[13]) ? 4'b0111 : 4'b0010;
										assign node1494 = (inp[9]) ? node1526 : node1495;
											assign node1495 = (inp[2]) ? node1513 : node1496;
												assign node1496 = (inp[10]) ? node1506 : node1497;
													assign node1497 = (inp[13]) ? node1501 : node1498;
														assign node1498 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node1501 = (inp[1]) ? node1503 : 4'b0011;
															assign node1503 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node1506 = (inp[13]) ? 4'b0111 : node1507;
														assign node1507 = (inp[0]) ? node1509 : 4'b0110;
															assign node1509 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node1513 = (inp[13]) ? node1515 : 4'b0011;
													assign node1515 = (inp[10]) ? node1523 : node1516;
														assign node1516 = (inp[0]) ? 4'b0110 : node1517;
															assign node1517 = (inp[1]) ? 4'b0111 : node1518;
																assign node1518 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1523 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node1526 = (inp[5]) ? node1538 : node1527;
												assign node1527 = (inp[0]) ? node1535 : node1528;
													assign node1528 = (inp[1]) ? node1532 : node1529;
														assign node1529 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node1532 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1535 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node1538 = (inp[1]) ? 4'b0110 : node1539;
													assign node1539 = (inp[2]) ? node1543 : node1540;
														assign node1540 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node1543 = (inp[10]) ? 4'b0010 : 4'b0111;
					assign node1547 = (inp[12]) ? node2237 : node1548;
						assign node1548 = (inp[4]) ? node1842 : node1549;
							assign node1549 = (inp[1]) ? node1723 : node1550;
								assign node1550 = (inp[2]) ? node1630 : node1551;
									assign node1551 = (inp[7]) ? node1593 : node1552;
										assign node1552 = (inp[15]) ? node1570 : node1553;
											assign node1553 = (inp[0]) ? node1563 : node1554;
												assign node1554 = (inp[10]) ? node1560 : node1555;
													assign node1555 = (inp[13]) ? node1557 : 4'b1000;
														assign node1557 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node1560 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node1563 = (inp[10]) ? node1565 : 4'b1001;
													assign node1565 = (inp[13]) ? node1567 : 4'b1000;
														assign node1567 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node1570 = (inp[11]) ? node1578 : node1571;
												assign node1571 = (inp[13]) ? 4'b1001 : node1572;
													assign node1572 = (inp[0]) ? node1574 : 4'b1001;
														assign node1574 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node1578 = (inp[5]) ? node1588 : node1579;
													assign node1579 = (inp[13]) ? node1585 : node1580;
														assign node1580 = (inp[9]) ? 4'b1001 : node1581;
															assign node1581 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node1585 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node1588 = (inp[10]) ? 4'b1000 : node1589;
														assign node1589 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node1593 = (inp[13]) ? node1607 : node1594;
											assign node1594 = (inp[5]) ? node1602 : node1595;
												assign node1595 = (inp[9]) ? node1597 : 4'b1001;
													assign node1597 = (inp[10]) ? node1599 : 4'b1000;
														assign node1599 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node1602 = (inp[9]) ? 4'b1001 : node1603;
													assign node1603 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node1607 = (inp[0]) ? node1621 : node1608;
												assign node1608 = (inp[15]) ? node1616 : node1609;
													assign node1609 = (inp[5]) ? node1613 : node1610;
														assign node1610 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node1613 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node1616 = (inp[5]) ? node1618 : 4'b1100;
														assign node1618 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node1621 = (inp[9]) ? node1623 : 4'b1100;
													assign node1623 = (inp[11]) ? node1627 : node1624;
														assign node1624 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node1627 = (inp[10]) ? 4'b1100 : 4'b1000;
									assign node1630 = (inp[7]) ? node1656 : node1631;
										assign node1631 = (inp[11]) ? node1641 : node1632;
											assign node1632 = (inp[5]) ? 4'b1101 : node1633;
												assign node1633 = (inp[13]) ? node1635 : 4'b1101;
													assign node1635 = (inp[10]) ? node1637 : 4'b1100;
														assign node1637 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node1641 = (inp[15]) ? node1651 : node1642;
												assign node1642 = (inp[5]) ? node1646 : node1643;
													assign node1643 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node1646 = (inp[13]) ? node1648 : 4'b1100;
														assign node1648 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node1651 = (inp[10]) ? node1653 : 4'b1101;
													assign node1653 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node1656 = (inp[11]) ? node1688 : node1657;
											assign node1657 = (inp[9]) ? node1671 : node1658;
												assign node1658 = (inp[10]) ? node1666 : node1659;
													assign node1659 = (inp[0]) ? 4'b1100 : node1660;
														assign node1660 = (inp[5]) ? node1662 : 4'b1000;
															assign node1662 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node1666 = (inp[5]) ? 4'b1100 : node1667;
														assign node1667 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node1671 = (inp[5]) ? node1679 : node1672;
													assign node1672 = (inp[15]) ? node1674 : 4'b1101;
														assign node1674 = (inp[13]) ? node1676 : 4'b1001;
															assign node1676 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node1679 = (inp[13]) ? node1683 : node1680;
														assign node1680 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node1683 = (inp[0]) ? node1685 : 4'b1101;
															assign node1685 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node1688 = (inp[13]) ? node1706 : node1689;
												assign node1689 = (inp[0]) ? node1697 : node1690;
													assign node1690 = (inp[10]) ? node1692 : 4'b1001;
														assign node1692 = (inp[5]) ? node1694 : 4'b1101;
															assign node1694 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node1697 = (inp[10]) ? node1703 : node1698;
														assign node1698 = (inp[15]) ? 4'b1000 : node1699;
															assign node1699 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node1703 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node1706 = (inp[10]) ? node1716 : node1707;
													assign node1707 = (inp[0]) ? node1709 : 4'b1000;
														assign node1709 = (inp[5]) ? node1713 : node1710;
															assign node1710 = (inp[9]) ? 4'b1001 : 4'b1100;
															assign node1713 = (inp[9]) ? 4'b1100 : 4'b1001;
													assign node1716 = (inp[0]) ? 4'b1000 : node1717;
														assign node1717 = (inp[15]) ? node1719 : 4'b1001;
															assign node1719 = (inp[5]) ? 4'b1100 : 4'b1001;
								assign node1723 = (inp[2]) ? node1771 : node1724;
									assign node1724 = (inp[7]) ? node1742 : node1725;
										assign node1725 = (inp[0]) ? 4'b1101 : node1726;
											assign node1726 = (inp[10]) ? node1734 : node1727;
												assign node1727 = (inp[11]) ? node1729 : 4'b1100;
													assign node1729 = (inp[5]) ? 4'b1101 : node1730;
														assign node1730 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node1734 = (inp[13]) ? 4'b1101 : node1735;
													assign node1735 = (inp[11]) ? node1737 : 4'b1101;
														assign node1737 = (inp[15]) ? 4'b1100 : 4'b1101;
										assign node1742 = (inp[0]) ? node1754 : node1743;
											assign node1743 = (inp[10]) ? node1749 : node1744;
												assign node1744 = (inp[13]) ? node1746 : 4'b1001;
													assign node1746 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node1749 = (inp[15]) ? 4'b1101 : node1750;
													assign node1750 = (inp[5]) ? 4'b1001 : 4'b1101;
											assign node1754 = (inp[5]) ? node1764 : node1755;
												assign node1755 = (inp[15]) ? node1759 : node1756;
													assign node1756 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node1759 = (inp[11]) ? 4'b1001 : node1760;
														assign node1760 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node1764 = (inp[15]) ? 4'b1100 : node1765;
													assign node1765 = (inp[9]) ? 4'b1000 : node1766;
														assign node1766 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node1771 = (inp[7]) ? node1801 : node1772;
										assign node1772 = (inp[15]) ? node1786 : node1773;
											assign node1773 = (inp[13]) ? node1779 : node1774;
												assign node1774 = (inp[0]) ? node1776 : 4'b1001;
													assign node1776 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node1779 = (inp[10]) ? node1783 : node1780;
													assign node1780 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node1783 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node1786 = (inp[5]) ? node1788 : 4'b1001;
												assign node1788 = (inp[13]) ? 4'b1001 : node1789;
													assign node1789 = (inp[11]) ? node1795 : node1790;
														assign node1790 = (inp[0]) ? node1792 : 4'b1001;
															assign node1792 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node1795 = (inp[10]) ? node1797 : 4'b1001;
															assign node1797 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node1801 = (inp[13]) ? node1827 : node1802;
											assign node1802 = (inp[11]) ? node1818 : node1803;
												assign node1803 = (inp[10]) ? node1807 : node1804;
													assign node1804 = (inp[0]) ? 4'b1001 : 4'b1101;
													assign node1807 = (inp[15]) ? node1813 : node1808;
														assign node1808 = (inp[5]) ? 4'b1101 : node1809;
															assign node1809 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node1813 = (inp[5]) ? 4'b1000 : node1814;
															assign node1814 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node1818 = (inp[0]) ? node1822 : node1819;
													assign node1819 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node1822 = (inp[5]) ? 4'b1001 : node1823;
														assign node1823 = (inp[15]) ? 4'b1101 : 4'b1001;
											assign node1827 = (inp[5]) ? node1837 : node1828;
												assign node1828 = (inp[15]) ? node1834 : node1829;
													assign node1829 = (inp[11]) ? 4'b1001 : node1830;
														assign node1830 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node1834 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node1837 = (inp[15]) ? node1839 : 4'b1100;
													assign node1839 = (inp[0]) ? 4'b1000 : 4'b1001;
							assign node1842 = (inp[15]) ? node2058 : node1843;
								assign node1843 = (inp[13]) ? node1963 : node1844;
									assign node1844 = (inp[9]) ? node1916 : node1845;
										assign node1845 = (inp[0]) ? node1879 : node1846;
											assign node1846 = (inp[10]) ? node1870 : node1847;
												assign node1847 = (inp[2]) ? node1859 : node1848;
													assign node1848 = (inp[1]) ? node1854 : node1849;
														assign node1849 = (inp[5]) ? node1851 : 4'b1010;
															assign node1851 = (inp[7]) ? 4'b1110 : 4'b1011;
														assign node1854 = (inp[7]) ? 4'b1110 : node1855;
															assign node1855 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node1859 = (inp[7]) ? node1861 : 4'b1111;
														assign node1861 = (inp[5]) ? node1867 : node1862;
															assign node1862 = (inp[11]) ? 4'b1010 : node1863;
																assign node1863 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node1867 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node1870 = (inp[5]) ? node1876 : node1871;
													assign node1871 = (inp[7]) ? node1873 : 4'b1011;
														assign node1873 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node1876 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node1879 = (inp[11]) ? node1891 : node1880;
												assign node1880 = (inp[5]) ? node1882 : 4'b1011;
													assign node1882 = (inp[2]) ? node1886 : node1883;
														assign node1883 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node1886 = (inp[7]) ? node1888 : 4'b1111;
															assign node1888 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node1891 = (inp[1]) ? node1903 : node1892;
													assign node1892 = (inp[7]) ? node1896 : node1893;
														assign node1893 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node1896 = (inp[2]) ? node1900 : node1897;
															assign node1897 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node1900 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node1903 = (inp[10]) ? node1909 : node1904;
														assign node1904 = (inp[2]) ? 4'b1110 : node1905;
															assign node1905 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node1909 = (inp[5]) ? node1911 : 4'b1010;
															assign node1911 = (inp[7]) ? node1913 : 4'b1010;
																assign node1913 = (inp[2]) ? 4'b1111 : 4'b1010;
										assign node1916 = (inp[2]) ? node1942 : node1917;
											assign node1917 = (inp[1]) ? node1931 : node1918;
												assign node1918 = (inp[5]) ? node1924 : node1919;
													assign node1919 = (inp[0]) ? node1921 : 4'b1010;
														assign node1921 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node1924 = (inp[7]) ? node1926 : 4'b1010;
														assign node1926 = (inp[10]) ? 4'b1111 : node1927;
															assign node1927 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node1931 = (inp[10]) ? node1937 : node1932;
													assign node1932 = (inp[0]) ? 4'b1111 : node1933;
														assign node1933 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node1937 = (inp[0]) ? 4'b1110 : node1938;
														assign node1938 = (inp[5]) ? 4'b1110 : 4'b1111;
											assign node1942 = (inp[1]) ? node1954 : node1943;
												assign node1943 = (inp[7]) ? node1949 : node1944;
													assign node1944 = (inp[10]) ? node1946 : 4'b1111;
														assign node1946 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node1949 = (inp[5]) ? 4'b1010 : node1950;
														assign node1950 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node1954 = (inp[7]) ? node1960 : node1955;
													assign node1955 = (inp[10]) ? node1957 : 4'b1010;
														assign node1957 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node1960 = (inp[0]) ? 4'b1111 : 4'b1011;
									assign node1963 = (inp[0]) ? node2011 : node1964;
										assign node1964 = (inp[7]) ? node1978 : node1965;
											assign node1965 = (inp[1]) ? node1971 : node1966;
												assign node1966 = (inp[2]) ? node1968 : 4'b1011;
													assign node1968 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node1971 = (inp[2]) ? 4'b1010 : node1972;
													assign node1972 = (inp[5]) ? 4'b1111 : node1973;
														assign node1973 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node1978 = (inp[9]) ? node2000 : node1979;
												assign node1979 = (inp[1]) ? node1987 : node1980;
													assign node1980 = (inp[11]) ? node1982 : 4'b1110;
														assign node1982 = (inp[10]) ? 4'b1010 : node1983;
															assign node1983 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node1987 = (inp[10]) ? node1995 : node1988;
														assign node1988 = (inp[2]) ? node1992 : node1989;
															assign node1989 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node1992 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node1995 = (inp[11]) ? node1997 : 4'b1011;
															assign node1997 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node2000 = (inp[1]) ? node2006 : node2001;
													assign node2001 = (inp[5]) ? 4'b1110 : node2002;
														assign node2002 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node2006 = (inp[2]) ? node2008 : 4'b1010;
														assign node2008 = (inp[11]) ? 4'b1010 : 4'b1111;
										assign node2011 = (inp[1]) ? node2033 : node2012;
											assign node2012 = (inp[7]) ? node2020 : node2013;
												assign node2013 = (inp[10]) ? 4'b1011 : node2014;
													assign node2014 = (inp[5]) ? 4'b1010 : node2015;
														assign node2015 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node2020 = (inp[5]) ? node2030 : node2021;
													assign node2021 = (inp[2]) ? 4'b1110 : node2022;
														assign node2022 = (inp[9]) ? node2026 : node2023;
															assign node2023 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node2026 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node2030 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node2033 = (inp[11]) ? node2045 : node2034;
												assign node2034 = (inp[2]) ? node2040 : node2035;
													assign node2035 = (inp[7]) ? node2037 : 4'b1110;
														assign node2037 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node2040 = (inp[5]) ? node2042 : 4'b1011;
														assign node2042 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node2045 = (inp[9]) ? node2053 : node2046;
													assign node2046 = (inp[2]) ? 4'b1111 : node2047;
														assign node2047 = (inp[5]) ? node2049 : 4'b1111;
															assign node2049 = (inp[7]) ? 4'b1011 : 4'b1111;
													assign node2053 = (inp[2]) ? 4'b1011 : node2054;
														assign node2054 = (inp[7]) ? 4'b1011 : 4'b1111;
								assign node2058 = (inp[5]) ? node2146 : node2059;
									assign node2059 = (inp[10]) ? node2105 : node2060;
										assign node2060 = (inp[0]) ? node2088 : node2061;
											assign node2061 = (inp[11]) ? node2077 : node2062;
												assign node2062 = (inp[7]) ? 4'b1010 : node2063;
													assign node2063 = (inp[13]) ? 4'b1110 : node2064;
														assign node2064 = (inp[9]) ? node2070 : node2065;
															assign node2065 = (inp[1]) ? 4'b1010 : node2066;
																assign node2066 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node2070 = (inp[1]) ? node2072 : 4'b1010;
																assign node2072 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node2077 = (inp[9]) ? node2083 : node2078;
													assign node2078 = (inp[1]) ? node2080 : 4'b1010;
														assign node2080 = (inp[7]) ? 4'b1010 : 4'b1110;
													assign node2083 = (inp[7]) ? node2085 : 4'b1111;
														assign node2085 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node2088 = (inp[2]) ? node2098 : node2089;
												assign node2089 = (inp[1]) ? node2095 : node2090;
													assign node2090 = (inp[13]) ? 4'b1011 : node2091;
														assign node2091 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node2095 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node2098 = (inp[1]) ? node2100 : 4'b1110;
													assign node2100 = (inp[11]) ? node2102 : 4'b1011;
														assign node2102 = (inp[13]) ? 4'b1011 : 4'b1010;
										assign node2105 = (inp[2]) ? node2131 : node2106;
											assign node2106 = (inp[1]) ? node2124 : node2107;
												assign node2107 = (inp[0]) ? node2119 : node2108;
													assign node2108 = (inp[9]) ? 4'b1011 : node2109;
														assign node2109 = (inp[13]) ? node2113 : node2110;
															assign node2110 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node2113 = (inp[7]) ? 4'b1011 : node2114;
																assign node2114 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node2119 = (inp[7]) ? node2121 : 4'b1010;
														assign node2121 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node2124 = (inp[11]) ? 4'b1111 : node2125;
													assign node2125 = (inp[0]) ? 4'b1110 : node2126;
														assign node2126 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node2131 = (inp[1]) ? 4'b1010 : node2132;
												assign node2132 = (inp[0]) ? node2134 : 4'b1110;
													assign node2134 = (inp[9]) ? node2140 : node2135;
														assign node2135 = (inp[7]) ? 4'b1111 : node2136;
															assign node2136 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node2140 = (inp[13]) ? node2142 : 4'b1110;
															assign node2142 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node2146 = (inp[13]) ? node2194 : node2147;
										assign node2147 = (inp[2]) ? node2165 : node2148;
											assign node2148 = (inp[1]) ? node2158 : node2149;
												assign node2149 = (inp[7]) ? node2153 : node2150;
													assign node2150 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node2153 = (inp[10]) ? 4'b1010 : node2154;
														assign node2154 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node2158 = (inp[7]) ? node2162 : node2159;
													assign node2159 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node2162 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node2165 = (inp[9]) ? node2173 : node2166;
												assign node2166 = (inp[7]) ? node2170 : node2167;
													assign node2167 = (inp[11]) ? 4'b1110 : 4'b1010;
													assign node2170 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node2173 = (inp[11]) ? node2187 : node2174;
													assign node2174 = (inp[1]) ? node2180 : node2175;
														assign node2175 = (inp[10]) ? 4'b1110 : node2176;
															assign node2176 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node2180 = (inp[7]) ? node2182 : 4'b1110;
															assign node2182 = (inp[0]) ? node2184 : 4'b1011;
																assign node2184 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node2187 = (inp[1]) ? node2191 : node2188;
														assign node2188 = (inp[7]) ? 4'b1111 : 4'b1011;
														assign node2191 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node2194 = (inp[1]) ? node2212 : node2195;
											assign node2195 = (inp[7]) ? node2203 : node2196;
												assign node2196 = (inp[2]) ? 4'b1011 : node2197;
													assign node2197 = (inp[10]) ? 4'b1110 : node2198;
														assign node2198 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node2203 = (inp[2]) ? 4'b1111 : node2204;
													assign node2204 = (inp[0]) ? 4'b1010 : node2205;
														assign node2205 = (inp[10]) ? node2207 : 4'b1011;
															assign node2207 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node2212 = (inp[10]) ? node2224 : node2213;
												assign node2213 = (inp[0]) ? node2219 : node2214;
													assign node2214 = (inp[11]) ? node2216 : 4'b1011;
														assign node2216 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node2219 = (inp[11]) ? node2221 : 4'b1010;
														assign node2221 = (inp[7]) ? 4'b1011 : 4'b1111;
												assign node2224 = (inp[2]) ? node2228 : node2225;
													assign node2225 = (inp[11]) ? 4'b1010 : 4'b1110;
													assign node2228 = (inp[7]) ? node2230 : 4'b1111;
														assign node2230 = (inp[0]) ? node2234 : node2231;
															assign node2231 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node2234 = (inp[11]) ? 4'b1010 : 4'b1011;
						assign node2237 = (inp[4]) ? node2579 : node2238;
							assign node2238 = (inp[10]) ? node2386 : node2239;
								assign node2239 = (inp[0]) ? node2309 : node2240;
									assign node2240 = (inp[2]) ? node2280 : node2241;
										assign node2241 = (inp[11]) ? node2261 : node2242;
											assign node2242 = (inp[5]) ? node2250 : node2243;
												assign node2243 = (inp[7]) ? node2247 : node2244;
													assign node2244 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node2247 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node2250 = (inp[1]) ? node2256 : node2251;
													assign node2251 = (inp[15]) ? node2253 : 4'b1111;
														assign node2253 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node2256 = (inp[7]) ? node2258 : 4'b1111;
														assign node2258 = (inp[15]) ? 4'b1111 : 4'b1011;
											assign node2261 = (inp[15]) ? node2271 : node2262;
												assign node2262 = (inp[1]) ? node2266 : node2263;
													assign node2263 = (inp[7]) ? 4'b1110 : 4'b1010;
													assign node2266 = (inp[5]) ? node2268 : 4'b1111;
														assign node2268 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node2271 = (inp[9]) ? node2275 : node2272;
													assign node2272 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node2275 = (inp[1]) ? 4'b1110 : node2276;
														assign node2276 = (inp[13]) ? 4'b1110 : 4'b1111;
										assign node2280 = (inp[1]) ? node2296 : node2281;
											assign node2281 = (inp[13]) ? node2291 : node2282;
												assign node2282 = (inp[15]) ? node2286 : node2283;
													assign node2283 = (inp[11]) ? 4'b1010 : 4'b1110;
													assign node2286 = (inp[5]) ? 4'b1110 : node2287;
														assign node2287 = (inp[9]) ? 4'b1110 : 4'b1011;
												assign node2291 = (inp[5]) ? node2293 : 4'b1110;
													assign node2293 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node2296 = (inp[13]) ? node2298 : 4'b1010;
												assign node2298 = (inp[5]) ? node2304 : node2299;
													assign node2299 = (inp[9]) ? node2301 : 4'b1110;
														assign node2301 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node2304 = (inp[11]) ? 4'b1010 : node2305;
														assign node2305 = (inp[15]) ? 4'b1011 : 4'b1010;
									assign node2309 = (inp[1]) ? node2343 : node2310;
										assign node2310 = (inp[2]) ? node2322 : node2311;
											assign node2311 = (inp[7]) ? node2319 : node2312;
												assign node2312 = (inp[13]) ? node2314 : 4'b1011;
													assign node2314 = (inp[11]) ? node2316 : 4'b1011;
														assign node2316 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node2319 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node2322 = (inp[7]) ? node2330 : node2323;
												assign node2323 = (inp[13]) ? node2325 : 4'b1111;
													assign node2325 = (inp[15]) ? node2327 : 4'b1111;
														assign node2327 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node2330 = (inp[9]) ? node2336 : node2331;
													assign node2331 = (inp[13]) ? node2333 : 4'b1111;
														assign node2333 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node2336 = (inp[15]) ? 4'b1010 : node2337;
														assign node2337 = (inp[13]) ? 4'b1110 : node2338;
															assign node2338 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node2343 = (inp[2]) ? node2367 : node2344;
											assign node2344 = (inp[7]) ? node2360 : node2345;
												assign node2345 = (inp[11]) ? node2347 : 4'b1110;
													assign node2347 = (inp[5]) ? node2353 : node2348;
														assign node2348 = (inp[13]) ? node2350 : 4'b1110;
															assign node2350 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node2353 = (inp[9]) ? node2355 : 4'b1111;
															assign node2355 = (inp[13]) ? 4'b1110 : node2356;
																assign node2356 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node2360 = (inp[15]) ? node2362 : 4'b1010;
													assign node2362 = (inp[5]) ? node2364 : 4'b1011;
														assign node2364 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node2367 = (inp[7]) ? node2371 : node2368;
												assign node2368 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node2371 = (inp[15]) ? node2379 : node2372;
													assign node2372 = (inp[5]) ? node2376 : node2373;
														assign node2373 = (inp[13]) ? 4'b1010 : 4'b1011;
														assign node2376 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node2379 = (inp[5]) ? node2383 : node2380;
														assign node2380 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node2383 = (inp[9]) ? 4'b1011 : 4'b1010;
								assign node2386 = (inp[7]) ? node2446 : node2387;
									assign node2387 = (inp[0]) ? node2417 : node2388;
										assign node2388 = (inp[13]) ? node2402 : node2389;
											assign node2389 = (inp[9]) ? node2395 : node2390;
												assign node2390 = (inp[1]) ? node2392 : 4'b1011;
													assign node2392 = (inp[2]) ? 4'b1011 : 4'b1110;
												assign node2395 = (inp[2]) ? node2399 : node2396;
													assign node2396 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node2399 = (inp[1]) ? 4'b1011 : 4'b1111;
											assign node2402 = (inp[11]) ? node2410 : node2403;
												assign node2403 = (inp[9]) ? node2405 : 4'b1110;
													assign node2405 = (inp[5]) ? 4'b1110 : node2406;
														assign node2406 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node2410 = (inp[1]) ? 4'b1011 : node2411;
													assign node2411 = (inp[2]) ? 4'b1111 : node2412;
														assign node2412 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node2417 = (inp[2]) ? node2433 : node2418;
											assign node2418 = (inp[1]) ? node2428 : node2419;
												assign node2419 = (inp[13]) ? node2421 : 4'b1010;
													assign node2421 = (inp[11]) ? node2425 : node2422;
														assign node2422 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node2425 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node2428 = (inp[11]) ? node2430 : 4'b1111;
													assign node2430 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node2433 = (inp[1]) ? node2441 : node2434;
												assign node2434 = (inp[13]) ? node2436 : 4'b1110;
													assign node2436 = (inp[11]) ? node2438 : 4'b1111;
														assign node2438 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node2441 = (inp[15]) ? 4'b1010 : node2442;
													assign node2442 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node2446 = (inp[13]) ? node2518 : node2447;
										assign node2447 = (inp[9]) ? node2495 : node2448;
											assign node2448 = (inp[1]) ? node2478 : node2449;
												assign node2449 = (inp[2]) ? node2465 : node2450;
													assign node2450 = (inp[15]) ? node2456 : node2451;
														assign node2451 = (inp[5]) ? 4'b1110 : node2452;
															assign node2452 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node2456 = (inp[5]) ? node2462 : node2457;
															assign node2457 = (inp[11]) ? node2459 : 4'b1111;
																assign node2459 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node2462 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node2465 = (inp[11]) ? node2475 : node2466;
														assign node2466 = (inp[0]) ? node2472 : node2467;
															assign node2467 = (inp[15]) ? 4'b1111 : node2468;
																assign node2468 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node2472 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node2475 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node2478 = (inp[11]) ? node2486 : node2479;
													assign node2479 = (inp[5]) ? node2481 : 4'b1110;
														assign node2481 = (inp[0]) ? 4'b1010 : node2482;
															assign node2482 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node2486 = (inp[5]) ? node2490 : node2487;
														assign node2487 = (inp[15]) ? 4'b1010 : 4'b1111;
														assign node2490 = (inp[0]) ? 4'b1111 : node2491;
															assign node2491 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node2495 = (inp[5]) ? node2513 : node2496;
												assign node2496 = (inp[1]) ? node2506 : node2497;
													assign node2497 = (inp[11]) ? node2503 : node2498;
														assign node2498 = (inp[2]) ? 4'b1011 : node2499;
															assign node2499 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node2503 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node2506 = (inp[15]) ? node2510 : node2507;
														assign node2507 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node2510 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node2513 = (inp[11]) ? node2515 : 4'b1011;
													assign node2515 = (inp[2]) ? 4'b1111 : 4'b1011;
										assign node2518 = (inp[11]) ? node2544 : node2519;
											assign node2519 = (inp[0]) ? node2537 : node2520;
												assign node2520 = (inp[5]) ? node2530 : node2521;
													assign node2521 = (inp[15]) ? node2527 : node2522;
														assign node2522 = (inp[1]) ? 4'b1111 : node2523;
															assign node2523 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node2527 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node2530 = (inp[2]) ? 4'b1011 : node2531;
														assign node2531 = (inp[9]) ? node2533 : 4'b1010;
															assign node2533 = (inp[15]) ? 4'b1110 : 4'b1010;
												assign node2537 = (inp[5]) ? node2539 : 4'b1110;
													assign node2539 = (inp[2]) ? node2541 : 4'b1011;
														assign node2541 = (inp[1]) ? 4'b1011 : 4'b1111;
											assign node2544 = (inp[9]) ? node2564 : node2545;
												assign node2545 = (inp[2]) ? node2551 : node2546;
													assign node2546 = (inp[0]) ? node2548 : 4'b1110;
														assign node2548 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node2551 = (inp[15]) ? node2555 : node2552;
														assign node2552 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node2555 = (inp[0]) ? node2559 : node2556;
															assign node2556 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node2559 = (inp[1]) ? node2561 : 4'b1110;
																assign node2561 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node2564 = (inp[0]) ? node2574 : node2565;
													assign node2565 = (inp[1]) ? node2567 : 4'b1010;
														assign node2567 = (inp[2]) ? 4'b1010 : node2568;
															assign node2568 = (inp[15]) ? node2570 : 4'b1011;
																assign node2570 = (inp[5]) ? 4'b1110 : 4'b1011;
													assign node2574 = (inp[1]) ? 4'b1010 : node2575;
														assign node2575 = (inp[2]) ? 4'b1111 : 4'b1110;
							assign node2579 = (inp[9]) ? node2771 : node2580;
								assign node2580 = (inp[10]) ? node2662 : node2581;
									assign node2581 = (inp[0]) ? node2621 : node2582;
										assign node2582 = (inp[5]) ? node2588 : node2583;
											assign node2583 = (inp[15]) ? node2585 : 4'b1000;
												assign node2585 = (inp[2]) ? 4'b1101 : 4'b1000;
											assign node2588 = (inp[11]) ? node2608 : node2589;
												assign node2589 = (inp[7]) ? node2599 : node2590;
													assign node2590 = (inp[15]) ? node2592 : 4'b1100;
														assign node2592 = (inp[1]) ? node2596 : node2593;
															assign node2593 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node2596 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node2599 = (inp[2]) ? node2605 : node2600;
														assign node2600 = (inp[13]) ? node2602 : 4'b1100;
															assign node2602 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node2605 = (inp[1]) ? 4'b1001 : 4'b1100;
												assign node2608 = (inp[1]) ? node2616 : node2609;
													assign node2609 = (inp[2]) ? node2613 : node2610;
														assign node2610 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node2613 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node2616 = (inp[2]) ? 4'b1000 : node2617;
														assign node2617 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node2621 = (inp[15]) ? node2645 : node2622;
											assign node2622 = (inp[2]) ? node2638 : node2623;
												assign node2623 = (inp[7]) ? node2635 : node2624;
													assign node2624 = (inp[11]) ? node2628 : node2625;
														assign node2625 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node2628 = (inp[1]) ? node2632 : node2629;
															assign node2629 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node2632 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node2635 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node2638 = (inp[1]) ? node2642 : node2639;
													assign node2639 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node2642 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node2645 = (inp[7]) ? node2653 : node2646;
												assign node2646 = (inp[11]) ? 4'b1100 : node2647;
													assign node2647 = (inp[2]) ? node2649 : 4'b1001;
														assign node2649 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node2653 = (inp[2]) ? node2657 : node2654;
													assign node2654 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node2657 = (inp[11]) ? 4'b1001 : node2658;
														assign node2658 = (inp[13]) ? 4'b1000 : 4'b1001;
									assign node2662 = (inp[13]) ? node2708 : node2663;
										assign node2663 = (inp[11]) ? node2679 : node2664;
											assign node2664 = (inp[5]) ? node2672 : node2665;
												assign node2665 = (inp[7]) ? node2669 : node2666;
													assign node2666 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node2669 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node2672 = (inp[0]) ? 4'b1001 : node2673;
													assign node2673 = (inp[2]) ? 4'b1100 : node2674;
														assign node2674 = (inp[1]) ? 4'b1101 : 4'b1001;
											assign node2679 = (inp[5]) ? node2691 : node2680;
												assign node2680 = (inp[0]) ? node2686 : node2681;
													assign node2681 = (inp[1]) ? node2683 : 4'b1000;
														assign node2683 = (inp[7]) ? 4'b1000 : 4'b1101;
													assign node2686 = (inp[7]) ? node2688 : 4'b1100;
														assign node2688 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node2691 = (inp[15]) ? node2703 : node2692;
													assign node2692 = (inp[0]) ? node2700 : node2693;
														assign node2693 = (inp[7]) ? node2695 : 4'b1101;
															assign node2695 = (inp[1]) ? node2697 : 4'b1000;
																assign node2697 = (inp[2]) ? 4'b1000 : 4'b1101;
														assign node2700 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node2703 = (inp[0]) ? node2705 : 4'b1000;
														assign node2705 = (inp[1]) ? 4'b1000 : 4'b1100;
										assign node2708 = (inp[0]) ? node2738 : node2709;
											assign node2709 = (inp[7]) ? node2733 : node2710;
												assign node2710 = (inp[5]) ? node2720 : node2711;
													assign node2711 = (inp[2]) ? 4'b1001 : node2712;
														assign node2712 = (inp[15]) ? node2716 : node2713;
															assign node2713 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node2716 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node2720 = (inp[11]) ? node2730 : node2721;
														assign node2721 = (inp[1]) ? node2725 : node2722;
															assign node2722 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node2725 = (inp[2]) ? node2727 : 4'b1101;
																assign node2727 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node2730 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node2733 = (inp[5]) ? 4'b1101 : node2734;
													assign node2734 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node2738 = (inp[15]) ? node2758 : node2739;
												assign node2739 = (inp[5]) ? node2747 : node2740;
													assign node2740 = (inp[11]) ? 4'b1000 : node2741;
														assign node2741 = (inp[1]) ? node2743 : 4'b1100;
															assign node2743 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node2747 = (inp[2]) ? node2753 : node2748;
														assign node2748 = (inp[1]) ? 4'b1100 : node2749;
															assign node2749 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node2753 = (inp[7]) ? 4'b1001 : node2754;
															assign node2754 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node2758 = (inp[1]) ? node2766 : node2759;
													assign node2759 = (inp[11]) ? 4'b1101 : node2760;
														assign node2760 = (inp[7]) ? node2762 : 4'b1000;
															assign node2762 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node2766 = (inp[11]) ? node2768 : 4'b1101;
														assign node2768 = (inp[5]) ? 4'b1000 : 4'b1001;
								assign node2771 = (inp[13]) ? node2851 : node2772;
									assign node2772 = (inp[5]) ? node2818 : node2773;
										assign node2773 = (inp[7]) ? node2797 : node2774;
											assign node2774 = (inp[0]) ? node2786 : node2775;
												assign node2775 = (inp[10]) ? node2779 : node2776;
													assign node2776 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node2779 = (inp[1]) ? 4'b1101 : node2780;
														assign node2780 = (inp[11]) ? 4'b1101 : node2781;
															assign node2781 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node2786 = (inp[15]) ? node2790 : node2787;
													assign node2787 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node2790 = (inp[1]) ? node2792 : 4'b1000;
														assign node2792 = (inp[2]) ? 4'b1001 : node2793;
															assign node2793 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node2797 = (inp[2]) ? node2809 : node2798;
												assign node2798 = (inp[10]) ? node2802 : node2799;
													assign node2799 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node2802 = (inp[0]) ? node2804 : 4'b1101;
														assign node2804 = (inp[1]) ? 4'b1001 : node2805;
															assign node2805 = (inp[11]) ? 4'b1101 : 4'b1001;
												assign node2809 = (inp[0]) ? node2815 : node2810;
													assign node2810 = (inp[1]) ? node2812 : 4'b1001;
														assign node2812 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node2815 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node2818 = (inp[10]) ? node2832 : node2819;
											assign node2819 = (inp[11]) ? node2827 : node2820;
												assign node2820 = (inp[0]) ? node2822 : 4'b1100;
													assign node2822 = (inp[15]) ? 4'b1101 : node2823;
														assign node2823 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node2827 = (inp[2]) ? 4'b1000 : node2828;
													assign node2828 = (inp[1]) ? 4'b1100 : 4'b1000;
											assign node2832 = (inp[2]) ? node2840 : node2833;
												assign node2833 = (inp[15]) ? node2837 : node2834;
													assign node2834 = (inp[0]) ? 4'b1100 : 4'b1000;
													assign node2837 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node2840 = (inp[1]) ? node2842 : 4'b1101;
													assign node2842 = (inp[0]) ? 4'b1000 : node2843;
														assign node2843 = (inp[11]) ? node2845 : 4'b1000;
															assign node2845 = (inp[15]) ? 4'b1001 : node2846;
																assign node2846 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node2851 = (inp[1]) ? node2889 : node2852;
										assign node2852 = (inp[2]) ? node2872 : node2853;
											assign node2853 = (inp[5]) ? node2867 : node2854;
												assign node2854 = (inp[11]) ? node2858 : node2855;
													assign node2855 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node2858 = (inp[7]) ? node2864 : node2859;
														assign node2859 = (inp[15]) ? 4'b1000 : node2860;
															assign node2860 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node2864 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node2867 = (inp[0]) ? node2869 : 4'b1001;
													assign node2869 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node2872 = (inp[5]) ? node2884 : node2873;
												assign node2873 = (inp[11]) ? node2879 : node2874;
													assign node2874 = (inp[7]) ? 4'b1000 : node2875;
														assign node2875 = (inp[0]) ? 4'b1001 : 4'b1101;
													assign node2879 = (inp[10]) ? 4'b1000 : node2880;
														assign node2880 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node2884 = (inp[0]) ? 4'b1100 : node2885;
													assign node2885 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node2889 = (inp[2]) ? node2911 : node2890;
											assign node2890 = (inp[7]) ? node2902 : node2891;
												assign node2891 = (inp[0]) ? node2893 : 4'b1101;
													assign node2893 = (inp[5]) ? node2897 : node2894;
														assign node2894 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node2897 = (inp[11]) ? node2899 : 4'b1101;
															assign node2899 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node2902 = (inp[5]) ? node2904 : 4'b1100;
													assign node2904 = (inp[11]) ? 4'b1100 : node2905;
														assign node2905 = (inp[0]) ? 4'b1101 : node2906;
															assign node2906 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node2911 = (inp[11]) ? node2919 : node2912;
												assign node2912 = (inp[5]) ? 4'b1000 : node2913;
													assign node2913 = (inp[7]) ? node2915 : 4'b1100;
														assign node2915 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node2919 = (inp[0]) ? 4'b1101 : 4'b1100;
				assign node2922 = (inp[10]) ? node4536 : node2923;
					assign node2923 = (inp[0]) ? node3745 : node2924;
						assign node2924 = (inp[8]) ? node3356 : node2925;
							assign node2925 = (inp[2]) ? node3151 : node2926;
								assign node2926 = (inp[13]) ? node3040 : node2927;
									assign node2927 = (inp[1]) ? node2989 : node2928;
										assign node2928 = (inp[5]) ? node2964 : node2929;
											assign node2929 = (inp[4]) ? node2949 : node2930;
												assign node2930 = (inp[11]) ? node2940 : node2931;
													assign node2931 = (inp[9]) ? node2937 : node2932;
														assign node2932 = (inp[15]) ? 4'b1011 : node2933;
															assign node2933 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node2937 = (inp[12]) ? 4'b1011 : 4'b1101;
													assign node2940 = (inp[7]) ? node2942 : 4'b1101;
														assign node2942 = (inp[12]) ? node2946 : node2943;
															assign node2943 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node2946 = (inp[15]) ? 4'b1010 : 4'b1100;
												assign node2949 = (inp[7]) ? node2957 : node2950;
													assign node2950 = (inp[15]) ? node2954 : node2951;
														assign node2951 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node2954 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node2957 = (inp[12]) ? node2959 : 4'b1011;
														assign node2959 = (inp[11]) ? node2961 : 4'b1000;
															assign node2961 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node2964 = (inp[7]) ? node2974 : node2965;
												assign node2965 = (inp[12]) ? node2971 : node2966;
													assign node2966 = (inp[15]) ? 4'b1111 : node2967;
														assign node2967 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node2971 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node2974 = (inp[11]) ? node2980 : node2975;
													assign node2975 = (inp[15]) ? node2977 : 4'b1111;
														assign node2977 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node2980 = (inp[9]) ? node2982 : 4'b1100;
														assign node2982 = (inp[12]) ? node2986 : node2983;
															assign node2983 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node2986 = (inp[4]) ? 4'b1101 : 4'b1110;
										assign node2989 = (inp[4]) ? node3017 : node2990;
											assign node2990 = (inp[15]) ? node3004 : node2991;
												assign node2991 = (inp[9]) ? node2995 : node2992;
													assign node2992 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node2995 = (inp[5]) ? node2999 : node2996;
														assign node2996 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node2999 = (inp[7]) ? node3001 : 4'b1010;
															assign node3001 = (inp[12]) ? 4'b1100 : 4'b1010;
												assign node3004 = (inp[9]) ? node3006 : 4'b1010;
													assign node3006 = (inp[7]) ? node3014 : node3007;
														assign node3007 = (inp[12]) ? 4'b1100 : node3008;
															assign node3008 = (inp[11]) ? 4'b1011 : node3009;
																assign node3009 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node3014 = (inp[12]) ? 4'b1011 : 4'b1101;
											assign node3017 = (inp[7]) ? node3025 : node3018;
												assign node3018 = (inp[12]) ? node3020 : 4'b1101;
													assign node3020 = (inp[11]) ? node3022 : 4'b1011;
														assign node3022 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node3025 = (inp[12]) ? node3033 : node3026;
													assign node3026 = (inp[9]) ? node3028 : 4'b1011;
														assign node3028 = (inp[15]) ? node3030 : 4'b1011;
															assign node3030 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node3033 = (inp[5]) ? 4'b1001 : node3034;
														assign node3034 = (inp[11]) ? 4'b1000 : node3035;
															assign node3035 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node3040 = (inp[7]) ? node3094 : node3041;
										assign node3041 = (inp[12]) ? node3065 : node3042;
											assign node3042 = (inp[4]) ? node3058 : node3043;
												assign node3043 = (inp[15]) ? node3047 : node3044;
													assign node3044 = (inp[9]) ? 4'b1101 : 4'b1000;
													assign node3047 = (inp[9]) ? node3053 : node3048;
														assign node3048 = (inp[11]) ? node3050 : 4'b1111;
															assign node3050 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node3053 = (inp[1]) ? node3055 : 4'b1010;
															assign node3055 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node3058 = (inp[5]) ? 4'b1100 : node3059;
													assign node3059 = (inp[11]) ? node3061 : 4'b1001;
														assign node3061 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node3065 = (inp[5]) ? node3081 : node3066;
												assign node3066 = (inp[9]) ? node3076 : node3067;
													assign node3067 = (inp[1]) ? node3071 : node3068;
														assign node3068 = (inp[15]) ? 4'b1111 : 4'b1010;
														assign node3071 = (inp[11]) ? 4'b1011 : node3072;
															assign node3072 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node3076 = (inp[4]) ? node3078 : 4'b1000;
														assign node3078 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node3081 = (inp[4]) ? node3091 : node3082;
													assign node3082 = (inp[11]) ? 4'b1110 : node3083;
														assign node3083 = (inp[1]) ? node3087 : node3084;
															assign node3084 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node3087 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node3091 = (inp[15]) ? 4'b1110 : 4'b1010;
										assign node3094 = (inp[5]) ? node3122 : node3095;
											assign node3095 = (inp[11]) ? node3115 : node3096;
												assign node3096 = (inp[4]) ? node3110 : node3097;
													assign node3097 = (inp[9]) ? node3107 : node3098;
														assign node3098 = (inp[15]) ? node3102 : node3099;
															assign node3099 = (inp[1]) ? 4'b1000 : 4'b1110;
															assign node3102 = (inp[12]) ? node3104 : 4'b1001;
																assign node3104 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node3107 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node3110 = (inp[12]) ? 4'b1101 : node3111;
														assign node3111 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node3115 = (inp[9]) ? 4'b1100 : node3116;
													assign node3116 = (inp[4]) ? node3118 : 4'b1111;
														assign node3118 = (inp[12]) ? 4'b1101 : 4'b1111;
											assign node3122 = (inp[1]) ? node3136 : node3123;
												assign node3123 = (inp[15]) ? node3125 : 4'b1011;
													assign node3125 = (inp[11]) ? node3127 : 4'b1001;
														assign node3127 = (inp[9]) ? node3129 : 4'b1000;
															assign node3129 = (inp[12]) ? node3133 : node3130;
																assign node3130 = (inp[4]) ? 4'b1010 : 4'b1001;
																assign node3133 = (inp[4]) ? 4'b1001 : 4'b1010;
												assign node3136 = (inp[12]) ? node3144 : node3137;
													assign node3137 = (inp[11]) ? node3141 : node3138;
														assign node3138 = (inp[4]) ? 4'b1110 : 4'b1001;
														assign node3141 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node3144 = (inp[4]) ? node3146 : 4'b1001;
														assign node3146 = (inp[11]) ? node3148 : 4'b1101;
															assign node3148 = (inp[15]) ? 4'b1100 : 4'b1101;
								assign node3151 = (inp[7]) ? node3267 : node3152;
									assign node3152 = (inp[12]) ? node3206 : node3153;
										assign node3153 = (inp[15]) ? node3179 : node3154;
											assign node3154 = (inp[13]) ? node3162 : node3155;
												assign node3155 = (inp[5]) ? node3157 : 4'b1101;
													assign node3157 = (inp[1]) ? 4'b1101 : node3158;
														assign node3158 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node3162 = (inp[11]) ? node3168 : node3163;
													assign node3163 = (inp[5]) ? node3165 : 4'b1001;
														assign node3165 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node3168 = (inp[4]) ? node3174 : node3169;
														assign node3169 = (inp[5]) ? node3171 : 4'b1001;
															assign node3171 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node3174 = (inp[5]) ? 4'b1000 : node3175;
															assign node3175 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node3179 = (inp[4]) ? node3193 : node3180;
												assign node3180 = (inp[9]) ? node3182 : 4'b1111;
													assign node3182 = (inp[5]) ? node3186 : node3183;
														assign node3183 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node3186 = (inp[11]) ? node3188 : 4'b1010;
															assign node3188 = (inp[1]) ? 4'b1110 : node3189;
																assign node3189 = (inp[13]) ? 4'b1110 : 4'b1011;
												assign node3193 = (inp[5]) ? node3201 : node3194;
													assign node3194 = (inp[13]) ? 4'b1100 : node3195;
														assign node3195 = (inp[9]) ? node3197 : 4'b1000;
															assign node3197 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3201 = (inp[9]) ? 4'b1101 : node3202;
														assign node3202 = (inp[11]) ? 4'b1001 : 4'b1100;
										assign node3206 = (inp[15]) ? node3236 : node3207;
											assign node3207 = (inp[9]) ? node3225 : node3208;
												assign node3208 = (inp[1]) ? node3218 : node3209;
													assign node3209 = (inp[4]) ? node3213 : node3210;
														assign node3210 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node3213 = (inp[5]) ? 4'b1111 : node3214;
															assign node3214 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node3218 = (inp[4]) ? node3220 : 4'b1110;
														assign node3220 = (inp[13]) ? 4'b1111 : node3221;
															assign node3221 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node3225 = (inp[4]) ? 4'b1011 : node3226;
													assign node3226 = (inp[1]) ? node3228 : 4'b1111;
														assign node3228 = (inp[11]) ? node3232 : node3229;
															assign node3229 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node3232 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node3236 = (inp[4]) ? node3252 : node3237;
												assign node3237 = (inp[5]) ? node3241 : node3238;
													assign node3238 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node3241 = (inp[11]) ? node3245 : node3242;
														assign node3242 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node3245 = (inp[13]) ? node3249 : node3246;
															assign node3246 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node3249 = (inp[1]) ? 4'b1100 : 4'b1001;
												assign node3252 = (inp[1]) ? node3260 : node3253;
													assign node3253 = (inp[13]) ? 4'b1011 : node3254;
														assign node3254 = (inp[9]) ? 4'b1111 : node3255;
															assign node3255 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node3260 = (inp[9]) ? node3262 : 4'b1010;
														assign node3262 = (inp[5]) ? 4'b1011 : node3263;
															assign node3263 = (inp[13]) ? 4'b1110 : 4'b1011;
									assign node3267 = (inp[12]) ? node3305 : node3268;
										assign node3268 = (inp[4]) ? node3282 : node3269;
											assign node3269 = (inp[15]) ? node3275 : node3270;
												assign node3270 = (inp[9]) ? node3272 : 4'b1110;
													assign node3272 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node3275 = (inp[13]) ? 4'b1100 : node3276;
													assign node3276 = (inp[1]) ? 4'b1101 : node3277;
														assign node3277 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node3282 = (inp[13]) ? node3298 : node3283;
												assign node3283 = (inp[11]) ? node3287 : node3284;
													assign node3284 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node3287 = (inp[1]) ? node3291 : node3288;
														assign node3288 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node3291 = (inp[5]) ? node3293 : 4'b1111;
															assign node3293 = (inp[9]) ? 4'b1111 : node3294;
																assign node3294 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node3298 = (inp[9]) ? node3302 : node3299;
													assign node3299 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node3302 = (inp[1]) ? 4'b1011 : 4'b1010;
										assign node3305 = (inp[4]) ? node3329 : node3306;
											assign node3306 = (inp[15]) ? node3320 : node3307;
												assign node3307 = (inp[5]) ? node3309 : 4'b1001;
													assign node3309 = (inp[13]) ? node3313 : node3310;
														assign node3310 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node3313 = (inp[1]) ? node3315 : 4'b1000;
															assign node3315 = (inp[9]) ? node3317 : 4'b1101;
																assign node3317 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node3320 = (inp[9]) ? 4'b1110 : node3321;
													assign node3321 = (inp[11]) ? node3325 : node3322;
														assign node3322 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node3325 = (inp[1]) ? 4'b1011 : 4'b1111;
											assign node3329 = (inp[5]) ? node3339 : node3330;
												assign node3330 = (inp[1]) ? 4'b1100 : node3331;
													assign node3331 = (inp[11]) ? 4'b1100 : node3332;
														assign node3332 = (inp[15]) ? 4'b1101 : node3333;
															assign node3333 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node3339 = (inp[11]) ? node3343 : node3340;
													assign node3340 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node3343 = (inp[13]) ? node3347 : node3344;
														assign node3344 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node3347 = (inp[1]) ? 4'b1000 : node3348;
															assign node3348 = (inp[9]) ? node3352 : node3349;
																assign node3349 = (inp[15]) ? 4'b1101 : 4'b1100;
																assign node3352 = (inp[15]) ? 4'b1100 : 4'b1101;
							assign node3356 = (inp[9]) ? node3544 : node3357;
								assign node3357 = (inp[11]) ? node3453 : node3358;
									assign node3358 = (inp[13]) ? node3402 : node3359;
										assign node3359 = (inp[7]) ? node3389 : node3360;
											assign node3360 = (inp[1]) ? node3380 : node3361;
												assign node3361 = (inp[5]) ? node3367 : node3362;
													assign node3362 = (inp[2]) ? 4'b1100 : node3363;
														assign node3363 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node3367 = (inp[12]) ? node3377 : node3368;
														assign node3368 = (inp[4]) ? node3372 : node3369;
															assign node3369 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node3372 = (inp[2]) ? 4'b1110 : node3373;
																assign node3373 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node3377 = (inp[15]) ? 4'b1101 : 4'b1001;
												assign node3380 = (inp[4]) ? 4'b1000 : node3381;
													assign node3381 = (inp[12]) ? node3383 : 4'b1001;
														assign node3383 = (inp[15]) ? 4'b1010 : node3384;
															assign node3384 = (inp[2]) ? 4'b1010 : 4'b1111;
											assign node3389 = (inp[12]) ? node3397 : node3390;
												assign node3390 = (inp[4]) ? node3392 : 4'b1101;
													assign node3392 = (inp[5]) ? 4'b1111 : node3393;
														assign node3393 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node3397 = (inp[15]) ? 4'b1010 : node3398;
													assign node3398 = (inp[2]) ? 4'b1100 : 4'b1001;
										assign node3402 = (inp[15]) ? node3424 : node3403;
											assign node3403 = (inp[5]) ? node3415 : node3404;
												assign node3404 = (inp[2]) ? node3410 : node3405;
													assign node3405 = (inp[12]) ? 4'b1010 : node3406;
														assign node3406 = (inp[4]) ? 4'b1010 : 4'b1000;
													assign node3410 = (inp[1]) ? 4'b1010 : node3411;
														assign node3411 = (inp[7]) ? 4'b1010 : 4'b1111;
												assign node3415 = (inp[7]) ? node3419 : node3416;
													assign node3416 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node3419 = (inp[1]) ? 4'b1010 : node3420;
														assign node3420 = (inp[4]) ? 4'b1010 : 4'b1111;
											assign node3424 = (inp[5]) ? node3440 : node3425;
												assign node3425 = (inp[4]) ? node3433 : node3426;
													assign node3426 = (inp[12]) ? node3430 : node3427;
														assign node3427 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node3430 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node3433 = (inp[2]) ? node3435 : 4'b1110;
														assign node3435 = (inp[1]) ? 4'b1101 : node3436;
															assign node3436 = (inp[7]) ? 4'b1111 : 4'b1011;
												assign node3440 = (inp[1]) ? node3442 : 4'b1010;
													assign node3442 = (inp[12]) ? node3448 : node3443;
														assign node3443 = (inp[2]) ? 4'b1100 : node3444;
															assign node3444 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node3448 = (inp[2]) ? node3450 : 4'b1111;
															assign node3450 = (inp[4]) ? 4'b1000 : 4'b1010;
									assign node3453 = (inp[4]) ? node3501 : node3454;
										assign node3454 = (inp[12]) ? node3476 : node3455;
											assign node3455 = (inp[15]) ? node3463 : node3456;
												assign node3456 = (inp[5]) ? 4'b1101 : node3457;
													assign node3457 = (inp[7]) ? 4'b1100 : node3458;
														assign node3458 = (inp[1]) ? 4'b1100 : 4'b1001;
												assign node3463 = (inp[5]) ? node3473 : node3464;
													assign node3464 = (inp[7]) ? node3470 : node3465;
														assign node3465 = (inp[1]) ? node3467 : 4'b1001;
															assign node3467 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node3470 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node3473 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node3476 = (inp[2]) ? node3488 : node3477;
												assign node3477 = (inp[1]) ? node3481 : node3478;
													assign node3478 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node3481 = (inp[5]) ? 4'b1111 : node3482;
														assign node3482 = (inp[7]) ? node3484 : 4'b1011;
															assign node3484 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node3488 = (inp[15]) ? node3494 : node3489;
													assign node3489 = (inp[7]) ? 4'b1110 : node3490;
														assign node3490 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node3494 = (inp[1]) ? node3496 : 4'b1110;
														assign node3496 = (inp[13]) ? 4'b1010 : node3497;
															assign node3497 = (inp[5]) ? 4'b1010 : 4'b1011;
										assign node3501 = (inp[12]) ? node3513 : node3502;
											assign node3502 = (inp[2]) ? node3510 : node3503;
												assign node3503 = (inp[13]) ? node3505 : 4'b1011;
													assign node3505 = (inp[15]) ? node3507 : 4'b1110;
														assign node3507 = (inp[1]) ? 4'b1110 : 4'b1010;
												assign node3510 = (inp[1]) ? 4'b1011 : 4'b1111;
											assign node3513 = (inp[5]) ? node3531 : node3514;
												assign node3514 = (inp[7]) ? node3524 : node3515;
													assign node3515 = (inp[13]) ? node3519 : node3516;
														assign node3516 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node3519 = (inp[1]) ? node3521 : 4'b1101;
															assign node3521 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node3524 = (inp[15]) ? 4'b1100 : node3525;
														assign node3525 = (inp[13]) ? node3527 : 4'b1000;
															assign node3527 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node3531 = (inp[2]) ? node3539 : node3532;
													assign node3532 = (inp[1]) ? 4'b1101 : node3533;
														assign node3533 = (inp[15]) ? node3535 : 4'b1001;
															assign node3535 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node3539 = (inp[1]) ? 4'b1000 : node3540;
														assign node3540 = (inp[13]) ? 4'b1001 : 4'b1000;
								assign node3544 = (inp[2]) ? node3654 : node3545;
									assign node3545 = (inp[1]) ? node3605 : node3546;
										assign node3546 = (inp[7]) ? node3578 : node3547;
											assign node3547 = (inp[13]) ? node3561 : node3548;
												assign node3548 = (inp[11]) ? node3556 : node3549;
													assign node3549 = (inp[4]) ? node3553 : node3550;
														assign node3550 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node3553 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node3556 = (inp[15]) ? 4'b1001 : node3557;
														assign node3557 = (inp[12]) ? 4'b1100 : 4'b1001;
												assign node3561 = (inp[4]) ? node3567 : node3562;
													assign node3562 = (inp[12]) ? 4'b1010 : node3563;
														assign node3563 = (inp[15]) ? 4'b1001 : 4'b1100;
													assign node3567 = (inp[12]) ? node3573 : node3568;
														assign node3568 = (inp[15]) ? node3570 : 4'b1010;
															assign node3570 = (inp[11]) ? 4'b1111 : 4'b1010;
														assign node3573 = (inp[15]) ? 4'b1100 : node3574;
															assign node3574 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node3578 = (inp[4]) ? node3592 : node3579;
												assign node3579 = (inp[12]) ? node3589 : node3580;
													assign node3580 = (inp[5]) ? 4'b1100 : node3581;
														assign node3581 = (inp[15]) ? node3585 : node3582;
															assign node3582 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node3585 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node3589 = (inp[15]) ? 4'b1010 : 4'b1111;
												assign node3592 = (inp[12]) ? 4'b1001 : node3593;
													assign node3593 = (inp[11]) ? node3595 : 4'b1010;
														assign node3595 = (inp[5]) ? node3599 : node3596;
															assign node3596 = (inp[13]) ? 4'b1011 : 4'b1010;
															assign node3599 = (inp[15]) ? 4'b1010 : node3600;
																assign node3600 = (inp[13]) ? 4'b1010 : 4'b1011;
										assign node3605 = (inp[7]) ? node3635 : node3606;
											assign node3606 = (inp[15]) ? node3622 : node3607;
												assign node3607 = (inp[13]) ? node3615 : node3608;
													assign node3608 = (inp[4]) ? node3612 : node3609;
														assign node3609 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node3612 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node3615 = (inp[11]) ? 4'b1111 : node3616;
														assign node3616 = (inp[4]) ? node3618 : 4'b1110;
															assign node3618 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node3622 = (inp[5]) ? node3632 : node3623;
													assign node3623 = (inp[4]) ? node3629 : node3624;
														assign node3624 = (inp[13]) ? 4'b1011 : node3625;
															assign node3625 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node3629 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node3632 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node3635 = (inp[4]) ? node3645 : node3636;
												assign node3636 = (inp[12]) ? node3640 : node3637;
													assign node3637 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node3640 = (inp[5]) ? 4'b1111 : node3641;
														assign node3641 = (inp[15]) ? 4'b1110 : 4'b1010;
												assign node3645 = (inp[12]) ? node3651 : node3646;
													assign node3646 = (inp[15]) ? node3648 : 4'b1110;
														assign node3648 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node3651 = (inp[13]) ? 4'b1100 : 4'b1101;
									assign node3654 = (inp[1]) ? node3698 : node3655;
										assign node3655 = (inp[7]) ? node3675 : node3656;
											assign node3656 = (inp[4]) ? node3666 : node3657;
												assign node3657 = (inp[12]) ? node3663 : node3658;
													assign node3658 = (inp[11]) ? node3660 : 4'b1100;
														assign node3660 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node3663 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node3666 = (inp[12]) ? node3668 : 4'b1010;
													assign node3668 = (inp[11]) ? node3670 : 4'b1100;
														assign node3670 = (inp[13]) ? 4'b1001 : node3671;
															assign node3671 = (inp[5]) ? 4'b1100 : 4'b1000;
											assign node3675 = (inp[4]) ? node3689 : node3676;
												assign node3676 = (inp[12]) ? node3680 : node3677;
													assign node3677 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node3680 = (inp[13]) ? node3684 : node3681;
														assign node3681 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node3684 = (inp[5]) ? 4'b1110 : node3685;
															assign node3685 = (inp[15]) ? 4'b1110 : 4'b1011;
												assign node3689 = (inp[12]) ? node3693 : node3690;
													assign node3690 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node3693 = (inp[15]) ? 4'b1100 : node3694;
														assign node3694 = (inp[13]) ? 4'b1101 : 4'b1100;
										assign node3698 = (inp[15]) ? node3722 : node3699;
											assign node3699 = (inp[13]) ? node3707 : node3700;
												assign node3700 = (inp[7]) ? node3704 : node3701;
													assign node3701 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node3704 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node3707 = (inp[11]) ? node3713 : node3708;
													assign node3708 = (inp[7]) ? 4'b1111 : node3709;
														assign node3709 = (inp[12]) ? 4'b1010 : 4'b1001;
													assign node3713 = (inp[7]) ? node3717 : node3714;
														assign node3714 = (inp[12]) ? 4'b1100 : 4'b1001;
														assign node3717 = (inp[5]) ? node3719 : 4'b1000;
															assign node3719 = (inp[4]) ? 4'b1010 : 4'b1000;
											assign node3722 = (inp[7]) ? node3736 : node3723;
												assign node3723 = (inp[5]) ? node3733 : node3724;
													assign node3724 = (inp[11]) ? node3730 : node3725;
														assign node3725 = (inp[12]) ? node3727 : 4'b1001;
															assign node3727 = (inp[4]) ? 4'b1101 : 4'b1110;
														assign node3730 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node3733 = (inp[12]) ? 4'b1010 : 4'b1001;
												assign node3736 = (inp[11]) ? 4'b1100 : node3737;
													assign node3737 = (inp[4]) ? node3741 : node3738;
														assign node3738 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node3741 = (inp[5]) ? 4'b1001 : 4'b1000;
						assign node3745 = (inp[8]) ? node4161 : node3746;
							assign node3746 = (inp[15]) ? node3948 : node3747;
								assign node3747 = (inp[4]) ? node3855 : node3748;
									assign node3748 = (inp[5]) ? node3804 : node3749;
										assign node3749 = (inp[1]) ? node3777 : node3750;
											assign node3750 = (inp[13]) ? node3766 : node3751;
												assign node3751 = (inp[2]) ? node3759 : node3752;
													assign node3752 = (inp[7]) ? node3756 : node3753;
														assign node3753 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node3756 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node3759 = (inp[9]) ? node3763 : node3760;
														assign node3760 = (inp[12]) ? 4'b1110 : 4'b1100;
														assign node3763 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node3766 = (inp[2]) ? node3774 : node3767;
													assign node3767 = (inp[9]) ? 4'b1000 : node3768;
														assign node3768 = (inp[7]) ? 4'b1110 : node3769;
															assign node3769 = (inp[12]) ? 4'b1110 : 4'b1100;
													assign node3774 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node3777 = (inp[7]) ? node3793 : node3778;
												assign node3778 = (inp[12]) ? node3788 : node3779;
													assign node3779 = (inp[11]) ? node3783 : node3780;
														assign node3780 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node3783 = (inp[9]) ? node3785 : 4'b1001;
															assign node3785 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node3788 = (inp[9]) ? 4'b1011 : node3789;
														assign node3789 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node3793 = (inp[12]) ? node3799 : node3794;
													assign node3794 = (inp[13]) ? node3796 : 4'b1011;
														assign node3796 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node3799 = (inp[13]) ? 4'b1100 : node3800;
														assign node3800 = (inp[2]) ? 4'b1000 : 4'b1100;
										assign node3804 = (inp[7]) ? node3832 : node3805;
											assign node3805 = (inp[12]) ? node3809 : node3806;
												assign node3806 = (inp[2]) ? 4'b1000 : 4'b1101;
												assign node3809 = (inp[11]) ? node3827 : node3810;
													assign node3810 = (inp[9]) ? node3818 : node3811;
														assign node3811 = (inp[1]) ? node3813 : 4'b1011;
															assign node3813 = (inp[2]) ? 4'b1011 : node3814;
																assign node3814 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node3818 = (inp[1]) ? node3822 : node3819;
															assign node3819 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node3822 = (inp[2]) ? 4'b1111 : node3823;
																assign node3823 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node3827 = (inp[13]) ? 4'b1011 : node3828;
														assign node3828 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node3832 = (inp[12]) ? node3852 : node3833;
												assign node3833 = (inp[9]) ? node3843 : node3834;
													assign node3834 = (inp[1]) ? node3838 : node3835;
														assign node3835 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node3838 = (inp[13]) ? 4'b1011 : node3839;
															assign node3839 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node3843 = (inp[2]) ? node3847 : node3844;
														assign node3844 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node3847 = (inp[13]) ? 4'b1111 : node3848;
															assign node3848 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node3852 = (inp[13]) ? 4'b1100 : 4'b1101;
									assign node3855 = (inp[11]) ? node3903 : node3856;
										assign node3856 = (inp[13]) ? node3872 : node3857;
											assign node3857 = (inp[2]) ? node3865 : node3858;
												assign node3858 = (inp[9]) ? node3860 : 4'b1010;
													assign node3860 = (inp[5]) ? 4'b1000 : node3861;
														assign node3861 = (inp[1]) ? 4'b1011 : 4'b1000;
												assign node3865 = (inp[12]) ? node3869 : node3866;
													assign node3866 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node3869 = (inp[9]) ? 4'b1000 : 4'b1100;
											assign node3872 = (inp[7]) ? node3888 : node3873;
												assign node3873 = (inp[12]) ? node3885 : node3874;
													assign node3874 = (inp[1]) ? node3882 : node3875;
														assign node3875 = (inp[2]) ? node3877 : 4'b1001;
															assign node3877 = (inp[5]) ? 4'b1100 : node3878;
																assign node3878 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node3882 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node3885 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node3888 = (inp[12]) ? node3894 : node3889;
													assign node3889 = (inp[9]) ? node3891 : 4'b1110;
														assign node3891 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node3894 = (inp[5]) ? node3900 : node3895;
														assign node3895 = (inp[9]) ? 4'b1101 : node3896;
															assign node3896 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node3900 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node3903 = (inp[1]) ? node3925 : node3904;
											assign node3904 = (inp[2]) ? node3916 : node3905;
												assign node3905 = (inp[5]) ? node3913 : node3906;
													assign node3906 = (inp[13]) ? 4'b1010 : node3907;
														assign node3907 = (inp[12]) ? 4'b1001 : node3908;
															assign node3908 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node3913 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node3916 = (inp[13]) ? node3922 : node3917;
													assign node3917 = (inp[9]) ? node3919 : 4'b1000;
														assign node3919 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node3922 = (inp[7]) ? 4'b1000 : 4'b1110;
											assign node3925 = (inp[12]) ? node3937 : node3926;
												assign node3926 = (inp[7]) ? node3932 : node3927;
													assign node3927 = (inp[5]) ? 4'b1101 : node3928;
														assign node3928 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node3932 = (inp[9]) ? node3934 : 4'b1110;
														assign node3934 = (inp[13]) ? 4'b1011 : 4'b1110;
												assign node3937 = (inp[7]) ? node3945 : node3938;
													assign node3938 = (inp[9]) ? node3942 : node3939;
														assign node3939 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node3942 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node3945 = (inp[9]) ? 4'b1001 : 4'b1000;
								assign node3948 = (inp[11]) ? node4048 : node3949;
									assign node3949 = (inp[13]) ? node4003 : node3950;
										assign node3950 = (inp[5]) ? node3978 : node3951;
											assign node3951 = (inp[7]) ? node3961 : node3952;
												assign node3952 = (inp[9]) ? node3954 : 4'b1100;
													assign node3954 = (inp[1]) ? 4'b1011 : node3955;
														assign node3955 = (inp[12]) ? 4'b1000 : node3956;
															assign node3956 = (inp[2]) ? 4'b1001 : 4'b1011;
												assign node3961 = (inp[2]) ? node3969 : node3962;
													assign node3962 = (inp[1]) ? 4'b1010 : node3963;
														assign node3963 = (inp[12]) ? 4'b1011 : node3964;
															assign node3964 = (inp[4]) ? 4'b1011 : 4'b1100;
													assign node3969 = (inp[4]) ? node3973 : node3970;
														assign node3970 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node3973 = (inp[12]) ? node3975 : 4'b1110;
															assign node3975 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node3978 = (inp[1]) ? node4000 : node3979;
												assign node3979 = (inp[2]) ? node3993 : node3980;
													assign node3980 = (inp[7]) ? node3988 : node3981;
														assign node3981 = (inp[4]) ? node3985 : node3982;
															assign node3982 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node3985 = (inp[12]) ? 4'b1011 : 4'b1000;
														assign node3988 = (inp[12]) ? 4'b1100 : node3989;
															assign node3989 = (inp[4]) ? 4'b1110 : 4'b1100;
													assign node3993 = (inp[7]) ? node3997 : node3994;
														assign node3994 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node3997 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node4000 = (inp[9]) ? 4'b1101 : 4'b1110;
										assign node4003 = (inp[4]) ? node4025 : node4004;
											assign node4004 = (inp[5]) ? node4014 : node4005;
												assign node4005 = (inp[2]) ? node4011 : node4006;
													assign node4006 = (inp[12]) ? node4008 : 4'b1001;
														assign node4008 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node4011 = (inp[12]) ? 4'b1010 : 4'b1000;
												assign node4014 = (inp[12]) ? node4020 : node4015;
													assign node4015 = (inp[7]) ? 4'b1000 : node4016;
														assign node4016 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node4020 = (inp[7]) ? 4'b1011 : node4021;
														assign node4021 = (inp[1]) ? 4'b1101 : 4'b1001;
											assign node4025 = (inp[2]) ? node4039 : node4026;
												assign node4026 = (inp[9]) ? node4034 : node4027;
													assign node4027 = (inp[12]) ? 4'b1110 : node4028;
														assign node4028 = (inp[7]) ? 4'b1110 : node4029;
															assign node4029 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node4034 = (inp[5]) ? node4036 : 4'b1001;
														assign node4036 = (inp[7]) ? 4'b1101 : 4'b1111;
												assign node4039 = (inp[5]) ? node4041 : 4'b1010;
													assign node4041 = (inp[1]) ? node4045 : node4042;
														assign node4042 = (inp[7]) ? 4'b1111 : 4'b1011;
														assign node4045 = (inp[12]) ? 4'b1010 : 4'b1011;
									assign node4048 = (inp[7]) ? node4098 : node4049;
										assign node4049 = (inp[5]) ? node4071 : node4050;
											assign node4050 = (inp[9]) ? node4062 : node4051;
												assign node4051 = (inp[13]) ? node4057 : node4052;
													assign node4052 = (inp[4]) ? node4054 : 4'b1110;
														assign node4054 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node4057 = (inp[12]) ? node4059 : 4'b1111;
														assign node4059 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node4062 = (inp[2]) ? node4066 : node4063;
													assign node4063 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node4066 = (inp[13]) ? node4068 : 4'b1001;
														assign node4068 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node4071 = (inp[1]) ? node4089 : node4072;
												assign node4072 = (inp[13]) ? node4080 : node4073;
													assign node4073 = (inp[9]) ? node4075 : 4'b1011;
														assign node4075 = (inp[12]) ? 4'b1010 : node4076;
															assign node4076 = (inp[2]) ? 4'b1010 : 4'b1000;
													assign node4080 = (inp[9]) ? 4'b1100 : node4081;
														assign node4081 = (inp[12]) ? node4085 : node4082;
															assign node4082 = (inp[4]) ? 4'b1000 : 4'b1110;
															assign node4085 = (inp[4]) ? 4'b1010 : 4'b1000;
												assign node4089 = (inp[2]) ? 4'b1000 : node4090;
													assign node4090 = (inp[9]) ? node4094 : node4091;
														assign node4091 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node4094 = (inp[12]) ? 4'b1101 : 4'b1010;
										assign node4098 = (inp[12]) ? node4120 : node4099;
											assign node4099 = (inp[4]) ? node4115 : node4100;
												assign node4100 = (inp[9]) ? node4108 : node4101;
													assign node4101 = (inp[5]) ? node4103 : 4'b1001;
														assign node4103 = (inp[2]) ? node4105 : 4'b1001;
															assign node4105 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node4108 = (inp[13]) ? 4'b1000 : node4109;
														assign node4109 = (inp[2]) ? 4'b1000 : node4110;
															assign node4110 = (inp[1]) ? 4'b1000 : 4'b1101;
												assign node4115 = (inp[1]) ? 4'b1010 : node4116;
													assign node4116 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node4120 = (inp[4]) ? node4132 : node4121;
												assign node4121 = (inp[5]) ? node4129 : node4122;
													assign node4122 = (inp[13]) ? node4126 : node4123;
														assign node4123 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node4126 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node4129 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node4132 = (inp[1]) ? node4150 : node4133;
													assign node4133 = (inp[5]) ? node4141 : node4134;
														assign node4134 = (inp[13]) ? node4138 : node4135;
															assign node4135 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node4138 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node4141 = (inp[13]) ? node4147 : node4142;
															assign node4142 = (inp[9]) ? node4144 : 4'b1101;
																assign node4144 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node4147 = (inp[9]) ? 4'b1101 : 4'b1000;
													assign node4150 = (inp[5]) ? node4156 : node4151;
														assign node4151 = (inp[2]) ? node4153 : 4'b1000;
															assign node4153 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node4156 = (inp[13]) ? 4'b1000 : node4157;
															assign node4157 = (inp[9]) ? 4'b1000 : 4'b1001;
							assign node4161 = (inp[13]) ? node4371 : node4162;
								assign node4162 = (inp[15]) ? node4284 : node4163;
									assign node4163 = (inp[7]) ? node4223 : node4164;
										assign node4164 = (inp[2]) ? node4194 : node4165;
											assign node4165 = (inp[5]) ? node4177 : node4166;
												assign node4166 = (inp[1]) ? node4170 : node4167;
													assign node4167 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node4170 = (inp[11]) ? node4172 : 4'b1101;
														assign node4172 = (inp[4]) ? 4'b1100 : node4173;
															assign node4173 = (inp[12]) ? 4'b1111 : 4'b1100;
												assign node4177 = (inp[1]) ? node4187 : node4178;
													assign node4178 = (inp[4]) ? node4182 : node4179;
														assign node4179 = (inp[12]) ? 4'b1011 : 4'b1101;
														assign node4182 = (inp[12]) ? node4184 : 4'b1111;
															assign node4184 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node4187 = (inp[12]) ? 4'b1001 : node4188;
														assign node4188 = (inp[4]) ? node4190 : 4'b1001;
															assign node4190 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node4194 = (inp[9]) ? node4206 : node4195;
												assign node4195 = (inp[1]) ? node4197 : 4'b1011;
													assign node4197 = (inp[12]) ? node4203 : node4198;
														assign node4198 = (inp[4]) ? 4'b1010 : node4199;
															assign node4199 = (inp[11]) ? 4'b1001 : 4'b1100;
														assign node4203 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node4206 = (inp[11]) ? node4218 : node4207;
													assign node4207 = (inp[4]) ? node4213 : node4208;
														assign node4208 = (inp[5]) ? node4210 : 4'b1101;
															assign node4210 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node4213 = (inp[12]) ? node4215 : 4'b1011;
															assign node4215 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node4218 = (inp[4]) ? 4'b1010 : node4219;
														assign node4219 = (inp[12]) ? 4'b1011 : 4'b1001;
										assign node4223 = (inp[11]) ? node4253 : node4224;
											assign node4224 = (inp[9]) ? node4238 : node4225;
												assign node4225 = (inp[1]) ? node4233 : node4226;
													assign node4226 = (inp[4]) ? node4230 : node4227;
														assign node4227 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node4230 = (inp[2]) ? 4'b1110 : 4'b1011;
													assign node4233 = (inp[12]) ? node4235 : 4'b1101;
														assign node4235 = (inp[2]) ? 4'b1001 : 4'b1011;
												assign node4238 = (inp[1]) ? node4248 : node4239;
													assign node4239 = (inp[2]) ? node4243 : node4240;
														assign node4240 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node4243 = (inp[4]) ? 4'b1110 : node4244;
															assign node4244 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node4248 = (inp[12]) ? 4'b1110 : node4249;
														assign node4249 = (inp[5]) ? 4'b1100 : 4'b1101;
											assign node4253 = (inp[2]) ? node4267 : node4254;
												assign node4254 = (inp[1]) ? node4264 : node4255;
													assign node4255 = (inp[5]) ? node4259 : node4256;
														assign node4256 = (inp[12]) ? 4'b1001 : 4'b1010;
														assign node4259 = (inp[4]) ? 4'b1010 : node4260;
															assign node4260 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node4264 = (inp[12]) ? 4'b1010 : 4'b1100;
												assign node4267 = (inp[1]) ? node4275 : node4268;
													assign node4268 = (inp[12]) ? node4272 : node4269;
														assign node4269 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node4272 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node4275 = (inp[4]) ? node4281 : node4276;
														assign node4276 = (inp[12]) ? node4278 : 4'b1001;
															assign node4278 = (inp[5]) ? 4'b1010 : 4'b1111;
														assign node4281 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node4284 = (inp[11]) ? node4322 : node4285;
										assign node4285 = (inp[1]) ? node4305 : node4286;
											assign node4286 = (inp[4]) ? node4302 : node4287;
												assign node4287 = (inp[12]) ? node4299 : node4288;
													assign node4288 = (inp[9]) ? 4'b1001 : node4289;
														assign node4289 = (inp[7]) ? node4291 : 4'b1100;
															assign node4291 = (inp[5]) ? node4295 : node4292;
																assign node4292 = (inp[2]) ? 4'b1100 : 4'b1001;
																assign node4295 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node4299 = (inp[2]) ? 4'b1110 : 4'b1011;
												assign node4302 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node4305 = (inp[12]) ? node4315 : node4306;
												assign node4306 = (inp[4]) ? node4310 : node4307;
													assign node4307 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node4310 = (inp[2]) ? 4'b1010 : node4311;
														assign node4311 = (inp[7]) ? 4'b1110 : 4'b1010;
												assign node4315 = (inp[4]) ? node4317 : 4'b1111;
													assign node4317 = (inp[2]) ? 4'b1000 : node4318;
														assign node4318 = (inp[5]) ? 4'b1100 : 4'b1001;
										assign node4322 = (inp[5]) ? node4346 : node4323;
											assign node4323 = (inp[4]) ? node4335 : node4324;
												assign node4324 = (inp[12]) ? node4328 : node4325;
													assign node4325 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node4328 = (inp[1]) ? 4'b1111 : node4329;
														assign node4329 = (inp[7]) ? node4331 : 4'b1011;
															assign node4331 = (inp[2]) ? 4'b1110 : 4'b1011;
												assign node4335 = (inp[12]) ? node4341 : node4336;
													assign node4336 = (inp[9]) ? node4338 : 4'b1111;
														assign node4338 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node4341 = (inp[7]) ? 4'b1101 : node4342;
														assign node4342 = (inp[9]) ? 4'b1100 : 4'b1001;
											assign node4346 = (inp[2]) ? node4358 : node4347;
												assign node4347 = (inp[1]) ? node4353 : node4348;
													assign node4348 = (inp[12]) ? 4'b1011 : node4349;
														assign node4349 = (inp[7]) ? 4'b1100 : 4'b1011;
													assign node4353 = (inp[7]) ? node4355 : 4'b1110;
														assign node4355 = (inp[12]) ? 4'b1110 : 4'b1111;
												assign node4358 = (inp[12]) ? node4368 : node4359;
													assign node4359 = (inp[4]) ? node4365 : node4360;
														assign node4360 = (inp[7]) ? node4362 : 4'b1000;
															assign node4362 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node4365 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node4368 = (inp[4]) ? 4'b1101 : 4'b1111;
								assign node4371 = (inp[7]) ? node4469 : node4372;
									assign node4372 = (inp[9]) ? node4424 : node4373;
										assign node4373 = (inp[12]) ? node4397 : node4374;
											assign node4374 = (inp[4]) ? node4384 : node4375;
												assign node4375 = (inp[11]) ? node4377 : 4'b1101;
													assign node4377 = (inp[2]) ? node4379 : 4'b1001;
														assign node4379 = (inp[5]) ? 4'b1100 : node4380;
															assign node4380 = (inp[1]) ? 4'b1001 : 4'b1100;
												assign node4384 = (inp[15]) ? node4392 : node4385;
													assign node4385 = (inp[1]) ? node4387 : 4'b1011;
														assign node4387 = (inp[2]) ? node4389 : 4'b1111;
															assign node4389 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node4392 = (inp[1]) ? 4'b1110 : node4393;
														assign node4393 = (inp[2]) ? 4'b1110 : 4'b1011;
											assign node4397 = (inp[4]) ? node4411 : node4398;
												assign node4398 = (inp[2]) ? node4406 : node4399;
													assign node4399 = (inp[11]) ? 4'b1110 : node4400;
														assign node4400 = (inp[1]) ? node4402 : 4'b1011;
															assign node4402 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node4406 = (inp[15]) ? 4'b1111 : node4407;
														assign node4407 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node4411 = (inp[11]) ? node4419 : node4412;
													assign node4412 = (inp[2]) ? 4'b1101 : node4413;
														assign node4413 = (inp[1]) ? 4'b1101 : node4414;
															assign node4414 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node4419 = (inp[1]) ? 4'b1001 : node4420;
														assign node4420 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node4424 = (inp[4]) ? node4446 : node4425;
											assign node4425 = (inp[12]) ? node4437 : node4426;
												assign node4426 = (inp[2]) ? node4432 : node4427;
													assign node4427 = (inp[15]) ? node4429 : 4'b1101;
														assign node4429 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node4432 = (inp[11]) ? 4'b1000 : node4433;
														assign node4433 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node4437 = (inp[15]) ? node4441 : node4438;
													assign node4438 = (inp[5]) ? 4'b1110 : 4'b1011;
													assign node4441 = (inp[2]) ? 4'b1111 : node4442;
														assign node4442 = (inp[5]) ? 4'b1010 : 4'b1110;
											assign node4446 = (inp[12]) ? node4460 : node4447;
												assign node4447 = (inp[11]) ? node4453 : node4448;
													assign node4448 = (inp[1]) ? node4450 : 4'b1111;
														assign node4450 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node4453 = (inp[5]) ? node4457 : node4454;
														assign node4454 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node4457 = (inp[15]) ? 4'b1011 : 4'b1111;
												assign node4460 = (inp[2]) ? node4464 : node4461;
													assign node4461 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node4464 = (inp[11]) ? 4'b1101 : node4465;
														assign node4465 = (inp[1]) ? 4'b1001 : 4'b1101;
									assign node4469 = (inp[1]) ? node4503 : node4470;
										assign node4470 = (inp[2]) ? node4484 : node4471;
											assign node4471 = (inp[15]) ? node4475 : node4472;
												assign node4472 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node4475 = (inp[12]) ? node4481 : node4476;
													assign node4476 = (inp[4]) ? node4478 : 4'b1100;
														assign node4478 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node4481 = (inp[4]) ? 4'b1001 : 4'b1011;
											assign node4484 = (inp[4]) ? node4494 : node4485;
												assign node4485 = (inp[12]) ? node4489 : node4486;
													assign node4486 = (inp[15]) ? 4'b1000 : 4'b1101;
													assign node4489 = (inp[5]) ? 4'b1111 : node4490;
														assign node4490 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node4494 = (inp[12]) ? node4500 : node4495;
													assign node4495 = (inp[11]) ? 4'b1110 : node4496;
														assign node4496 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node4500 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node4503 = (inp[2]) ? node4521 : node4504;
											assign node4504 = (inp[4]) ? node4518 : node4505;
												assign node4505 = (inp[12]) ? node4513 : node4506;
													assign node4506 = (inp[15]) ? 4'b1001 : node4507;
														assign node4507 = (inp[5]) ? node4509 : 4'b1101;
															assign node4509 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node4513 = (inp[5]) ? 4'b1110 : node4514;
														assign node4514 = (inp[15]) ? 4'b1111 : 4'b1011;
												assign node4518 = (inp[12]) ? 4'b1101 : 4'b1111;
											assign node4521 = (inp[9]) ? node4529 : node4522;
												assign node4522 = (inp[4]) ? node4526 : node4523;
													assign node4523 = (inp[5]) ? 4'b1011 : 4'b1000;
													assign node4526 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node4529 = (inp[12]) ? node4533 : node4530;
													assign node4530 = (inp[15]) ? 4'b1101 : 4'b1000;
													assign node4533 = (inp[11]) ? 4'b1111 : 4'b1110;
					assign node4536 = (inp[0]) ? node5314 : node4537;
						assign node4537 = (inp[8]) ? node4967 : node4538;
							assign node4538 = (inp[1]) ? node4758 : node4539;
								assign node4539 = (inp[9]) ? node4653 : node4540;
									assign node4540 = (inp[12]) ? node4588 : node4541;
										assign node4541 = (inp[7]) ? node4565 : node4542;
											assign node4542 = (inp[15]) ? node4556 : node4543;
												assign node4543 = (inp[2]) ? 4'b1000 : node4544;
													assign node4544 = (inp[11]) ? node4550 : node4545;
														assign node4545 = (inp[13]) ? 4'b1001 : node4546;
															assign node4546 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node4550 = (inp[13]) ? 4'b1001 : node4551;
															assign node4551 = (inp[5]) ? 4'b1100 : 4'b1000;
												assign node4556 = (inp[4]) ? node4560 : node4557;
													assign node4557 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node4560 = (inp[13]) ? 4'b1100 : node4561;
														assign node4561 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node4565 = (inp[15]) ? node4577 : node4566;
												assign node4566 = (inp[5]) ? node4572 : node4567;
													assign node4567 = (inp[2]) ? node4569 : 4'b1110;
														assign node4569 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node4572 = (inp[2]) ? node4574 : 4'b1010;
														assign node4574 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node4577 = (inp[4]) ? node4581 : node4578;
													assign node4578 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node4581 = (inp[11]) ? node4583 : 4'b1011;
														assign node4583 = (inp[5]) ? 4'b1110 : node4584;
															assign node4584 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node4588 = (inp[7]) ? node4630 : node4589;
											assign node4589 = (inp[5]) ? node4607 : node4590;
												assign node4590 = (inp[15]) ? node4596 : node4591;
													assign node4591 = (inp[13]) ? node4593 : 4'b1010;
														assign node4593 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node4596 = (inp[4]) ? node4600 : node4597;
														assign node4597 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node4600 = (inp[13]) ? node4604 : node4601;
															assign node4601 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node4604 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node4607 = (inp[11]) ? node4621 : node4608;
													assign node4608 = (inp[13]) ? node4616 : node4609;
														assign node4609 = (inp[15]) ? 4'b1110 : node4610;
															assign node4610 = (inp[2]) ? node4612 : 4'b1110;
																assign node4612 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node4616 = (inp[15]) ? 4'b1001 : node4617;
															assign node4617 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node4621 = (inp[2]) ? 4'b1011 : node4622;
														assign node4622 = (inp[4]) ? node4624 : 4'b1111;
															assign node4624 = (inp[13]) ? node4626 : 4'b1111;
																assign node4626 = (inp[15]) ? 4'b1111 : 4'b1010;
											assign node4630 = (inp[4]) ? node4640 : node4631;
												assign node4631 = (inp[15]) ? node4633 : 4'b1000;
													assign node4633 = (inp[11]) ? node4637 : node4634;
														assign node4634 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node4637 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node4640 = (inp[11]) ? node4646 : node4641;
													assign node4641 = (inp[2]) ? 4'b1101 : node4642;
														assign node4642 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node4646 = (inp[2]) ? 4'b1001 : node4647;
														assign node4647 = (inp[13]) ? node4649 : 4'b1101;
															assign node4649 = (inp[15]) ? 4'b1101 : 4'b1001;
									assign node4653 = (inp[13]) ? node4701 : node4654;
										assign node4654 = (inp[7]) ? node4680 : node4655;
											assign node4655 = (inp[12]) ? node4669 : node4656;
												assign node4656 = (inp[4]) ? node4662 : node4657;
													assign node4657 = (inp[2]) ? 4'b1100 : node4658;
														assign node4658 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node4662 = (inp[5]) ? 4'b1100 : node4663;
														assign node4663 = (inp[11]) ? 4'b1001 : node4664;
															assign node4664 = (inp[2]) ? 4'b1101 : 4'b1000;
												assign node4669 = (inp[11]) ? node4675 : node4670;
													assign node4670 = (inp[5]) ? node4672 : 4'b1010;
														assign node4672 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node4675 = (inp[2]) ? 4'b1011 : node4676;
														assign node4676 = (inp[5]) ? 4'b1110 : 4'b1111;
											assign node4680 = (inp[2]) ? node4690 : node4681;
												assign node4681 = (inp[5]) ? 4'b1110 : node4682;
													assign node4682 = (inp[15]) ? node4684 : 4'b1000;
														assign node4684 = (inp[11]) ? 4'b1010 : node4685;
															assign node4685 = (inp[4]) ? 4'b1010 : 4'b1100;
												assign node4690 = (inp[15]) ? node4698 : node4691;
													assign node4691 = (inp[11]) ? 4'b1100 : node4692;
														assign node4692 = (inp[5]) ? node4694 : 4'b1001;
															assign node4694 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node4698 = (inp[11]) ? 4'b1000 : 4'b1110;
										assign node4701 = (inp[2]) ? node4727 : node4702;
											assign node4702 = (inp[5]) ? node4716 : node4703;
												assign node4703 = (inp[11]) ? node4709 : node4704;
													assign node4704 = (inp[7]) ? node4706 : 4'b1110;
														assign node4706 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node4709 = (inp[4]) ? node4713 : node4710;
														assign node4710 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node4713 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node4716 = (inp[12]) ? node4724 : node4717;
													assign node4717 = (inp[11]) ? 4'b1011 : node4718;
														assign node4718 = (inp[4]) ? 4'b1001 : node4719;
															assign node4719 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node4724 = (inp[15]) ? 4'b1000 : 4'b1001;
											assign node4727 = (inp[5]) ? node4741 : node4728;
												assign node4728 = (inp[4]) ? node4736 : node4729;
													assign node4729 = (inp[15]) ? node4733 : node4730;
														assign node4730 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node4733 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node4736 = (inp[12]) ? 4'b1011 : node4737;
														assign node4737 = (inp[15]) ? 4'b1100 : 4'b1010;
												assign node4741 = (inp[4]) ? node4751 : node4742;
													assign node4742 = (inp[7]) ? node4746 : node4743;
														assign node4743 = (inp[12]) ? 4'b1000 : 4'b1101;
														assign node4746 = (inp[15]) ? node4748 : 4'b1110;
															assign node4748 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node4751 = (inp[7]) ? node4753 : 4'b1110;
														assign node4753 = (inp[12]) ? node4755 : 4'b1110;
															assign node4755 = (inp[15]) ? 4'b1101 : 4'b1100;
								assign node4758 = (inp[7]) ? node4862 : node4759;
									assign node4759 = (inp[12]) ? node4805 : node4760;
										assign node4760 = (inp[15]) ? node4784 : node4761;
											assign node4761 = (inp[9]) ? node4775 : node4762;
												assign node4762 = (inp[13]) ? node4770 : node4763;
													assign node4763 = (inp[2]) ? node4765 : 4'b1001;
														assign node4765 = (inp[5]) ? node4767 : 4'b1101;
															assign node4767 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node4770 = (inp[4]) ? node4772 : 4'b1101;
														assign node4772 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node4775 = (inp[11]) ? node4781 : node4776;
													assign node4776 = (inp[2]) ? node4778 : 4'b1000;
														assign node4778 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node4781 = (inp[5]) ? 4'b1100 : 4'b1101;
											assign node4784 = (inp[4]) ? node4794 : node4785;
												assign node4785 = (inp[2]) ? node4789 : node4786;
													assign node4786 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node4789 = (inp[13]) ? 4'b1011 : node4790;
														assign node4790 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node4794 = (inp[2]) ? node4798 : node4795;
													assign node4795 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node4798 = (inp[13]) ? node4802 : node4799;
														assign node4799 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node4802 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node4805 = (inp[15]) ? node4843 : node4806;
											assign node4806 = (inp[9]) ? node4824 : node4807;
												assign node4807 = (inp[11]) ? node4813 : node4808;
													assign node4808 = (inp[5]) ? node4810 : 4'b1110;
														assign node4810 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node4813 = (inp[5]) ? node4815 : 4'b1010;
														assign node4815 = (inp[2]) ? node4817 : 4'b1110;
															assign node4817 = (inp[4]) ? node4821 : node4818;
																assign node4818 = (inp[13]) ? 4'b1011 : 4'b1110;
																assign node4821 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node4824 = (inp[5]) ? node4830 : node4825;
													assign node4825 = (inp[2]) ? node4827 : 4'b1111;
														assign node4827 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node4830 = (inp[2]) ? node4838 : node4831;
														assign node4831 = (inp[11]) ? node4835 : node4832;
															assign node4832 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node4835 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node4838 = (inp[4]) ? 4'b1111 : node4839;
															assign node4839 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node4843 = (inp[4]) ? node4855 : node4844;
												assign node4844 = (inp[2]) ? node4852 : node4845;
													assign node4845 = (inp[13]) ? node4849 : node4846;
														assign node4846 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node4849 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node4852 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node4855 = (inp[11]) ? node4857 : 4'b1010;
													assign node4857 = (inp[5]) ? 4'b1111 : node4858;
														assign node4858 = (inp[2]) ? 4'b1111 : 4'b1010;
									assign node4862 = (inp[12]) ? node4912 : node4863;
										assign node4863 = (inp[15]) ? node4885 : node4864;
											assign node4864 = (inp[9]) ? node4874 : node4865;
												assign node4865 = (inp[11]) ? node4871 : node4866;
													assign node4866 = (inp[2]) ? 4'b1110 : node4867;
														assign node4867 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node4871 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node4874 = (inp[11]) ? node4876 : 4'b1010;
													assign node4876 = (inp[5]) ? node4878 : 4'b1010;
														assign node4878 = (inp[4]) ? 4'b1011 : node4879;
															assign node4879 = (inp[13]) ? node4881 : 4'b1111;
																assign node4881 = (inp[2]) ? 4'b1010 : 4'b1111;
											assign node4885 = (inp[4]) ? node4903 : node4886;
												assign node4886 = (inp[13]) ? node4890 : node4887;
													assign node4887 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node4890 = (inp[9]) ? 4'b1001 : node4891;
														assign node4891 = (inp[2]) ? node4895 : node4892;
															assign node4892 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node4895 = (inp[5]) ? node4899 : node4896;
																assign node4896 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node4899 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node4903 = (inp[11]) ? node4909 : node4904;
													assign node4904 = (inp[13]) ? node4906 : 4'b1011;
														assign node4906 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node4909 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node4912 = (inp[15]) ? node4942 : node4913;
											assign node4913 = (inp[13]) ? node4931 : node4914;
												assign node4914 = (inp[2]) ? node4924 : node4915;
													assign node4915 = (inp[4]) ? node4919 : node4916;
														assign node4916 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node4919 = (inp[9]) ? 4'b1001 : node4920;
															assign node4920 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node4924 = (inp[4]) ? 4'b1101 : node4925;
														assign node4925 = (inp[9]) ? node4927 : 4'b1001;
															assign node4927 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4931 = (inp[9]) ? node4939 : node4932;
													assign node4932 = (inp[2]) ? node4936 : node4933;
														assign node4933 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node4936 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node4939 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node4942 = (inp[4]) ? node4958 : node4943;
												assign node4943 = (inp[5]) ? node4951 : node4944;
													assign node4944 = (inp[2]) ? node4948 : node4945;
														assign node4945 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node4948 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node4951 = (inp[2]) ? node4955 : node4952;
														assign node4952 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node4955 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node4958 = (inp[11]) ? node4962 : node4959;
													assign node4959 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node4962 = (inp[2]) ? node4964 : 4'b1001;
														assign node4964 = (inp[9]) ? 4'b1001 : 4'b1000;
							assign node4967 = (inp[7]) ? node5171 : node4968;
								assign node4968 = (inp[5]) ? node5074 : node4969;
									assign node4969 = (inp[2]) ? node5029 : node4970;
										assign node4970 = (inp[11]) ? node4994 : node4971;
											assign node4971 = (inp[15]) ? node4983 : node4972;
												assign node4972 = (inp[1]) ? node4980 : node4973;
													assign node4973 = (inp[12]) ? node4977 : node4974;
														assign node4974 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node4977 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node4980 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node4983 = (inp[1]) ? node4989 : node4984;
													assign node4984 = (inp[13]) ? 4'b1110 : node4985;
														assign node4985 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node4989 = (inp[4]) ? node4991 : 4'b1101;
														assign node4991 = (inp[12]) ? 4'b1001 : 4'b1010;
											assign node4994 = (inp[13]) ? node5010 : node4995;
												assign node4995 = (inp[12]) ? node5003 : node4996;
													assign node4996 = (inp[4]) ? node5000 : node4997;
														assign node4997 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node5000 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node5003 = (inp[4]) ? node5005 : 4'b1111;
														assign node5005 = (inp[15]) ? node5007 : 4'b1001;
															assign node5007 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node5010 = (inp[9]) ? node5022 : node5011;
													assign node5011 = (inp[12]) ? node5017 : node5012;
														assign node5012 = (inp[15]) ? 4'b1100 : node5013;
															assign node5013 = (inp[1]) ? 4'b1111 : 4'b1001;
														assign node5017 = (inp[15]) ? node5019 : 4'b1100;
															assign node5019 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node5022 = (inp[12]) ? node5024 : 4'b1000;
														assign node5024 = (inp[15]) ? node5026 : 4'b1100;
															assign node5026 = (inp[1]) ? 4'b1000 : 4'b1100;
										assign node5029 = (inp[11]) ? node5055 : node5030;
											assign node5030 = (inp[4]) ? node5038 : node5031;
												assign node5031 = (inp[12]) ? node5033 : 4'b1000;
													assign node5033 = (inp[13]) ? 4'b1011 : node5034;
														assign node5034 = (inp[15]) ? 4'b1111 : 4'b1011;
												assign node5038 = (inp[12]) ? node5048 : node5039;
													assign node5039 = (inp[9]) ? node5045 : node5040;
														assign node5040 = (inp[15]) ? node5042 : 4'b1011;
															assign node5042 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node5045 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node5048 = (inp[9]) ? node5050 : 4'b1101;
														assign node5050 = (inp[15]) ? node5052 : 4'b1000;
															assign node5052 = (inp[1]) ? 4'b1101 : 4'b1001;
											assign node5055 = (inp[1]) ? node5067 : node5056;
												assign node5056 = (inp[15]) ? node5062 : node5057;
													assign node5057 = (inp[12]) ? node5059 : 4'b1101;
														assign node5059 = (inp[4]) ? 4'b1101 : 4'b1111;
													assign node5062 = (inp[4]) ? 4'b1010 : node5063;
														assign node5063 = (inp[12]) ? 4'b1011 : 4'b1101;
												assign node5067 = (inp[12]) ? node5069 : 4'b1001;
													assign node5069 = (inp[13]) ? 4'b1110 : node5070;
														assign node5070 = (inp[4]) ? 4'b1000 : 4'b1010;
									assign node5074 = (inp[11]) ? node5138 : node5075;
										assign node5075 = (inp[1]) ? node5109 : node5076;
											assign node5076 = (inp[2]) ? node5092 : node5077;
												assign node5077 = (inp[15]) ? node5085 : node5078;
													assign node5078 = (inp[12]) ? node5082 : node5079;
														assign node5079 = (inp[4]) ? 4'b1111 : 4'b1101;
														assign node5082 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node5085 = (inp[12]) ? node5089 : node5086;
														assign node5086 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node5089 = (inp[13]) ? 4'b1000 : 4'b1011;
												assign node5092 = (inp[13]) ? node5100 : node5093;
													assign node5093 = (inp[4]) ? node5097 : node5094;
														assign node5094 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node5097 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node5100 = (inp[15]) ? node5104 : node5101;
														assign node5101 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node5104 = (inp[4]) ? 4'b1111 : node5105;
															assign node5105 = (inp[12]) ? 4'b1111 : 4'b1101;
											assign node5109 = (inp[12]) ? node5119 : node5110;
												assign node5110 = (inp[4]) ? 4'b1010 : node5111;
													assign node5111 = (inp[15]) ? node5115 : node5112;
														assign node5112 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node5115 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node5119 = (inp[4]) ? node5133 : node5120;
													assign node5120 = (inp[2]) ? node5124 : node5121;
														assign node5121 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node5124 = (inp[9]) ? node5126 : 4'b1010;
															assign node5126 = (inp[13]) ? node5130 : node5127;
																assign node5127 = (inp[15]) ? 4'b1010 : 4'b1011;
																assign node5130 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node5133 = (inp[13]) ? 4'b1001 : node5134;
														assign node5134 = (inp[2]) ? 4'b1000 : 4'b1100;
										assign node5138 = (inp[12]) ? node5154 : node5139;
											assign node5139 = (inp[4]) ? node5147 : node5140;
												assign node5140 = (inp[9]) ? 4'b1000 : node5141;
													assign node5141 = (inp[2]) ? 4'b1101 : node5142;
														assign node5142 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node5147 = (inp[1]) ? node5149 : 4'b1011;
													assign node5149 = (inp[2]) ? 4'b1111 : node5150;
														assign node5150 = (inp[15]) ? 4'b1111 : 4'b1010;
											assign node5154 = (inp[4]) ? node5164 : node5155;
												assign node5155 = (inp[1]) ? node5161 : node5156;
													assign node5156 = (inp[2]) ? node5158 : 4'b1011;
														assign node5158 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node5161 = (inp[2]) ? 4'b1011 : 4'b1110;
												assign node5164 = (inp[15]) ? 4'b1001 : node5165;
													assign node5165 = (inp[13]) ? 4'b1100 : node5166;
														assign node5166 = (inp[1]) ? 4'b1100 : 4'b1101;
								assign node5171 = (inp[1]) ? node5243 : node5172;
									assign node5172 = (inp[2]) ? node5210 : node5173;
										assign node5173 = (inp[5]) ? node5197 : node5174;
											assign node5174 = (inp[12]) ? node5186 : node5175;
												assign node5175 = (inp[4]) ? 4'b1011 : node5176;
													assign node5176 = (inp[9]) ? 4'b1001 : node5177;
														assign node5177 = (inp[11]) ? node5179 : 4'b1001;
															assign node5179 = (inp[13]) ? 4'b1000 : node5180;
																assign node5180 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node5186 = (inp[4]) ? node5192 : node5187;
													assign node5187 = (inp[15]) ? node5189 : 4'b1111;
														assign node5189 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node5192 = (inp[11]) ? node5194 : 4'b1000;
														assign node5194 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node5197 = (inp[9]) ? node5205 : node5198;
												assign node5198 = (inp[12]) ? node5202 : node5199;
													assign node5199 = (inp[4]) ? 4'b1010 : 4'b1000;
													assign node5202 = (inp[4]) ? 4'b1000 : 4'b1011;
												assign node5205 = (inp[13]) ? 4'b1000 : node5206;
													assign node5206 = (inp[4]) ? 4'b1001 : 4'b1000;
										assign node5210 = (inp[15]) ? node5226 : node5211;
											assign node5211 = (inp[12]) ? node5221 : node5212;
												assign node5212 = (inp[4]) ? 4'b1110 : node5213;
													assign node5213 = (inp[9]) ? node5217 : node5214;
														assign node5214 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node5217 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node5221 = (inp[13]) ? node5223 : 4'b1101;
													assign node5223 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node5226 = (inp[5]) ? node5236 : node5227;
												assign node5227 = (inp[4]) ? node5231 : node5228;
													assign node5228 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node5231 = (inp[12]) ? node5233 : 4'b1111;
														assign node5233 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node5236 = (inp[12]) ? node5240 : node5237;
													assign node5237 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node5240 = (inp[4]) ? 4'b1101 : 4'b1111;
									assign node5243 = (inp[2]) ? node5275 : node5244;
										assign node5244 = (inp[5]) ? node5264 : node5245;
											assign node5245 = (inp[15]) ? node5251 : node5246;
												assign node5246 = (inp[4]) ? node5248 : 4'b1011;
													assign node5248 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node5251 = (inp[13]) ? node5261 : node5252;
													assign node5252 = (inp[11]) ? 4'b1111 : node5253;
														assign node5253 = (inp[4]) ? node5257 : node5254;
															assign node5254 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node5257 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node5261 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node5264 = (inp[4]) ? node5272 : node5265;
												assign node5265 = (inp[11]) ? node5269 : node5266;
													assign node5266 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node5269 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node5272 = (inp[12]) ? 4'b1101 : 4'b1111;
										assign node5275 = (inp[4]) ? node5291 : node5276;
											assign node5276 = (inp[12]) ? node5282 : node5277;
												assign node5277 = (inp[9]) ? node5279 : 4'b1101;
													assign node5279 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node5282 = (inp[15]) ? node5288 : node5283;
													assign node5283 = (inp[5]) ? 4'b1011 : node5284;
														assign node5284 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node5288 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node5291 = (inp[12]) ? node5301 : node5292;
												assign node5292 = (inp[13]) ? 4'b1011 : node5293;
													assign node5293 = (inp[15]) ? node5297 : node5294;
														assign node5294 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node5297 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node5301 = (inp[13]) ? 4'b1001 : node5302;
													assign node5302 = (inp[5]) ? node5308 : node5303;
														assign node5303 = (inp[9]) ? 4'b1001 : node5304;
															assign node5304 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node5308 = (inp[15]) ? node5310 : 4'b1000;
															assign node5310 = (inp[9]) ? 4'b1000 : 4'b1001;
						assign node5314 = (inp[8]) ? node5740 : node5315;
							assign node5315 = (inp[9]) ? node5535 : node5316;
								assign node5316 = (inp[7]) ? node5424 : node5317;
									assign node5317 = (inp[12]) ? node5365 : node5318;
										assign node5318 = (inp[4]) ? node5342 : node5319;
											assign node5319 = (inp[15]) ? node5329 : node5320;
												assign node5320 = (inp[2]) ? node5324 : node5321;
													assign node5321 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5324 = (inp[13]) ? node5326 : 4'b1100;
														assign node5326 = (inp[5]) ? 4'b1100 : 4'b1000;
												assign node5329 = (inp[2]) ? node5333 : node5330;
													assign node5330 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node5333 = (inp[1]) ? 4'b1010 : node5334;
														assign node5334 = (inp[13]) ? node5338 : node5335;
															assign node5335 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node5338 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node5342 = (inp[5]) ? node5352 : node5343;
												assign node5343 = (inp[11]) ? node5345 : 4'b1001;
													assign node5345 = (inp[13]) ? 4'b1100 : node5346;
														assign node5346 = (inp[15]) ? node5348 : 4'b1001;
															assign node5348 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node5352 = (inp[2]) ? node5362 : node5353;
													assign node5353 = (inp[1]) ? 4'b1000 : node5354;
														assign node5354 = (inp[11]) ? node5358 : node5355;
															assign node5355 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node5358 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node5362 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node5365 = (inp[4]) ? node5393 : node5366;
											assign node5366 = (inp[15]) ? node5380 : node5367;
												assign node5367 = (inp[13]) ? node5371 : node5368;
													assign node5368 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node5371 = (inp[2]) ? node5375 : node5372;
														assign node5372 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node5375 = (inp[1]) ? node5377 : 4'b1010;
															assign node5377 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node5380 = (inp[2]) ? node5388 : node5381;
													assign node5381 = (inp[13]) ? 4'b1000 : node5382;
														assign node5382 = (inp[1]) ? 4'b1101 : node5383;
															assign node5383 = (inp[5]) ? 4'b1000 : 4'b1101;
													assign node5388 = (inp[13]) ? 4'b1101 : node5389;
														assign node5389 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node5393 = (inp[15]) ? node5409 : node5394;
												assign node5394 = (inp[1]) ? node5402 : node5395;
													assign node5395 = (inp[2]) ? node5399 : node5396;
														assign node5396 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node5399 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node5402 = (inp[5]) ? node5406 : node5403;
														assign node5403 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node5406 = (inp[11]) ? 4'b1011 : 4'b1111;
												assign node5409 = (inp[5]) ? node5413 : node5410;
													assign node5410 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node5413 = (inp[13]) ? node5419 : node5414;
														assign node5414 = (inp[2]) ? 4'b1110 : node5415;
															assign node5415 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node5419 = (inp[2]) ? node5421 : 4'b1111;
															assign node5421 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node5424 = (inp[12]) ? node5474 : node5425;
										assign node5425 = (inp[15]) ? node5447 : node5426;
											assign node5426 = (inp[4]) ? node5438 : node5427;
												assign node5427 = (inp[1]) ? node5429 : 4'b1011;
													assign node5429 = (inp[5]) ? node5433 : node5430;
														assign node5430 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node5433 = (inp[11]) ? 4'b1011 : node5434;
															assign node5434 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node5438 = (inp[5]) ? node5444 : node5439;
													assign node5439 = (inp[1]) ? node5441 : 4'b1011;
														assign node5441 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node5444 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node5447 = (inp[4]) ? node5465 : node5448;
												assign node5448 = (inp[11]) ? node5456 : node5449;
													assign node5449 = (inp[5]) ? 4'b1101 : node5450;
														assign node5450 = (inp[2]) ? node5452 : 4'b1101;
															assign node5452 = (inp[1]) ? 4'b1000 : 4'b1101;
													assign node5456 = (inp[13]) ? node5460 : node5457;
														assign node5457 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node5460 = (inp[5]) ? 4'b1000 : node5461;
															assign node5461 = (inp[1]) ? 4'b1101 : 4'b1000;
												assign node5465 = (inp[5]) ? node5469 : node5466;
													assign node5466 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node5469 = (inp[1]) ? 4'b1111 : node5470;
														assign node5470 = (inp[11]) ? 4'b1010 : 4'b1110;
										assign node5474 = (inp[15]) ? node5510 : node5475;
											assign node5475 = (inp[1]) ? node5491 : node5476;
												assign node5476 = (inp[11]) ? node5484 : node5477;
													assign node5477 = (inp[4]) ? node5481 : node5478;
														assign node5478 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node5481 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node5484 = (inp[2]) ? node5486 : 4'b1101;
														assign node5486 = (inp[5]) ? 4'b1101 : node5487;
															assign node5487 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node5491 = (inp[2]) ? node5493 : 4'b1001;
													assign node5493 = (inp[5]) ? node5503 : node5494;
														assign node5494 = (inp[13]) ? node5500 : node5495;
															assign node5495 = (inp[4]) ? node5497 : 4'b1000;
																assign node5497 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node5500 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node5503 = (inp[13]) ? node5507 : node5504;
															assign node5504 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node5507 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node5510 = (inp[4]) ? node5524 : node5511;
												assign node5511 = (inp[2]) ? node5515 : node5512;
													assign node5512 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node5515 = (inp[11]) ? node5519 : node5516;
														assign node5516 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node5519 = (inp[1]) ? node5521 : 4'b1010;
															assign node5521 = (inp[5]) ? 4'b1111 : 4'b1011;
												assign node5524 = (inp[13]) ? node5532 : node5525;
													assign node5525 = (inp[11]) ? 4'b1000 : node5526;
														assign node5526 = (inp[5]) ? node5528 : 4'b1100;
															assign node5528 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node5532 = (inp[1]) ? 4'b1101 : 4'b1100;
								assign node5535 = (inp[13]) ? node5641 : node5536;
									assign node5536 = (inp[1]) ? node5582 : node5537;
										assign node5537 = (inp[4]) ? node5563 : node5538;
											assign node5538 = (inp[7]) ? node5550 : node5539;
												assign node5539 = (inp[2]) ? node5543 : node5540;
													assign node5540 = (inp[11]) ? 4'b1000 : 4'b1100;
													assign node5543 = (inp[5]) ? node5547 : node5544;
														assign node5544 = (inp[12]) ? 4'b1001 : 4'b1110;
														assign node5547 = (inp[11]) ? 4'b1001 : 4'b1101;
												assign node5550 = (inp[15]) ? node5554 : node5551;
													assign node5551 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node5554 = (inp[12]) ? node5558 : node5555;
														assign node5555 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node5558 = (inp[11]) ? node5560 : 4'b1011;
															assign node5560 = (inp[2]) ? 4'b1011 : 4'b1110;
											assign node5563 = (inp[12]) ? node5571 : node5564;
												assign node5564 = (inp[2]) ? node5568 : node5565;
													assign node5565 = (inp[5]) ? 4'b1111 : 4'b1010;
													assign node5568 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node5571 = (inp[7]) ? node5577 : node5572;
													assign node5572 = (inp[11]) ? 4'b1111 : node5573;
														assign node5573 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node5577 = (inp[15]) ? node5579 : 4'b1000;
														assign node5579 = (inp[11]) ? 4'b1001 : 4'b1101;
										assign node5582 = (inp[2]) ? node5612 : node5583;
											assign node5583 = (inp[12]) ? node5601 : node5584;
												assign node5584 = (inp[15]) ? node5590 : node5585;
													assign node5585 = (inp[7]) ? 4'b1010 : node5586;
														assign node5586 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node5590 = (inp[7]) ? node5596 : node5591;
														assign node5591 = (inp[5]) ? 4'b1011 : node5592;
															assign node5592 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node5596 = (inp[5]) ? 4'b1100 : node5597;
															assign node5597 = (inp[4]) ? 4'b1011 : 4'b1001;
												assign node5601 = (inp[7]) ? node5607 : node5602;
													assign node5602 = (inp[5]) ? node5604 : 4'b1110;
														assign node5604 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node5607 = (inp[15]) ? node5609 : 4'b1101;
														assign node5609 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node5612 = (inp[12]) ? node5624 : node5613;
												assign node5613 = (inp[7]) ? node5619 : node5614;
													assign node5614 = (inp[15]) ? node5616 : 4'b1101;
														assign node5616 = (inp[4]) ? 4'b1000 : 4'b1111;
													assign node5619 = (inp[11]) ? 4'b1110 : node5620;
														assign node5620 = (inp[4]) ? 4'b1111 : 4'b1100;
												assign node5624 = (inp[7]) ? node5632 : node5625;
													assign node5625 = (inp[15]) ? 4'b1000 : node5626;
														assign node5626 = (inp[5]) ? node5628 : 4'b1111;
															assign node5628 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node5632 = (inp[4]) ? node5636 : node5633;
														assign node5633 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node5636 = (inp[15]) ? 4'b1100 : node5637;
															assign node5637 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node5641 = (inp[2]) ? node5691 : node5642;
										assign node5642 = (inp[11]) ? node5664 : node5643;
											assign node5643 = (inp[5]) ? node5657 : node5644;
												assign node5644 = (inp[7]) ? node5654 : node5645;
													assign node5645 = (inp[12]) ? node5649 : node5646;
														assign node5646 = (inp[1]) ? 4'b1110 : 4'b1000;
														assign node5649 = (inp[15]) ? node5651 : 4'b1110;
															assign node5651 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node5654 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node5657 = (inp[4]) ? node5659 : 4'b1111;
													assign node5659 = (inp[15]) ? 4'b1110 : node5660;
														assign node5660 = (inp[7]) ? 4'b1110 : 4'b1101;
											assign node5664 = (inp[5]) ? node5676 : node5665;
												assign node5665 = (inp[12]) ? node5669 : node5666;
													assign node5666 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node5669 = (inp[7]) ? node5673 : node5670;
														assign node5670 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node5673 = (inp[15]) ? 4'b1110 : 4'b1101;
												assign node5676 = (inp[12]) ? node5680 : node5677;
													assign node5677 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node5680 = (inp[7]) ? node5682 : 4'b1001;
														assign node5682 = (inp[15]) ? node5688 : node5683;
															assign node5683 = (inp[1]) ? 4'b1001 : node5684;
																assign node5684 = (inp[4]) ? 4'b1001 : 4'b1100;
															assign node5688 = (inp[1]) ? 4'b1100 : 4'b1000;
										assign node5691 = (inp[1]) ? node5717 : node5692;
											assign node5692 = (inp[12]) ? node5710 : node5693;
												assign node5693 = (inp[5]) ? node5703 : node5694;
													assign node5694 = (inp[4]) ? node5698 : node5695;
														assign node5695 = (inp[15]) ? 4'b1100 : 4'b1011;
														assign node5698 = (inp[7]) ? node5700 : 4'b1000;
															assign node5700 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node5703 = (inp[4]) ? node5705 : 4'b1110;
														assign node5705 = (inp[7]) ? 4'b1111 : node5706;
															assign node5706 = (inp[15]) ? 4'b1000 : 4'b1101;
												assign node5710 = (inp[11]) ? node5712 : 4'b1001;
													assign node5712 = (inp[5]) ? node5714 : 4'b1011;
														assign node5714 = (inp[15]) ? 4'b1010 : 4'b1111;
											assign node5717 = (inp[15]) ? node5729 : node5718;
												assign node5718 = (inp[12]) ? node5724 : node5719;
													assign node5719 = (inp[11]) ? 4'b1010 : node5720;
														assign node5720 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node5724 = (inp[11]) ? 4'b1100 : node5725;
														assign node5725 = (inp[7]) ? 4'b1000 : 4'b1010;
												assign node5729 = (inp[12]) ? node5735 : node5730;
													assign node5730 = (inp[11]) ? 4'b1100 : node5731;
														assign node5731 = (inp[4]) ? 4'b1010 : 4'b1100;
													assign node5735 = (inp[7]) ? node5737 : 4'b1010;
														assign node5737 = (inp[4]) ? 4'b1000 : 4'b1010;
							assign node5740 = (inp[7]) ? node5922 : node5741;
								assign node5741 = (inp[2]) ? node5829 : node5742;
									assign node5742 = (inp[1]) ? node5788 : node5743;
										assign node5743 = (inp[15]) ? node5765 : node5744;
											assign node5744 = (inp[5]) ? node5756 : node5745;
												assign node5745 = (inp[12]) ? node5753 : node5746;
													assign node5746 = (inp[4]) ? 4'b1010 : node5747;
														assign node5747 = (inp[11]) ? node5749 : 4'b1000;
															assign node5749 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node5753 = (inp[13]) ? 4'b1001 : 4'b1011;
												assign node5756 = (inp[12]) ? node5762 : node5757;
													assign node5757 = (inp[9]) ? 4'b1101 : node5758;
														assign node5758 = (inp[11]) ? 4'b1100 : 4'b1110;
													assign node5762 = (inp[4]) ? 4'b1101 : 4'b1010;
											assign node5765 = (inp[5]) ? node5773 : node5766;
												assign node5766 = (inp[13]) ? 4'b1111 : node5767;
													assign node5767 = (inp[12]) ? node5769 : 4'b1000;
														assign node5769 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node5773 = (inp[9]) ? node5777 : node5774;
													assign node5774 = (inp[12]) ? 4'b1001 : 4'b1011;
													assign node5777 = (inp[13]) ? node5779 : 4'b1010;
														assign node5779 = (inp[12]) ? node5785 : node5780;
															assign node5780 = (inp[4]) ? 4'b1010 : node5781;
																assign node5781 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node5785 = (inp[11]) ? 4'b1011 : 4'b1001;
										assign node5788 = (inp[13]) ? node5804 : node5789;
											assign node5789 = (inp[4]) ? node5797 : node5790;
												assign node5790 = (inp[12]) ? node5792 : 4'b1100;
													assign node5792 = (inp[5]) ? 4'b1110 : node5793;
														assign node5793 = (inp[15]) ? 4'b1011 : 4'b1110;
												assign node5797 = (inp[12]) ? node5799 : 4'b1111;
													assign node5799 = (inp[5]) ? node5801 : 4'b1101;
														assign node5801 = (inp[9]) ? 4'b1000 : 4'b1101;
											assign node5804 = (inp[4]) ? node5816 : node5805;
												assign node5805 = (inp[12]) ? node5813 : node5806;
													assign node5806 = (inp[11]) ? 4'b1101 : node5807;
														assign node5807 = (inp[5]) ? node5809 : 4'b1100;
															assign node5809 = (inp[9]) ? 4'b1001 : 4'b1100;
													assign node5813 = (inp[9]) ? 4'b1011 : 4'b1110;
												assign node5816 = (inp[12]) ? node5820 : node5817;
													assign node5817 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node5820 = (inp[11]) ? 4'b1000 : node5821;
														assign node5821 = (inp[9]) ? 4'b1100 : node5822;
															assign node5822 = (inp[15]) ? node5824 : 4'b1100;
																assign node5824 = (inp[5]) ? 4'b1100 : 4'b1000;
									assign node5829 = (inp[1]) ? node5875 : node5830;
										assign node5830 = (inp[15]) ? node5854 : node5831;
											assign node5831 = (inp[5]) ? node5845 : node5832;
												assign node5832 = (inp[13]) ? node5838 : node5833;
													assign node5833 = (inp[11]) ? node5835 : 4'b1100;
														assign node5835 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node5838 = (inp[4]) ? node5842 : node5839;
														assign node5839 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node5842 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node5845 = (inp[12]) ? node5851 : node5846;
													assign node5846 = (inp[4]) ? 4'b1010 : node5847;
														assign node5847 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node5851 = (inp[4]) ? 4'b1001 : 4'b1111;
											assign node5854 = (inp[5]) ? node5864 : node5855;
												assign node5855 = (inp[12]) ? node5859 : node5856;
													assign node5856 = (inp[11]) ? 4'b1101 : 4'b1011;
													assign node5859 = (inp[4]) ? node5861 : 4'b1010;
														assign node5861 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node5864 = (inp[13]) ? node5870 : node5865;
													assign node5865 = (inp[4]) ? node5867 : 4'b1101;
														assign node5867 = (inp[12]) ? 4'b1101 : 4'b1110;
													assign node5870 = (inp[12]) ? 4'b1100 : node5871;
														assign node5871 = (inp[11]) ? 4'b1100 : 4'b1110;
										assign node5875 = (inp[5]) ? node5903 : node5876;
											assign node5876 = (inp[15]) ? node5892 : node5877;
												assign node5877 = (inp[9]) ? node5885 : node5878;
													assign node5878 = (inp[12]) ? node5882 : node5879;
														assign node5879 = (inp[13]) ? 4'b1010 : 4'b1000;
														assign node5882 = (inp[11]) ? 4'b1011 : 4'b1001;
													assign node5885 = (inp[13]) ? node5887 : 4'b1001;
														assign node5887 = (inp[11]) ? 4'b1001 : node5888;
															assign node5888 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node5892 = (inp[12]) ? node5898 : node5893;
													assign node5893 = (inp[4]) ? 4'b1110 : node5894;
														assign node5894 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5898 = (inp[4]) ? 4'b1101 : node5899;
														assign node5899 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node5903 = (inp[15]) ? node5915 : node5904;
												assign node5904 = (inp[12]) ? node5912 : node5905;
													assign node5905 = (inp[4]) ? node5907 : 4'b1100;
														assign node5907 = (inp[11]) ? 4'b1110 : node5908;
															assign node5908 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node5912 = (inp[13]) ? 4'b1011 : 4'b1010;
												assign node5915 = (inp[4]) ? node5919 : node5916;
													assign node5916 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5919 = (inp[12]) ? 4'b1000 : 4'b1011;
								assign node5922 = (inp[13]) ? node6008 : node5923;
									assign node5923 = (inp[5]) ? node5971 : node5924;
										assign node5924 = (inp[15]) ? node5944 : node5925;
											assign node5925 = (inp[2]) ? node5935 : node5926;
												assign node5926 = (inp[1]) ? node5932 : node5927;
													assign node5927 = (inp[12]) ? 4'b1110 : node5928;
														assign node5928 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node5932 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node5935 = (inp[4]) ? node5939 : node5936;
													assign node5936 = (inp[1]) ? 4'b1110 : 4'b1100;
													assign node5939 = (inp[1]) ? node5941 : 4'b1100;
														assign node5941 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node5944 = (inp[11]) ? node5958 : node5945;
												assign node5945 = (inp[2]) ? node5951 : node5946;
													assign node5946 = (inp[12]) ? 4'b1110 : node5947;
														assign node5947 = (inp[4]) ? 4'b1111 : 4'b1101;
													assign node5951 = (inp[4]) ? node5955 : node5952;
														assign node5952 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node5955 = (inp[12]) ? 4'b1101 : 4'b1110;
												assign node5958 = (inp[2]) ? node5966 : node5959;
													assign node5959 = (inp[1]) ? 4'b1100 : node5960;
														assign node5960 = (inp[12]) ? 4'b1010 : node5961;
															assign node5961 = (inp[9]) ? 4'b1010 : 4'b1000;
													assign node5966 = (inp[12]) ? 4'b1111 : node5967;
														assign node5967 = (inp[9]) ? 4'b1010 : 4'b1100;
										assign node5971 = (inp[12]) ? node5989 : node5972;
											assign node5972 = (inp[4]) ? node5978 : node5973;
												assign node5973 = (inp[11]) ? 4'b1000 : node5974;
													assign node5974 = (inp[2]) ? 4'b1000 : 4'b1101;
												assign node5978 = (inp[15]) ? node5982 : node5979;
													assign node5979 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node5982 = (inp[9]) ? 4'b1110 : node5983;
														assign node5983 = (inp[1]) ? 4'b1111 : node5984;
															assign node5984 = (inp[2]) ? 4'b1111 : 4'b1010;
											assign node5989 = (inp[4]) ? node5995 : node5990;
												assign node5990 = (inp[2]) ? 4'b1010 : node5991;
													assign node5991 = (inp[11]) ? 4'b1011 : 4'b1111;
												assign node5995 = (inp[11]) ? node6001 : node5996;
													assign node5996 = (inp[1]) ? node5998 : 4'b1101;
														assign node5998 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node6001 = (inp[1]) ? node6003 : 4'b1000;
														assign node6003 = (inp[15]) ? 4'b1000 : node6004;
															assign node6004 = (inp[2]) ? 4'b1001 : 4'b1101;
									assign node6008 = (inp[11]) ? node6064 : node6009;
										assign node6009 = (inp[5]) ? node6041 : node6010;
											assign node6010 = (inp[9]) ? node6024 : node6011;
												assign node6011 = (inp[2]) ? node6013 : 4'b1110;
													assign node6013 = (inp[1]) ? node6019 : node6014;
														assign node6014 = (inp[12]) ? node6016 : 4'b1101;
															assign node6016 = (inp[4]) ? 4'b1101 : 4'b1010;
														assign node6019 = (inp[4]) ? 4'b1010 : node6020;
															assign node6020 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node6024 = (inp[4]) ? node6034 : node6025;
													assign node6025 = (inp[12]) ? node6031 : node6026;
														assign node6026 = (inp[1]) ? node6028 : 4'b1100;
															assign node6028 = (inp[15]) ? 4'b1001 : 4'b1100;
														assign node6031 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node6034 = (inp[2]) ? node6038 : node6035;
														assign node6035 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node6038 = (inp[1]) ? 4'b1000 : 4'b1100;
											assign node6041 = (inp[15]) ? node6047 : node6042;
												assign node6042 = (inp[2]) ? 4'b1010 : node6043;
													assign node6043 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node6047 = (inp[1]) ? node6053 : node6048;
													assign node6048 = (inp[2]) ? node6050 : 4'b1010;
														assign node6050 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node6053 = (inp[4]) ? node6059 : node6054;
														assign node6054 = (inp[12]) ? 4'b1010 : node6055;
															assign node6055 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node6059 = (inp[2]) ? 4'b1010 : node6060;
															assign node6060 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node6064 = (inp[4]) ? node6090 : node6065;
											assign node6065 = (inp[12]) ? node6081 : node6066;
												assign node6066 = (inp[15]) ? node6074 : node6067;
													assign node6067 = (inp[2]) ? node6071 : node6068;
														assign node6068 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6071 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node6074 = (inp[9]) ? node6076 : 4'b1100;
														assign node6076 = (inp[1]) ? 4'b1001 : node6077;
															assign node6077 = (inp[5]) ? 4'b1001 : 4'b1100;
												assign node6081 = (inp[9]) ? node6085 : node6082;
													assign node6082 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node6085 = (inp[2]) ? node6087 : 4'b1010;
														assign node6087 = (inp[1]) ? 4'b1010 : 4'b1110;
											assign node6090 = (inp[1]) ? node6098 : node6091;
												assign node6091 = (inp[2]) ? node6095 : node6092;
													assign node6092 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node6095 = (inp[12]) ? 4'b1100 : 4'b1111;
												assign node6098 = (inp[2]) ? 4'b1010 : 4'b1110;
			assign node6101 = (inp[14]) ? node8609 : node6102;
				assign node6102 = (inp[8]) ? node7404 : node6103;
					assign node6103 = (inp[13]) ? node6761 : node6104;
						assign node6104 = (inp[5]) ? node6432 : node6105;
							assign node6105 = (inp[12]) ? node6247 : node6106;
								assign node6106 = (inp[15]) ? node6146 : node6107;
									assign node6107 = (inp[7]) ? node6123 : node6108;
										assign node6108 = (inp[9]) ? node6114 : node6109;
											assign node6109 = (inp[11]) ? node6111 : 4'b1000;
												assign node6111 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node6114 = (inp[11]) ? node6120 : node6115;
												assign node6115 = (inp[1]) ? 4'b1001 : node6116;
													assign node6116 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node6120 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node6123 = (inp[9]) ? node6137 : node6124;
											assign node6124 = (inp[11]) ? node6132 : node6125;
												assign node6125 = (inp[2]) ? node6127 : 4'b1010;
													assign node6127 = (inp[1]) ? node6129 : 4'b1011;
														assign node6129 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node6132 = (inp[2]) ? node6134 : 4'b1011;
													assign node6134 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node6137 = (inp[11]) ? node6143 : node6138;
												assign node6138 = (inp[2]) ? node6140 : 4'b1011;
													assign node6140 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node6143 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node6146 = (inp[7]) ? node6204 : node6147;
										assign node6147 = (inp[4]) ? node6183 : node6148;
											assign node6148 = (inp[10]) ? node6166 : node6149;
												assign node6149 = (inp[0]) ? node6157 : node6150;
													assign node6150 = (inp[2]) ? node6152 : 4'b1010;
														assign node6152 = (inp[11]) ? 4'b1010 : node6153;
															assign node6153 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node6157 = (inp[1]) ? 4'b1011 : node6158;
														assign node6158 = (inp[2]) ? node6162 : node6159;
															assign node6159 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node6162 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node6166 = (inp[9]) ? node6172 : node6167;
													assign node6167 = (inp[1]) ? node6169 : 4'b1011;
														assign node6169 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node6172 = (inp[2]) ? node6174 : 4'b1010;
														assign node6174 = (inp[1]) ? 4'b1011 : node6175;
															assign node6175 = (inp[0]) ? node6179 : node6176;
																assign node6176 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node6179 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node6183 = (inp[1]) ? node6197 : node6184;
												assign node6184 = (inp[2]) ? node6190 : node6185;
													assign node6185 = (inp[11]) ? node6187 : 4'b1011;
														assign node6187 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node6190 = (inp[0]) ? 4'b1010 : node6191;
														assign node6191 = (inp[9]) ? 4'b1010 : node6192;
															assign node6192 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node6197 = (inp[2]) ? 4'b1110 : node6198;
													assign node6198 = (inp[0]) ? 4'b1111 : node6199;
														assign node6199 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node6204 = (inp[4]) ? node6224 : node6205;
											assign node6205 = (inp[1]) ? node6215 : node6206;
												assign node6206 = (inp[10]) ? node6208 : 4'b1101;
													assign node6208 = (inp[9]) ? node6210 : 4'b1101;
														assign node6210 = (inp[11]) ? 4'b1100 : node6211;
															assign node6211 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6215 = (inp[0]) ? 4'b1000 : node6216;
													assign node6216 = (inp[10]) ? node6218 : 4'b1000;
														assign node6218 = (inp[2]) ? node6220 : 4'b1001;
															assign node6220 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node6224 = (inp[2]) ? node6236 : node6225;
												assign node6225 = (inp[0]) ? 4'b1000 : node6226;
													assign node6226 = (inp[10]) ? 4'b1001 : node6227;
														assign node6227 = (inp[1]) ? node6229 : 4'b1001;
															assign node6229 = (inp[11]) ? node6231 : 4'b1000;
																assign node6231 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node6236 = (inp[10]) ? 4'b1001 : node6237;
													assign node6237 = (inp[1]) ? 4'b1001 : node6238;
														assign node6238 = (inp[0]) ? 4'b1000 : node6239;
															assign node6239 = (inp[9]) ? node6241 : 4'b1001;
																assign node6241 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node6247 = (inp[15]) ? node6347 : node6248;
									assign node6248 = (inp[7]) ? node6306 : node6249;
										assign node6249 = (inp[0]) ? node6277 : node6250;
											assign node6250 = (inp[11]) ? node6262 : node6251;
												assign node6251 = (inp[1]) ? node6257 : node6252;
													assign node6252 = (inp[4]) ? 4'b1100 : node6253;
														assign node6253 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node6257 = (inp[9]) ? 4'b1000 : node6258;
														assign node6258 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node6262 = (inp[9]) ? node6272 : node6263;
													assign node6263 = (inp[2]) ? node6267 : node6264;
														assign node6264 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node6267 = (inp[10]) ? 4'b1100 : node6268;
															assign node6268 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node6272 = (inp[10]) ? node6274 : 4'b1101;
														assign node6274 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node6277 = (inp[2]) ? node6289 : node6278;
												assign node6278 = (inp[1]) ? node6280 : 4'b1101;
													assign node6280 = (inp[4]) ? node6286 : node6281;
														assign node6281 = (inp[9]) ? node6283 : 4'b1100;
															assign node6283 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node6286 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node6289 = (inp[4]) ? node6297 : node6290;
													assign node6290 = (inp[1]) ? 4'b1101 : node6291;
														assign node6291 = (inp[10]) ? node6293 : 4'b1001;
															assign node6293 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node6297 = (inp[1]) ? node6303 : node6298;
														assign node6298 = (inp[11]) ? node6300 : 4'b1101;
															assign node6300 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6303 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node6306 = (inp[9]) ? node6324 : node6307;
											assign node6307 = (inp[0]) ? node6319 : node6308;
												assign node6308 = (inp[1]) ? node6314 : node6309;
													assign node6309 = (inp[2]) ? node6311 : 4'b1011;
														assign node6311 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node6314 = (inp[11]) ? node6316 : 4'b1010;
														assign node6316 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node6319 = (inp[2]) ? 4'b1110 : node6320;
													assign node6320 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node6324 = (inp[0]) ? node6336 : node6325;
												assign node6325 = (inp[10]) ? node6327 : 4'b1110;
													assign node6327 = (inp[1]) ? node6331 : node6328;
														assign node6328 = (inp[11]) ? 4'b1110 : 4'b1010;
														assign node6331 = (inp[4]) ? 4'b1011 : node6332;
															assign node6332 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node6336 = (inp[11]) ? node6342 : node6337;
													assign node6337 = (inp[4]) ? node6339 : 4'b1111;
														assign node6339 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node6342 = (inp[2]) ? 4'b1110 : node6343;
														assign node6343 = (inp[4]) ? 4'b1111 : 4'b1011;
									assign node6347 = (inp[7]) ? node6393 : node6348;
										assign node6348 = (inp[4]) ? node6380 : node6349;
											assign node6349 = (inp[1]) ? node6359 : node6350;
												assign node6350 = (inp[0]) ? 4'b1010 : node6351;
													assign node6351 = (inp[10]) ? node6353 : 4'b1011;
														assign node6353 = (inp[9]) ? 4'b1011 : node6354;
															assign node6354 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node6359 = (inp[9]) ? node6373 : node6360;
													assign node6360 = (inp[0]) ? 4'b1111 : node6361;
														assign node6361 = (inp[10]) ? node6367 : node6362;
															assign node6362 = (inp[11]) ? 4'b1110 : node6363;
																assign node6363 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node6367 = (inp[11]) ? node6369 : 4'b1111;
																assign node6369 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node6373 = (inp[0]) ? 4'b1110 : node6374;
														assign node6374 = (inp[2]) ? 4'b1111 : node6375;
															assign node6375 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node6380 = (inp[10]) ? node6388 : node6381;
												assign node6381 = (inp[9]) ? 4'b1011 : node6382;
													assign node6382 = (inp[2]) ? node6384 : 4'b1011;
														assign node6384 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node6388 = (inp[0]) ? node6390 : 4'b1010;
													assign node6390 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node6393 = (inp[1]) ? node6419 : node6394;
											assign node6394 = (inp[4]) ? node6404 : node6395;
												assign node6395 = (inp[2]) ? 4'b1001 : node6396;
													assign node6396 = (inp[11]) ? node6400 : node6397;
														assign node6397 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node6400 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node6404 = (inp[0]) ? node6414 : node6405;
													assign node6405 = (inp[9]) ? node6407 : 4'b1101;
														assign node6407 = (inp[2]) ? node6411 : node6408;
															assign node6408 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node6411 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node6414 = (inp[9]) ? 4'b1100 : node6415;
														assign node6415 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node6419 = (inp[4]) ? node6421 : 4'b1001;
												assign node6421 = (inp[11]) ? node6427 : node6422;
													assign node6422 = (inp[9]) ? 4'b1000 : node6423;
														assign node6423 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node6427 = (inp[10]) ? node6429 : 4'b1001;
														assign node6429 = (inp[9]) ? 4'b1001 : 4'b1000;
							assign node6432 = (inp[12]) ? node6594 : node6433;
								assign node6433 = (inp[15]) ? node6499 : node6434;
									assign node6434 = (inp[7]) ? node6466 : node6435;
										assign node6435 = (inp[4]) ? node6457 : node6436;
											assign node6436 = (inp[11]) ? node6450 : node6437;
												assign node6437 = (inp[9]) ? node6443 : node6438;
													assign node6438 = (inp[0]) ? node6440 : 4'b1100;
														assign node6440 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6443 = (inp[1]) ? node6445 : 4'b1101;
														assign node6445 = (inp[2]) ? node6447 : 4'b1101;
															assign node6447 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6450 = (inp[9]) ? 4'b1100 : node6451;
													assign node6451 = (inp[0]) ? node6453 : 4'b1101;
														assign node6453 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node6457 = (inp[2]) ? node6461 : node6458;
												assign node6458 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node6461 = (inp[9]) ? node6463 : 4'b1100;
													assign node6463 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node6466 = (inp[1]) ? node6478 : node6467;
											assign node6467 = (inp[0]) ? 4'b1111 : node6468;
												assign node6468 = (inp[10]) ? 4'b1110 : node6469;
													assign node6469 = (inp[2]) ? node6471 : 4'b1111;
														assign node6471 = (inp[11]) ? 4'b1110 : node6472;
															assign node6472 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node6478 = (inp[4]) ? node6490 : node6479;
												assign node6479 = (inp[9]) ? node6483 : node6480;
													assign node6480 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node6483 = (inp[11]) ? 4'b1111 : node6484;
														assign node6484 = (inp[2]) ? node6486 : 4'b1110;
															assign node6486 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node6490 = (inp[2]) ? 4'b1110 : node6491;
													assign node6491 = (inp[10]) ? node6493 : 4'b1111;
														assign node6493 = (inp[9]) ? 4'b1110 : node6494;
															assign node6494 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node6499 = (inp[7]) ? node6551 : node6500;
										assign node6500 = (inp[4]) ? node6528 : node6501;
											assign node6501 = (inp[1]) ? node6517 : node6502;
												assign node6502 = (inp[10]) ? node6512 : node6503;
													assign node6503 = (inp[0]) ? 4'b1110 : node6504;
														assign node6504 = (inp[11]) ? node6508 : node6505;
															assign node6505 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node6508 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node6512 = (inp[11]) ? node6514 : 4'b1111;
														assign node6514 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node6517 = (inp[2]) ? node6523 : node6518;
													assign node6518 = (inp[10]) ? node6520 : 4'b1111;
														assign node6520 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6523 = (inp[0]) ? node6525 : 4'b1110;
														assign node6525 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node6528 = (inp[1]) ? node6544 : node6529;
												assign node6529 = (inp[0]) ? node6537 : node6530;
													assign node6530 = (inp[2]) ? node6532 : 4'b1110;
														assign node6532 = (inp[11]) ? 4'b1111 : node6533;
															assign node6533 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6537 = (inp[2]) ? 4'b1110 : node6538;
														assign node6538 = (inp[9]) ? node6540 : 4'b1110;
															assign node6540 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node6544 = (inp[0]) ? 4'b1011 : node6545;
													assign node6545 = (inp[11]) ? node6547 : 4'b1010;
														assign node6547 = (inp[9]) ? 4'b1011 : 4'b1010;
										assign node6551 = (inp[4]) ? node6573 : node6552;
											assign node6552 = (inp[1]) ? node6566 : node6553;
												assign node6553 = (inp[0]) ? node6561 : node6554;
													assign node6554 = (inp[11]) ? 4'b1001 : node6555;
														assign node6555 = (inp[9]) ? 4'b1001 : node6556;
															assign node6556 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node6561 = (inp[11]) ? node6563 : 4'b1001;
														assign node6563 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6566 = (inp[11]) ? 4'b1101 : node6567;
													assign node6567 = (inp[9]) ? 4'b1101 : node6568;
														assign node6568 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node6573 = (inp[0]) ? node6587 : node6574;
												assign node6574 = (inp[10]) ? node6580 : node6575;
													assign node6575 = (inp[9]) ? 4'b1100 : node6576;
														assign node6576 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node6580 = (inp[2]) ? 4'b1101 : node6581;
														assign node6581 = (inp[11]) ? node6583 : 4'b1100;
															assign node6583 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node6587 = (inp[9]) ? 4'b1101 : node6588;
													assign node6588 = (inp[1]) ? 4'b1101 : node6589;
														assign node6589 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node6594 = (inp[15]) ? node6682 : node6595;
									assign node6595 = (inp[7]) ? node6643 : node6596;
										assign node6596 = (inp[10]) ? node6620 : node6597;
											assign node6597 = (inp[11]) ? node6605 : node6598;
												assign node6598 = (inp[1]) ? node6602 : node6599;
													assign node6599 = (inp[4]) ? 4'b1001 : 4'b1100;
													assign node6602 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6605 = (inp[9]) ? node6613 : node6606;
													assign node6606 = (inp[0]) ? 4'b1101 : node6607;
														assign node6607 = (inp[1]) ? 4'b1000 : node6608;
															assign node6608 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node6613 = (inp[2]) ? node6615 : 4'b1100;
														assign node6615 = (inp[0]) ? 4'b1101 : node6616;
															assign node6616 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node6620 = (inp[11]) ? node6630 : node6621;
												assign node6621 = (inp[2]) ? node6623 : 4'b1101;
													assign node6623 = (inp[4]) ? node6627 : node6624;
														assign node6624 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node6627 = (inp[1]) ? 4'b1100 : 4'b1001;
												assign node6630 = (inp[4]) ? node6636 : node6631;
													assign node6631 = (inp[1]) ? node6633 : 4'b1100;
														assign node6633 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node6636 = (inp[1]) ? node6638 : 4'b1001;
														assign node6638 = (inp[2]) ? 4'b1101 : node6639;
															assign node6639 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node6643 = (inp[1]) ? node6669 : node6644;
											assign node6644 = (inp[4]) ? node6656 : node6645;
												assign node6645 = (inp[0]) ? 4'b1111 : node6646;
													assign node6646 = (inp[10]) ? node6648 : 4'b1110;
														assign node6648 = (inp[2]) ? node6650 : 4'b1111;
															assign node6650 = (inp[11]) ? node6652 : 4'b1110;
																assign node6652 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node6656 = (inp[9]) ? node6660 : node6657;
													assign node6657 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6660 = (inp[11]) ? node6664 : node6661;
														assign node6661 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node6664 = (inp[10]) ? node6666 : 4'b1010;
															assign node6666 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node6669 = (inp[4]) ? node6675 : node6670;
												assign node6670 = (inp[11]) ? 4'b1010 : node6671;
													assign node6671 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node6675 = (inp[9]) ? node6677 : 4'b1110;
													assign node6677 = (inp[0]) ? node6679 : 4'b1110;
														assign node6679 = (inp[10]) ? 4'b1111 : 4'b1110;
									assign node6682 = (inp[7]) ? node6730 : node6683;
										assign node6683 = (inp[4]) ? node6705 : node6684;
											assign node6684 = (inp[1]) ? node6698 : node6685;
												assign node6685 = (inp[0]) ? node6693 : node6686;
													assign node6686 = (inp[10]) ? 4'b1110 : node6687;
														assign node6687 = (inp[2]) ? node6689 : 4'b1110;
															assign node6689 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node6693 = (inp[11]) ? 4'b1111 : node6694;
														assign node6694 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node6698 = (inp[9]) ? node6702 : node6699;
													assign node6699 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node6702 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node6705 = (inp[1]) ? node6719 : node6706;
												assign node6706 = (inp[0]) ? node6710 : node6707;
													assign node6707 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6710 = (inp[2]) ? 4'b1110 : node6711;
														assign node6711 = (inp[11]) ? node6715 : node6712;
															assign node6712 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node6715 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node6719 = (inp[11]) ? node6725 : node6720;
													assign node6720 = (inp[2]) ? node6722 : 4'b1110;
														assign node6722 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6725 = (inp[10]) ? node6727 : 4'b1111;
														assign node6727 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node6730 = (inp[1]) ? node6748 : node6731;
											assign node6731 = (inp[4]) ? node6741 : node6732;
												assign node6732 = (inp[10]) ? node6738 : node6733;
													assign node6733 = (inp[2]) ? node6735 : 4'b1100;
														assign node6735 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node6738 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6741 = (inp[0]) ? node6743 : 4'b1000;
													assign node6743 = (inp[10]) ? node6745 : 4'b1001;
														assign node6745 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node6748 = (inp[9]) ? 4'b1101 : node6749;
												assign node6749 = (inp[4]) ? node6751 : 4'b1101;
													assign node6751 = (inp[10]) ? node6753 : 4'b1100;
														assign node6753 = (inp[2]) ? 4'b1101 : node6754;
															assign node6754 = (inp[11]) ? 4'b1100 : node6755;
																assign node6755 = (inp[0]) ? 4'b1101 : 4'b1100;
						assign node6761 = (inp[5]) ? node7059 : node6762;
							assign node6762 = (inp[12]) ? node6884 : node6763;
								assign node6763 = (inp[15]) ? node6823 : node6764;
									assign node6764 = (inp[7]) ? node6794 : node6765;
										assign node6765 = (inp[9]) ? node6779 : node6766;
											assign node6766 = (inp[11]) ? node6774 : node6767;
												assign node6767 = (inp[2]) ? node6769 : 4'b1100;
													assign node6769 = (inp[0]) ? 4'b1101 : node6770;
														assign node6770 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node6774 = (inp[2]) ? node6776 : 4'b1101;
													assign node6776 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node6779 = (inp[11]) ? node6785 : node6780;
												assign node6780 = (inp[1]) ? 4'b1101 : node6781;
													assign node6781 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node6785 = (inp[2]) ? node6787 : 4'b1100;
													assign node6787 = (inp[10]) ? 4'b1101 : node6788;
														assign node6788 = (inp[0]) ? 4'b1100 : node6789;
															assign node6789 = (inp[4]) ? 4'b1101 : 4'b1100;
										assign node6794 = (inp[1]) ? node6808 : node6795;
											assign node6795 = (inp[2]) ? node6803 : node6796;
												assign node6796 = (inp[11]) ? node6800 : node6797;
													assign node6797 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node6800 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node6803 = (inp[11]) ? 4'b1111 : node6804;
													assign node6804 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node6808 = (inp[11]) ? node6814 : node6809;
												assign node6809 = (inp[9]) ? 4'b1111 : node6810;
													assign node6810 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node6814 = (inp[9]) ? 4'b1110 : node6815;
													assign node6815 = (inp[2]) ? node6817 : 4'b1111;
														assign node6817 = (inp[4]) ? 4'b1111 : node6818;
															assign node6818 = (inp[10]) ? 4'b1111 : 4'b1110;
									assign node6823 = (inp[7]) ? node6855 : node6824;
										assign node6824 = (inp[1]) ? node6838 : node6825;
											assign node6825 = (inp[9]) ? node6829 : node6826;
												assign node6826 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node6829 = (inp[2]) ? node6833 : node6830;
													assign node6830 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node6833 = (inp[11]) ? node6835 : 4'b1111;
														assign node6835 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node6838 = (inp[4]) ? node6844 : node6839;
												assign node6839 = (inp[10]) ? node6841 : 4'b1110;
													assign node6841 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node6844 = (inp[9]) ? node6850 : node6845;
													assign node6845 = (inp[2]) ? node6847 : 4'b1010;
														assign node6847 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node6850 = (inp[11]) ? node6852 : 4'b1011;
														assign node6852 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node6855 = (inp[10]) ? node6863 : node6856;
											assign node6856 = (inp[9]) ? 4'b1100 : node6857;
												assign node6857 = (inp[11]) ? 4'b1101 : node6858;
													assign node6858 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node6863 = (inp[11]) ? node6875 : node6864;
												assign node6864 = (inp[4]) ? node6868 : node6865;
													assign node6865 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node6868 = (inp[1]) ? 4'b1101 : node6869;
														assign node6869 = (inp[0]) ? 4'b1100 : node6870;
															assign node6870 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node6875 = (inp[9]) ? node6879 : node6876;
													assign node6876 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node6879 = (inp[4]) ? node6881 : 4'b1100;
														assign node6881 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node6884 = (inp[15]) ? node6976 : node6885;
									assign node6885 = (inp[7]) ? node6927 : node6886;
										assign node6886 = (inp[9]) ? node6906 : node6887;
											assign node6887 = (inp[4]) ? node6895 : node6888;
												assign node6888 = (inp[1]) ? node6890 : 4'b1101;
													assign node6890 = (inp[0]) ? 4'b1001 : node6891;
														assign node6891 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node6895 = (inp[1]) ? node6899 : node6896;
													assign node6896 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node6899 = (inp[10]) ? 4'b1101 : node6900;
														assign node6900 = (inp[2]) ? 4'b1101 : node6901;
															assign node6901 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node6906 = (inp[1]) ? node6922 : node6907;
												assign node6907 = (inp[4]) ? node6913 : node6908;
													assign node6908 = (inp[2]) ? 4'b1101 : node6909;
														assign node6909 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6913 = (inp[10]) ? 4'b1000 : node6914;
														assign node6914 = (inp[0]) ? node6916 : 4'b1000;
															assign node6916 = (inp[2]) ? 4'b1001 : node6917;
																assign node6917 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6922 = (inp[4]) ? node6924 : 4'b1000;
													assign node6924 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node6927 = (inp[2]) ? node6955 : node6928;
											assign node6928 = (inp[9]) ? node6944 : node6929;
												assign node6929 = (inp[10]) ? node6941 : node6930;
													assign node6930 = (inp[11]) ? node6934 : node6931;
														assign node6931 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node6934 = (inp[1]) ? node6938 : node6935;
															assign node6935 = (inp[0]) ? 4'b1110 : 4'b1010;
															assign node6938 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node6941 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node6944 = (inp[0]) ? 4'b1010 : node6945;
													assign node6945 = (inp[10]) ? node6951 : node6946;
														assign node6946 = (inp[1]) ? 4'b1110 : node6947;
															assign node6947 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node6951 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node6955 = (inp[0]) ? node6969 : node6956;
												assign node6956 = (inp[1]) ? node6964 : node6957;
													assign node6957 = (inp[4]) ? 4'b1011 : node6958;
														assign node6958 = (inp[11]) ? 4'b1111 : node6959;
															assign node6959 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node6964 = (inp[4]) ? 4'b1110 : node6965;
														assign node6965 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node6969 = (inp[1]) ? node6973 : node6970;
													assign node6970 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node6973 = (inp[4]) ? 4'b1111 : 4'b1011;
									assign node6976 = (inp[7]) ? node7014 : node6977;
										assign node6977 = (inp[1]) ? node6991 : node6978;
											assign node6978 = (inp[10]) ? node6984 : node6979;
												assign node6979 = (inp[9]) ? 4'b1110 : node6980;
													assign node6980 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node6984 = (inp[11]) ? node6986 : 4'b1111;
													assign node6986 = (inp[9]) ? 4'b1111 : node6987;
														assign node6987 = (inp[4]) ? 4'b1110 : 4'b1111;
											assign node6991 = (inp[4]) ? node7005 : node6992;
												assign node6992 = (inp[11]) ? node6998 : node6993;
													assign node6993 = (inp[9]) ? 4'b1010 : node6994;
														assign node6994 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node6998 = (inp[0]) ? node7000 : 4'b1011;
														assign node7000 = (inp[9]) ? 4'b1010 : node7001;
															assign node7001 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node7005 = (inp[2]) ? node7011 : node7006;
													assign node7006 = (inp[0]) ? 4'b1111 : node7007;
														assign node7007 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node7011 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node7014 = (inp[1]) ? node7034 : node7015;
											assign node7015 = (inp[4]) ? node7023 : node7016;
												assign node7016 = (inp[2]) ? node7018 : 4'b1101;
													assign node7018 = (inp[0]) ? 4'b1100 : node7019;
														assign node7019 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node7023 = (inp[2]) ? 4'b1001 : node7024;
													assign node7024 = (inp[9]) ? node7026 : 4'b1000;
														assign node7026 = (inp[10]) ? 4'b1001 : node7027;
															assign node7027 = (inp[11]) ? node7029 : 4'b1000;
																assign node7029 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node7034 = (inp[4]) ? node7044 : node7035;
												assign node7035 = (inp[2]) ? node7041 : node7036;
													assign node7036 = (inp[10]) ? 4'b1100 : node7037;
														assign node7037 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node7041 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node7044 = (inp[2]) ? node7050 : node7045;
													assign node7045 = (inp[11]) ? 4'b1101 : node7046;
														assign node7046 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node7050 = (inp[11]) ? 4'b1100 : node7051;
														assign node7051 = (inp[10]) ? node7055 : node7052;
															assign node7052 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7055 = (inp[0]) ? 4'b1100 : 4'b1101;
							assign node7059 = (inp[12]) ? node7247 : node7060;
								assign node7060 = (inp[15]) ? node7150 : node7061;
									assign node7061 = (inp[7]) ? node7099 : node7062;
										assign node7062 = (inp[1]) ? node7084 : node7063;
											assign node7063 = (inp[10]) ? node7079 : node7064;
												assign node7064 = (inp[11]) ? node7070 : node7065;
													assign node7065 = (inp[4]) ? node7067 : 4'b1001;
														assign node7067 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7070 = (inp[9]) ? node7072 : 4'b1000;
														assign node7072 = (inp[4]) ? node7076 : node7073;
															assign node7073 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node7076 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node7079 = (inp[2]) ? node7081 : 4'b1001;
													assign node7081 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node7084 = (inp[10]) ? node7086 : 4'b1000;
												assign node7086 = (inp[2]) ? node7094 : node7087;
													assign node7087 = (inp[11]) ? node7089 : 4'b1000;
														assign node7089 = (inp[4]) ? 4'b1000 : node7090;
															assign node7090 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7094 = (inp[9]) ? node7096 : 4'b1001;
														assign node7096 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node7099 = (inp[10]) ? node7125 : node7100;
											assign node7100 = (inp[11]) ? node7114 : node7101;
												assign node7101 = (inp[1]) ? node7105 : node7102;
													assign node7102 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node7105 = (inp[2]) ? node7109 : node7106;
														assign node7106 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node7109 = (inp[9]) ? 4'b1011 : node7110;
															assign node7110 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node7114 = (inp[9]) ? node7122 : node7115;
													assign node7115 = (inp[0]) ? 4'b1011 : node7116;
														assign node7116 = (inp[4]) ? 4'b1011 : node7117;
															assign node7117 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node7122 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node7125 = (inp[4]) ? node7135 : node7126;
												assign node7126 = (inp[11]) ? 4'b1010 : node7127;
													assign node7127 = (inp[9]) ? node7129 : 4'b1010;
														assign node7129 = (inp[0]) ? 4'b1011 : node7130;
															assign node7130 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node7135 = (inp[9]) ? node7145 : node7136;
													assign node7136 = (inp[2]) ? node7140 : node7137;
														assign node7137 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node7140 = (inp[0]) ? 4'b1010 : node7141;
															assign node7141 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node7145 = (inp[0]) ? 4'b1011 : node7146;
														assign node7146 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node7150 = (inp[7]) ? node7204 : node7151;
										assign node7151 = (inp[4]) ? node7183 : node7152;
											assign node7152 = (inp[2]) ? node7174 : node7153;
												assign node7153 = (inp[11]) ? node7169 : node7154;
													assign node7154 = (inp[10]) ? node7164 : node7155;
														assign node7155 = (inp[1]) ? 4'b1011 : node7156;
															assign node7156 = (inp[9]) ? node7160 : node7157;
																assign node7157 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node7160 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7164 = (inp[1]) ? 4'b1010 : node7165;
															assign node7165 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node7169 = (inp[9]) ? 4'b1010 : node7170;
														assign node7170 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node7174 = (inp[10]) ? node7178 : node7175;
													assign node7175 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node7178 = (inp[0]) ? 4'b1011 : node7179;
														assign node7179 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node7183 = (inp[1]) ? node7193 : node7184;
												assign node7184 = (inp[2]) ? 4'b1011 : node7185;
													assign node7185 = (inp[0]) ? node7189 : node7186;
														assign node7186 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node7189 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node7193 = (inp[9]) ? node7201 : node7194;
													assign node7194 = (inp[0]) ? node7196 : 4'b1111;
														assign node7196 = (inp[11]) ? node7198 : 4'b1111;
															assign node7198 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node7201 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node7204 = (inp[4]) ? node7228 : node7205;
											assign node7205 = (inp[1]) ? node7215 : node7206;
												assign node7206 = (inp[10]) ? node7208 : 4'b1100;
													assign node7208 = (inp[11]) ? node7212 : node7209;
														assign node7209 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node7212 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node7215 = (inp[10]) ? node7217 : 4'b1001;
													assign node7217 = (inp[9]) ? 4'b1000 : node7218;
														assign node7218 = (inp[2]) ? 4'b1001 : node7219;
															assign node7219 = (inp[0]) ? node7223 : node7220;
																assign node7220 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node7223 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node7228 = (inp[9]) ? node7234 : node7229;
												assign node7229 = (inp[2]) ? 4'b1001 : node7230;
													assign node7230 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node7234 = (inp[1]) ? node7242 : node7235;
													assign node7235 = (inp[11]) ? node7239 : node7236;
														assign node7236 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node7239 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node7242 = (inp[2]) ? node7244 : 4'b1000;
														assign node7244 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node7247 = (inp[15]) ? node7317 : node7248;
									assign node7248 = (inp[7]) ? node7284 : node7249;
										assign node7249 = (inp[0]) ? node7267 : node7250;
											assign node7250 = (inp[10]) ? node7258 : node7251;
												assign node7251 = (inp[1]) ? node7255 : node7252;
													assign node7252 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7255 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node7258 = (inp[11]) ? node7260 : 4'b1101;
													assign node7260 = (inp[9]) ? node7262 : 4'b1100;
														assign node7262 = (inp[1]) ? node7264 : 4'b1101;
															assign node7264 = (inp[4]) ? 4'b1000 : 4'b1101;
											assign node7267 = (inp[4]) ? node7277 : node7268;
												assign node7268 = (inp[1]) ? node7274 : node7269;
													assign node7269 = (inp[9]) ? 4'b1001 : node7270;
														assign node7270 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node7274 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node7277 = (inp[1]) ? node7279 : 4'b1101;
													assign node7279 = (inp[2]) ? node7281 : 4'b1001;
														assign node7281 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node7284 = (inp[11]) ? node7302 : node7285;
											assign node7285 = (inp[10]) ? node7291 : node7286;
												assign node7286 = (inp[2]) ? 4'b1110 : node7287;
													assign node7287 = (inp[1]) ? 4'b1011 : 4'b1110;
												assign node7291 = (inp[2]) ? node7295 : node7292;
													assign node7292 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node7295 = (inp[4]) ? node7299 : node7296;
														assign node7296 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node7299 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node7302 = (inp[10]) ? node7308 : node7303;
												assign node7303 = (inp[2]) ? node7305 : 4'b1111;
													assign node7305 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node7308 = (inp[4]) ? node7314 : node7309;
													assign node7309 = (inp[0]) ? node7311 : 4'b1010;
														assign node7311 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node7314 = (inp[1]) ? 4'b1010 : 4'b1111;
									assign node7317 = (inp[7]) ? node7349 : node7318;
										assign node7318 = (inp[1]) ? node7326 : node7319;
											assign node7319 = (inp[11]) ? node7323 : node7320;
												assign node7320 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node7323 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node7326 = (inp[4]) ? node7346 : node7327;
												assign node7327 = (inp[2]) ? node7337 : node7328;
													assign node7328 = (inp[10]) ? 4'b1110 : node7329;
														assign node7329 = (inp[0]) ? 4'b1110 : node7330;
															assign node7330 = (inp[9]) ? 4'b1111 : node7331;
																assign node7331 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node7337 = (inp[11]) ? 4'b1111 : node7338;
														assign node7338 = (inp[10]) ? node7342 : node7339;
															assign node7339 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node7342 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node7346 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node7349 = (inp[1]) ? node7373 : node7350;
											assign node7350 = (inp[4]) ? node7370 : node7351;
												assign node7351 = (inp[0]) ? node7363 : node7352;
													assign node7352 = (inp[2]) ? 4'b1000 : node7353;
														assign node7353 = (inp[10]) ? node7357 : node7354;
															assign node7354 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node7357 = (inp[9]) ? 4'b1001 : node7358;
																assign node7358 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node7363 = (inp[2]) ? 4'b1001 : node7364;
														assign node7364 = (inp[9]) ? node7366 : 4'b1000;
															assign node7366 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node7370 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node7373 = (inp[2]) ? node7383 : node7374;
												assign node7374 = (inp[10]) ? node7376 : 4'b1000;
													assign node7376 = (inp[0]) ? node7378 : 4'b1000;
														assign node7378 = (inp[9]) ? 4'b1001 : node7379;
															assign node7379 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node7383 = (inp[10]) ? node7393 : node7384;
													assign node7384 = (inp[4]) ? node7386 : 4'b1000;
														assign node7386 = (inp[11]) ? node7390 : node7387;
															assign node7387 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node7390 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7393 = (inp[4]) ? node7399 : node7394;
														assign node7394 = (inp[9]) ? node7396 : 4'b1001;
															assign node7396 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7399 = (inp[0]) ? 4'b1000 : node7400;
															assign node7400 = (inp[11]) ? 4'b1000 : 4'b1001;
					assign node7404 = (inp[4]) ? node8014 : node7405;
						assign node7405 = (inp[15]) ? node7735 : node7406;
							assign node7406 = (inp[2]) ? node7562 : node7407;
								assign node7407 = (inp[9]) ? node7483 : node7408;
									assign node7408 = (inp[1]) ? node7444 : node7409;
										assign node7409 = (inp[5]) ? node7423 : node7410;
											assign node7410 = (inp[7]) ? node7418 : node7411;
												assign node7411 = (inp[0]) ? node7415 : node7412;
													assign node7412 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node7415 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node7418 = (inp[12]) ? node7420 : 4'b0001;
													assign node7420 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node7423 = (inp[7]) ? node7437 : node7424;
												assign node7424 = (inp[12]) ? node7432 : node7425;
													assign node7425 = (inp[10]) ? 4'b0101 : node7426;
														assign node7426 = (inp[13]) ? 4'b0100 : node7427;
															assign node7427 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node7432 = (inp[13]) ? 4'b0100 : node7433;
														assign node7433 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node7437 = (inp[12]) ? node7439 : 4'b0100;
													assign node7439 = (inp[13]) ? node7441 : 4'b0001;
														assign node7441 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node7444 = (inp[10]) ? node7464 : node7445;
											assign node7445 = (inp[11]) ? node7453 : node7446;
												assign node7446 = (inp[7]) ? 4'b0001 : node7447;
													assign node7447 = (inp[5]) ? 4'b0001 : node7448;
														assign node7448 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node7453 = (inp[7]) ? node7457 : node7454;
													assign node7454 = (inp[5]) ? 4'b0001 : 4'b0100;
													assign node7457 = (inp[5]) ? node7461 : node7458;
														assign node7458 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node7461 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node7464 = (inp[0]) ? node7476 : node7465;
												assign node7465 = (inp[7]) ? node7471 : node7466;
													assign node7466 = (inp[11]) ? 4'b0100 : node7467;
														assign node7467 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node7471 = (inp[5]) ? node7473 : 4'b0101;
														assign node7473 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node7476 = (inp[11]) ? node7480 : node7477;
													assign node7477 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node7480 = (inp[12]) ? 4'b0101 : 4'b0100;
									assign node7483 = (inp[12]) ? node7519 : node7484;
										assign node7484 = (inp[11]) ? node7504 : node7485;
											assign node7485 = (inp[7]) ? node7495 : node7486;
												assign node7486 = (inp[10]) ? 4'b0001 : node7487;
													assign node7487 = (inp[1]) ? node7489 : 4'b0001;
														assign node7489 = (inp[13]) ? node7491 : 4'b0000;
															assign node7491 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node7495 = (inp[5]) ? node7501 : node7496;
													assign node7496 = (inp[0]) ? node7498 : 4'b0000;
														assign node7498 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node7501 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node7504 = (inp[5]) ? node7512 : node7505;
												assign node7505 = (inp[1]) ? node7509 : node7506;
													assign node7506 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node7509 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node7512 = (inp[1]) ? 4'b0001 : node7513;
													assign node7513 = (inp[7]) ? 4'b0101 : node7514;
														assign node7514 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node7519 = (inp[1]) ? node7545 : node7520;
											assign node7520 = (inp[10]) ? node7528 : node7521;
												assign node7521 = (inp[0]) ? 4'b0000 : node7522;
													assign node7522 = (inp[11]) ? node7524 : 4'b0100;
														assign node7524 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node7528 = (inp[11]) ? node7538 : node7529;
													assign node7529 = (inp[0]) ? node7535 : node7530;
														assign node7530 = (inp[5]) ? 4'b0000 : node7531;
															assign node7531 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node7535 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node7538 = (inp[7]) ? 4'b0101 : node7539;
														assign node7539 = (inp[5]) ? node7541 : 4'b0000;
															assign node7541 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node7545 = (inp[0]) ? node7553 : node7546;
												assign node7546 = (inp[10]) ? node7550 : node7547;
													assign node7547 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node7550 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node7553 = (inp[10]) ? node7559 : node7554;
													assign node7554 = (inp[13]) ? 4'b0101 : node7555;
														assign node7555 = (inp[7]) ? 4'b0000 : 4'b0101;
													assign node7559 = (inp[13]) ? 4'b0000 : 4'b0100;
								assign node7562 = (inp[0]) ? node7646 : node7563;
									assign node7563 = (inp[11]) ? node7599 : node7564;
										assign node7564 = (inp[13]) ? node7586 : node7565;
											assign node7565 = (inp[7]) ? node7573 : node7566;
												assign node7566 = (inp[1]) ? node7568 : 4'b0100;
													assign node7568 = (inp[5]) ? 4'b0001 : node7569;
														assign node7569 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node7573 = (inp[12]) ? node7577 : node7574;
													assign node7574 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node7577 = (inp[9]) ? node7581 : node7578;
														assign node7578 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node7581 = (inp[5]) ? node7583 : 4'b0000;
															assign node7583 = (inp[10]) ? 4'b0101 : 4'b0000;
											assign node7586 = (inp[1]) ? node7592 : node7587;
												assign node7587 = (inp[5]) ? 4'b0101 : node7588;
													assign node7588 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node7592 = (inp[7]) ? node7596 : node7593;
													assign node7593 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node7596 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node7599 = (inp[13]) ? node7619 : node7600;
											assign node7600 = (inp[10]) ? node7610 : node7601;
												assign node7601 = (inp[12]) ? node7603 : 4'b0001;
													assign node7603 = (inp[7]) ? node7605 : 4'b0001;
														assign node7605 = (inp[1]) ? node7607 : 4'b0100;
															assign node7607 = (inp[5]) ? 4'b0100 : 4'b0001;
												assign node7610 = (inp[9]) ? node7612 : 4'b0101;
													assign node7612 = (inp[1]) ? 4'b0100 : node7613;
														assign node7613 = (inp[5]) ? node7615 : 4'b0001;
															assign node7615 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node7619 = (inp[5]) ? node7635 : node7620;
												assign node7620 = (inp[9]) ? node7626 : node7621;
													assign node7621 = (inp[1]) ? 4'b0100 : node7622;
														assign node7622 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node7626 = (inp[12]) ? node7630 : node7627;
														assign node7627 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7630 = (inp[1]) ? 4'b0000 : node7631;
															assign node7631 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node7635 = (inp[10]) ? 4'b0001 : node7636;
													assign node7636 = (inp[7]) ? node7640 : node7637;
														assign node7637 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node7640 = (inp[1]) ? 4'b0101 : node7641;
															assign node7641 = (inp[12]) ? 4'b0000 : 4'b0101;
									assign node7646 = (inp[5]) ? node7696 : node7647;
										assign node7647 = (inp[1]) ? node7677 : node7648;
											assign node7648 = (inp[7]) ? node7670 : node7649;
												assign node7649 = (inp[9]) ? node7659 : node7650;
													assign node7650 = (inp[12]) ? 4'b0001 : node7651;
														assign node7651 = (inp[10]) ? node7655 : node7652;
															assign node7652 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node7655 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node7659 = (inp[12]) ? node7665 : node7660;
														assign node7660 = (inp[10]) ? node7662 : 4'b0000;
															assign node7662 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node7665 = (inp[10]) ? 4'b0000 : node7666;
															assign node7666 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node7670 = (inp[12]) ? node7674 : node7671;
													assign node7671 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node7674 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node7677 = (inp[10]) ? node7685 : node7678;
												assign node7678 = (inp[12]) ? 4'b0101 : node7679;
													assign node7679 = (inp[13]) ? node7681 : 4'b0101;
														assign node7681 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node7685 = (inp[12]) ? node7691 : node7686;
													assign node7686 = (inp[11]) ? node7688 : 4'b0101;
														assign node7688 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node7691 = (inp[7]) ? node7693 : 4'b0100;
														assign node7693 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node7696 = (inp[1]) ? node7716 : node7697;
											assign node7697 = (inp[11]) ? node7701 : node7698;
												assign node7698 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7701 = (inp[12]) ? node7711 : node7702;
													assign node7702 = (inp[9]) ? node7706 : node7703;
														assign node7703 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node7706 = (inp[10]) ? 4'b0100 : node7707;
															assign node7707 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node7711 = (inp[9]) ? node7713 : 4'b0001;
														assign node7713 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node7716 = (inp[12]) ? node7726 : node7717;
												assign node7717 = (inp[13]) ? node7723 : node7718;
													assign node7718 = (inp[11]) ? 4'b0000 : node7719;
														assign node7719 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node7723 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node7726 = (inp[7]) ? node7730 : node7727;
													assign node7727 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node7730 = (inp[11]) ? 4'b0100 : node7731;
														assign node7731 = (inp[13]) ? 4'b0101 : 4'b0100;
							assign node7735 = (inp[0]) ? node7871 : node7736;
								assign node7736 = (inp[7]) ? node7810 : node7737;
									assign node7737 = (inp[11]) ? node7769 : node7738;
										assign node7738 = (inp[13]) ? node7754 : node7739;
											assign node7739 = (inp[1]) ? node7743 : node7740;
												assign node7740 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node7743 = (inp[5]) ? 4'b0011 : node7744;
													assign node7744 = (inp[10]) ? node7748 : node7745;
														assign node7745 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node7748 = (inp[2]) ? 4'b0110 : node7749;
															assign node7749 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node7754 = (inp[12]) ? node7766 : node7755;
												assign node7755 = (inp[9]) ? node7761 : node7756;
													assign node7756 = (inp[5]) ? node7758 : 4'b0110;
														assign node7758 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node7761 = (inp[2]) ? node7763 : 4'b0110;
														assign node7763 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node7766 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node7769 = (inp[10]) ? node7797 : node7770;
											assign node7770 = (inp[13]) ? node7780 : node7771;
												assign node7771 = (inp[1]) ? node7773 : 4'b0111;
													assign node7773 = (inp[5]) ? node7777 : node7774;
														assign node7774 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node7777 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node7780 = (inp[12]) ? node7792 : node7781;
													assign node7781 = (inp[1]) ? node7787 : node7782;
														assign node7782 = (inp[5]) ? node7784 : 4'b0010;
															assign node7784 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node7787 = (inp[5]) ? node7789 : 4'b0111;
															assign node7789 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node7792 = (inp[5]) ? 4'b0110 : node7793;
														assign node7793 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node7797 = (inp[2]) ? node7805 : node7798;
												assign node7798 = (inp[9]) ? node7802 : node7799;
													assign node7799 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node7802 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node7805 = (inp[5]) ? 4'b0111 : node7806;
													assign node7806 = (inp[1]) ? 4'b0111 : 4'b0011;
									assign node7810 = (inp[12]) ? node7834 : node7811;
										assign node7811 = (inp[11]) ? node7829 : node7812;
											assign node7812 = (inp[10]) ? node7822 : node7813;
												assign node7813 = (inp[13]) ? node7815 : 4'b0110;
													assign node7815 = (inp[9]) ? 4'b0110 : node7816;
														assign node7816 = (inp[5]) ? 4'b0011 : node7817;
															assign node7817 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node7822 = (inp[5]) ? node7824 : 4'b0011;
													assign node7824 = (inp[1]) ? 4'b0110 : node7825;
														assign node7825 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node7829 = (inp[2]) ? node7831 : 4'b0010;
												assign node7831 = (inp[5]) ? 4'b0111 : 4'b0010;
										assign node7834 = (inp[9]) ? node7856 : node7835;
											assign node7835 = (inp[11]) ? node7845 : node7836;
												assign node7836 = (inp[5]) ? node7842 : node7837;
													assign node7837 = (inp[1]) ? 4'b0110 : node7838;
														assign node7838 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node7842 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node7845 = (inp[10]) ? node7849 : node7846;
													assign node7846 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node7849 = (inp[13]) ? node7851 : 4'b0011;
														assign node7851 = (inp[5]) ? node7853 : 4'b0111;
															assign node7853 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node7856 = (inp[11]) ? node7866 : node7857;
												assign node7857 = (inp[2]) ? 4'b0111 : node7858;
													assign node7858 = (inp[1]) ? node7862 : node7859;
														assign node7859 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node7862 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node7866 = (inp[2]) ? node7868 : 4'b0110;
													assign node7868 = (inp[1]) ? 4'b0110 : 4'b0010;
								assign node7871 = (inp[11]) ? node7933 : node7872;
									assign node7872 = (inp[1]) ? node7902 : node7873;
										assign node7873 = (inp[5]) ? node7891 : node7874;
											assign node7874 = (inp[12]) ? node7882 : node7875;
												assign node7875 = (inp[7]) ? 4'b0111 : node7876;
													assign node7876 = (inp[13]) ? node7878 : 4'b0011;
														assign node7878 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node7882 = (inp[7]) ? node7888 : node7883;
													assign node7883 = (inp[13]) ? node7885 : 4'b0011;
														assign node7885 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node7888 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node7891 = (inp[13]) ? node7897 : node7892;
												assign node7892 = (inp[7]) ? node7894 : 4'b0111;
													assign node7894 = (inp[12]) ? 4'b0111 : 4'b0010;
												assign node7897 = (inp[12]) ? node7899 : 4'b0010;
													assign node7899 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node7902 = (inp[13]) ? node7922 : node7903;
											assign node7903 = (inp[9]) ? node7907 : node7904;
												assign node7904 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node7907 = (inp[10]) ? node7917 : node7908;
													assign node7908 = (inp[7]) ? 4'b0111 : node7909;
														assign node7909 = (inp[5]) ? 4'b0010 : node7910;
															assign node7910 = (inp[2]) ? 4'b0110 : node7911;
																assign node7911 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node7917 = (inp[12]) ? node7919 : 4'b0010;
														assign node7919 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node7922 = (inp[7]) ? node7930 : node7923;
												assign node7923 = (inp[5]) ? node7927 : node7924;
													assign node7924 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node7927 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node7930 = (inp[2]) ? 4'b0111 : 4'b0011;
									assign node7933 = (inp[2]) ? node7971 : node7934;
										assign node7934 = (inp[5]) ? node7948 : node7935;
											assign node7935 = (inp[1]) ? node7943 : node7936;
												assign node7936 = (inp[10]) ? node7938 : 4'b0110;
													assign node7938 = (inp[9]) ? 4'b0011 : node7939;
														assign node7939 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node7943 = (inp[7]) ? 4'b0110 : node7944;
													assign node7944 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node7948 = (inp[1]) ? node7960 : node7949;
												assign node7949 = (inp[13]) ? node7955 : node7950;
													assign node7950 = (inp[12]) ? 4'b0110 : node7951;
														assign node7951 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node7955 = (inp[7]) ? node7957 : 4'b0111;
														assign node7957 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node7960 = (inp[7]) ? node7968 : node7961;
													assign node7961 = (inp[13]) ? node7965 : node7962;
														assign node7962 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node7965 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node7968 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node7971 = (inp[10]) ? node7991 : node7972;
											assign node7972 = (inp[13]) ? node7982 : node7973;
												assign node7973 = (inp[5]) ? node7977 : node7974;
													assign node7974 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node7977 = (inp[1]) ? 4'b0010 : node7978;
														assign node7978 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node7982 = (inp[1]) ? node7986 : node7983;
													assign node7983 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node7986 = (inp[5]) ? node7988 : 4'b0110;
														assign node7988 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node7991 = (inp[12]) ? node8003 : node7992;
												assign node7992 = (inp[13]) ? node7998 : node7993;
													assign node7993 = (inp[9]) ? 4'b0110 : node7994;
														assign node7994 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node7998 = (inp[7]) ? node8000 : 4'b0011;
														assign node8000 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node8003 = (inp[5]) ? node8011 : node8004;
													assign node8004 = (inp[1]) ? node8006 : 4'b0010;
														assign node8006 = (inp[7]) ? 4'b0110 : node8007;
															assign node8007 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node8011 = (inp[1]) ? 4'b0010 : 4'b0110;
						assign node8014 = (inp[15]) ? node8340 : node8015;
							assign node8015 = (inp[7]) ? node8181 : node8016;
								assign node8016 = (inp[1]) ? node8080 : node8017;
									assign node8017 = (inp[2]) ? node8041 : node8018;
										assign node8018 = (inp[13]) ? node8030 : node8019;
											assign node8019 = (inp[11]) ? 4'b0111 : node8020;
												assign node8020 = (inp[0]) ? 4'b0010 : node8021;
													assign node8021 = (inp[9]) ? node8023 : 4'b0110;
														assign node8023 = (inp[10]) ? 4'b0110 : node8024;
															assign node8024 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node8030 = (inp[5]) ? node8036 : node8031;
												assign node8031 = (inp[10]) ? node8033 : 4'b0111;
													assign node8033 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node8036 = (inp[12]) ? 4'b0010 : node8037;
													assign node8037 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node8041 = (inp[13]) ? node8061 : node8042;
											assign node8042 = (inp[5]) ? node8052 : node8043;
												assign node8043 = (inp[12]) ? 4'b0111 : node8044;
													assign node8044 = (inp[11]) ? node8048 : node8045;
														assign node8045 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node8048 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node8052 = (inp[12]) ? node8058 : node8053;
													assign node8053 = (inp[0]) ? 4'b0110 : node8054;
														assign node8054 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node8058 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node8061 = (inp[10]) ? node8071 : node8062;
												assign node8062 = (inp[12]) ? node8068 : node8063;
													assign node8063 = (inp[9]) ? 4'b0110 : node8064;
														assign node8064 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node8068 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node8071 = (inp[9]) ? node8073 : 4'b0010;
													assign node8073 = (inp[0]) ? node8075 : 4'b0111;
														assign node8075 = (inp[11]) ? node8077 : 4'b0111;
															assign node8077 = (inp[12]) ? 4'b0110 : 4'b0010;
									assign node8080 = (inp[9]) ? node8124 : node8081;
										assign node8081 = (inp[5]) ? node8107 : node8082;
											assign node8082 = (inp[12]) ? node8098 : node8083;
												assign node8083 = (inp[11]) ? node8093 : node8084;
													assign node8084 = (inp[0]) ? node8090 : node8085;
														assign node8085 = (inp[2]) ? node8087 : 4'b0110;
															assign node8087 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node8090 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node8093 = (inp[2]) ? 4'b0111 : node8094;
														assign node8094 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node8098 = (inp[13]) ? 4'b0011 : node8099;
													assign node8099 = (inp[11]) ? node8103 : node8100;
														assign node8100 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node8103 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node8107 = (inp[12]) ? node8117 : node8108;
												assign node8108 = (inp[0]) ? node8114 : node8109;
													assign node8109 = (inp[11]) ? 4'b0010 : node8110;
														assign node8110 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node8114 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node8117 = (inp[11]) ? 4'b0111 : node8118;
													assign node8118 = (inp[13]) ? 4'b0110 : node8119;
														assign node8119 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node8124 = (inp[10]) ? node8156 : node8125;
											assign node8125 = (inp[2]) ? node8143 : node8126;
												assign node8126 = (inp[13]) ? node8138 : node8127;
													assign node8127 = (inp[12]) ? 4'b0010 : node8128;
														assign node8128 = (inp[5]) ? node8130 : 4'b0111;
															assign node8130 = (inp[0]) ? node8134 : node8131;
																assign node8131 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node8134 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node8138 = (inp[0]) ? 4'b0111 : node8139;
														assign node8139 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node8143 = (inp[11]) ? node8153 : node8144;
													assign node8144 = (inp[5]) ? node8148 : node8145;
														assign node8145 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node8148 = (inp[0]) ? 4'b0011 : node8149;
															assign node8149 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node8153 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node8156 = (inp[11]) ? node8176 : node8157;
												assign node8157 = (inp[13]) ? node8169 : node8158;
													assign node8158 = (inp[5]) ? node8162 : node8159;
														assign node8159 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node8162 = (inp[12]) ? 4'b0110 : node8163;
															assign node8163 = (inp[2]) ? node8165 : 4'b0011;
																assign node8165 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node8169 = (inp[0]) ? node8171 : 4'b0110;
														assign node8171 = (inp[12]) ? node8173 : 4'b0010;
															assign node8173 = (inp[5]) ? 4'b0111 : 4'b0010;
												assign node8176 = (inp[0]) ? node8178 : 4'b0010;
													assign node8178 = (inp[5]) ? 4'b0110 : 4'b0011;
								assign node8181 = (inp[9]) ? node8269 : node8182;
									assign node8182 = (inp[11]) ? node8236 : node8183;
										assign node8183 = (inp[12]) ? node8211 : node8184;
											assign node8184 = (inp[1]) ? node8202 : node8185;
												assign node8185 = (inp[5]) ? node8191 : node8186;
													assign node8186 = (inp[0]) ? 4'b0011 : node8187;
														assign node8187 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node8191 = (inp[10]) ? node8193 : 4'b0110;
														assign node8193 = (inp[2]) ? 4'b0111 : node8194;
															assign node8194 = (inp[0]) ? node8198 : node8195;
																assign node8195 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node8198 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node8202 = (inp[5]) ? node8206 : node8203;
													assign node8203 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node8206 = (inp[0]) ? 4'b0011 : node8207;
														assign node8207 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node8211 = (inp[1]) ? node8225 : node8212;
												assign node8212 = (inp[5]) ? node8222 : node8213;
													assign node8213 = (inp[10]) ? node8215 : 4'b0011;
														assign node8215 = (inp[0]) ? 4'b0010 : node8216;
															assign node8216 = (inp[2]) ? node8218 : 4'b0011;
																assign node8218 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node8222 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node8225 = (inp[5]) ? node8231 : node8226;
													assign node8226 = (inp[13]) ? 4'b0110 : node8227;
														assign node8227 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node8231 = (inp[10]) ? node8233 : 4'b0010;
														assign node8233 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node8236 = (inp[0]) ? node8248 : node8237;
											assign node8237 = (inp[5]) ? node8245 : node8238;
												assign node8238 = (inp[1]) ? node8242 : node8239;
													assign node8239 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node8242 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node8245 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node8248 = (inp[2]) ? node8256 : node8249;
												assign node8249 = (inp[5]) ? node8253 : node8250;
													assign node8250 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node8253 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node8256 = (inp[12]) ? node8264 : node8257;
													assign node8257 = (inp[13]) ? node8261 : node8258;
														assign node8258 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node8261 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node8264 = (inp[5]) ? 4'b0110 : node8265;
														assign node8265 = (inp[10]) ? 4'b0111 : 4'b0011;
									assign node8269 = (inp[1]) ? node8313 : node8270;
										assign node8270 = (inp[5]) ? node8300 : node8271;
											assign node8271 = (inp[12]) ? node8291 : node8272;
												assign node8272 = (inp[11]) ? node8282 : node8273;
													assign node8273 = (inp[2]) ? node8275 : 4'b0011;
														assign node8275 = (inp[13]) ? node8279 : node8276;
															assign node8276 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node8279 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node8282 = (inp[10]) ? 4'b0010 : node8283;
														assign node8283 = (inp[0]) ? node8285 : 4'b0011;
															assign node8285 = (inp[2]) ? node8287 : 4'b0010;
																assign node8287 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node8291 = (inp[0]) ? node8293 : 4'b0010;
													assign node8293 = (inp[11]) ? 4'b0011 : node8294;
														assign node8294 = (inp[10]) ? 4'b0010 : node8295;
															assign node8295 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node8300 = (inp[13]) ? 4'b0110 : node8301;
												assign node8301 = (inp[10]) ? node8303 : 4'b0111;
													assign node8303 = (inp[0]) ? 4'b0110 : node8304;
														assign node8304 = (inp[11]) ? node8308 : node8305;
															assign node8305 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node8308 = (inp[12]) ? 4'b0111 : 4'b0110;
										assign node8313 = (inp[5]) ? node8323 : node8314;
											assign node8314 = (inp[11]) ? 4'b0111 : node8315;
												assign node8315 = (inp[10]) ? 4'b0111 : node8316;
													assign node8316 = (inp[13]) ? node8318 : 4'b0110;
														assign node8318 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node8323 = (inp[0]) ? node8335 : node8324;
												assign node8324 = (inp[11]) ? node8330 : node8325;
													assign node8325 = (inp[10]) ? node8327 : 4'b0010;
														assign node8327 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node8330 = (inp[13]) ? 4'b0011 : node8331;
														assign node8331 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node8335 = (inp[11]) ? node8337 : 4'b0011;
													assign node8337 = (inp[13]) ? 4'b0010 : 4'b0011;
							assign node8340 = (inp[11]) ? node8484 : node8341;
								assign node8341 = (inp[0]) ? node8411 : node8342;
									assign node8342 = (inp[1]) ? node8372 : node8343;
										assign node8343 = (inp[5]) ? node8359 : node8344;
											assign node8344 = (inp[7]) ? node8352 : node8345;
												assign node8345 = (inp[12]) ? 4'b0000 : node8346;
													assign node8346 = (inp[13]) ? 4'b0101 : node8347;
														assign node8347 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node8352 = (inp[12]) ? 4'b0001 : node8353;
													assign node8353 = (inp[10]) ? node8355 : 4'b0000;
														assign node8355 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node8359 = (inp[7]) ? node8369 : node8360;
												assign node8360 = (inp[12]) ? node8364 : node8361;
													assign node8361 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node8364 = (inp[10]) ? node8366 : 4'b0100;
														assign node8366 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node8369 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node8372 = (inp[7]) ? node8398 : node8373;
											assign node8373 = (inp[2]) ? node8383 : node8374;
												assign node8374 = (inp[5]) ? node8380 : node8375;
													assign node8375 = (inp[12]) ? node8377 : 4'b0000;
														assign node8377 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node8380 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node8383 = (inp[9]) ? node8391 : node8384;
													assign node8384 = (inp[10]) ? 4'b0101 : node8385;
														assign node8385 = (inp[12]) ? node8387 : 4'b0000;
															assign node8387 = (inp[5]) ? 4'b0000 : 4'b0101;
													assign node8391 = (inp[5]) ? node8393 : 4'b0000;
														assign node8393 = (inp[12]) ? 4'b0000 : node8394;
															assign node8394 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node8398 = (inp[5]) ? node8404 : node8399;
												assign node8399 = (inp[13]) ? 4'b0100 : node8400;
													assign node8400 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node8404 = (inp[10]) ? 4'b0000 : node8405;
													assign node8405 = (inp[9]) ? 4'b0000 : node8406;
														assign node8406 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node8411 = (inp[13]) ? node8463 : node8412;
										assign node8412 = (inp[5]) ? node8442 : node8413;
											assign node8413 = (inp[9]) ? node8433 : node8414;
												assign node8414 = (inp[12]) ? node8428 : node8415;
													assign node8415 = (inp[2]) ? node8421 : node8416;
														assign node8416 = (inp[1]) ? node8418 : 4'b0001;
															assign node8418 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node8421 = (inp[1]) ? node8425 : node8422;
															assign node8422 = (inp[7]) ? 4'b0001 : 4'b0100;
															assign node8425 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node8428 = (inp[7]) ? 4'b0100 : node8429;
														assign node8429 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node8433 = (inp[1]) ? node8437 : node8434;
													assign node8434 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node8437 = (inp[7]) ? 4'b0101 : node8438;
														assign node8438 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node8442 = (inp[12]) ? node8458 : node8443;
												assign node8443 = (inp[9]) ? node8453 : node8444;
													assign node8444 = (inp[7]) ? node8448 : node8445;
														assign node8445 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node8448 = (inp[1]) ? 4'b0001 : node8449;
															assign node8449 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node8453 = (inp[7]) ? 4'b0000 : node8454;
														assign node8454 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node8458 = (inp[2]) ? node8460 : 4'b0000;
													assign node8460 = (inp[1]) ? 4'b0001 : 4'b0101;
										assign node8463 = (inp[5]) ? node8479 : node8464;
											assign node8464 = (inp[7]) ? node8476 : node8465;
												assign node8465 = (inp[9]) ? node8471 : node8466;
													assign node8466 = (inp[2]) ? node8468 : 4'b0001;
														assign node8468 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node8471 = (inp[1]) ? 4'b0100 : node8472;
														assign node8472 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node8476 = (inp[1]) ? 4'b0101 : 4'b0001;
											assign node8479 = (inp[1]) ? 4'b0001 : node8480;
												assign node8480 = (inp[12]) ? 4'b0101 : 4'b0001;
								assign node8484 = (inp[0]) ? node8536 : node8485;
									assign node8485 = (inp[2]) ? node8519 : node8486;
										assign node8486 = (inp[13]) ? node8504 : node8487;
											assign node8487 = (inp[1]) ? node8495 : node8488;
												assign node8488 = (inp[12]) ? node8490 : 4'b0101;
													assign node8490 = (inp[5]) ? 4'b0100 : node8491;
														assign node8491 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node8495 = (inp[5]) ? node8499 : node8496;
													assign node8496 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node8499 = (inp[12]) ? 4'b0000 : node8500;
														assign node8500 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node8504 = (inp[9]) ? node8514 : node8505;
												assign node8505 = (inp[10]) ? node8507 : 4'b0100;
													assign node8507 = (inp[7]) ? 4'b0001 : node8508;
														assign node8508 = (inp[12]) ? node8510 : 4'b0100;
															assign node8510 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node8514 = (inp[1]) ? 4'b0001 : node8515;
													assign node8515 = (inp[5]) ? 4'b0101 : 4'b0000;
										assign node8519 = (inp[1]) ? node8529 : node8520;
											assign node8520 = (inp[12]) ? 4'b0101 : node8521;
												assign node8521 = (inp[13]) ? 4'b0100 : node8522;
													assign node8522 = (inp[9]) ? 4'b0001 : node8523;
														assign node8523 = (inp[10]) ? 4'b0100 : 4'b0001;
											assign node8529 = (inp[5]) ? 4'b0001 : node8530;
												assign node8530 = (inp[7]) ? 4'b0101 : node8531;
													assign node8531 = (inp[12]) ? 4'b0100 : 4'b0001;
									assign node8536 = (inp[2]) ? node8580 : node8537;
										assign node8537 = (inp[13]) ? node8559 : node8538;
											assign node8538 = (inp[9]) ? node8546 : node8539;
												assign node8539 = (inp[1]) ? node8543 : node8540;
													assign node8540 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node8543 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node8546 = (inp[12]) ? node8550 : node8547;
													assign node8547 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node8550 = (inp[5]) ? node8556 : node8551;
														assign node8551 = (inp[1]) ? node8553 : 4'b0001;
															assign node8553 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node8556 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node8559 = (inp[10]) ? node8569 : node8560;
												assign node8560 = (inp[1]) ? node8564 : node8561;
													assign node8561 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node8564 = (inp[7]) ? 4'b0100 : node8565;
														assign node8565 = (inp[12]) ? 4'b0000 : 4'b0101;
												assign node8569 = (inp[1]) ? 4'b0000 : node8570;
													assign node8570 = (inp[5]) ? node8576 : node8571;
														assign node8571 = (inp[12]) ? node8573 : 4'b0000;
															assign node8573 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node8576 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node8580 = (inp[1]) ? node8600 : node8581;
											assign node8581 = (inp[5]) ? node8593 : node8582;
												assign node8582 = (inp[13]) ? node8588 : node8583;
													assign node8583 = (inp[7]) ? 4'b0000 : node8584;
														assign node8584 = (inp[12]) ? 4'b0000 : 4'b0101;
													assign node8588 = (inp[12]) ? node8590 : 4'b0001;
														assign node8590 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node8593 = (inp[10]) ? node8597 : node8594;
													assign node8594 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node8597 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node8600 = (inp[5]) ? node8606 : node8601;
												assign node8601 = (inp[7]) ? 4'b0100 : node8602;
													assign node8602 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node8606 = (inp[7]) ? 4'b0000 : 4'b0100;
				assign node8609 = (inp[4]) ? node9759 : node8610;
					assign node8610 = (inp[8]) ? node9236 : node8611;
						assign node8611 = (inp[7]) ? node8959 : node8612;
							assign node8612 = (inp[10]) ? node8770 : node8613;
								assign node8613 = (inp[12]) ? node8685 : node8614;
									assign node8614 = (inp[13]) ? node8652 : node8615;
										assign node8615 = (inp[1]) ? node8641 : node8616;
											assign node8616 = (inp[5]) ? node8622 : node8617;
												assign node8617 = (inp[9]) ? 4'b0001 : node8618;
													assign node8618 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node8622 = (inp[9]) ? node8628 : node8623;
													assign node8623 = (inp[11]) ? 4'b0001 : node8624;
														assign node8624 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node8628 = (inp[11]) ? node8636 : node8629;
														assign node8629 = (inp[0]) ? node8633 : node8630;
															assign node8630 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node8633 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node8636 = (inp[2]) ? node8638 : 4'b0001;
															assign node8638 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node8641 = (inp[15]) ? node8647 : node8642;
												assign node8642 = (inp[2]) ? node8644 : 4'b0000;
													assign node8644 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node8647 = (inp[2]) ? 4'b0100 : node8648;
													assign node8648 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node8652 = (inp[15]) ? node8666 : node8653;
											assign node8653 = (inp[5]) ? node8659 : node8654;
												assign node8654 = (inp[9]) ? 4'b0100 : node8655;
													assign node8655 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node8659 = (inp[11]) ? 4'b0101 : node8660;
													assign node8660 = (inp[2]) ? 4'b0100 : node8661;
														assign node8661 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node8666 = (inp[1]) ? node8674 : node8667;
												assign node8667 = (inp[0]) ? node8669 : 4'b0100;
													assign node8669 = (inp[2]) ? node8671 : 4'b0100;
														assign node8671 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node8674 = (inp[9]) ? 4'b0001 : node8675;
													assign node8675 = (inp[2]) ? node8681 : node8676;
														assign node8676 = (inp[5]) ? node8678 : 4'b0000;
															assign node8678 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node8681 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node8685 = (inp[13]) ? node8737 : node8686;
										assign node8686 = (inp[1]) ? node8712 : node8687;
											assign node8687 = (inp[9]) ? node8701 : node8688;
												assign node8688 = (inp[15]) ? node8690 : 4'b0101;
													assign node8690 = (inp[0]) ? node8692 : 4'b0101;
														assign node8692 = (inp[11]) ? node8698 : node8693;
															assign node8693 = (inp[5]) ? 4'b0100 : node8694;
																assign node8694 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node8698 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node8701 = (inp[2]) ? node8707 : node8702;
													assign node8702 = (inp[0]) ? node8704 : 4'b0101;
														assign node8704 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node8707 = (inp[5]) ? node8709 : 4'b0100;
														assign node8709 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node8712 = (inp[15]) ? node8726 : node8713;
												assign node8713 = (inp[0]) ? node8721 : node8714;
													assign node8714 = (inp[9]) ? node8718 : node8715;
														assign node8715 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node8718 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node8721 = (inp[11]) ? 4'b0100 : node8722;
														assign node8722 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node8726 = (inp[0]) ? node8728 : 4'b0000;
													assign node8728 = (inp[11]) ? node8730 : 4'b0001;
														assign node8730 = (inp[5]) ? node8734 : node8731;
															assign node8731 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node8734 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node8737 = (inp[1]) ? node8751 : node8738;
											assign node8738 = (inp[0]) ? 4'b0000 : node8739;
												assign node8739 = (inp[5]) ? node8741 : 4'b0001;
													assign node8741 = (inp[15]) ? node8743 : 4'b0001;
														assign node8743 = (inp[11]) ? node8747 : node8744;
															assign node8744 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node8747 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node8751 = (inp[15]) ? node8759 : node8752;
												assign node8752 = (inp[0]) ? 4'b0001 : node8753;
													assign node8753 = (inp[5]) ? 4'b0000 : node8754;
														assign node8754 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node8759 = (inp[0]) ? 4'b0101 : node8760;
													assign node8760 = (inp[5]) ? 4'b0101 : node8761;
														assign node8761 = (inp[11]) ? node8765 : node8762;
															assign node8762 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node8765 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node8770 = (inp[0]) ? node8866 : node8771;
									assign node8771 = (inp[9]) ? node8811 : node8772;
										assign node8772 = (inp[2]) ? node8794 : node8773;
											assign node8773 = (inp[12]) ? node8783 : node8774;
												assign node8774 = (inp[5]) ? node8778 : node8775;
													assign node8775 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node8778 = (inp[1]) ? node8780 : 4'b0101;
														assign node8780 = (inp[13]) ? 4'b0000 : 4'b0101;
												assign node8783 = (inp[5]) ? node8789 : node8784;
													assign node8784 = (inp[1]) ? node8786 : 4'b0001;
														assign node8786 = (inp[11]) ? 4'b0001 : 4'b0101;
													assign node8789 = (inp[1]) ? node8791 : 4'b0000;
														assign node8791 = (inp[15]) ? 4'b0101 : 4'b0000;
											assign node8794 = (inp[15]) ? node8802 : node8795;
												assign node8795 = (inp[12]) ? node8799 : node8796;
													assign node8796 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node8799 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node8802 = (inp[5]) ? node8804 : 4'b0001;
													assign node8804 = (inp[12]) ? 4'b0001 : node8805;
														assign node8805 = (inp[11]) ? 4'b0100 : node8806;
															assign node8806 = (inp[13]) ? 4'b0100 : 4'b0001;
										assign node8811 = (inp[2]) ? node8835 : node8812;
											assign node8812 = (inp[12]) ? node8826 : node8813;
												assign node8813 = (inp[15]) ? node8817 : node8814;
													assign node8814 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node8817 = (inp[5]) ? node8821 : node8818;
														assign node8818 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node8821 = (inp[11]) ? node8823 : 4'b0100;
															assign node8823 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node8826 = (inp[13]) ? node8830 : node8827;
													assign node8827 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node8830 = (inp[1]) ? node8832 : 4'b0000;
														assign node8832 = (inp[11]) ? 4'b0100 : 4'b0000;
											assign node8835 = (inp[1]) ? node8851 : node8836;
												assign node8836 = (inp[13]) ? node8840 : node8837;
													assign node8837 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node8840 = (inp[12]) ? node8842 : 4'b0100;
														assign node8842 = (inp[11]) ? node8844 : 4'b0000;
															assign node8844 = (inp[15]) ? node8848 : node8845;
																assign node8845 = (inp[5]) ? 4'b0001 : 4'b0000;
																assign node8848 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node8851 = (inp[12]) ? node8861 : node8852;
													assign node8852 = (inp[11]) ? node8858 : node8853;
														assign node8853 = (inp[13]) ? 4'b0100 : node8854;
															assign node8854 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node8858 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node8861 = (inp[15]) ? node8863 : 4'b0101;
														assign node8863 = (inp[5]) ? 4'b0101 : 4'b0000;
									assign node8866 = (inp[5]) ? node8914 : node8867;
										assign node8867 = (inp[2]) ? node8895 : node8868;
											assign node8868 = (inp[12]) ? node8882 : node8869;
												assign node8869 = (inp[13]) ? node8875 : node8870;
													assign node8870 = (inp[9]) ? 4'b0001 : node8871;
														assign node8871 = (inp[1]) ? 4'b0101 : 4'b0000;
													assign node8875 = (inp[15]) ? node8877 : 4'b0101;
														assign node8877 = (inp[1]) ? node8879 : 4'b0101;
															assign node8879 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node8882 = (inp[13]) ? node8888 : node8883;
													assign node8883 = (inp[9]) ? 4'b0100 : node8884;
														assign node8884 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node8888 = (inp[15]) ? node8892 : node8889;
														assign node8889 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node8892 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node8895 = (inp[9]) ? node8905 : node8896;
												assign node8896 = (inp[15]) ? 4'b0001 : node8897;
													assign node8897 = (inp[11]) ? node8899 : 4'b0101;
														assign node8899 = (inp[13]) ? node8901 : 4'b0001;
															assign node8901 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node8905 = (inp[11]) ? 4'b0000 : node8906;
													assign node8906 = (inp[13]) ? node8910 : node8907;
														assign node8907 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node8910 = (inp[15]) ? 4'b0101 : 4'b0001;
										assign node8914 = (inp[15]) ? node8940 : node8915;
											assign node8915 = (inp[2]) ? node8927 : node8916;
												assign node8916 = (inp[13]) ? node8922 : node8917;
													assign node8917 = (inp[12]) ? 4'b0100 : node8918;
														assign node8918 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node8922 = (inp[9]) ? node8924 : 4'b0000;
														assign node8924 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node8927 = (inp[9]) ? node8935 : node8928;
													assign node8928 = (inp[12]) ? node8932 : node8929;
														assign node8929 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node8932 = (inp[1]) ? 4'b0101 : 4'b0000;
													assign node8935 = (inp[12]) ? node8937 : 4'b0001;
														assign node8937 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node8940 = (inp[13]) ? node8954 : node8941;
												assign node8941 = (inp[12]) ? node8945 : node8942;
													assign node8942 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node8945 = (inp[1]) ? node8947 : 4'b0100;
														assign node8947 = (inp[2]) ? node8951 : node8948;
															assign node8948 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node8951 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node8954 = (inp[1]) ? node8956 : 4'b0100;
													assign node8956 = (inp[12]) ? 4'b0101 : 4'b0001;
							assign node8959 = (inp[13]) ? node9123 : node8960;
								assign node8960 = (inp[12]) ? node9036 : node8961;
									assign node8961 = (inp[15]) ? node8991 : node8962;
										assign node8962 = (inp[0]) ? node8984 : node8963;
											assign node8963 = (inp[11]) ? node8979 : node8964;
												assign node8964 = (inp[5]) ? node8972 : node8965;
													assign node8965 = (inp[1]) ? 4'b0010 : node8966;
														assign node8966 = (inp[9]) ? 4'b0011 : node8967;
															assign node8967 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node8972 = (inp[1]) ? 4'b0011 : node8973;
														assign node8973 = (inp[2]) ? 4'b0010 : node8974;
															assign node8974 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node8979 = (inp[5]) ? 4'b0010 : node8980;
													assign node8980 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node8984 = (inp[2]) ? node8988 : node8985;
												assign node8985 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node8988 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node8991 = (inp[1]) ? node9013 : node8992;
											assign node8992 = (inp[5]) ? node9008 : node8993;
												assign node8993 = (inp[10]) ? node9003 : node8994;
													assign node8994 = (inp[0]) ? 4'b0110 : node8995;
														assign node8995 = (inp[11]) ? 4'b0111 : node8996;
															assign node8996 = (inp[2]) ? node8998 : 4'b0110;
																assign node8998 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node9003 = (inp[9]) ? 4'b0111 : node9004;
														assign node9004 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node9008 = (inp[2]) ? node9010 : 4'b0110;
													assign node9010 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node9013 = (inp[2]) ? node9031 : node9014;
												assign node9014 = (inp[10]) ? node9026 : node9015;
													assign node9015 = (inp[11]) ? node9017 : 4'b0010;
														assign node9017 = (inp[5]) ? node9019 : 4'b0010;
															assign node9019 = (inp[9]) ? node9023 : node9020;
																assign node9020 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node9023 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node9026 = (inp[5]) ? node9028 : 4'b0011;
														assign node9028 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node9031 = (inp[9]) ? node9033 : 4'b0010;
													assign node9033 = (inp[0]) ? 4'b0011 : 4'b0010;
									assign node9036 = (inp[1]) ? node9082 : node9037;
										assign node9037 = (inp[15]) ? node9049 : node9038;
											assign node9038 = (inp[9]) ? 4'b0110 : node9039;
												assign node9039 = (inp[10]) ? node9045 : node9040;
													assign node9040 = (inp[2]) ? 4'b0111 : node9041;
														assign node9041 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node9045 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node9049 = (inp[5]) ? node9063 : node9050;
												assign node9050 = (inp[11]) ? node9058 : node9051;
													assign node9051 = (inp[2]) ? node9055 : node9052;
														assign node9052 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node9055 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node9058 = (inp[10]) ? 4'b0010 : node9059;
														assign node9059 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node9063 = (inp[9]) ? node9073 : node9064;
													assign node9064 = (inp[11]) ? node9066 : 4'b0010;
														assign node9066 = (inp[2]) ? node9070 : node9067;
															assign node9067 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node9070 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node9073 = (inp[11]) ? node9075 : 4'b0011;
														assign node9075 = (inp[0]) ? node9079 : node9076;
															assign node9076 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node9079 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node9082 = (inp[10]) ? node9098 : node9083;
											assign node9083 = (inp[5]) ? node9085 : 4'b0110;
												assign node9085 = (inp[15]) ? node9091 : node9086;
													assign node9086 = (inp[9]) ? node9088 : 4'b0111;
														assign node9088 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node9091 = (inp[2]) ? node9095 : node9092;
														assign node9092 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node9095 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node9098 = (inp[0]) ? node9116 : node9099;
												assign node9099 = (inp[11]) ? node9107 : node9100;
													assign node9100 = (inp[5]) ? node9102 : 4'b0110;
														assign node9102 = (inp[2]) ? 4'b0111 : node9103;
															assign node9103 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node9107 = (inp[9]) ? node9109 : 4'b0111;
														assign node9109 = (inp[5]) ? node9111 : 4'b0110;
															assign node9111 = (inp[2]) ? 4'b0111 : node9112;
																assign node9112 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node9116 = (inp[9]) ? 4'b0111 : node9117;
													assign node9117 = (inp[15]) ? node9119 : 4'b0111;
														assign node9119 = (inp[11]) ? 4'b0110 : 4'b0111;
								assign node9123 = (inp[12]) ? node9187 : node9124;
									assign node9124 = (inp[1]) ? node9154 : node9125;
										assign node9125 = (inp[15]) ? node9143 : node9126;
											assign node9126 = (inp[11]) ? node9132 : node9127;
												assign node9127 = (inp[2]) ? 4'b0110 : node9128;
													assign node9128 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node9132 = (inp[2]) ? 4'b0111 : node9133;
													assign node9133 = (inp[5]) ? node9137 : node9134;
														assign node9134 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node9137 = (inp[0]) ? 4'b0111 : node9138;
															assign node9138 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node9143 = (inp[9]) ? node9151 : node9144;
												assign node9144 = (inp[10]) ? 4'b0010 : node9145;
													assign node9145 = (inp[11]) ? node9147 : 4'b0011;
														assign node9147 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node9151 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node9154 = (inp[15]) ? node9174 : node9155;
											assign node9155 = (inp[11]) ? node9167 : node9156;
												assign node9156 = (inp[9]) ? 4'b0111 : node9157;
													assign node9157 = (inp[2]) ? node9161 : node9158;
														assign node9158 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node9161 = (inp[0]) ? 4'b0111 : node9162;
															assign node9162 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node9167 = (inp[5]) ? node9169 : 4'b0110;
													assign node9169 = (inp[2]) ? node9171 : 4'b0111;
														assign node9171 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node9174 = (inp[2]) ? node9182 : node9175;
												assign node9175 = (inp[9]) ? node9179 : node9176;
													assign node9176 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node9179 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node9182 = (inp[9]) ? 4'b0110 : node9183;
													assign node9183 = (inp[0]) ? 4'b0111 : 4'b0110;
									assign node9187 = (inp[15]) ? node9205 : node9188;
										assign node9188 = (inp[9]) ? node9196 : node9189;
											assign node9189 = (inp[11]) ? node9191 : 4'b0011;
												assign node9191 = (inp[5]) ? node9193 : 4'b0010;
													assign node9193 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node9196 = (inp[11]) ? 4'b0010 : node9197;
												assign node9197 = (inp[1]) ? node9199 : 4'b0010;
													assign node9199 = (inp[2]) ? node9201 : 4'b0011;
														assign node9201 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node9205 = (inp[1]) ? node9227 : node9206;
											assign node9206 = (inp[0]) ? node9216 : node9207;
												assign node9207 = (inp[5]) ? 4'b0111 : node9208;
													assign node9208 = (inp[10]) ? 4'b0111 : node9209;
														assign node9209 = (inp[9]) ? node9211 : 4'b0110;
															assign node9211 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node9216 = (inp[11]) ? node9222 : node9217;
													assign node9217 = (inp[9]) ? 4'b0111 : node9218;
														assign node9218 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node9222 = (inp[5]) ? 4'b0110 : node9223;
														assign node9223 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node9227 = (inp[10]) ? 4'b0010 : node9228;
												assign node9228 = (inp[11]) ? 4'b0011 : node9229;
													assign node9229 = (inp[0]) ? node9231 : 4'b0011;
														assign node9231 = (inp[2]) ? 4'b0011 : 4'b0010;
						assign node9236 = (inp[15]) ? node9540 : node9237;
							assign node9237 = (inp[10]) ? node9407 : node9238;
								assign node9238 = (inp[2]) ? node9324 : node9239;
									assign node9239 = (inp[0]) ? node9281 : node9240;
										assign node9240 = (inp[9]) ? node9260 : node9241;
											assign node9241 = (inp[1]) ? node9253 : node9242;
												assign node9242 = (inp[12]) ? node9246 : node9243;
													assign node9243 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node9246 = (inp[13]) ? node9248 : 4'b0110;
														assign node9248 = (inp[5]) ? 4'b0111 : node9249;
															assign node9249 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node9253 = (inp[12]) ? node9255 : 4'b0110;
													assign node9255 = (inp[13]) ? 4'b0010 : node9256;
														assign node9256 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node9260 = (inp[13]) ? node9272 : node9261;
												assign node9261 = (inp[7]) ? 4'b0110 : node9262;
													assign node9262 = (inp[5]) ? node9266 : node9263;
														assign node9263 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node9266 = (inp[11]) ? 4'b0010 : node9267;
															assign node9267 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node9272 = (inp[1]) ? node9278 : node9273;
													assign node9273 = (inp[7]) ? 4'b0111 : node9274;
														assign node9274 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node9278 = (inp[12]) ? 4'b0010 : 4'b0111;
										assign node9281 = (inp[5]) ? node9297 : node9282;
											assign node9282 = (inp[7]) ? node9290 : node9283;
												assign node9283 = (inp[1]) ? node9287 : node9284;
													assign node9284 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node9287 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node9290 = (inp[12]) ? node9294 : node9291;
													assign node9291 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node9294 = (inp[1]) ? 4'b0011 : 4'b0110;
											assign node9297 = (inp[11]) ? node9315 : node9298;
												assign node9298 = (inp[13]) ? node9308 : node9299;
													assign node9299 = (inp[7]) ? node9305 : node9300;
														assign node9300 = (inp[1]) ? node9302 : 4'b0011;
															assign node9302 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node9305 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node9308 = (inp[7]) ? 4'b0011 : node9309;
														assign node9309 = (inp[12]) ? node9311 : 4'b0110;
															assign node9311 = (inp[1]) ? 4'b0011 : 4'b0110;
												assign node9315 = (inp[12]) ? node9317 : 4'b0010;
													assign node9317 = (inp[1]) ? node9321 : node9318;
														assign node9318 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node9321 = (inp[13]) ? 4'b0011 : 4'b0010;
									assign node9324 = (inp[0]) ? node9370 : node9325;
										assign node9325 = (inp[5]) ? node9349 : node9326;
											assign node9326 = (inp[13]) ? node9342 : node9327;
												assign node9327 = (inp[11]) ? node9337 : node9328;
													assign node9328 = (inp[7]) ? node9330 : 4'b0111;
														assign node9330 = (inp[9]) ? 4'b0111 : node9331;
															assign node9331 = (inp[12]) ? 4'b0011 : node9332;
																assign node9332 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node9337 = (inp[9]) ? node9339 : 4'b0011;
														assign node9339 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node9342 = (inp[9]) ? 4'b0011 : node9343;
													assign node9343 = (inp[11]) ? node9345 : 4'b0011;
														assign node9345 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node9349 = (inp[7]) ? node9363 : node9350;
												assign node9350 = (inp[13]) ? node9360 : node9351;
													assign node9351 = (inp[9]) ? node9353 : 4'b0011;
														assign node9353 = (inp[1]) ? node9357 : node9354;
															assign node9354 = (inp[11]) ? 4'b0111 : 4'b0011;
															assign node9357 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node9360 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node9363 = (inp[13]) ? 4'b0011 : node9364;
													assign node9364 = (inp[1]) ? node9366 : 4'b0010;
														assign node9366 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node9370 = (inp[5]) ? node9380 : node9371;
											assign node9371 = (inp[1]) ? node9377 : node9372;
												assign node9372 = (inp[12]) ? node9374 : 4'b0010;
													assign node9374 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node9377 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node9380 = (inp[11]) ? node9400 : node9381;
												assign node9381 = (inp[12]) ? node9393 : node9382;
													assign node9382 = (inp[1]) ? node9388 : node9383;
														assign node9383 = (inp[13]) ? node9385 : 4'b0010;
															assign node9385 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node9388 = (inp[7]) ? node9390 : 4'b0110;
															assign node9390 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node9393 = (inp[1]) ? 4'b0011 : node9394;
														assign node9394 = (inp[7]) ? 4'b0110 : node9395;
															assign node9395 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node9400 = (inp[13]) ? node9402 : 4'b0011;
													assign node9402 = (inp[1]) ? 4'b0010 : node9403;
														assign node9403 = (inp[7]) ? 4'b0010 : 4'b0011;
								assign node9407 = (inp[7]) ? node9481 : node9408;
									assign node9408 = (inp[9]) ? node9456 : node9409;
										assign node9409 = (inp[1]) ? node9431 : node9410;
											assign node9410 = (inp[12]) ? node9422 : node9411;
												assign node9411 = (inp[5]) ? node9413 : 4'b0010;
													assign node9413 = (inp[2]) ? node9415 : 4'b0010;
														assign node9415 = (inp[0]) ? node9419 : node9416;
															assign node9416 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node9419 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node9422 = (inp[11]) ? 4'b0110 : node9423;
													assign node9423 = (inp[2]) ? node9425 : 4'b0111;
														assign node9425 = (inp[0]) ? 4'b0111 : node9426;
															assign node9426 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node9431 = (inp[12]) ? node9447 : node9432;
												assign node9432 = (inp[11]) ? 4'b0111 : node9433;
													assign node9433 = (inp[5]) ? node9437 : node9434;
														assign node9434 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node9437 = (inp[13]) ? 4'b0111 : node9438;
															assign node9438 = (inp[0]) ? node9442 : node9439;
																assign node9439 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node9442 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node9447 = (inp[0]) ? node9449 : 4'b0010;
													assign node9449 = (inp[11]) ? node9451 : 4'b0011;
														assign node9451 = (inp[2]) ? 4'b0011 : node9452;
															assign node9452 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node9456 = (inp[1]) ? node9474 : node9457;
											assign node9457 = (inp[12]) ? node9461 : node9458;
												assign node9458 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node9461 = (inp[0]) ? node9463 : 4'b0110;
													assign node9463 = (inp[11]) ? node9469 : node9464;
														assign node9464 = (inp[2]) ? node9466 : 4'b0111;
															assign node9466 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node9469 = (inp[2]) ? node9471 : 4'b0110;
															assign node9471 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node9474 = (inp[12]) ? node9476 : 4'b0110;
												assign node9476 = (inp[0]) ? 4'b0010 : node9477;
													assign node9477 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node9481 = (inp[1]) ? node9511 : node9482;
										assign node9482 = (inp[12]) ? node9502 : node9483;
											assign node9483 = (inp[13]) ? node9497 : node9484;
												assign node9484 = (inp[5]) ? node9492 : node9485;
													assign node9485 = (inp[0]) ? node9489 : node9486;
														assign node9486 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node9489 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node9492 = (inp[11]) ? node9494 : 4'b0010;
														assign node9494 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node9497 = (inp[9]) ? node9499 : 4'b0011;
													assign node9499 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node9502 = (inp[5]) ? node9506 : node9503;
												assign node9503 = (inp[13]) ? 4'b0111 : 4'b0110;
												assign node9506 = (inp[2]) ? 4'b0111 : node9507;
													assign node9507 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node9511 = (inp[12]) ? node9527 : node9512;
											assign node9512 = (inp[11]) ? node9522 : node9513;
												assign node9513 = (inp[9]) ? 4'b0111 : node9514;
													assign node9514 = (inp[13]) ? node9516 : 4'b0111;
														assign node9516 = (inp[0]) ? 4'b0110 : node9517;
															assign node9517 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node9522 = (inp[0]) ? 4'b0110 : node9523;
													assign node9523 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node9527 = (inp[2]) ? node9535 : node9528;
												assign node9528 = (inp[0]) ? node9532 : node9529;
													assign node9529 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node9532 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node9535 = (inp[0]) ? 4'b0010 : node9536;
													assign node9536 = (inp[11]) ? 4'b0011 : 4'b0010;
							assign node9540 = (inp[2]) ? node9616 : node9541;
								assign node9541 = (inp[0]) ? node9577 : node9542;
									assign node9542 = (inp[1]) ? node9560 : node9543;
										assign node9543 = (inp[12]) ? node9553 : node9544;
											assign node9544 = (inp[13]) ? node9546 : 4'b0010;
												assign node9546 = (inp[7]) ? node9550 : node9547;
													assign node9547 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node9550 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node9553 = (inp[5]) ? 4'b0110 : node9554;
												assign node9554 = (inp[13]) ? node9556 : 4'b0111;
													assign node9556 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node9560 = (inp[12]) ? node9572 : node9561;
											assign node9561 = (inp[13]) ? 4'b0110 : node9562;
												assign node9562 = (inp[10]) ? node9566 : node9563;
													assign node9563 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node9566 = (inp[11]) ? 4'b0110 : node9567;
														assign node9567 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node9572 = (inp[5]) ? 4'b0010 : node9573;
												assign node9573 = (inp[13]) ? 4'b0010 : 4'b0011;
									assign node9577 = (inp[5]) ? node9605 : node9578;
										assign node9578 = (inp[12]) ? node9586 : node9579;
											assign node9579 = (inp[1]) ? node9581 : 4'b0011;
												assign node9581 = (inp[7]) ? node9583 : 4'b0111;
													assign node9583 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node9586 = (inp[1]) ? node9596 : node9587;
												assign node9587 = (inp[9]) ? node9589 : 4'b0111;
													assign node9589 = (inp[11]) ? 4'b0111 : node9590;
														assign node9590 = (inp[7]) ? 4'b0110 : node9591;
															assign node9591 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node9596 = (inp[11]) ? node9600 : node9597;
													assign node9597 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node9600 = (inp[13]) ? 4'b0011 : node9601;
														assign node9601 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node9605 = (inp[1]) ? node9609 : node9606;
											assign node9606 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node9609 = (inp[12]) ? 4'b0011 : node9610;
												assign node9610 = (inp[7]) ? 4'b0111 : node9611;
													assign node9611 = (inp[10]) ? 4'b0111 : 4'b0110;
								assign node9616 = (inp[0]) ? node9684 : node9617;
									assign node9617 = (inp[5]) ? node9659 : node9618;
										assign node9618 = (inp[12]) ? node9630 : node9619;
											assign node9619 = (inp[1]) ? node9625 : node9620;
												assign node9620 = (inp[7]) ? 4'b0011 : node9621;
													assign node9621 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node9625 = (inp[7]) ? node9627 : 4'b0111;
													assign node9627 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node9630 = (inp[1]) ? node9642 : node9631;
												assign node9631 = (inp[11]) ? 4'b0110 : node9632;
													assign node9632 = (inp[9]) ? node9636 : node9633;
														assign node9633 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node9636 = (inp[10]) ? 4'b0110 : node9637;
															assign node9637 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node9642 = (inp[10]) ? node9648 : node9643;
													assign node9643 = (inp[7]) ? 4'b0011 : node9644;
														assign node9644 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node9648 = (inp[11]) ? node9654 : node9649;
														assign node9649 = (inp[7]) ? 4'b0011 : node9650;
															assign node9650 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node9654 = (inp[13]) ? node9656 : 4'b0010;
															assign node9656 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node9659 = (inp[11]) ? node9671 : node9660;
											assign node9660 = (inp[7]) ? 4'b0111 : node9661;
												assign node9661 = (inp[13]) ? node9667 : node9662;
													assign node9662 = (inp[1]) ? 4'b0110 : node9663;
														assign node9663 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node9667 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node9671 = (inp[12]) ? node9681 : node9672;
												assign node9672 = (inp[1]) ? node9678 : node9673;
													assign node9673 = (inp[7]) ? node9675 : 4'b0011;
														assign node9675 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node9678 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node9681 = (inp[1]) ? 4'b0011 : 4'b0111;
									assign node9684 = (inp[10]) ? node9718 : node9685;
										assign node9685 = (inp[9]) ? node9695 : node9686;
											assign node9686 = (inp[13]) ? 4'b0110 : node9687;
												assign node9687 = (inp[1]) ? node9691 : node9688;
													assign node9688 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node9691 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node9695 = (inp[7]) ? node9705 : node9696;
												assign node9696 = (inp[11]) ? node9700 : node9697;
													assign node9697 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node9700 = (inp[13]) ? node9702 : 4'b0010;
														assign node9702 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node9705 = (inp[11]) ? node9713 : node9706;
													assign node9706 = (inp[13]) ? node9708 : 4'b0010;
														assign node9708 = (inp[1]) ? node9710 : 4'b0110;
															assign node9710 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node9713 = (inp[1]) ? node9715 : 4'b0110;
														assign node9715 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node9718 = (inp[7]) ? node9732 : node9719;
											assign node9719 = (inp[1]) ? node9725 : node9720;
												assign node9720 = (inp[12]) ? node9722 : 4'b0010;
													assign node9722 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node9725 = (inp[12]) ? 4'b0010 : node9726;
													assign node9726 = (inp[5]) ? node9728 : 4'b0110;
														assign node9728 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node9732 = (inp[5]) ? node9738 : node9733;
												assign node9733 = (inp[13]) ? 4'b0010 : node9734;
													assign node9734 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node9738 = (inp[9]) ? node9748 : node9739;
													assign node9739 = (inp[13]) ? node9741 : 4'b0110;
														assign node9741 = (inp[12]) ? node9745 : node9742;
															assign node9742 = (inp[11]) ? 4'b0110 : 4'b0011;
															assign node9745 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node9748 = (inp[13]) ? node9756 : node9749;
														assign node9749 = (inp[1]) ? node9753 : node9750;
															assign node9750 = (inp[11]) ? 4'b0110 : 4'b0010;
															assign node9753 = (inp[11]) ? 4'b0010 : 4'b0110;
														assign node9756 = (inp[1]) ? 4'b0010 : 4'b0011;
					assign node9759 = (inp[8]) ? node10253 : node9760;
						assign node9760 = (inp[7]) ? node10038 : node9761;
							assign node9761 = (inp[0]) ? node9909 : node9762;
								assign node9762 = (inp[11]) ? node9844 : node9763;
									assign node9763 = (inp[15]) ? node9801 : node9764;
										assign node9764 = (inp[13]) ? node9786 : node9765;
											assign node9765 = (inp[1]) ? node9773 : node9766;
												assign node9766 = (inp[5]) ? node9770 : node9767;
													assign node9767 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node9770 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node9773 = (inp[2]) ? node9781 : node9774;
													assign node9774 = (inp[10]) ? node9776 : 4'b0010;
														assign node9776 = (inp[5]) ? node9778 : 4'b0010;
															assign node9778 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node9781 = (inp[10]) ? node9783 : 4'b0011;
														assign node9783 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node9786 = (inp[9]) ? node9794 : node9787;
												assign node9787 = (inp[5]) ? node9789 : 4'b0110;
													assign node9789 = (inp[12]) ? node9791 : 4'b0111;
														assign node9791 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node9794 = (inp[5]) ? node9796 : 4'b0111;
													assign node9796 = (inp[12]) ? node9798 : 4'b0110;
														assign node9798 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node9801 = (inp[13]) ? node9823 : node9802;
											assign node9802 = (inp[12]) ? node9814 : node9803;
												assign node9803 = (inp[10]) ? node9805 : 4'b0111;
													assign node9805 = (inp[2]) ? node9807 : 4'b0110;
														assign node9807 = (inp[1]) ? node9811 : node9808;
															assign node9808 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node9811 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node9814 = (inp[10]) ? 4'b0111 : node9815;
													assign node9815 = (inp[1]) ? 4'b0111 : node9816;
														assign node9816 = (inp[9]) ? node9818 : 4'b0110;
															assign node9818 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node9823 = (inp[12]) ? node9837 : node9824;
												assign node9824 = (inp[9]) ? node9830 : node9825;
													assign node9825 = (inp[1]) ? node9827 : 4'b0011;
														assign node9827 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node9830 = (inp[2]) ? 4'b0010 : node9831;
														assign node9831 = (inp[1]) ? node9833 : 4'b0011;
															assign node9833 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node9837 = (inp[9]) ? 4'b0011 : node9838;
													assign node9838 = (inp[1]) ? 4'b0011 : node9839;
														assign node9839 = (inp[5]) ? 4'b0011 : 4'b0010;
									assign node9844 = (inp[13]) ? node9862 : node9845;
										assign node9845 = (inp[15]) ? 4'b0111 : node9846;
											assign node9846 = (inp[1]) ? node9854 : node9847;
												assign node9847 = (inp[5]) ? node9851 : node9848;
													assign node9848 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node9851 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node9854 = (inp[10]) ? node9856 : 4'b0011;
													assign node9856 = (inp[9]) ? node9858 : 4'b0011;
														assign node9858 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node9862 = (inp[15]) ? node9878 : node9863;
											assign node9863 = (inp[5]) ? node9869 : node9864;
												assign node9864 = (inp[12]) ? node9866 : 4'b0111;
													assign node9866 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node9869 = (inp[10]) ? node9875 : node9870;
													assign node9870 = (inp[1]) ? 4'b0110 : node9871;
														assign node9871 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node9875 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node9878 = (inp[1]) ? node9888 : node9879;
												assign node9879 = (inp[5]) ? 4'b0011 : node9880;
													assign node9880 = (inp[2]) ? 4'b0011 : node9881;
														assign node9881 = (inp[9]) ? 4'b0010 : node9882;
															assign node9882 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node9888 = (inp[9]) ? node9900 : node9889;
													assign node9889 = (inp[2]) ? node9891 : 4'b0011;
														assign node9891 = (inp[10]) ? node9897 : node9892;
															assign node9892 = (inp[12]) ? node9894 : 4'b0011;
																assign node9894 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node9897 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node9900 = (inp[10]) ? 4'b0010 : node9901;
														assign node9901 = (inp[2]) ? 4'b0011 : node9902;
															assign node9902 = (inp[5]) ? 4'b0010 : node9903;
																assign node9903 = (inp[12]) ? 4'b0010 : 4'b0011;
								assign node9909 = (inp[13]) ? node9981 : node9910;
									assign node9910 = (inp[15]) ? node9944 : node9911;
										assign node9911 = (inp[10]) ? node9923 : node9912;
											assign node9912 = (inp[5]) ? 4'b0010 : node9913;
												assign node9913 = (inp[1]) ? 4'b0010 : node9914;
													assign node9914 = (inp[12]) ? node9918 : node9915;
														assign node9915 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node9918 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node9923 = (inp[2]) ? node9937 : node9924;
												assign node9924 = (inp[5]) ? node9928 : node9925;
													assign node9925 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node9928 = (inp[1]) ? 4'b0011 : node9929;
														assign node9929 = (inp[12]) ? node9933 : node9930;
															assign node9930 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node9933 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node9937 = (inp[12]) ? 4'b0010 : node9938;
													assign node9938 = (inp[5]) ? node9940 : 4'b0011;
														assign node9940 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node9944 = (inp[2]) ? node9968 : node9945;
											assign node9945 = (inp[12]) ? node9955 : node9946;
												assign node9946 = (inp[5]) ? 4'b0111 : node9947;
													assign node9947 = (inp[1]) ? node9951 : node9948;
														assign node9948 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node9951 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node9955 = (inp[5]) ? node9961 : node9956;
													assign node9956 = (inp[10]) ? 4'b0111 : node9957;
														assign node9957 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node9961 = (inp[11]) ? node9963 : 4'b0111;
														assign node9963 = (inp[1]) ? 4'b0110 : node9964;
															assign node9964 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node9968 = (inp[5]) ? node9970 : 4'b0110;
												assign node9970 = (inp[1]) ? node9976 : node9971;
													assign node9971 = (inp[12]) ? 4'b0110 : node9972;
														assign node9972 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node9976 = (inp[10]) ? 4'b0111 : node9977;
														assign node9977 = (inp[12]) ? 4'b0111 : 4'b0110;
									assign node9981 = (inp[15]) ? node9999 : node9982;
										assign node9982 = (inp[11]) ? node9988 : node9983;
											assign node9983 = (inp[9]) ? node9985 : 4'b0111;
												assign node9985 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node9988 = (inp[12]) ? 4'b0111 : node9989;
												assign node9989 = (inp[2]) ? node9991 : 4'b0110;
													assign node9991 = (inp[1]) ? 4'b0111 : node9992;
														assign node9992 = (inp[9]) ? 4'b0111 : node9993;
															assign node9993 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node9999 = (inp[11]) ? node10009 : node10000;
											assign node10000 = (inp[10]) ? 4'b0010 : node10001;
												assign node10001 = (inp[9]) ? node10005 : node10002;
													assign node10002 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node10005 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node10009 = (inp[1]) ? node10033 : node10010;
												assign node10010 = (inp[12]) ? node10022 : node10011;
													assign node10011 = (inp[10]) ? node10017 : node10012;
														assign node10012 = (inp[9]) ? 4'b0011 : node10013;
															assign node10013 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node10017 = (inp[5]) ? node10019 : 4'b0011;
															assign node10019 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node10022 = (inp[2]) ? node10028 : node10023;
														assign node10023 = (inp[5]) ? node10025 : 4'b0010;
															assign node10025 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node10028 = (inp[9]) ? node10030 : 4'b0011;
															assign node10030 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node10033 = (inp[2]) ? 4'b0010 : node10034;
													assign node10034 = (inp[9]) ? 4'b0011 : 4'b0010;
							assign node10038 = (inp[11]) ? node10178 : node10039;
								assign node10039 = (inp[10]) ? node10085 : node10040;
									assign node10040 = (inp[1]) ? node10070 : node10041;
										assign node10041 = (inp[13]) ? node10053 : node10042;
											assign node10042 = (inp[9]) ? node10044 : 4'b0000;
												assign node10044 = (inp[2]) ? node10046 : 4'b0001;
													assign node10046 = (inp[12]) ? node10048 : 4'b0001;
														assign node10048 = (inp[0]) ? node10050 : 4'b0000;
															assign node10050 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node10053 = (inp[0]) ? node10063 : node10054;
												assign node10054 = (inp[9]) ? node10056 : 4'b0100;
													assign node10056 = (inp[2]) ? node10058 : 4'b0100;
														assign node10058 = (inp[12]) ? 4'b0101 : node10059;
															assign node10059 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node10063 = (inp[9]) ? node10067 : node10064;
													assign node10064 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node10067 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node10070 = (inp[13]) ? node10078 : node10071;
											assign node10071 = (inp[12]) ? node10073 : 4'b0101;
												assign node10073 = (inp[9]) ? node10075 : 4'b0100;
													assign node10075 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node10078 = (inp[9]) ? node10082 : node10079;
												assign node10079 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node10082 = (inp[0]) ? 4'b0000 : 4'b0001;
									assign node10085 = (inp[5]) ? node10127 : node10086;
										assign node10086 = (inp[12]) ? node10106 : node10087;
											assign node10087 = (inp[13]) ? node10103 : node10088;
												assign node10088 = (inp[1]) ? node10090 : 4'b0000;
													assign node10090 = (inp[2]) ? node10098 : node10091;
														assign node10091 = (inp[15]) ? node10095 : node10092;
															assign node10092 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node10095 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node10098 = (inp[9]) ? node10100 : 4'b0100;
															assign node10100 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node10103 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node10106 = (inp[15]) ? node10112 : node10107;
												assign node10107 = (inp[1]) ? node10109 : 4'b0001;
													assign node10109 = (inp[0]) ? 4'b0100 : 4'b0001;
												assign node10112 = (inp[13]) ? node10118 : node10113;
													assign node10113 = (inp[1]) ? 4'b0100 : node10114;
														assign node10114 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node10118 = (inp[2]) ? 4'b0100 : node10119;
														assign node10119 = (inp[0]) ? node10123 : node10120;
															assign node10120 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node10123 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node10127 = (inp[15]) ? node10145 : node10128;
											assign node10128 = (inp[2]) ? node10138 : node10129;
												assign node10129 = (inp[13]) ? node10133 : node10130;
													assign node10130 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node10133 = (inp[9]) ? 4'b0100 : node10134;
														assign node10134 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node10138 = (inp[9]) ? node10142 : node10139;
													assign node10139 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node10142 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node10145 = (inp[9]) ? node10163 : node10146;
												assign node10146 = (inp[0]) ? node10152 : node10147;
													assign node10147 = (inp[12]) ? node10149 : 4'b0000;
														assign node10149 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node10152 = (inp[2]) ? node10158 : node10153;
														assign node10153 = (inp[1]) ? node10155 : 4'b0100;
															assign node10155 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node10158 = (inp[13]) ? 4'b0001 : node10159;
															assign node10159 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node10163 = (inp[1]) ? node10173 : node10164;
													assign node10164 = (inp[13]) ? node10168 : node10165;
														assign node10165 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node10168 = (inp[12]) ? node10170 : 4'b0101;
															assign node10170 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node10173 = (inp[13]) ? node10175 : 4'b0100;
														assign node10175 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node10178 = (inp[9]) ? node10216 : node10179;
									assign node10179 = (inp[0]) ? node10199 : node10180;
										assign node10180 = (inp[13]) ? node10188 : node10181;
											assign node10181 = (inp[1]) ? node10185 : node10182;
												assign node10182 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node10185 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node10188 = (inp[1]) ? 4'b0000 : node10189;
												assign node10189 = (inp[10]) ? node10191 : 4'b0100;
													assign node10191 = (inp[15]) ? node10195 : node10192;
														assign node10192 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node10195 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node10199 = (inp[13]) ? node10211 : node10200;
											assign node10200 = (inp[1]) ? node10208 : node10201;
												assign node10201 = (inp[5]) ? node10203 : 4'b0000;
													assign node10203 = (inp[15]) ? node10205 : 4'b0001;
														assign node10205 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node10208 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node10211 = (inp[1]) ? 4'b0001 : node10212;
												assign node10212 = (inp[12]) ? 4'b0101 : 4'b0100;
									assign node10216 = (inp[0]) ? node10230 : node10217;
										assign node10217 = (inp[13]) ? node10225 : node10218;
											assign node10218 = (inp[1]) ? node10222 : node10219;
												assign node10219 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node10222 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node10225 = (inp[1]) ? 4'b0001 : node10226;
												assign node10226 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node10230 = (inp[13]) ? node10248 : node10231;
											assign node10231 = (inp[1]) ? node10245 : node10232;
												assign node10232 = (inp[2]) ? node10242 : node10233;
													assign node10233 = (inp[5]) ? 4'b0001 : node10234;
														assign node10234 = (inp[15]) ? node10238 : node10235;
															assign node10235 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node10238 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node10242 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node10245 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node10248 = (inp[1]) ? 4'b0000 : node10249;
												assign node10249 = (inp[12]) ? 4'b0100 : 4'b0101;
						assign node10253 = (inp[1]) ? node10381 : node10254;
							assign node10254 = (inp[15]) ? node10310 : node10255;
								assign node10255 = (inp[7]) ? node10279 : node10256;
									assign node10256 = (inp[0]) ? node10268 : node10257;
										assign node10257 = (inp[5]) ? node10263 : node10258;
											assign node10258 = (inp[12]) ? node10260 : 4'b0000;
												assign node10260 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node10263 = (inp[13]) ? node10265 : 4'b0001;
												assign node10265 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node10268 = (inp[5]) ? node10274 : node10269;
											assign node10269 = (inp[10]) ? 4'b0001 : node10270;
												assign node10270 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node10274 = (inp[12]) ? node10276 : 4'b0000;
												assign node10276 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node10279 = (inp[5]) ? node10295 : node10280;
										assign node10280 = (inp[10]) ? node10288 : node10281;
											assign node10281 = (inp[2]) ? 4'b0101 : node10282;
												assign node10282 = (inp[0]) ? node10284 : 4'b0101;
													assign node10284 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node10288 = (inp[12]) ? node10292 : node10289;
												assign node10289 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node10292 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node10295 = (inp[10]) ? node10303 : node10296;
											assign node10296 = (inp[0]) ? node10300 : node10297;
												assign node10297 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node10300 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node10303 = (inp[12]) ? node10307 : node10304;
												assign node10304 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node10307 = (inp[0]) ? 4'b0100 : 4'b0101;
								assign node10310 = (inp[13]) ? node10334 : node10311;
									assign node10311 = (inp[12]) ? node10323 : node10312;
										assign node10312 = (inp[0]) ? node10318 : node10313;
											assign node10313 = (inp[5]) ? node10315 : 4'b0100;
												assign node10315 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node10318 = (inp[7]) ? 4'b0101 : node10319;
												assign node10319 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node10323 = (inp[0]) ? node10329 : node10324;
											assign node10324 = (inp[5]) ? 4'b0101 : node10325;
												assign node10325 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node10329 = (inp[5]) ? 4'b0100 : node10330;
												assign node10330 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node10334 = (inp[2]) ? node10352 : node10335;
										assign node10335 = (inp[0]) ? node10341 : node10336;
											assign node10336 = (inp[12]) ? 4'b0101 : node10337;
												assign node10337 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node10341 = (inp[12]) ? node10347 : node10342;
												assign node10342 = (inp[5]) ? 4'b0101 : node10343;
													assign node10343 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node10347 = (inp[5]) ? 4'b0100 : node10348;
													assign node10348 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node10352 = (inp[12]) ? node10362 : node10353;
											assign node10353 = (inp[0]) ? node10359 : node10354;
												assign node10354 = (inp[5]) ? 4'b0100 : node10355;
													assign node10355 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node10359 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node10362 = (inp[9]) ? node10374 : node10363;
												assign node10363 = (inp[7]) ? node10371 : node10364;
													assign node10364 = (inp[5]) ? node10368 : node10365;
														assign node10365 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node10368 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node10371 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node10374 = (inp[7]) ? 4'b0101 : node10375;
													assign node10375 = (inp[10]) ? 4'b0101 : node10376;
														assign node10376 = (inp[0]) ? 4'b0101 : 4'b0100;
							assign node10381 = (inp[15]) ? node10459 : node10382;
								assign node10382 = (inp[7]) ? node10406 : node10383;
									assign node10383 = (inp[5]) ? node10395 : node10384;
										assign node10384 = (inp[0]) ? node10390 : node10385;
											assign node10385 = (inp[13]) ? 4'b0100 : node10386;
												assign node10386 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node10390 = (inp[12]) ? node10392 : 4'b0101;
												assign node10392 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node10395 = (inp[0]) ? node10401 : node10396;
											assign node10396 = (inp[13]) ? 4'b0101 : node10397;
												assign node10397 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node10401 = (inp[12]) ? node10403 : 4'b0100;
												assign node10403 = (inp[13]) ? 4'b0100 : 4'b0101;
									assign node10406 = (inp[11]) ? node10432 : node10407;
										assign node10407 = (inp[10]) ? node10415 : node10408;
											assign node10408 = (inp[0]) ? node10412 : node10409;
												assign node10409 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node10412 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node10415 = (inp[9]) ? node10427 : node10416;
												assign node10416 = (inp[5]) ? node10422 : node10417;
													assign node10417 = (inp[2]) ? node10419 : 4'b0001;
														assign node10419 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node10422 = (inp[13]) ? 4'b0001 : node10423;
														assign node10423 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node10427 = (inp[0]) ? node10429 : 4'b0001;
													assign node10429 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node10432 = (inp[12]) ? node10454 : node10433;
											assign node10433 = (inp[10]) ? node10445 : node10434;
												assign node10434 = (inp[9]) ? node10436 : 4'b0001;
													assign node10436 = (inp[2]) ? node10440 : node10437;
														assign node10437 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node10440 = (inp[13]) ? node10442 : 4'b0000;
															assign node10442 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node10445 = (inp[5]) ? node10449 : node10446;
													assign node10446 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node10449 = (inp[2]) ? node10451 : 4'b0000;
														assign node10451 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node10454 = (inp[13]) ? 4'b0000 : node10455;
												assign node10455 = (inp[5]) ? 4'b0001 : 4'b0000;
								assign node10459 = (inp[0]) ? node10473 : node10460;
									assign node10460 = (inp[7]) ? 4'b0001 : node10461;
										assign node10461 = (inp[12]) ? node10469 : node10462;
											assign node10462 = (inp[13]) ? node10466 : node10463;
												assign node10463 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node10466 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node10469 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node10473 = (inp[7]) ? 4'b0000 : node10474;
										assign node10474 = (inp[5]) ? node10480 : node10475;
											assign node10475 = (inp[12]) ? 4'b0001 : node10476;
												assign node10476 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node10480 = (inp[13]) ? 4'b0000 : node10481;
												assign node10481 = (inp[12]) ? 4'b0000 : 4'b0001;
		assign node10486 = (inp[8]) ? node15542 : node10487;
			assign node10487 = (inp[14]) ? node13195 : node10488;
				assign node10488 = (inp[7]) ? node11828 : node10489;
					assign node10489 = (inp[15]) ? node11177 : node10490;
						assign node10490 = (inp[6]) ? node10878 : node10491;
							assign node10491 = (inp[0]) ? node10687 : node10492;
								assign node10492 = (inp[9]) ? node10570 : node10493;
									assign node10493 = (inp[4]) ? node10527 : node10494;
										assign node10494 = (inp[12]) ? node10518 : node10495;
											assign node10495 = (inp[13]) ? node10505 : node10496;
												assign node10496 = (inp[10]) ? node10500 : node10497;
													assign node10497 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node10500 = (inp[2]) ? 4'b1101 : node10501;
														assign node10501 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node10505 = (inp[10]) ? node10513 : node10506;
													assign node10506 = (inp[2]) ? node10510 : node10507;
														assign node10507 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node10510 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node10513 = (inp[5]) ? 4'b1000 : node10514;
														assign node10514 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node10518 = (inp[5]) ? 4'b1011 : node10519;
												assign node10519 = (inp[2]) ? node10521 : 4'b1111;
													assign node10521 = (inp[1]) ? 4'b1111 : node10522;
														assign node10522 = (inp[13]) ? 4'b1010 : 4'b1111;
										assign node10527 = (inp[12]) ? node10545 : node10528;
											assign node10528 = (inp[2]) ? node10536 : node10529;
												assign node10529 = (inp[13]) ? node10531 : 4'b1011;
													assign node10531 = (inp[5]) ? 4'b1110 : node10532;
														assign node10532 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node10536 = (inp[11]) ? node10542 : node10537;
													assign node10537 = (inp[1]) ? 4'b1010 : node10538;
														assign node10538 = (inp[13]) ? 4'b1010 : 4'b1111;
													assign node10542 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node10545 = (inp[2]) ? node10561 : node10546;
												assign node10546 = (inp[13]) ? node10556 : node10547;
													assign node10547 = (inp[1]) ? node10553 : node10548;
														assign node10548 = (inp[5]) ? node10550 : 4'b1100;
															assign node10550 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node10553 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node10556 = (inp[10]) ? node10558 : 4'b1001;
														assign node10558 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node10561 = (inp[13]) ? node10567 : node10562;
													assign node10562 = (inp[1]) ? 4'b1000 : node10563;
														assign node10563 = (inp[11]) ? 4'b1000 : 4'b1100;
													assign node10567 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node10570 = (inp[10]) ? node10638 : node10571;
										assign node10571 = (inp[5]) ? node10603 : node10572;
											assign node10572 = (inp[12]) ? node10586 : node10573;
												assign node10573 = (inp[4]) ? node10579 : node10574;
													assign node10574 = (inp[13]) ? 4'b1100 : node10575;
														assign node10575 = (inp[11]) ? 4'b1101 : 4'b1001;
													assign node10579 = (inp[1]) ? node10581 : 4'b1011;
														assign node10581 = (inp[13]) ? 4'b1111 : node10582;
															assign node10582 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node10586 = (inp[4]) ? node10596 : node10587;
													assign node10587 = (inp[2]) ? 4'b1010 : node10588;
														assign node10588 = (inp[1]) ? node10592 : node10589;
															assign node10589 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node10592 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node10596 = (inp[2]) ? node10600 : node10597;
														assign node10597 = (inp[11]) ? 4'b1101 : 4'b1001;
														assign node10600 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node10603 = (inp[1]) ? node10621 : node10604;
												assign node10604 = (inp[13]) ? node10612 : node10605;
													assign node10605 = (inp[2]) ? node10609 : node10606;
														assign node10606 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node10609 = (inp[11]) ? 4'b1101 : 4'b1110;
													assign node10612 = (inp[2]) ? node10618 : node10613;
														assign node10613 = (inp[4]) ? 4'b1100 : node10614;
															assign node10614 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10618 = (inp[11]) ? 4'b1010 : 4'b1000;
												assign node10621 = (inp[11]) ? node10633 : node10622;
													assign node10622 = (inp[13]) ? node10628 : node10623;
														assign node10623 = (inp[2]) ? node10625 : 4'b1010;
															assign node10625 = (inp[12]) ? 4'b1110 : 4'b1111;
														assign node10628 = (inp[12]) ? 4'b1111 : node10629;
															assign node10629 = (inp[4]) ? 4'b1110 : 4'b1100;
													assign node10633 = (inp[2]) ? 4'b1100 : node10634;
														assign node10634 = (inp[12]) ? 4'b1101 : 4'b1111;
										assign node10638 = (inp[1]) ? node10656 : node10639;
											assign node10639 = (inp[11]) ? node10649 : node10640;
												assign node10640 = (inp[12]) ? node10642 : 4'b1010;
													assign node10642 = (inp[4]) ? node10646 : node10643;
														assign node10643 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node10646 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node10649 = (inp[4]) ? 4'b1111 : node10650;
													assign node10650 = (inp[5]) ? 4'b1101 : node10651;
														assign node10651 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node10656 = (inp[13]) ? node10678 : node10657;
												assign node10657 = (inp[2]) ? node10669 : node10658;
													assign node10658 = (inp[5]) ? node10664 : node10659;
														assign node10659 = (inp[11]) ? 4'b1100 : node10660;
															assign node10660 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node10664 = (inp[12]) ? 4'b1100 : node10665;
															assign node10665 = (inp[4]) ? 4'b1011 : 4'b1000;
													assign node10669 = (inp[12]) ? node10675 : node10670;
														assign node10670 = (inp[4]) ? 4'b1010 : node10671;
															assign node10671 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10675 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node10678 = (inp[5]) ? node10684 : node10679;
													assign node10679 = (inp[12]) ? node10681 : 4'b1001;
														assign node10681 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node10684 = (inp[2]) ? 4'b1011 : 4'b1001;
								assign node10687 = (inp[4]) ? node10781 : node10688;
									assign node10688 = (inp[12]) ? node10720 : node10689;
										assign node10689 = (inp[1]) ? node10695 : node10690;
											assign node10690 = (inp[2]) ? node10692 : 4'b1000;
												assign node10692 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node10695 = (inp[5]) ? node10705 : node10696;
												assign node10696 = (inp[9]) ? node10700 : node10697;
													assign node10697 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node10700 = (inp[13]) ? 4'b1101 : node10701;
														assign node10701 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node10705 = (inp[2]) ? node10713 : node10706;
													assign node10706 = (inp[13]) ? node10708 : 4'b1000;
														assign node10708 = (inp[9]) ? 4'b1100 : node10709;
															assign node10709 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node10713 = (inp[13]) ? node10717 : node10714;
														assign node10714 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node10717 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node10720 = (inp[2]) ? node10752 : node10721;
											assign node10721 = (inp[9]) ? node10739 : node10722;
												assign node10722 = (inp[5]) ? node10736 : node10723;
													assign node10723 = (inp[11]) ? node10727 : node10724;
														assign node10724 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node10727 = (inp[10]) ? node10731 : node10728;
															assign node10728 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node10731 = (inp[13]) ? 4'b1011 : node10732;
																assign node10732 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node10736 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node10739 = (inp[13]) ? node10749 : node10740;
													assign node10740 = (inp[1]) ? node10746 : node10741;
														assign node10741 = (inp[11]) ? node10743 : 4'b1010;
															assign node10743 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node10746 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node10749 = (inp[11]) ? 4'b1010 : 4'b1110;
											assign node10752 = (inp[13]) ? node10770 : node10753;
												assign node10753 = (inp[11]) ? node10761 : node10754;
													assign node10754 = (inp[10]) ? 4'b1110 : node10755;
														assign node10755 = (inp[9]) ? 4'b1110 : node10756;
															assign node10756 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node10761 = (inp[10]) ? node10767 : node10762;
														assign node10762 = (inp[9]) ? node10764 : 4'b1111;
															assign node10764 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node10767 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node10770 = (inp[9]) ? node10778 : node10771;
													assign node10771 = (inp[11]) ? node10773 : 4'b1010;
														assign node10773 = (inp[5]) ? 4'b1011 : node10774;
															assign node10774 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node10778 = (inp[1]) ? 4'b1111 : 4'b1011;
									assign node10781 = (inp[12]) ? node10833 : node10782;
										assign node10782 = (inp[13]) ? node10812 : node10783;
											assign node10783 = (inp[11]) ? node10803 : node10784;
												assign node10784 = (inp[10]) ? node10796 : node10785;
													assign node10785 = (inp[2]) ? node10791 : node10786;
														assign node10786 = (inp[1]) ? node10788 : 4'b1010;
															assign node10788 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node10791 = (inp[1]) ? node10793 : 4'b1111;
															assign node10793 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node10796 = (inp[2]) ? node10798 : 4'b1111;
														assign node10798 = (inp[5]) ? 4'b1110 : node10799;
															assign node10799 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node10803 = (inp[2]) ? 4'b1111 : node10804;
													assign node10804 = (inp[5]) ? node10808 : node10805;
														assign node10805 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node10808 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node10812 = (inp[2]) ? node10824 : node10813;
												assign node10813 = (inp[1]) ? node10819 : node10814;
													assign node10814 = (inp[5]) ? 4'b1111 : node10815;
														assign node10815 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node10819 = (inp[5]) ? 4'b1110 : node10820;
														assign node10820 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node10824 = (inp[5]) ? node10828 : node10825;
													assign node10825 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node10828 = (inp[1]) ? node10830 : 4'b1010;
														assign node10830 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node10833 = (inp[10]) ? node10863 : node10834;
											assign node10834 = (inp[5]) ? node10854 : node10835;
												assign node10835 = (inp[1]) ? node10847 : node10836;
													assign node10836 = (inp[2]) ? node10844 : node10837;
														assign node10837 = (inp[13]) ? 4'b1001 : node10838;
															assign node10838 = (inp[9]) ? 4'b1100 : node10839;
																assign node10839 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10844 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node10847 = (inp[11]) ? node10849 : 4'b1000;
														assign node10849 = (inp[13]) ? 4'b1101 : node10850;
															assign node10850 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node10854 = (inp[9]) ? node10856 : 4'b1100;
													assign node10856 = (inp[2]) ? node10858 : 4'b1100;
														assign node10858 = (inp[1]) ? 4'b1000 : node10859;
															assign node10859 = (inp[13]) ? 4'b1000 : 4'b1100;
											assign node10863 = (inp[11]) ? node10873 : node10864;
												assign node10864 = (inp[5]) ? 4'b1101 : node10865;
													assign node10865 = (inp[9]) ? node10867 : 4'b1001;
														assign node10867 = (inp[2]) ? node10869 : 4'b1000;
															assign node10869 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node10873 = (inp[13]) ? 4'b1101 : node10874;
													assign node10874 = (inp[9]) ? 4'b1001 : 4'b1101;
							assign node10878 = (inp[12]) ? node11028 : node10879;
								assign node10879 = (inp[13]) ? node10973 : node10880;
									assign node10880 = (inp[5]) ? node10928 : node10881;
										assign node10881 = (inp[1]) ? node10911 : node10882;
											assign node10882 = (inp[2]) ? node10898 : node10883;
												assign node10883 = (inp[10]) ? node10891 : node10884;
													assign node10884 = (inp[4]) ? node10888 : node10885;
														assign node10885 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node10888 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node10891 = (inp[11]) ? node10893 : 4'b1001;
														assign node10893 = (inp[0]) ? 4'b1001 : node10894;
															assign node10894 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node10898 = (inp[4]) ? 4'b1000 : node10899;
													assign node10899 = (inp[0]) ? node10901 : 4'b1000;
														assign node10901 = (inp[10]) ? 4'b1000 : node10902;
															assign node10902 = (inp[9]) ? node10906 : node10903;
																assign node10903 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node10906 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node10911 = (inp[4]) ? node10919 : node10912;
												assign node10912 = (inp[2]) ? node10914 : 4'b1100;
													assign node10914 = (inp[9]) ? node10916 : 4'b1101;
														assign node10916 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node10919 = (inp[11]) ? 4'b1000 : node10920;
													assign node10920 = (inp[9]) ? node10922 : 4'b1000;
														assign node10922 = (inp[0]) ? node10924 : 4'b1001;
															assign node10924 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node10928 = (inp[1]) ? node10954 : node10929;
											assign node10929 = (inp[9]) ? node10935 : node10930;
												assign node10930 = (inp[11]) ? node10932 : 4'b1100;
													assign node10932 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node10935 = (inp[10]) ? node10949 : node10936;
													assign node10936 = (inp[4]) ? 4'b1100 : node10937;
														assign node10937 = (inp[11]) ? node10943 : node10938;
															assign node10938 = (inp[2]) ? 4'b1101 : node10939;
																assign node10939 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node10943 = (inp[0]) ? node10945 : 4'b1100;
																assign node10945 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node10949 = (inp[0]) ? 4'b1101 : node10950;
														assign node10950 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node10954 = (inp[4]) ? node10966 : node10955;
												assign node10955 = (inp[10]) ? 4'b1000 : node10956;
													assign node10956 = (inp[9]) ? node10962 : node10957;
														assign node10957 = (inp[11]) ? node10959 : 4'b1000;
															assign node10959 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node10962 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node10966 = (inp[0]) ? node10970 : node10967;
													assign node10967 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node10970 = (inp[10]) ? 4'b1100 : 4'b1101;
									assign node10973 = (inp[5]) ? node10999 : node10974;
										assign node10974 = (inp[4]) ? node10986 : node10975;
											assign node10975 = (inp[1]) ? node10979 : node10976;
												assign node10976 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node10979 = (inp[2]) ? 4'b1001 : node10980;
													assign node10980 = (inp[11]) ? node10982 : 4'b1000;
														assign node10982 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node10986 = (inp[0]) ? node10988 : 4'b1100;
												assign node10988 = (inp[9]) ? node10994 : node10989;
													assign node10989 = (inp[11]) ? node10991 : 4'b1100;
														assign node10991 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node10994 = (inp[11]) ? node10996 : 4'b1101;
														assign node10996 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node10999 = (inp[1]) ? node11015 : node11000;
											assign node11000 = (inp[10]) ? node11008 : node11001;
												assign node11001 = (inp[2]) ? 4'b1001 : node11002;
													assign node11002 = (inp[9]) ? node11004 : 4'b1000;
														assign node11004 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node11008 = (inp[9]) ? 4'b1000 : node11009;
													assign node11009 = (inp[11]) ? node11011 : 4'b1001;
														assign node11011 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node11015 = (inp[4]) ? node11021 : node11016;
												assign node11016 = (inp[9]) ? 4'b1100 : node11017;
													assign node11017 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node11021 = (inp[9]) ? 4'b1001 : node11022;
													assign node11022 = (inp[10]) ? 4'b1000 : node11023;
														assign node11023 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node11028 = (inp[5]) ? node11104 : node11029;
									assign node11029 = (inp[13]) ? node11071 : node11030;
										assign node11030 = (inp[4]) ? node11052 : node11031;
											assign node11031 = (inp[10]) ? node11045 : node11032;
												assign node11032 = (inp[11]) ? node11040 : node11033;
													assign node11033 = (inp[0]) ? 4'b1000 : node11034;
														assign node11034 = (inp[9]) ? node11036 : 4'b1000;
															assign node11036 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node11040 = (inp[1]) ? 4'b1001 : node11041;
														assign node11041 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node11045 = (inp[11]) ? node11047 : 4'b1001;
													assign node11047 = (inp[1]) ? node11049 : 4'b1000;
														assign node11049 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node11052 = (inp[1]) ? node11066 : node11053;
												assign node11053 = (inp[0]) ? node11055 : 4'b1000;
													assign node11055 = (inp[9]) ? 4'b1001 : node11056;
														assign node11056 = (inp[10]) ? node11060 : node11057;
															assign node11057 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node11060 = (inp[2]) ? 4'b1001 : node11061;
																assign node11061 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node11066 = (inp[9]) ? node11068 : 4'b1101;
													assign node11068 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node11071 = (inp[1]) ? node11093 : node11072;
											assign node11072 = (inp[2]) ? node11080 : node11073;
												assign node11073 = (inp[4]) ? node11075 : 4'b1100;
													assign node11075 = (inp[9]) ? node11077 : 4'b1101;
														assign node11077 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node11080 = (inp[4]) ? node11090 : node11081;
													assign node11081 = (inp[10]) ? node11083 : 4'b1101;
														assign node11083 = (inp[0]) ? node11087 : node11084;
															assign node11084 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node11087 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node11090 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node11093 = (inp[4]) ? node11099 : node11094;
												assign node11094 = (inp[9]) ? 4'b1101 : node11095;
													assign node11095 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node11099 = (inp[9]) ? 4'b1000 : node11100;
													assign node11100 = (inp[2]) ? 4'b1001 : 4'b1000;
									assign node11104 = (inp[13]) ? node11144 : node11105;
										assign node11105 = (inp[1]) ? node11125 : node11106;
											assign node11106 = (inp[2]) ? node11118 : node11107;
												assign node11107 = (inp[4]) ? node11109 : 4'b1101;
													assign node11109 = (inp[0]) ? 4'b1101 : node11110;
														assign node11110 = (inp[11]) ? node11114 : node11111;
															assign node11111 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node11114 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node11118 = (inp[4]) ? 4'b1101 : node11119;
													assign node11119 = (inp[10]) ? node11121 : 4'b1100;
														assign node11121 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node11125 = (inp[4]) ? node11131 : node11126;
												assign node11126 = (inp[9]) ? node11128 : 4'b1101;
													assign node11128 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node11131 = (inp[9]) ? node11135 : node11132;
													assign node11132 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11135 = (inp[0]) ? node11137 : 4'b1000;
														assign node11137 = (inp[10]) ? node11139 : 4'b1000;
															assign node11139 = (inp[2]) ? node11141 : 4'b1001;
																assign node11141 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node11144 = (inp[4]) ? node11162 : node11145;
											assign node11145 = (inp[1]) ? node11157 : node11146;
												assign node11146 = (inp[2]) ? node11152 : node11147;
													assign node11147 = (inp[11]) ? node11149 : 4'b1000;
														assign node11149 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node11152 = (inp[11]) ? node11154 : 4'b1001;
														assign node11154 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node11157 = (inp[2]) ? 4'b1000 : node11158;
													assign node11158 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node11162 = (inp[1]) ? 4'b1101 : node11163;
												assign node11163 = (inp[2]) ? node11171 : node11164;
													assign node11164 = (inp[11]) ? node11166 : 4'b1001;
														assign node11166 = (inp[0]) ? 4'b1001 : node11167;
															assign node11167 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node11171 = (inp[9]) ? node11173 : 4'b1000;
														assign node11173 = (inp[0]) ? 4'b1000 : 4'b1001;
						assign node11177 = (inp[6]) ? node11519 : node11178;
							assign node11178 = (inp[12]) ? node11372 : node11179;
								assign node11179 = (inp[10]) ? node11287 : node11180;
									assign node11180 = (inp[9]) ? node11238 : node11181;
										assign node11181 = (inp[2]) ? node11199 : node11182;
											assign node11182 = (inp[4]) ? node11188 : node11183;
												assign node11183 = (inp[13]) ? node11185 : 4'b1000;
													assign node11185 = (inp[1]) ? 4'b1000 : 4'b1101;
												assign node11188 = (inp[13]) ? node11194 : node11189;
													assign node11189 = (inp[1]) ? node11191 : 4'b1100;
														assign node11191 = (inp[0]) ? 4'b1001 : 4'b1100;
													assign node11194 = (inp[1]) ? node11196 : 4'b1000;
														assign node11196 = (inp[5]) ? 4'b1001 : 4'b1100;
											assign node11199 = (inp[13]) ? node11221 : node11200;
												assign node11200 = (inp[5]) ? node11210 : node11201;
													assign node11201 = (inp[4]) ? node11205 : node11202;
														assign node11202 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node11205 = (inp[1]) ? node11207 : 4'b1001;
															assign node11207 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node11210 = (inp[4]) ? 4'b1000 : node11211;
														assign node11211 = (inp[11]) ? 4'b1101 : node11212;
															assign node11212 = (inp[0]) ? node11216 : node11213;
																assign node11213 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node11216 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node11221 = (inp[4]) ? node11227 : node11222;
													assign node11222 = (inp[5]) ? node11224 : 4'b1100;
														assign node11224 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node11227 = (inp[1]) ? node11231 : node11228;
														assign node11228 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node11231 = (inp[5]) ? node11233 : 4'b1000;
															assign node11233 = (inp[0]) ? 4'b1100 : node11234;
																assign node11234 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node11238 = (inp[0]) ? node11262 : node11239;
											assign node11239 = (inp[1]) ? node11251 : node11240;
												assign node11240 = (inp[5]) ? node11246 : node11241;
													assign node11241 = (inp[2]) ? 4'b1101 : node11242;
														assign node11242 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node11246 = (inp[11]) ? node11248 : 4'b1001;
														assign node11248 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node11251 = (inp[4]) ? node11259 : node11252;
													assign node11252 = (inp[11]) ? 4'b1100 : node11253;
														assign node11253 = (inp[2]) ? node11255 : 4'b1101;
															assign node11255 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node11259 = (inp[11]) ? 4'b1001 : 4'b1101;
											assign node11262 = (inp[1]) ? node11276 : node11263;
												assign node11263 = (inp[13]) ? node11271 : node11264;
													assign node11264 = (inp[4]) ? 4'b1101 : node11265;
														assign node11265 = (inp[11]) ? 4'b1101 : node11266;
															assign node11266 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node11271 = (inp[11]) ? 4'b1100 : node11272;
														assign node11272 = (inp[5]) ? 4'b1100 : 4'b1000;
												assign node11276 = (inp[4]) ? node11284 : node11277;
													assign node11277 = (inp[5]) ? 4'b1101 : node11278;
														assign node11278 = (inp[2]) ? node11280 : 4'b1001;
															assign node11280 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node11284 = (inp[13]) ? 4'b1101 : 4'b1000;
									assign node11287 = (inp[9]) ? node11329 : node11288;
										assign node11288 = (inp[0]) ? node11304 : node11289;
											assign node11289 = (inp[1]) ? node11297 : node11290;
												assign node11290 = (inp[4]) ? node11292 : 4'b1001;
													assign node11292 = (inp[2]) ? 4'b1100 : node11293;
														assign node11293 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node11297 = (inp[4]) ? node11301 : node11298;
													assign node11298 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node11301 = (inp[13]) ? 4'b1001 : 4'b1000;
											assign node11304 = (inp[2]) ? node11314 : node11305;
												assign node11305 = (inp[4]) ? 4'b1001 : node11306;
													assign node11306 = (inp[1]) ? node11308 : 4'b1100;
														assign node11308 = (inp[13]) ? 4'b1101 : node11309;
															assign node11309 = (inp[5]) ? 4'b1001 : 4'b1101;
												assign node11314 = (inp[11]) ? node11320 : node11315;
													assign node11315 = (inp[4]) ? 4'b1000 : node11316;
														assign node11316 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node11320 = (inp[4]) ? 4'b1101 : node11321;
														assign node11321 = (inp[1]) ? node11325 : node11322;
															assign node11322 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node11325 = (inp[13]) ? 4'b1101 : 4'b1000;
										assign node11329 = (inp[4]) ? node11359 : node11330;
											assign node11330 = (inp[5]) ? node11344 : node11331;
												assign node11331 = (inp[11]) ? node11341 : node11332;
													assign node11332 = (inp[13]) ? node11338 : node11333;
														assign node11333 = (inp[0]) ? 4'b1001 : node11334;
															assign node11334 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node11338 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node11341 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node11344 = (inp[0]) ? node11350 : node11345;
													assign node11345 = (inp[2]) ? 4'b1000 : node11346;
														assign node11346 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node11350 = (inp[13]) ? 4'b1001 : node11351;
														assign node11351 = (inp[2]) ? 4'b1100 : node11352;
															assign node11352 = (inp[11]) ? node11354 : 4'b1000;
																assign node11354 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node11359 = (inp[0]) ? node11365 : node11360;
												assign node11360 = (inp[13]) ? 4'b1101 : node11361;
													assign node11361 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node11365 = (inp[1]) ? 4'b1100 : node11366;
													assign node11366 = (inp[13]) ? 4'b1000 : node11367;
														assign node11367 = (inp[2]) ? 4'b1000 : 4'b1100;
								assign node11372 = (inp[0]) ? node11450 : node11373;
									assign node11373 = (inp[2]) ? node11413 : node11374;
										assign node11374 = (inp[10]) ? node11392 : node11375;
											assign node11375 = (inp[5]) ? 4'b1010 : node11376;
												assign node11376 = (inp[9]) ? node11388 : node11377;
													assign node11377 = (inp[4]) ? node11383 : node11378;
														assign node11378 = (inp[11]) ? 4'b1010 : node11379;
															assign node11379 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node11383 = (inp[1]) ? node11385 : 4'b1110;
															assign node11385 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node11388 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node11392 = (inp[4]) ? node11402 : node11393;
												assign node11393 = (inp[9]) ? node11395 : 4'b1011;
													assign node11395 = (inp[11]) ? node11397 : 4'b1011;
														assign node11397 = (inp[5]) ? node11399 : 4'b1010;
															assign node11399 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node11402 = (inp[1]) ? node11406 : node11403;
													assign node11403 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node11406 = (inp[5]) ? node11410 : node11407;
														assign node11407 = (inp[13]) ? 4'b1011 : 4'b1110;
														assign node11410 = (inp[9]) ? 4'b1011 : 4'b1110;
										assign node11413 = (inp[13]) ? node11433 : node11414;
											assign node11414 = (inp[1]) ? node11424 : node11415;
												assign node11415 = (inp[4]) ? node11417 : 4'b1110;
													assign node11417 = (inp[5]) ? node11419 : 4'b1111;
														assign node11419 = (inp[10]) ? node11421 : 4'b1110;
															assign node11421 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node11424 = (inp[5]) ? 4'b1111 : node11425;
													assign node11425 = (inp[4]) ? node11427 : 4'b1010;
														assign node11427 = (inp[9]) ? 4'b1011 : node11428;
															assign node11428 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node11433 = (inp[1]) ? node11443 : node11434;
												assign node11434 = (inp[11]) ? node11438 : node11435;
													assign node11435 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node11438 = (inp[9]) ? 4'b1011 : node11439;
														assign node11439 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node11443 = (inp[5]) ? 4'b1010 : node11444;
													assign node11444 = (inp[10]) ? 4'b1111 : node11445;
														assign node11445 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node11450 = (inp[2]) ? node11484 : node11451;
										assign node11451 = (inp[13]) ? node11469 : node11452;
											assign node11452 = (inp[5]) ? node11462 : node11453;
												assign node11453 = (inp[1]) ? node11457 : node11454;
													assign node11454 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node11457 = (inp[4]) ? 4'b1111 : node11458;
														assign node11458 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node11462 = (inp[9]) ? node11466 : node11463;
													assign node11463 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11466 = (inp[4]) ? 4'b1011 : 4'b1010;
											assign node11469 = (inp[1]) ? node11479 : node11470;
												assign node11470 = (inp[5]) ? node11476 : node11471;
													assign node11471 = (inp[10]) ? node11473 : 4'b1110;
														assign node11473 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node11476 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node11479 = (inp[5]) ? node11481 : 4'b1011;
													assign node11481 = (inp[10]) ? 4'b1111 : 4'b1110;
										assign node11484 = (inp[13]) ? node11504 : node11485;
											assign node11485 = (inp[5]) ? node11493 : node11486;
												assign node11486 = (inp[1]) ? node11488 : 4'b1110;
													assign node11488 = (inp[11]) ? 4'b1010 : node11489;
														assign node11489 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node11493 = (inp[4]) ? node11495 : 4'b1110;
													assign node11495 = (inp[1]) ? node11497 : 4'b1111;
														assign node11497 = (inp[9]) ? node11499 : 4'b1110;
															assign node11499 = (inp[11]) ? 4'b1110 : node11500;
																assign node11500 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node11504 = (inp[1]) ? node11510 : node11505;
												assign node11505 = (inp[4]) ? node11507 : 4'b1011;
													assign node11507 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node11510 = (inp[5]) ? node11516 : node11511;
													assign node11511 = (inp[11]) ? node11513 : 4'b1110;
														assign node11513 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node11516 = (inp[11]) ? 4'b1010 : 4'b1011;
							assign node11519 = (inp[11]) ? node11673 : node11520;
								assign node11520 = (inp[13]) ? node11602 : node11521;
									assign node11521 = (inp[5]) ? node11561 : node11522;
										assign node11522 = (inp[12]) ? node11548 : node11523;
											assign node11523 = (inp[10]) ? node11539 : node11524;
												assign node11524 = (inp[0]) ? node11532 : node11525;
													assign node11525 = (inp[1]) ? node11529 : node11526;
														assign node11526 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node11529 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node11532 = (inp[9]) ? node11536 : node11533;
														assign node11533 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node11536 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node11539 = (inp[2]) ? node11541 : 4'b1010;
													assign node11541 = (inp[1]) ? node11543 : 4'b1110;
														assign node11543 = (inp[9]) ? 4'b1011 : node11544;
															assign node11544 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node11548 = (inp[4]) ? 4'b1010 : node11549;
												assign node11549 = (inp[0]) ? node11551 : 4'b1010;
													assign node11551 = (inp[1]) ? node11557 : node11552;
														assign node11552 = (inp[2]) ? 4'b1010 : node11553;
															assign node11553 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node11557 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node11561 = (inp[12]) ? node11581 : node11562;
											assign node11562 = (inp[0]) ? node11572 : node11563;
												assign node11563 = (inp[4]) ? node11569 : node11564;
													assign node11564 = (inp[1]) ? node11566 : 4'b1110;
														assign node11566 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node11569 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node11572 = (inp[1]) ? node11578 : node11573;
													assign node11573 = (inp[9]) ? 4'b1110 : node11574;
														assign node11574 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node11578 = (inp[4]) ? 4'b1110 : 4'b1011;
											assign node11581 = (inp[9]) ? node11587 : node11582;
												assign node11582 = (inp[2]) ? 4'b1110 : node11583;
													assign node11583 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node11587 = (inp[2]) ? 4'b1111 : node11588;
													assign node11588 = (inp[10]) ? node11594 : node11589;
														assign node11589 = (inp[1]) ? 4'b1110 : node11590;
															assign node11590 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node11594 = (inp[4]) ? node11598 : node11595;
															assign node11595 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node11598 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node11602 = (inp[5]) ? node11642 : node11603;
										assign node11603 = (inp[9]) ? node11627 : node11604;
											assign node11604 = (inp[12]) ? node11614 : node11605;
												assign node11605 = (inp[1]) ? node11609 : node11606;
													assign node11606 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11609 = (inp[4]) ? 4'b1110 : node11610;
														assign node11610 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node11614 = (inp[0]) ? 4'b1111 : node11615;
													assign node11615 = (inp[1]) ? node11621 : node11616;
														assign node11616 = (inp[4]) ? 4'b1110 : node11617;
															assign node11617 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node11621 = (inp[10]) ? 4'b1111 : node11622;
															assign node11622 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node11627 = (inp[0]) ? node11637 : node11628;
												assign node11628 = (inp[4]) ? 4'b1111 : node11629;
													assign node11629 = (inp[2]) ? 4'b1111 : node11630;
														assign node11630 = (inp[12]) ? 4'b1110 : node11631;
															assign node11631 = (inp[1]) ? 4'b1011 : 4'b1110;
												assign node11637 = (inp[12]) ? 4'b1110 : node11638;
													assign node11638 = (inp[2]) ? 4'b1110 : 4'b1010;
										assign node11642 = (inp[12]) ? node11660 : node11643;
											assign node11643 = (inp[4]) ? node11653 : node11644;
												assign node11644 = (inp[1]) ? node11650 : node11645;
													assign node11645 = (inp[9]) ? node11647 : 4'b1011;
														assign node11647 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node11650 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node11653 = (inp[1]) ? 4'b1010 : node11654;
													assign node11654 = (inp[9]) ? node11656 : 4'b1110;
														assign node11656 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node11660 = (inp[1]) ? node11666 : node11661;
												assign node11661 = (inp[2]) ? node11663 : 4'b1011;
													assign node11663 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node11666 = (inp[10]) ? node11668 : 4'b1010;
													assign node11668 = (inp[2]) ? 4'b1011 : node11669;
														assign node11669 = (inp[0]) ? 4'b1010 : 4'b1011;
								assign node11673 = (inp[12]) ? node11759 : node11674;
									assign node11674 = (inp[9]) ? node11722 : node11675;
										assign node11675 = (inp[1]) ? node11703 : node11676;
											assign node11676 = (inp[10]) ? node11692 : node11677;
												assign node11677 = (inp[4]) ? node11685 : node11678;
													assign node11678 = (inp[0]) ? node11680 : 4'b1111;
														assign node11680 = (inp[5]) ? node11682 : 4'b1110;
															assign node11682 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node11685 = (inp[2]) ? 4'b1111 : node11686;
														assign node11686 = (inp[5]) ? node11688 : 4'b1011;
															assign node11688 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node11692 = (inp[2]) ? node11700 : node11693;
													assign node11693 = (inp[13]) ? node11697 : node11694;
														assign node11694 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node11697 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node11700 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node11703 = (inp[10]) ? node11717 : node11704;
												assign node11704 = (inp[5]) ? node11710 : node11705;
													assign node11705 = (inp[13]) ? 4'b1011 : node11706;
														assign node11706 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11710 = (inp[0]) ? node11712 : 4'b1010;
														assign node11712 = (inp[2]) ? 4'b1111 : node11713;
															assign node11713 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node11717 = (inp[4]) ? 4'b1110 : node11718;
													assign node11718 = (inp[5]) ? 4'b1010 : 4'b1111;
										assign node11722 = (inp[10]) ? node11730 : node11723;
											assign node11723 = (inp[2]) ? 4'b1010 : node11724;
												assign node11724 = (inp[0]) ? 4'b1110 : node11725;
													assign node11725 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node11730 = (inp[4]) ? node11746 : node11731;
												assign node11731 = (inp[5]) ? node11741 : node11732;
													assign node11732 = (inp[1]) ? node11738 : node11733;
														assign node11733 = (inp[13]) ? 4'b1111 : node11734;
															assign node11734 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node11738 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node11741 = (inp[0]) ? 4'b1010 : node11742;
														assign node11742 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node11746 = (inp[13]) ? node11750 : node11747;
													assign node11747 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node11750 = (inp[2]) ? node11756 : node11751;
														assign node11751 = (inp[0]) ? 4'b1011 : node11752;
															assign node11752 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node11756 = (inp[0]) ? 4'b1111 : 4'b1011;
									assign node11759 = (inp[9]) ? node11795 : node11760;
										assign node11760 = (inp[2]) ? node11782 : node11761;
											assign node11761 = (inp[13]) ? node11771 : node11762;
												assign node11762 = (inp[5]) ? node11768 : node11763;
													assign node11763 = (inp[10]) ? 4'b1011 : node11764;
														assign node11764 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node11768 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node11771 = (inp[5]) ? node11777 : node11772;
													assign node11772 = (inp[4]) ? node11774 : 4'b1110;
														assign node11774 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node11777 = (inp[4]) ? node11779 : 4'b1011;
														assign node11779 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node11782 = (inp[5]) ? node11792 : node11783;
												assign node11783 = (inp[13]) ? node11787 : node11784;
													assign node11784 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node11787 = (inp[0]) ? 4'b1110 : node11788;
														assign node11788 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node11792 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node11795 = (inp[0]) ? node11811 : node11796;
											assign node11796 = (inp[2]) ? node11806 : node11797;
												assign node11797 = (inp[13]) ? node11801 : node11798;
													assign node11798 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node11801 = (inp[5]) ? 4'b1011 : node11802;
														assign node11802 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node11806 = (inp[13]) ? node11808 : 4'b1110;
													assign node11808 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node11811 = (inp[2]) ? node11821 : node11812;
												assign node11812 = (inp[4]) ? node11818 : node11813;
													assign node11813 = (inp[13]) ? node11815 : 4'b1111;
														assign node11815 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node11818 = (inp[13]) ? 4'b1111 : 4'b1110;
												assign node11821 = (inp[5]) ? node11825 : node11822;
													assign node11822 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node11825 = (inp[1]) ? 4'b1110 : 4'b1010;
					assign node11828 = (inp[15]) ? node12512 : node11829;
						assign node11829 = (inp[6]) ? node12219 : node11830;
							assign node11830 = (inp[13]) ? node12008 : node11831;
								assign node11831 = (inp[1]) ? node11907 : node11832;
									assign node11832 = (inp[2]) ? node11860 : node11833;
										assign node11833 = (inp[9]) ? node11843 : node11834;
											assign node11834 = (inp[0]) ? node11838 : node11835;
												assign node11835 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node11838 = (inp[12]) ? 4'b1100 : node11839;
													assign node11839 = (inp[10]) ? 4'b1100 : 4'b1011;
											assign node11843 = (inp[11]) ? node11851 : node11844;
												assign node11844 = (inp[10]) ? 4'b1101 : node11845;
													assign node11845 = (inp[4]) ? 4'b1011 : node11846;
														assign node11846 = (inp[12]) ? 4'b1100 : 4'b1111;
												assign node11851 = (inp[10]) ? node11857 : node11852;
													assign node11852 = (inp[12]) ? 4'b1010 : node11853;
														assign node11853 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node11857 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node11860 = (inp[11]) ? node11884 : node11861;
											assign node11861 = (inp[9]) ? node11875 : node11862;
												assign node11862 = (inp[10]) ? node11870 : node11863;
													assign node11863 = (inp[12]) ? node11867 : node11864;
														assign node11864 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node11867 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node11870 = (inp[12]) ? 4'b1001 : node11871;
														assign node11871 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node11875 = (inp[10]) ? node11881 : node11876;
													assign node11876 = (inp[12]) ? node11878 : 4'b1000;
														assign node11878 = (inp[0]) ? 4'b1000 : 4'b1110;
													assign node11881 = (inp[4]) ? 4'b1001 : 4'b1111;
											assign node11884 = (inp[10]) ? node11890 : node11885;
												assign node11885 = (inp[4]) ? 4'b1001 : node11886;
													assign node11886 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node11890 = (inp[12]) ? node11902 : node11891;
													assign node11891 = (inp[4]) ? node11895 : node11892;
														assign node11892 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node11895 = (inp[0]) ? 4'b1000 : node11896;
															assign node11896 = (inp[9]) ? 4'b1000 : node11897;
																assign node11897 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node11902 = (inp[9]) ? node11904 : 4'b1000;
														assign node11904 = (inp[5]) ? 4'b1000 : 4'b1001;
									assign node11907 = (inp[2]) ? node11963 : node11908;
										assign node11908 = (inp[4]) ? node11936 : node11909;
											assign node11909 = (inp[12]) ? node11923 : node11910;
												assign node11910 = (inp[9]) ? node11918 : node11911;
													assign node11911 = (inp[10]) ? node11915 : node11912;
														assign node11912 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node11915 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node11918 = (inp[10]) ? 4'b1010 : node11919;
														assign node11919 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node11923 = (inp[5]) ? node11931 : node11924;
													assign node11924 = (inp[0]) ? 4'b1001 : node11925;
														assign node11925 = (inp[9]) ? 4'b1000 : node11926;
															assign node11926 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node11931 = (inp[0]) ? node11933 : 4'b1100;
														assign node11933 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node11936 = (inp[12]) ? node11948 : node11937;
												assign node11937 = (inp[5]) ? node11943 : node11938;
													assign node11938 = (inp[11]) ? 4'b1000 : node11939;
														assign node11939 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node11943 = (inp[11]) ? 4'b1100 : node11944;
														assign node11944 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node11948 = (inp[5]) ? node11958 : node11949;
													assign node11949 = (inp[11]) ? node11955 : node11950;
														assign node11950 = (inp[10]) ? node11952 : 4'b1110;
															assign node11952 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node11955 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node11958 = (inp[9]) ? node11960 : 4'b1011;
														assign node11960 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node11963 = (inp[5]) ? node11985 : node11964;
											assign node11964 = (inp[11]) ? node11980 : node11965;
												assign node11965 = (inp[12]) ? node11971 : node11966;
													assign node11966 = (inp[0]) ? node11968 : 4'b1100;
														assign node11968 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node11971 = (inp[4]) ? node11977 : node11972;
														assign node11972 = (inp[0]) ? 4'b1101 : node11973;
															assign node11973 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node11977 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node11980 = (inp[4]) ? 4'b1100 : node11981;
													assign node11981 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node11985 = (inp[10]) ? node11995 : node11986;
												assign node11986 = (inp[12]) ? node11992 : node11987;
													assign node11987 = (inp[9]) ? node11989 : 4'b1000;
														assign node11989 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11992 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node11995 = (inp[4]) ? node12003 : node11996;
													assign node11996 = (inp[11]) ? node11998 : 4'b1000;
														assign node11998 = (inp[0]) ? node12000 : 4'b1110;
															assign node12000 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12003 = (inp[12]) ? 4'b1110 : node12004;
														assign node12004 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node12008 = (inp[12]) ? node12120 : node12009;
									assign node12009 = (inp[4]) ? node12081 : node12010;
										assign node12010 = (inp[2]) ? node12048 : node12011;
											assign node12011 = (inp[5]) ? node12029 : node12012;
												assign node12012 = (inp[10]) ? node12020 : node12013;
													assign node12013 = (inp[11]) ? node12017 : node12014;
														assign node12014 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12017 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12020 = (inp[1]) ? node12026 : node12021;
														assign node12021 = (inp[11]) ? node12023 : 4'b1111;
															assign node12023 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node12026 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12029 = (inp[1]) ? node12043 : node12030;
													assign node12030 = (inp[11]) ? node12038 : node12031;
														assign node12031 = (inp[10]) ? node12033 : 4'b1010;
															assign node12033 = (inp[9]) ? 4'b1011 : node12034;
																assign node12034 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12038 = (inp[10]) ? 4'b1010 : node12039;
															assign node12039 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12043 = (inp[9]) ? node12045 : 4'b1111;
														assign node12045 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node12048 = (inp[5]) ? node12064 : node12049;
												assign node12049 = (inp[9]) ? node12053 : node12050;
													assign node12050 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node12053 = (inp[0]) ? 4'b1011 : node12054;
														assign node12054 = (inp[11]) ? node12058 : node12055;
															assign node12055 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node12058 = (inp[10]) ? 4'b1010 : node12059;
																assign node12059 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node12064 = (inp[1]) ? node12072 : node12065;
													assign node12065 = (inp[9]) ? node12069 : node12066;
														assign node12066 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node12069 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node12072 = (inp[10]) ? 4'b1010 : node12073;
														assign node12073 = (inp[9]) ? 4'b1011 : node12074;
															assign node12074 = (inp[11]) ? node12076 : 4'b1010;
																assign node12076 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node12081 = (inp[2]) ? node12105 : node12082;
											assign node12082 = (inp[5]) ? node12092 : node12083;
												assign node12083 = (inp[1]) ? node12089 : node12084;
													assign node12084 = (inp[9]) ? 4'b1001 : node12085;
														assign node12085 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node12089 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node12092 = (inp[0]) ? node12100 : node12093;
													assign node12093 = (inp[1]) ? 4'b1000 : node12094;
														assign node12094 = (inp[10]) ? 4'b1001 : node12095;
															assign node12095 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node12100 = (inp[1]) ? 4'b1001 : node12101;
														assign node12101 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node12105 = (inp[5]) ? node12113 : node12106;
												assign node12106 = (inp[1]) ? node12108 : 4'b1100;
													assign node12108 = (inp[11]) ? node12110 : 4'b1000;
														assign node12110 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node12113 = (inp[9]) ? node12115 : 4'b1100;
													assign node12115 = (inp[1]) ? node12117 : 4'b1101;
														assign node12117 = (inp[0]) ? 4'b1101 : 4'b1100;
									assign node12120 = (inp[4]) ? node12174 : node12121;
										assign node12121 = (inp[2]) ? node12153 : node12122;
											assign node12122 = (inp[5]) ? node12138 : node12123;
												assign node12123 = (inp[1]) ? node12131 : node12124;
													assign node12124 = (inp[0]) ? node12126 : 4'b1000;
														assign node12126 = (inp[10]) ? 4'b1001 : node12127;
															assign node12127 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node12131 = (inp[10]) ? 4'b1101 : node12132;
														assign node12132 = (inp[9]) ? node12134 : 4'b1100;
															assign node12134 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node12138 = (inp[11]) ? 4'b1001 : node12139;
													assign node12139 = (inp[9]) ? node12147 : node12140;
														assign node12140 = (inp[10]) ? node12142 : 4'b1000;
															assign node12142 = (inp[1]) ? node12144 : 4'b1001;
																assign node12144 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node12147 = (inp[0]) ? node12149 : 4'b1001;
															assign node12149 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node12153 = (inp[5]) ? node12163 : node12154;
												assign node12154 = (inp[1]) ? node12158 : node12155;
													assign node12155 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node12158 = (inp[9]) ? 4'b1001 : node12159;
														assign node12159 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node12163 = (inp[11]) ? node12165 : 4'b1101;
													assign node12165 = (inp[1]) ? node12167 : 4'b1100;
														assign node12167 = (inp[0]) ? 4'b1101 : node12168;
															assign node12168 = (inp[9]) ? node12170 : 4'b1100;
																assign node12170 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node12174 = (inp[2]) ? node12198 : node12175;
											assign node12175 = (inp[5]) ? node12187 : node12176;
												assign node12176 = (inp[1]) ? node12182 : node12177;
													assign node12177 = (inp[10]) ? 4'b1110 : node12178;
														assign node12178 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node12182 = (inp[9]) ? node12184 : 4'b1011;
														assign node12184 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node12187 = (inp[9]) ? node12193 : node12188;
													assign node12188 = (inp[0]) ? node12190 : 4'b1111;
														assign node12190 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node12193 = (inp[10]) ? 4'b1110 : node12194;
														assign node12194 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node12198 = (inp[5]) ? node12206 : node12199;
												assign node12199 = (inp[11]) ? node12203 : node12200;
													assign node12200 = (inp[0]) ? 4'b1111 : 4'b1011;
													assign node12203 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node12206 = (inp[0]) ? node12208 : 4'b1011;
													assign node12208 = (inp[9]) ? node12214 : node12209;
														assign node12209 = (inp[1]) ? 4'b1010 : node12210;
															assign node12210 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node12214 = (inp[1]) ? node12216 : 4'b1011;
															assign node12216 = (inp[11]) ? 4'b1010 : 4'b1011;
							assign node12219 = (inp[5]) ? node12377 : node12220;
								assign node12220 = (inp[13]) ? node12300 : node12221;
									assign node12221 = (inp[1]) ? node12275 : node12222;
										assign node12222 = (inp[2]) ? node12242 : node12223;
											assign node12223 = (inp[10]) ? node12237 : node12224;
												assign node12224 = (inp[4]) ? node12230 : node12225;
													assign node12225 = (inp[0]) ? node12227 : 4'b1010;
														assign node12227 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12230 = (inp[12]) ? 4'b1011 : node12231;
														assign node12231 = (inp[9]) ? node12233 : 4'b1110;
															assign node12233 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12237 = (inp[12]) ? node12239 : 4'b1011;
													assign node12239 = (inp[0]) ? 4'b1011 : 4'b1111;
											assign node12242 = (inp[9]) ? node12262 : node12243;
												assign node12243 = (inp[0]) ? node12253 : node12244;
													assign node12244 = (inp[10]) ? node12246 : 4'b1011;
														assign node12246 = (inp[4]) ? node12250 : node12247;
															assign node12247 = (inp[12]) ? 4'b1110 : 4'b1011;
															assign node12250 = (inp[12]) ? 4'b1011 : 4'b1110;
													assign node12253 = (inp[10]) ? node12259 : node12254;
														assign node12254 = (inp[11]) ? 4'b1110 : node12255;
															assign node12255 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node12259 = (inp[4]) ? 4'b1111 : 4'b1010;
												assign node12262 = (inp[12]) ? node12266 : node12263;
													assign node12263 = (inp[4]) ? 4'b1111 : 4'b1010;
													assign node12266 = (inp[4]) ? 4'b1010 : node12267;
														assign node12267 = (inp[11]) ? node12271 : node12268;
															assign node12268 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12271 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node12275 = (inp[12]) ? node12291 : node12276;
											assign node12276 = (inp[10]) ? node12282 : node12277;
												assign node12277 = (inp[9]) ? node12279 : 4'b1011;
													assign node12279 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node12282 = (inp[2]) ? node12288 : node12283;
													assign node12283 = (inp[4]) ? 4'b1010 : node12284;
														assign node12284 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node12288 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node12291 = (inp[0]) ? node12297 : node12292;
												assign node12292 = (inp[11]) ? 4'b1010 : node12293;
													assign node12293 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node12297 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node12300 = (inp[1]) ? node12340 : node12301;
										assign node12301 = (inp[0]) ? node12319 : node12302;
											assign node12302 = (inp[2]) ? node12310 : node12303;
												assign node12303 = (inp[9]) ? node12305 : 4'b1111;
													assign node12305 = (inp[12]) ? 4'b1010 : node12306;
														assign node12306 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12310 = (inp[9]) ? 4'b1111 : node12311;
													assign node12311 = (inp[10]) ? node12315 : node12312;
														assign node12312 = (inp[11]) ? 4'b1011 : 4'b1111;
														assign node12315 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node12319 = (inp[2]) ? node12329 : node12320;
												assign node12320 = (inp[11]) ? node12322 : 4'b1010;
													assign node12322 = (inp[9]) ? node12324 : 4'b1011;
														assign node12324 = (inp[12]) ? 4'b1011 : node12325;
															assign node12325 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node12329 = (inp[4]) ? node12333 : node12330;
													assign node12330 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node12333 = (inp[10]) ? node12335 : 4'b1111;
														assign node12335 = (inp[9]) ? node12337 : 4'b1110;
															assign node12337 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node12340 = (inp[10]) ? node12358 : node12341;
											assign node12341 = (inp[4]) ? node12349 : node12342;
												assign node12342 = (inp[11]) ? node12344 : 4'b1110;
													assign node12344 = (inp[9]) ? node12346 : 4'b1110;
														assign node12346 = (inp[12]) ? 4'b1110 : 4'b1111;
												assign node12349 = (inp[9]) ? node12353 : node12350;
													assign node12350 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12353 = (inp[11]) ? 4'b1110 : node12354;
														assign node12354 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node12358 = (inp[4]) ? node12370 : node12359;
												assign node12359 = (inp[0]) ? 4'b1111 : node12360;
													assign node12360 = (inp[12]) ? node12366 : node12361;
														assign node12361 = (inp[11]) ? node12363 : 4'b1110;
															assign node12363 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node12366 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node12370 = (inp[12]) ? 4'b1111 : node12371;
													assign node12371 = (inp[0]) ? node12373 : 4'b1111;
														assign node12373 = (inp[2]) ? 4'b1110 : 4'b1111;
								assign node12377 = (inp[13]) ? node12439 : node12378;
									assign node12378 = (inp[1]) ? node12424 : node12379;
										assign node12379 = (inp[11]) ? node12405 : node12380;
											assign node12380 = (inp[10]) ? node12394 : node12381;
												assign node12381 = (inp[9]) ? node12389 : node12382;
													assign node12382 = (inp[12]) ? node12386 : node12383;
														assign node12383 = (inp[0]) ? 4'b1011 : 4'b1111;
														assign node12386 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node12389 = (inp[2]) ? node12391 : 4'b1111;
														assign node12391 = (inp[12]) ? 4'b1011 : 4'b1110;
												assign node12394 = (inp[12]) ? node12402 : node12395;
													assign node12395 = (inp[4]) ? 4'b1011 : node12396;
														assign node12396 = (inp[9]) ? 4'b1110 : node12397;
															assign node12397 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node12402 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node12405 = (inp[2]) ? node12417 : node12406;
												assign node12406 = (inp[12]) ? node12412 : node12407;
													assign node12407 = (inp[10]) ? 4'b1010 : node12408;
														assign node12408 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12412 = (inp[0]) ? 4'b1011 : node12413;
														assign node12413 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node12417 = (inp[9]) ? node12419 : 4'b1111;
													assign node12419 = (inp[12]) ? 4'b1010 : node12420;
														assign node12420 = (inp[0]) ? 4'b1111 : 4'b1011;
										assign node12424 = (inp[2]) ? node12434 : node12425;
											assign node12425 = (inp[11]) ? node12427 : 4'b1110;
												assign node12427 = (inp[12]) ? 4'b1111 : node12428;
													assign node12428 = (inp[0]) ? 4'b1110 : node12429;
														assign node12429 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node12434 = (inp[11]) ? node12436 : 4'b1111;
												assign node12436 = (inp[9]) ? 4'b1111 : 4'b1110;
									assign node12439 = (inp[1]) ? node12477 : node12440;
										assign node12440 = (inp[12]) ? node12460 : node12441;
											assign node12441 = (inp[4]) ? node12453 : node12442;
												assign node12442 = (inp[9]) ? node12448 : node12443;
													assign node12443 = (inp[11]) ? node12445 : 4'b1010;
														assign node12445 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node12448 = (inp[11]) ? 4'b1010 : node12449;
														assign node12449 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node12453 = (inp[9]) ? node12455 : 4'b1110;
													assign node12455 = (inp[11]) ? node12457 : 4'b1111;
														assign node12457 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node12460 = (inp[4]) ? node12464 : node12461;
												assign node12461 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node12464 = (inp[11]) ? node12474 : node12465;
													assign node12465 = (inp[9]) ? node12471 : node12466;
														assign node12466 = (inp[2]) ? node12468 : 4'b1011;
															assign node12468 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12471 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12474 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node12477 = (inp[4]) ? node12497 : node12478;
											assign node12478 = (inp[10]) ? node12488 : node12479;
												assign node12479 = (inp[11]) ? node12481 : 4'b1010;
													assign node12481 = (inp[9]) ? node12483 : 4'b1011;
														assign node12483 = (inp[12]) ? node12485 : 4'b1011;
															assign node12485 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node12488 = (inp[11]) ? node12492 : node12489;
													assign node12489 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12492 = (inp[9]) ? 4'b1010 : node12493;
														assign node12493 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node12497 = (inp[10]) ? node12503 : node12498;
												assign node12498 = (inp[12]) ? 4'b1010 : node12499;
													assign node12499 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node12503 = (inp[12]) ? 4'b1011 : node12504;
													assign node12504 = (inp[9]) ? node12508 : node12505;
														assign node12505 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12508 = (inp[0]) ? 4'b1010 : 4'b1011;
						assign node12512 = (inp[6]) ? node12834 : node12513;
							assign node12513 = (inp[12]) ? node12687 : node12514;
								assign node12514 = (inp[13]) ? node12610 : node12515;
									assign node12515 = (inp[2]) ? node12561 : node12516;
										assign node12516 = (inp[4]) ? node12540 : node12517;
											assign node12517 = (inp[5]) ? node12531 : node12518;
												assign node12518 = (inp[11]) ? 4'b1110 : node12519;
													assign node12519 = (inp[9]) ? node12525 : node12520;
														assign node12520 = (inp[0]) ? 4'b1111 : node12521;
															assign node12521 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node12525 = (inp[10]) ? node12527 : 4'b1110;
															assign node12527 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node12531 = (inp[1]) ? node12535 : node12532;
													assign node12532 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12535 = (inp[10]) ? node12537 : 4'b1111;
														assign node12537 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node12540 = (inp[5]) ? node12552 : node12541;
												assign node12541 = (inp[0]) ? node12547 : node12542;
													assign node12542 = (inp[9]) ? 4'b1010 : node12543;
														assign node12543 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node12547 = (inp[10]) ? node12549 : 4'b1011;
														assign node12549 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node12552 = (inp[1]) ? node12556 : node12553;
													assign node12553 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node12556 = (inp[9]) ? node12558 : 4'b1010;
														assign node12558 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node12561 = (inp[11]) ? node12589 : node12562;
											assign node12562 = (inp[5]) ? node12574 : node12563;
												assign node12563 = (inp[4]) ? node12569 : node12564;
													assign node12564 = (inp[1]) ? 4'b1010 : node12565;
														assign node12565 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12569 = (inp[1]) ? 4'b1110 : node12570;
														assign node12570 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node12574 = (inp[0]) ? node12584 : node12575;
													assign node12575 = (inp[4]) ? 4'b1011 : node12576;
														assign node12576 = (inp[1]) ? 4'b1011 : node12577;
															assign node12577 = (inp[10]) ? node12579 : 4'b1110;
																assign node12579 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node12584 = (inp[4]) ? node12586 : 4'b1111;
														assign node12586 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node12589 = (inp[10]) ? node12607 : node12590;
												assign node12590 = (inp[4]) ? node12598 : node12591;
													assign node12591 = (inp[1]) ? 4'b1010 : node12592;
														assign node12592 = (inp[9]) ? node12594 : 4'b1111;
															assign node12594 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node12598 = (inp[9]) ? 4'b1111 : node12599;
														assign node12599 = (inp[1]) ? node12601 : 4'b1111;
															assign node12601 = (inp[0]) ? 4'b1110 : node12602;
																assign node12602 = (inp[5]) ? 4'b1110 : 4'b1111;
												assign node12607 = (inp[9]) ? 4'b1011 : 4'b1111;
									assign node12610 = (inp[2]) ? node12650 : node12611;
										assign node12611 = (inp[0]) ? node12635 : node12612;
											assign node12612 = (inp[10]) ? node12622 : node12613;
												assign node12613 = (inp[1]) ? node12619 : node12614;
													assign node12614 = (inp[11]) ? 4'b1110 : node12615;
														assign node12615 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node12619 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node12622 = (inp[4]) ? node12630 : node12623;
													assign node12623 = (inp[5]) ? 4'b1111 : node12624;
														assign node12624 = (inp[9]) ? 4'b1011 : node12625;
															assign node12625 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node12630 = (inp[5]) ? node12632 : 4'b1110;
														assign node12632 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node12635 = (inp[4]) ? node12645 : node12636;
												assign node12636 = (inp[5]) ? node12642 : node12637;
													assign node12637 = (inp[11]) ? 4'b1010 : node12638;
														assign node12638 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12642 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node12645 = (inp[9]) ? node12647 : 4'b1110;
													assign node12647 = (inp[5]) ? 4'b1011 : 4'b1111;
										assign node12650 = (inp[4]) ? node12668 : node12651;
											assign node12651 = (inp[1]) ? node12655 : node12652;
												assign node12652 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node12655 = (inp[9]) ? node12657 : 4'b1111;
													assign node12657 = (inp[10]) ? node12659 : 4'b1111;
														assign node12659 = (inp[11]) ? 4'b1111 : node12660;
															assign node12660 = (inp[5]) ? node12664 : node12661;
																assign node12661 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node12664 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node12668 = (inp[9]) ? node12680 : node12669;
												assign node12669 = (inp[1]) ? node12671 : 4'b1011;
													assign node12671 = (inp[10]) ? 4'b1011 : node12672;
														assign node12672 = (inp[11]) ? node12674 : 4'b1010;
															assign node12674 = (inp[0]) ? 4'b1010 : node12675;
																assign node12675 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node12680 = (inp[10]) ? node12682 : 4'b1011;
													assign node12682 = (inp[1]) ? 4'b1010 : node12683;
														assign node12683 = (inp[11]) ? 4'b1111 : 4'b1011;
								assign node12687 = (inp[9]) ? node12755 : node12688;
									assign node12688 = (inp[0]) ? node12724 : node12689;
										assign node12689 = (inp[10]) ? node12711 : node12690;
											assign node12690 = (inp[5]) ? node12702 : node12691;
												assign node12691 = (inp[11]) ? node12697 : node12692;
													assign node12692 = (inp[4]) ? node12694 : 4'b1100;
														assign node12694 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12697 = (inp[2]) ? 4'b1101 : node12698;
														assign node12698 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node12702 = (inp[2]) ? node12708 : node12703;
													assign node12703 = (inp[11]) ? node12705 : 4'b1101;
														assign node12705 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node12708 = (inp[13]) ? 4'b1000 : 4'b1100;
											assign node12711 = (inp[11]) ? node12717 : node12712;
												assign node12712 = (inp[2]) ? 4'b1001 : node12713;
													assign node12713 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node12717 = (inp[13]) ? node12721 : node12718;
													assign node12718 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12721 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node12724 = (inp[10]) ? node12732 : node12725;
											assign node12725 = (inp[5]) ? node12727 : 4'b1100;
												assign node12727 = (inp[2]) ? 4'b1001 : node12728;
													assign node12728 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node12732 = (inp[5]) ? node12746 : node12733;
												assign node12733 = (inp[2]) ? node12739 : node12734;
													assign node12734 = (inp[4]) ? 4'b1000 : node12735;
														assign node12735 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node12739 = (inp[1]) ? node12743 : node12740;
														assign node12740 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node12743 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node12746 = (inp[13]) ? node12750 : node12747;
													assign node12747 = (inp[2]) ? 4'b1100 : 4'b1001;
													assign node12750 = (inp[2]) ? 4'b1001 : node12751;
														assign node12751 = (inp[4]) ? 4'b1101 : 4'b1100;
									assign node12755 = (inp[10]) ? node12799 : node12756;
										assign node12756 = (inp[2]) ? node12780 : node12757;
											assign node12757 = (inp[13]) ? node12767 : node12758;
												assign node12758 = (inp[5]) ? node12762 : node12759;
													assign node12759 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node12762 = (inp[4]) ? 4'b1000 : node12763;
														assign node12763 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node12767 = (inp[1]) ? node12773 : node12768;
													assign node12768 = (inp[11]) ? node12770 : 4'b1101;
														assign node12770 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node12773 = (inp[5]) ? node12777 : node12774;
														assign node12774 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node12777 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node12780 = (inp[13]) ? node12788 : node12781;
												assign node12781 = (inp[5]) ? 4'b1101 : node12782;
													assign node12782 = (inp[1]) ? node12784 : 4'b1101;
														assign node12784 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node12788 = (inp[11]) ? node12794 : node12789;
													assign node12789 = (inp[5]) ? 4'b1000 : node12790;
														assign node12790 = (inp[1]) ? 4'b1101 : 4'b1000;
													assign node12794 = (inp[1]) ? 4'b1001 : node12795;
														assign node12795 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node12799 = (inp[1]) ? node12819 : node12800;
											assign node12800 = (inp[2]) ? node12812 : node12801;
												assign node12801 = (inp[13]) ? node12807 : node12802;
													assign node12802 = (inp[4]) ? 4'b1001 : node12803;
														assign node12803 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node12807 = (inp[0]) ? 4'b1101 : node12808;
														assign node12808 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node12812 = (inp[13]) ? node12814 : 4'b1100;
													assign node12814 = (inp[0]) ? node12816 : 4'b1000;
														assign node12816 = (inp[5]) ? 4'b1001 : 4'b1000;
											assign node12819 = (inp[13]) ? node12829 : node12820;
												assign node12820 = (inp[5]) ? node12822 : 4'b1000;
													assign node12822 = (inp[0]) ? node12826 : node12823;
														assign node12823 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node12826 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node12829 = (inp[5]) ? node12831 : 4'b1100;
													assign node12831 = (inp[2]) ? 4'b1000 : 4'b1100;
							assign node12834 = (inp[1]) ? node13014 : node12835;
								assign node12835 = (inp[0]) ? node12943 : node12836;
									assign node12836 = (inp[2]) ? node12870 : node12837;
										assign node12837 = (inp[4]) ? node12855 : node12838;
											assign node12838 = (inp[5]) ? node12848 : node12839;
												assign node12839 = (inp[13]) ? node12845 : node12840;
													assign node12840 = (inp[11]) ? 4'b1001 : node12841;
														assign node12841 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node12845 = (inp[12]) ? 4'b1101 : 4'b1100;
												assign node12848 = (inp[13]) ? node12850 : 4'b1100;
													assign node12850 = (inp[9]) ? node12852 : 4'b1000;
														assign node12852 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node12855 = (inp[11]) ? node12865 : node12856;
												assign node12856 = (inp[10]) ? 4'b1100 : node12857;
													assign node12857 = (inp[13]) ? node12859 : 4'b1101;
														assign node12859 = (inp[12]) ? node12861 : 4'b1001;
															assign node12861 = (inp[9]) ? 4'b1100 : 4'b1001;
												assign node12865 = (inp[12]) ? 4'b1001 : node12866;
													assign node12866 = (inp[5]) ? 4'b1001 : 4'b1101;
										assign node12870 = (inp[12]) ? node12902 : node12871;
											assign node12871 = (inp[13]) ? node12885 : node12872;
												assign node12872 = (inp[10]) ? node12880 : node12873;
													assign node12873 = (inp[5]) ? node12875 : 4'b1101;
														assign node12875 = (inp[9]) ? node12877 : 4'b1100;
															assign node12877 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node12880 = (inp[4]) ? node12882 : 4'b1001;
														assign node12882 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node12885 = (inp[4]) ? node12895 : node12886;
													assign node12886 = (inp[5]) ? node12892 : node12887;
														assign node12887 = (inp[9]) ? 4'b1100 : node12888;
															assign node12888 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12892 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12895 = (inp[5]) ? 4'b1100 : node12896;
														assign node12896 = (inp[11]) ? 4'b1000 : node12897;
															assign node12897 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node12902 = (inp[11]) ? node12924 : node12903;
												assign node12903 = (inp[10]) ? node12915 : node12904;
													assign node12904 = (inp[9]) ? node12912 : node12905;
														assign node12905 = (inp[4]) ? node12907 : 4'b1001;
															assign node12907 = (inp[5]) ? 4'b1100 : node12908;
																assign node12908 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node12912 = (inp[5]) ? 4'b1001 : 4'b1100;
													assign node12915 = (inp[13]) ? node12919 : node12916;
														assign node12916 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node12919 = (inp[9]) ? node12921 : 4'b1100;
															assign node12921 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node12924 = (inp[4]) ? node12936 : node12925;
													assign node12925 = (inp[5]) ? node12931 : node12926;
														assign node12926 = (inp[13]) ? node12928 : 4'b1000;
															assign node12928 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node12931 = (inp[9]) ? 4'b1000 : node12932;
															assign node12932 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node12936 = (inp[5]) ? node12940 : node12937;
														assign node12937 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node12940 = (inp[13]) ? 4'b1000 : 4'b1100;
									assign node12943 = (inp[5]) ? node12981 : node12944;
										assign node12944 = (inp[13]) ? node12966 : node12945;
											assign node12945 = (inp[4]) ? node12963 : node12946;
												assign node12946 = (inp[10]) ? node12954 : node12947;
													assign node12947 = (inp[2]) ? node12949 : 4'b1000;
														assign node12949 = (inp[11]) ? 4'b1000 : node12950;
															assign node12950 = (inp[12]) ? 4'b1001 : 4'b1000;
													assign node12954 = (inp[12]) ? node12958 : node12955;
														assign node12955 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12958 = (inp[11]) ? 4'b1000 : node12959;
															assign node12959 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node12963 = (inp[2]) ? 4'b1001 : 4'b1100;
											assign node12966 = (inp[12]) ? node12972 : node12967;
												assign node12967 = (inp[2]) ? node12969 : 4'b1000;
													assign node12969 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node12972 = (inp[10]) ? 4'b1101 : node12973;
													assign node12973 = (inp[9]) ? node12977 : node12974;
														assign node12974 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12977 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node12981 = (inp[13]) ? node13003 : node12982;
											assign node12982 = (inp[12]) ? node12988 : node12983;
												assign node12983 = (inp[4]) ? 4'b1001 : node12984;
													assign node12984 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node12988 = (inp[11]) ? node12992 : node12989;
													assign node12989 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node12992 = (inp[2]) ? node13000 : node12993;
														assign node12993 = (inp[10]) ? node12995 : 4'b1100;
															assign node12995 = (inp[9]) ? 4'b1101 : node12996;
																assign node12996 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node13000 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node13003 = (inp[12]) ? node13011 : node13004;
												assign node13004 = (inp[4]) ? node13006 : 4'b1001;
													assign node13006 = (inp[11]) ? node13008 : 4'b1101;
														assign node13008 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node13011 = (inp[10]) ? 4'b1001 : 4'b1000;
								assign node13014 = (inp[2]) ? node13102 : node13015;
									assign node13015 = (inp[4]) ? node13063 : node13016;
										assign node13016 = (inp[9]) ? node13034 : node13017;
											assign node13017 = (inp[13]) ? node13029 : node13018;
												assign node13018 = (inp[11]) ? 4'b1001 : node13019;
													assign node13019 = (inp[0]) ? 4'b1000 : node13020;
														assign node13020 = (inp[5]) ? node13024 : node13021;
															assign node13021 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node13024 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node13029 = (inp[11]) ? 4'b1101 : node13030;
													assign node13030 = (inp[12]) ? 4'b1001 : 4'b1101;
											assign node13034 = (inp[13]) ? node13046 : node13035;
												assign node13035 = (inp[11]) ? node13039 : node13036;
													assign node13036 = (inp[0]) ? 4'b1001 : 4'b1100;
													assign node13039 = (inp[12]) ? node13043 : node13040;
														assign node13040 = (inp[0]) ? 4'b1100 : 4'b1000;
														assign node13043 = (inp[5]) ? 4'b1100 : 4'b1000;
												assign node13046 = (inp[5]) ? node13056 : node13047;
													assign node13047 = (inp[12]) ? 4'b1101 : node13048;
														assign node13048 = (inp[0]) ? node13052 : node13049;
															assign node13049 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13052 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node13056 = (inp[12]) ? node13060 : node13057;
														assign node13057 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13060 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node13063 = (inp[0]) ? node13079 : node13064;
											assign node13064 = (inp[13]) ? node13070 : node13065;
												assign node13065 = (inp[5]) ? 4'b1101 : node13066;
													assign node13066 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node13070 = (inp[5]) ? 4'b1000 : node13071;
													assign node13071 = (inp[12]) ? 4'b1100 : node13072;
														assign node13072 = (inp[11]) ? 4'b1100 : node13073;
															assign node13073 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node13079 = (inp[13]) ? node13091 : node13080;
												assign node13080 = (inp[5]) ? node13084 : node13081;
													assign node13081 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node13084 = (inp[10]) ? 4'b1100 : node13085;
														assign node13085 = (inp[11]) ? node13087 : 4'b1101;
															assign node13087 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node13091 = (inp[5]) ? node13095 : node13092;
													assign node13092 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13095 = (inp[10]) ? node13097 : 4'b1000;
														assign node13097 = (inp[11]) ? node13099 : 4'b1001;
															assign node13099 = (inp[9]) ? 4'b1000 : 4'b1001;
									assign node13102 = (inp[13]) ? node13140 : node13103;
										assign node13103 = (inp[5]) ? node13127 : node13104;
											assign node13104 = (inp[4]) ? node13114 : node13105;
												assign node13105 = (inp[12]) ? node13109 : node13106;
													assign node13106 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node13109 = (inp[11]) ? 4'b1000 : node13110;
														assign node13110 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node13114 = (inp[9]) ? node13120 : node13115;
													assign node13115 = (inp[0]) ? 4'b1000 : node13116;
														assign node13116 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node13120 = (inp[12]) ? node13122 : 4'b1001;
														assign node13122 = (inp[10]) ? 4'b1000 : node13123;
															assign node13123 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node13127 = (inp[4]) ? node13135 : node13128;
												assign node13128 = (inp[12]) ? node13130 : 4'b1000;
													assign node13130 = (inp[9]) ? 4'b1101 : node13131;
														assign node13131 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node13135 = (inp[9]) ? 4'b1100 : node13136;
													assign node13136 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node13140 = (inp[5]) ? node13154 : node13141;
											assign node13141 = (inp[4]) ? node13149 : node13142;
												assign node13142 = (inp[12]) ? 4'b1100 : node13143;
													assign node13143 = (inp[11]) ? 4'b1001 : node13144;
														assign node13144 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node13149 = (inp[0]) ? 4'b1101 : node13150;
													assign node13150 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node13154 = (inp[4]) ? node13172 : node13155;
												assign node13155 = (inp[12]) ? node13163 : node13156;
													assign node13156 = (inp[9]) ? node13160 : node13157;
														assign node13157 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node13160 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13163 = (inp[0]) ? node13165 : 4'b1001;
														assign node13165 = (inp[9]) ? node13169 : node13166;
															assign node13166 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node13169 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node13172 = (inp[10]) ? node13190 : node13173;
													assign node13173 = (inp[12]) ? node13179 : node13174;
														assign node13174 = (inp[0]) ? 4'b1001 : node13175;
															assign node13175 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node13179 = (inp[0]) ? node13185 : node13180;
															assign node13180 = (inp[9]) ? 4'b1001 : node13181;
																assign node13181 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13185 = (inp[11]) ? 4'b1000 : node13186;
																assign node13186 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13190 = (inp[12]) ? 4'b1000 : node13191;
														assign node13191 = (inp[0]) ? 4'b1001 : 4'b1000;
				assign node13195 = (inp[7]) ? node14391 : node13196;
					assign node13196 = (inp[6]) ? node13878 : node13197;
						assign node13197 = (inp[12]) ? node13519 : node13198;
							assign node13198 = (inp[4]) ? node13362 : node13199;
								assign node13199 = (inp[15]) ? node13289 : node13200;
									assign node13200 = (inp[9]) ? node13236 : node13201;
										assign node13201 = (inp[5]) ? node13225 : node13202;
											assign node13202 = (inp[2]) ? node13210 : node13203;
												assign node13203 = (inp[13]) ? node13207 : node13204;
													assign node13204 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node13207 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node13210 = (inp[11]) ? node13220 : node13211;
													assign node13211 = (inp[10]) ? node13213 : 4'b0111;
														assign node13213 = (inp[13]) ? 4'b0010 : node13214;
															assign node13214 = (inp[0]) ? node13216 : 4'b0010;
																assign node13216 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node13220 = (inp[13]) ? 4'b0010 : node13221;
														assign node13221 = (inp[10]) ? 4'b0111 : 4'b0010;
											assign node13225 = (inp[1]) ? 4'b0110 : node13226;
												assign node13226 = (inp[10]) ? node13232 : node13227;
													assign node13227 = (inp[11]) ? 4'b0111 : node13228;
														assign node13228 = (inp[0]) ? 4'b0111 : 4'b0011;
													assign node13232 = (inp[0]) ? 4'b0011 : 4'b0110;
										assign node13236 = (inp[1]) ? node13270 : node13237;
											assign node13237 = (inp[11]) ? node13251 : node13238;
												assign node13238 = (inp[5]) ? node13246 : node13239;
													assign node13239 = (inp[13]) ? 4'b0010 : node13240;
														assign node13240 = (inp[2]) ? 4'b0111 : node13241;
															assign node13241 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node13246 = (inp[10]) ? node13248 : 4'b0110;
														assign node13248 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node13251 = (inp[10]) ? node13261 : node13252;
													assign node13252 = (inp[5]) ? node13254 : 4'b0010;
														assign node13254 = (inp[0]) ? 4'b0011 : node13255;
															assign node13255 = (inp[13]) ? 4'b0011 : node13256;
																assign node13256 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node13261 = (inp[5]) ? node13265 : node13262;
														assign node13262 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node13265 = (inp[2]) ? node13267 : 4'b0010;
															assign node13267 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node13270 = (inp[10]) ? node13276 : node13271;
												assign node13271 = (inp[11]) ? 4'b0110 : node13272;
													assign node13272 = (inp[0]) ? 4'b0110 : 4'b0010;
												assign node13276 = (inp[0]) ? node13284 : node13277;
													assign node13277 = (inp[2]) ? node13281 : node13278;
														assign node13278 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node13281 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node13284 = (inp[5]) ? 4'b0111 : node13285;
														assign node13285 = (inp[11]) ? 4'b0110 : 4'b0111;
									assign node13289 = (inp[11]) ? node13317 : node13290;
										assign node13290 = (inp[10]) ? node13302 : node13291;
											assign node13291 = (inp[5]) ? node13293 : 4'b0101;
												assign node13293 = (inp[2]) ? node13297 : node13294;
													assign node13294 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node13297 = (inp[0]) ? node13299 : 4'b0101;
														assign node13299 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node13302 = (inp[9]) ? node13312 : node13303;
												assign node13303 = (inp[1]) ? node13309 : node13304;
													assign node13304 = (inp[2]) ? 4'b0000 : node13305;
														assign node13305 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node13309 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node13312 = (inp[2]) ? node13314 : 4'b0100;
													assign node13314 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node13317 = (inp[0]) ? node13337 : node13318;
											assign node13318 = (inp[13]) ? node13326 : node13319;
												assign node13319 = (inp[10]) ? node13321 : 4'b0000;
													assign node13321 = (inp[1]) ? node13323 : 4'b0001;
														assign node13323 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node13326 = (inp[2]) ? node13332 : node13327;
													assign node13327 = (inp[5]) ? node13329 : 4'b0101;
														assign node13329 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node13332 = (inp[9]) ? node13334 : 4'b0001;
														assign node13334 = (inp[5]) ? 4'b0100 : 4'b0001;
											assign node13337 = (inp[2]) ? node13351 : node13338;
												assign node13338 = (inp[9]) ? node13346 : node13339;
													assign node13339 = (inp[13]) ? node13341 : 4'b0100;
														assign node13341 = (inp[5]) ? node13343 : 4'b0100;
															assign node13343 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node13346 = (inp[13]) ? node13348 : 4'b0001;
														assign node13348 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node13351 = (inp[5]) ? 4'b0101 : node13352;
													assign node13352 = (inp[13]) ? node13356 : node13353;
														assign node13353 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node13356 = (inp[1]) ? node13358 : 4'b0001;
															assign node13358 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node13362 = (inp[2]) ? node13450 : node13363;
									assign node13363 = (inp[13]) ? node13405 : node13364;
										assign node13364 = (inp[15]) ? node13388 : node13365;
											assign node13365 = (inp[5]) ? node13379 : node13366;
												assign node13366 = (inp[1]) ? node13374 : node13367;
													assign node13367 = (inp[10]) ? node13369 : 4'b0000;
														assign node13369 = (inp[9]) ? 4'b0001 : node13370;
															assign node13370 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node13374 = (inp[0]) ? node13376 : 4'b0001;
														assign node13376 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node13379 = (inp[1]) ? node13383 : node13380;
													assign node13380 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node13383 = (inp[0]) ? node13385 : 4'b0101;
														assign node13385 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node13388 = (inp[0]) ? node13398 : node13389;
												assign node13389 = (inp[11]) ? node13391 : 4'b0101;
													assign node13391 = (inp[9]) ? 4'b0101 : node13392;
														assign node13392 = (inp[10]) ? 4'b0100 : node13393;
															assign node13393 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node13398 = (inp[1]) ? node13402 : node13399;
													assign node13399 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node13402 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node13405 = (inp[15]) ? node13427 : node13406;
											assign node13406 = (inp[1]) ? node13420 : node13407;
												assign node13407 = (inp[10]) ? node13413 : node13408;
													assign node13408 = (inp[9]) ? node13410 : 4'b0100;
														assign node13410 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node13413 = (inp[5]) ? node13415 : 4'b0101;
														assign node13415 = (inp[0]) ? node13417 : 4'b0100;
															assign node13417 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node13420 = (inp[5]) ? node13424 : node13421;
													assign node13421 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node13424 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node13427 = (inp[5]) ? node13441 : node13428;
												assign node13428 = (inp[0]) ? node13436 : node13429;
													assign node13429 = (inp[10]) ? 4'b0001 : node13430;
														assign node13430 = (inp[11]) ? node13432 : 4'b0000;
															assign node13432 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node13436 = (inp[10]) ? 4'b0000 : node13437;
														assign node13437 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node13441 = (inp[1]) ? node13445 : node13442;
													assign node13442 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node13445 = (inp[11]) ? node13447 : 4'b0100;
														assign node13447 = (inp[0]) ? 4'b0101 : 4'b0100;
									assign node13450 = (inp[15]) ? node13478 : node13451;
										assign node13451 = (inp[13]) ? node13471 : node13452;
											assign node13452 = (inp[1]) ? node13462 : node13453;
												assign node13453 = (inp[11]) ? node13455 : 4'b0101;
													assign node13455 = (inp[0]) ? node13459 : node13456;
														assign node13456 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node13459 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node13462 = (inp[5]) ? node13468 : node13463;
													assign node13463 = (inp[9]) ? 4'b0100 : node13464;
														assign node13464 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node13468 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node13471 = (inp[5]) ? node13475 : node13472;
												assign node13472 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node13475 = (inp[1]) ? 4'b0101 : 4'b0001;
										assign node13478 = (inp[13]) ? node13494 : node13479;
											assign node13479 = (inp[1]) ? node13487 : node13480;
												assign node13480 = (inp[0]) ? node13482 : 4'b0000;
													assign node13482 = (inp[10]) ? node13484 : 4'b0000;
														assign node13484 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node13487 = (inp[5]) ? node13489 : 4'b0001;
													assign node13489 = (inp[10]) ? 4'b0100 : node13490;
														assign node13490 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node13494 = (inp[5]) ? node13512 : node13495;
												assign node13495 = (inp[11]) ? node13505 : node13496;
													assign node13496 = (inp[9]) ? node13498 : 4'b0100;
														assign node13498 = (inp[0]) ? 4'b0101 : node13499;
															assign node13499 = (inp[1]) ? 4'b0100 : node13500;
																assign node13500 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node13505 = (inp[0]) ? node13507 : 4'b0101;
														assign node13507 = (inp[9]) ? 4'b0101 : node13508;
															assign node13508 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node13512 = (inp[1]) ? 4'b0000 : node13513;
													assign node13513 = (inp[10]) ? node13515 : 4'b0100;
														assign node13515 = (inp[9]) ? 4'b0100 : 4'b0101;
							assign node13519 = (inp[4]) ? node13699 : node13520;
								assign node13520 = (inp[15]) ? node13608 : node13521;
									assign node13521 = (inp[10]) ? node13569 : node13522;
										assign node13522 = (inp[0]) ? node13546 : node13523;
											assign node13523 = (inp[9]) ? node13533 : node13524;
												assign node13524 = (inp[1]) ? node13526 : 4'b0000;
													assign node13526 = (inp[13]) ? node13528 : 4'b0001;
														assign node13528 = (inp[2]) ? node13530 : 4'b0100;
															assign node13530 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node13533 = (inp[5]) ? node13543 : node13534;
													assign node13534 = (inp[2]) ? 4'b0100 : node13535;
														assign node13535 = (inp[1]) ? node13539 : node13536;
															assign node13536 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node13539 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node13543 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node13546 = (inp[5]) ? node13556 : node13547;
												assign node13547 = (inp[13]) ? node13551 : node13548;
													assign node13548 = (inp[11]) ? 4'b0000 : 4'b0100;
													assign node13551 = (inp[1]) ? node13553 : 4'b0100;
														assign node13553 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node13556 = (inp[2]) ? node13562 : node13557;
													assign node13557 = (inp[11]) ? 4'b0100 : node13558;
														assign node13558 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node13562 = (inp[13]) ? node13566 : node13563;
														assign node13563 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node13566 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node13569 = (inp[13]) ? node13585 : node13570;
											assign node13570 = (inp[2]) ? node13580 : node13571;
												assign node13571 = (inp[5]) ? node13575 : node13572;
													assign node13572 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node13575 = (inp[9]) ? node13577 : 4'b0001;
														assign node13577 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node13580 = (inp[5]) ? 4'b0100 : node13581;
													assign node13581 = (inp[1]) ? 4'b0101 : 4'b0001;
											assign node13585 = (inp[11]) ? node13595 : node13586;
												assign node13586 = (inp[5]) ? node13592 : node13587;
													assign node13587 = (inp[1]) ? node13589 : 4'b0001;
														assign node13589 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node13592 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node13595 = (inp[0]) ? node13605 : node13596;
													assign node13596 = (inp[1]) ? node13602 : node13597;
														assign node13597 = (inp[2]) ? node13599 : 4'b0000;
															assign node13599 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node13602 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node13605 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node13608 = (inp[1]) ? node13670 : node13609;
										assign node13609 = (inp[9]) ? node13639 : node13610;
											assign node13610 = (inp[2]) ? node13626 : node13611;
												assign node13611 = (inp[0]) ? node13619 : node13612;
													assign node13612 = (inp[13]) ? 4'b0111 : node13613;
														assign node13613 = (inp[11]) ? 4'b0111 : node13614;
															assign node13614 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node13619 = (inp[10]) ? node13623 : node13620;
														assign node13620 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node13623 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node13626 = (inp[0]) ? node13634 : node13627;
													assign node13627 = (inp[13]) ? node13631 : node13628;
														assign node13628 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node13631 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node13634 = (inp[10]) ? node13636 : 4'b0010;
														assign node13636 = (inp[11]) ? 4'b0111 : 4'b0011;
											assign node13639 = (inp[5]) ? node13655 : node13640;
												assign node13640 = (inp[13]) ? node13648 : node13641;
													assign node13641 = (inp[2]) ? node13645 : node13642;
														assign node13642 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node13645 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node13648 = (inp[10]) ? node13650 : 4'b0010;
														assign node13650 = (inp[0]) ? 4'b0011 : node13651;
															assign node13651 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node13655 = (inp[0]) ? node13659 : node13656;
													assign node13656 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node13659 = (inp[10]) ? node13665 : node13660;
														assign node13660 = (inp[13]) ? node13662 : 4'b0011;
															assign node13662 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node13665 = (inp[2]) ? 4'b0110 : node13666;
															assign node13666 = (inp[13]) ? 4'b0111 : 4'b0011;
										assign node13670 = (inp[13]) ? node13690 : node13671;
											assign node13671 = (inp[2]) ? node13685 : node13672;
												assign node13672 = (inp[0]) ? 4'b0011 : node13673;
													assign node13673 = (inp[5]) ? node13675 : 4'b0010;
														assign node13675 = (inp[11]) ? 4'b0011 : node13676;
															assign node13676 = (inp[10]) ? node13680 : node13677;
																assign node13677 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node13680 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node13685 = (inp[0]) ? 4'b0111 : node13686;
													assign node13686 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node13690 = (inp[2]) ? 4'b0011 : node13691;
												assign node13691 = (inp[11]) ? 4'b0111 : node13692;
													assign node13692 = (inp[10]) ? 4'b0111 : node13693;
														assign node13693 = (inp[5]) ? 4'b0110 : 4'b0111;
								assign node13699 = (inp[11]) ? node13773 : node13700;
									assign node13700 = (inp[1]) ? node13738 : node13701;
										assign node13701 = (inp[2]) ? node13725 : node13702;
											assign node13702 = (inp[5]) ? node13712 : node13703;
												assign node13703 = (inp[9]) ? node13709 : node13704;
													assign node13704 = (inp[13]) ? 4'b0110 : node13705;
														assign node13705 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node13709 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node13712 = (inp[0]) ? node13718 : node13713;
													assign node13713 = (inp[13]) ? 4'b0110 : node13714;
														assign node13714 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node13718 = (inp[15]) ? node13720 : 4'b0110;
														assign node13720 = (inp[9]) ? node13722 : 4'b0110;
															assign node13722 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node13725 = (inp[10]) ? node13727 : 4'b0111;
												assign node13727 = (inp[15]) ? node13729 : 4'b0110;
													assign node13729 = (inp[9]) ? node13731 : 4'b0111;
														assign node13731 = (inp[13]) ? node13735 : node13732;
															assign node13732 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node13735 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node13738 = (inp[13]) ? node13758 : node13739;
											assign node13739 = (inp[15]) ? node13749 : node13740;
												assign node13740 = (inp[2]) ? node13744 : node13741;
													assign node13741 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node13744 = (inp[5]) ? node13746 : 4'b0010;
														assign node13746 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node13749 = (inp[2]) ? node13751 : 4'b0010;
													assign node13751 = (inp[10]) ? node13753 : 4'b0111;
														assign node13753 = (inp[9]) ? node13755 : 4'b0111;
															assign node13755 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node13758 = (inp[9]) ? node13766 : node13759;
												assign node13759 = (inp[5]) ? node13763 : node13760;
													assign node13760 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node13763 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node13766 = (inp[5]) ? node13768 : 4'b0111;
													assign node13768 = (inp[2]) ? 4'b0011 : node13769;
														assign node13769 = (inp[15]) ? 4'b0111 : 4'b0011;
									assign node13773 = (inp[9]) ? node13821 : node13774;
										assign node13774 = (inp[2]) ? node13804 : node13775;
											assign node13775 = (inp[10]) ? node13791 : node13776;
												assign node13776 = (inp[5]) ? node13786 : node13777;
													assign node13777 = (inp[15]) ? 4'b0111 : node13778;
														assign node13778 = (inp[0]) ? node13780 : 4'b0111;
															assign node13780 = (inp[1]) ? 4'b0110 : node13781;
																assign node13781 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node13786 = (inp[0]) ? node13788 : 4'b0110;
														assign node13788 = (inp[15]) ? 4'b0010 : 4'b0110;
												assign node13791 = (inp[0]) ? node13799 : node13792;
													assign node13792 = (inp[15]) ? 4'b0011 : node13793;
														assign node13793 = (inp[13]) ? 4'b0111 : node13794;
															assign node13794 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node13799 = (inp[5]) ? 4'b0011 : node13800;
														assign node13800 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node13804 = (inp[13]) ? node13816 : node13805;
												assign node13805 = (inp[15]) ? node13813 : node13806;
													assign node13806 = (inp[1]) ? node13808 : 4'b0110;
														assign node13808 = (inp[5]) ? 4'b0011 : node13809;
															assign node13809 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node13813 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node13816 = (inp[1]) ? node13818 : 4'b0010;
													assign node13818 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node13821 = (inp[0]) ? node13851 : node13822;
											assign node13822 = (inp[10]) ? node13838 : node13823;
												assign node13823 = (inp[5]) ? node13833 : node13824;
													assign node13824 = (inp[13]) ? node13830 : node13825;
														assign node13825 = (inp[1]) ? node13827 : 4'b0110;
															assign node13827 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node13830 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node13833 = (inp[1]) ? 4'b0111 : node13834;
														assign node13834 = (inp[13]) ? 4'b0111 : 4'b0010;
												assign node13838 = (inp[1]) ? node13844 : node13839;
													assign node13839 = (inp[5]) ? node13841 : 4'b0010;
														assign node13841 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node13844 = (inp[5]) ? node13846 : 4'b0111;
														assign node13846 = (inp[2]) ? node13848 : 4'b0110;
															assign node13848 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node13851 = (inp[2]) ? node13865 : node13852;
												assign node13852 = (inp[5]) ? node13854 : 4'b0010;
													assign node13854 = (inp[1]) ? node13858 : node13855;
														assign node13855 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node13858 = (inp[10]) ? 4'b0110 : node13859;
															assign node13859 = (inp[15]) ? 4'b0011 : node13860;
																assign node13860 = (inp[13]) ? 4'b0011 : 4'b0110;
												assign node13865 = (inp[1]) ? node13873 : node13866;
													assign node13866 = (inp[13]) ? 4'b0110 : node13867;
														assign node13867 = (inp[10]) ? 4'b0111 : node13868;
															assign node13868 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node13873 = (inp[15]) ? 4'b0110 : node13874;
														assign node13874 = (inp[13]) ? 4'b0111 : 4'b0011;
						assign node13878 = (inp[9]) ? node14138 : node13879;
							assign node13879 = (inp[5]) ? node14013 : node13880;
								assign node13880 = (inp[4]) ? node13972 : node13881;
									assign node13881 = (inp[11]) ? node13925 : node13882;
										assign node13882 = (inp[0]) ? node13910 : node13883;
											assign node13883 = (inp[2]) ? node13897 : node13884;
												assign node13884 = (inp[13]) ? node13894 : node13885;
													assign node13885 = (inp[10]) ? node13887 : 4'b0110;
														assign node13887 = (inp[12]) ? 4'b0110 : node13888;
															assign node13888 = (inp[15]) ? 4'b0011 : node13889;
																assign node13889 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node13894 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node13897 = (inp[15]) ? node13901 : node13898;
													assign node13898 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node13901 = (inp[12]) ? node13907 : node13902;
														assign node13902 = (inp[13]) ? 4'b0110 : node13903;
															assign node13903 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node13907 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node13910 = (inp[2]) ? node13922 : node13911;
												assign node13911 = (inp[13]) ? node13919 : node13912;
													assign node13912 = (inp[12]) ? 4'b0111 : node13913;
														assign node13913 = (inp[1]) ? node13915 : 4'b0011;
															assign node13915 = (inp[15]) ? 4'b0010 : 4'b0111;
													assign node13919 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node13922 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node13925 = (inp[15]) ? node13945 : node13926;
											assign node13926 = (inp[1]) ? node13938 : node13927;
												assign node13927 = (inp[13]) ? node13933 : node13928;
													assign node13928 = (inp[2]) ? 4'b0111 : node13929;
														assign node13929 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node13933 = (inp[12]) ? node13935 : 4'b0110;
														assign node13935 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node13938 = (inp[13]) ? 4'b0111 : node13939;
													assign node13939 = (inp[2]) ? node13941 : 4'b0110;
														assign node13941 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node13945 = (inp[12]) ? node13957 : node13946;
												assign node13946 = (inp[13]) ? node13954 : node13947;
													assign node13947 = (inp[1]) ? node13949 : 4'b0011;
														assign node13949 = (inp[2]) ? 4'b0010 : node13950;
															assign node13950 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node13954 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node13957 = (inp[13]) ? node13967 : node13958;
													assign node13958 = (inp[1]) ? node13962 : node13959;
														assign node13959 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node13962 = (inp[2]) ? node13964 : 4'b0111;
															assign node13964 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node13967 = (inp[0]) ? node13969 : 4'b0010;
														assign node13969 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node13972 = (inp[12]) ? node13998 : node13973;
										assign node13973 = (inp[15]) ? node13981 : node13974;
											assign node13974 = (inp[13]) ? node13976 : 4'b0010;
												assign node13976 = (inp[0]) ? 4'b0110 : node13977;
													assign node13977 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node13981 = (inp[13]) ? node13987 : node13982;
												assign node13982 = (inp[11]) ? 4'b0111 : node13983;
													assign node13983 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node13987 = (inp[10]) ? node13993 : node13988;
													assign node13988 = (inp[0]) ? 4'b0011 : node13989;
														assign node13989 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node13993 = (inp[11]) ? node13995 : 4'b0010;
														assign node13995 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node13998 = (inp[15]) ? node14010 : node13999;
											assign node13999 = (inp[13]) ? node14005 : node14000;
												assign node14000 = (inp[1]) ? node14002 : 4'b0010;
													assign node14002 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node14005 = (inp[0]) ? 4'b0110 : node14006;
													assign node14006 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node14010 = (inp[13]) ? 4'b0010 : 4'b0110;
								assign node14013 = (inp[4]) ? node14095 : node14014;
									assign node14014 = (inp[2]) ? node14050 : node14015;
										assign node14015 = (inp[13]) ? node14031 : node14016;
											assign node14016 = (inp[11]) ? node14026 : node14017;
												assign node14017 = (inp[0]) ? node14019 : 4'b0010;
													assign node14019 = (inp[15]) ? 4'b0010 : node14020;
														assign node14020 = (inp[12]) ? node14022 : 4'b0110;
															assign node14022 = (inp[1]) ? 4'b0011 : 4'b0110;
												assign node14026 = (inp[12]) ? 4'b0110 : node14027;
													assign node14027 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node14031 = (inp[12]) ? node14043 : node14032;
												assign node14032 = (inp[10]) ? node14036 : node14033;
													assign node14033 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node14036 = (inp[0]) ? node14040 : node14037;
														assign node14037 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node14040 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node14043 = (inp[1]) ? node14047 : node14044;
													assign node14044 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node14047 = (inp[15]) ? 4'b0010 : 4'b0110;
										assign node14050 = (inp[11]) ? node14078 : node14051;
											assign node14051 = (inp[13]) ? node14059 : node14052;
												assign node14052 = (inp[10]) ? 4'b0011 : node14053;
													assign node14053 = (inp[1]) ? node14055 : 4'b0111;
														assign node14055 = (inp[0]) ? 4'b0111 : 4'b0011;
												assign node14059 = (inp[0]) ? node14065 : node14060;
													assign node14060 = (inp[12]) ? node14062 : 4'b0010;
														assign node14062 = (inp[1]) ? 4'b0111 : 4'b0010;
													assign node14065 = (inp[12]) ? node14073 : node14066;
														assign node14066 = (inp[10]) ? node14068 : 4'b0111;
															assign node14068 = (inp[15]) ? node14070 : 4'b0111;
																assign node14070 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node14073 = (inp[1]) ? 4'b0111 : node14074;
															assign node14074 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node14078 = (inp[12]) ? node14092 : node14079;
												assign node14079 = (inp[13]) ? node14085 : node14080;
													assign node14080 = (inp[15]) ? 4'b0010 : node14081;
														assign node14081 = (inp[0]) ? 4'b0111 : 4'b0011;
													assign node14085 = (inp[1]) ? 4'b0111 : node14086;
														assign node14086 = (inp[15]) ? 4'b0110 : node14087;
															assign node14087 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node14092 = (inp[15]) ? 4'b0011 : 4'b0010;
									assign node14095 = (inp[12]) ? node14125 : node14096;
										assign node14096 = (inp[0]) ? node14114 : node14097;
											assign node14097 = (inp[1]) ? node14107 : node14098;
												assign node14098 = (inp[11]) ? node14100 : 4'b0011;
													assign node14100 = (inp[2]) ? 4'b0111 : node14101;
														assign node14101 = (inp[10]) ? node14103 : 4'b0011;
															assign node14103 = (inp[15]) ? 4'b0111 : 4'b0011;
												assign node14107 = (inp[11]) ? node14109 : 4'b0110;
													assign node14109 = (inp[13]) ? node14111 : 4'b0011;
														assign node14111 = (inp[15]) ? 4'b0010 : 4'b0110;
											assign node14114 = (inp[1]) ? node14120 : node14115;
												assign node14115 = (inp[15]) ? node14117 : 4'b0111;
													assign node14117 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node14120 = (inp[13]) ? node14122 : 4'b0111;
													assign node14122 = (inp[11]) ? 4'b0011 : 4'b0111;
										assign node14125 = (inp[15]) ? node14135 : node14126;
											assign node14126 = (inp[13]) ? node14132 : node14127;
												assign node14127 = (inp[11]) ? node14129 : 4'b0011;
													assign node14129 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node14132 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node14135 = (inp[13]) ? 4'b0011 : 4'b0111;
							assign node14138 = (inp[5]) ? node14270 : node14139;
								assign node14139 = (inp[4]) ? node14229 : node14140;
									assign node14140 = (inp[1]) ? node14198 : node14141;
										assign node14141 = (inp[11]) ? node14163 : node14142;
											assign node14142 = (inp[10]) ? node14160 : node14143;
												assign node14143 = (inp[2]) ? node14149 : node14144;
													assign node14144 = (inp[0]) ? 4'b0011 : node14145;
														assign node14145 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node14149 = (inp[0]) ? node14155 : node14150;
														assign node14150 = (inp[12]) ? 4'b0110 : node14151;
															assign node14151 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node14155 = (inp[12]) ? 4'b0111 : node14156;
															assign node14156 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node14160 = (inp[15]) ? 4'b0110 : 4'b0111;
											assign node14163 = (inp[2]) ? node14181 : node14164;
												assign node14164 = (inp[0]) ? node14176 : node14165;
													assign node14165 = (inp[10]) ? node14167 : 4'b0111;
														assign node14167 = (inp[13]) ? node14171 : node14168;
															assign node14168 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node14171 = (inp[12]) ? node14173 : 4'b0111;
																assign node14173 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node14176 = (inp[15]) ? 4'b0010 : node14177;
														assign node14177 = (inp[13]) ? 4'b0111 : 4'b0010;
												assign node14181 = (inp[10]) ? node14187 : node14182;
													assign node14182 = (inp[0]) ? node14184 : 4'b0010;
														assign node14184 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node14187 = (inp[0]) ? node14193 : node14188;
														assign node14188 = (inp[13]) ? 4'b0011 : node14189;
															assign node14189 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node14193 = (inp[15]) ? 4'b0111 : node14194;
															assign node14194 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node14198 = (inp[2]) ? node14210 : node14199;
											assign node14199 = (inp[0]) ? node14205 : node14200;
												assign node14200 = (inp[10]) ? 4'b0111 : node14201;
													assign node14201 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node14205 = (inp[10]) ? node14207 : 4'b0110;
													assign node14207 = (inp[11]) ? 4'b0011 : 4'b0110;
											assign node14210 = (inp[12]) ? node14220 : node14211;
												assign node14211 = (inp[0]) ? node14213 : 4'b0011;
													assign node14213 = (inp[15]) ? node14217 : node14214;
														assign node14214 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node14217 = (inp[13]) ? 4'b0110 : 4'b0010;
												assign node14220 = (inp[0]) ? node14222 : 4'b0110;
													assign node14222 = (inp[10]) ? 4'b0011 : node14223;
														assign node14223 = (inp[11]) ? node14225 : 4'b0111;
															assign node14225 = (inp[15]) ? 4'b0111 : 4'b0011;
									assign node14229 = (inp[12]) ? node14255 : node14230;
										assign node14230 = (inp[15]) ? node14242 : node14231;
											assign node14231 = (inp[13]) ? node14237 : node14232;
												assign node14232 = (inp[2]) ? 4'b0011 : node14233;
													assign node14233 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node14237 = (inp[0]) ? 4'b0111 : node14238;
													assign node14238 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node14242 = (inp[13]) ? node14252 : node14243;
												assign node14243 = (inp[2]) ? node14247 : node14244;
													assign node14244 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node14247 = (inp[10]) ? node14249 : 4'b0110;
														assign node14249 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node14252 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node14255 = (inp[15]) ? node14267 : node14256;
											assign node14256 = (inp[13]) ? node14262 : node14257;
												assign node14257 = (inp[1]) ? node14259 : 4'b0011;
													assign node14259 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node14262 = (inp[10]) ? 4'b0111 : node14263;
													assign node14263 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node14267 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node14270 = (inp[4]) ? node14328 : node14271;
									assign node14271 = (inp[2]) ? node14297 : node14272;
										assign node14272 = (inp[12]) ? node14286 : node14273;
											assign node14273 = (inp[13]) ? node14281 : node14274;
												assign node14274 = (inp[15]) ? node14278 : node14275;
													assign node14275 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node14278 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node14281 = (inp[0]) ? 4'b0111 : node14282;
													assign node14282 = (inp[15]) ? 4'b0110 : 4'b0010;
											assign node14286 = (inp[15]) ? node14294 : node14287;
												assign node14287 = (inp[0]) ? node14289 : 4'b0011;
													assign node14289 = (inp[13]) ? 4'b0010 : node14290;
														assign node14290 = (inp[1]) ? 4'b0010 : 4'b0111;
												assign node14294 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node14297 = (inp[15]) ? node14315 : node14298;
											assign node14298 = (inp[13]) ? node14306 : node14299;
												assign node14299 = (inp[1]) ? node14303 : node14300;
													assign node14300 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node14303 = (inp[12]) ? 4'b0011 : 4'b0110;
												assign node14306 = (inp[1]) ? node14312 : node14307;
													assign node14307 = (inp[12]) ? 4'b0011 : node14308;
														assign node14308 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node14312 = (inp[12]) ? 4'b0110 : 4'b0011;
											assign node14315 = (inp[12]) ? node14325 : node14316;
												assign node14316 = (inp[13]) ? node14320 : node14317;
													assign node14317 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node14320 = (inp[0]) ? node14322 : 4'b0110;
														assign node14322 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node14325 = (inp[13]) ? 4'b0010 : 4'b0110;
									assign node14328 = (inp[12]) ? node14376 : node14329;
										assign node14329 = (inp[11]) ? node14347 : node14330;
											assign node14330 = (inp[15]) ? node14338 : node14331;
												assign node14331 = (inp[13]) ? 4'b0110 : node14332;
													assign node14332 = (inp[1]) ? 4'b0010 : node14333;
														assign node14333 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node14338 = (inp[13]) ? node14342 : node14339;
													assign node14339 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node14342 = (inp[2]) ? node14344 : 4'b0011;
														assign node14344 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node14347 = (inp[10]) ? node14365 : node14348;
												assign node14348 = (inp[2]) ? node14354 : node14349;
													assign node14349 = (inp[1]) ? 4'b0110 : node14350;
														assign node14350 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node14354 = (inp[1]) ? node14362 : node14355;
														assign node14355 = (inp[0]) ? node14357 : 4'b0110;
															assign node14357 = (inp[13]) ? 4'b0110 : node14358;
																assign node14358 = (inp[15]) ? 4'b0111 : 4'b0011;
														assign node14362 = (inp[15]) ? 4'b0011 : 4'b0111;
												assign node14365 = (inp[0]) ? node14373 : node14366;
													assign node14366 = (inp[1]) ? 4'b0111 : node14367;
														assign node14367 = (inp[15]) ? 4'b0110 : node14368;
															assign node14368 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node14373 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node14376 = (inp[15]) ? node14388 : node14377;
											assign node14377 = (inp[13]) ? node14383 : node14378;
												assign node14378 = (inp[0]) ? node14380 : 4'b0010;
													assign node14380 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node14383 = (inp[0]) ? 4'b0110 : node14384;
													assign node14384 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node14388 = (inp[13]) ? 4'b0010 : 4'b0110;
					assign node14391 = (inp[6]) ? node15147 : node14392;
						assign node14392 = (inp[12]) ? node14810 : node14393;
							assign node14393 = (inp[15]) ? node14595 : node14394;
								assign node14394 = (inp[4]) ? node14516 : node14395;
									assign node14395 = (inp[10]) ? node14455 : node14396;
										assign node14396 = (inp[13]) ? node14424 : node14397;
											assign node14397 = (inp[2]) ? node14415 : node14398;
												assign node14398 = (inp[1]) ? node14406 : node14399;
													assign node14399 = (inp[11]) ? node14403 : node14400;
														assign node14400 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node14403 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node14406 = (inp[11]) ? node14410 : node14407;
														assign node14407 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node14410 = (inp[9]) ? node14412 : 4'b0001;
															assign node14412 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node14415 = (inp[1]) ? node14421 : node14416;
													assign node14416 = (inp[5]) ? 4'b0101 : node14417;
														assign node14417 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node14421 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node14424 = (inp[2]) ? node14442 : node14425;
												assign node14425 = (inp[1]) ? node14431 : node14426;
													assign node14426 = (inp[5]) ? node14428 : 4'b0001;
														assign node14428 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node14431 = (inp[9]) ? node14433 : 4'b0100;
														assign node14433 = (inp[5]) ? node14439 : node14434;
															assign node14434 = (inp[0]) ? 4'b0101 : node14435;
																assign node14435 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node14439 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node14442 = (inp[11]) ? node14446 : node14443;
													assign node14443 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node14446 = (inp[0]) ? node14452 : node14447;
														assign node14447 = (inp[1]) ? node14449 : 4'b0001;
															assign node14449 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node14452 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node14455 = (inp[1]) ? node14477 : node14456;
											assign node14456 = (inp[9]) ? node14466 : node14457;
												assign node14457 = (inp[0]) ? 4'b0100 : node14458;
													assign node14458 = (inp[5]) ? 4'b0000 : node14459;
														assign node14459 = (inp[11]) ? 4'b0100 : node14460;
															assign node14460 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node14466 = (inp[11]) ? node14472 : node14467;
													assign node14467 = (inp[2]) ? node14469 : 4'b0101;
														assign node14469 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node14472 = (inp[0]) ? 4'b0000 : node14473;
														assign node14473 = (inp[5]) ? 4'b0101 : 4'b0000;
											assign node14477 = (inp[0]) ? node14497 : node14478;
												assign node14478 = (inp[9]) ? node14490 : node14479;
													assign node14479 = (inp[5]) ? node14485 : node14480;
														assign node14480 = (inp[13]) ? 4'b0001 : node14481;
															assign node14481 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node14485 = (inp[2]) ? 4'b0000 : node14486;
															assign node14486 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node14490 = (inp[13]) ? node14494 : node14491;
														assign node14491 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node14494 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node14497 = (inp[11]) ? node14511 : node14498;
													assign node14498 = (inp[5]) ? node14506 : node14499;
														assign node14499 = (inp[13]) ? node14503 : node14500;
															assign node14500 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node14503 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node14506 = (inp[2]) ? node14508 : 4'b0000;
															assign node14508 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node14511 = (inp[5]) ? 4'b0001 : node14512;
														assign node14512 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node14516 = (inp[10]) ? node14552 : node14517;
										assign node14517 = (inp[9]) ? node14535 : node14518;
											assign node14518 = (inp[2]) ? node14528 : node14519;
												assign node14519 = (inp[13]) ? node14523 : node14520;
													assign node14520 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node14523 = (inp[5]) ? 4'b0110 : node14524;
														assign node14524 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node14528 = (inp[11]) ? 4'b0011 : node14529;
													assign node14529 = (inp[1]) ? node14531 : 4'b0010;
														assign node14531 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node14535 = (inp[11]) ? node14543 : node14536;
												assign node14536 = (inp[5]) ? 4'b0011 : node14537;
													assign node14537 = (inp[0]) ? 4'b0010 : node14538;
														assign node14538 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node14543 = (inp[13]) ? node14547 : node14544;
													assign node14544 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node14547 = (inp[2]) ? 4'b0011 : node14548;
														assign node14548 = (inp[0]) ? 4'b0111 : 4'b0011;
										assign node14552 = (inp[11]) ? node14576 : node14553;
											assign node14553 = (inp[5]) ? node14565 : node14554;
												assign node14554 = (inp[0]) ? node14560 : node14555;
													assign node14555 = (inp[9]) ? 4'b0110 : node14556;
														assign node14556 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node14560 = (inp[13]) ? 4'b0110 : node14561;
														assign node14561 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node14565 = (inp[0]) ? node14569 : node14566;
													assign node14566 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node14569 = (inp[13]) ? node14573 : node14570;
														assign node14570 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node14573 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node14576 = (inp[2]) ? node14584 : node14577;
												assign node14577 = (inp[13]) ? 4'b0110 : node14578;
													assign node14578 = (inp[1]) ? 4'b0010 : node14579;
														assign node14579 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node14584 = (inp[0]) ? node14588 : node14585;
													assign node14585 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node14588 = (inp[5]) ? node14592 : node14589;
														assign node14589 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node14592 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node14595 = (inp[0]) ? node14705 : node14596;
									assign node14596 = (inp[11]) ? node14648 : node14597;
										assign node14597 = (inp[13]) ? node14629 : node14598;
											assign node14598 = (inp[9]) ? node14608 : node14599;
												assign node14599 = (inp[4]) ? node14603 : node14600;
													assign node14600 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node14603 = (inp[2]) ? node14605 : 4'b0110;
														assign node14605 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node14608 = (inp[4]) ? node14622 : node14609;
													assign node14609 = (inp[5]) ? node14619 : node14610;
														assign node14610 = (inp[1]) ? node14616 : node14611;
															assign node14611 = (inp[2]) ? node14613 : 4'b0011;
																assign node14613 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node14616 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node14619 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node14622 = (inp[5]) ? node14624 : 4'b0111;
														assign node14624 = (inp[10]) ? node14626 : 4'b0011;
															assign node14626 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node14629 = (inp[9]) ? node14637 : node14630;
												assign node14630 = (inp[4]) ? node14634 : node14631;
													assign node14631 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node14634 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node14637 = (inp[2]) ? node14639 : 4'b0010;
													assign node14639 = (inp[5]) ? node14641 : 4'b0110;
														assign node14641 = (inp[4]) ? node14643 : 4'b0110;
															assign node14643 = (inp[1]) ? 4'b0010 : node14644;
																assign node14644 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node14648 = (inp[4]) ? node14680 : node14649;
											assign node14649 = (inp[1]) ? node14671 : node14650;
												assign node14650 = (inp[2]) ? node14660 : node14651;
													assign node14651 = (inp[5]) ? node14655 : node14652;
														assign node14652 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node14655 = (inp[9]) ? 4'b0110 : node14656;
															assign node14656 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node14660 = (inp[9]) ? node14662 : 4'b0111;
														assign node14662 = (inp[5]) ? node14666 : node14663;
															assign node14663 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node14666 = (inp[13]) ? node14668 : 4'b0011;
																assign node14668 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node14671 = (inp[9]) ? node14677 : node14672;
													assign node14672 = (inp[10]) ? node14674 : 4'b0010;
														assign node14674 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node14677 = (inp[10]) ? 4'b0010 : 4'b0111;
											assign node14680 = (inp[13]) ? node14694 : node14681;
												assign node14681 = (inp[2]) ? 4'b0011 : node14682;
													assign node14682 = (inp[9]) ? node14688 : node14683;
														assign node14683 = (inp[1]) ? 4'b0010 : node14684;
															assign node14684 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node14688 = (inp[10]) ? node14690 : 4'b0011;
															assign node14690 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node14694 = (inp[5]) ? 4'b0111 : node14695;
													assign node14695 = (inp[9]) ? node14701 : node14696;
														assign node14696 = (inp[2]) ? 4'b0110 : node14697;
															assign node14697 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node14701 = (inp[10]) ? 4'b0010 : 4'b0011;
									assign node14705 = (inp[11]) ? node14767 : node14706;
										assign node14706 = (inp[5]) ? node14730 : node14707;
											assign node14707 = (inp[10]) ? node14721 : node14708;
												assign node14708 = (inp[4]) ? node14712 : node14709;
													assign node14709 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node14712 = (inp[9]) ? node14714 : 4'b0011;
														assign node14714 = (inp[13]) ? node14718 : node14715;
															assign node14715 = (inp[1]) ? 4'b0010 : 4'b0111;
															assign node14718 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node14721 = (inp[9]) ? 4'b0110 : node14722;
													assign node14722 = (inp[13]) ? 4'b0110 : node14723;
														assign node14723 = (inp[1]) ? node14725 : 4'b0111;
															assign node14725 = (inp[2]) ? 4'b0010 : 4'b0111;
											assign node14730 = (inp[4]) ? node14748 : node14731;
												assign node14731 = (inp[2]) ? node14737 : node14732;
													assign node14732 = (inp[10]) ? 4'b0011 : node14733;
														assign node14733 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node14737 = (inp[13]) ? node14745 : node14738;
														assign node14738 = (inp[1]) ? 4'b0010 : node14739;
															assign node14739 = (inp[9]) ? node14741 : 4'b0011;
																assign node14741 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node14745 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node14748 = (inp[9]) ? node14754 : node14749;
													assign node14749 = (inp[2]) ? 4'b0010 : node14750;
														assign node14750 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node14754 = (inp[10]) ? 4'b0010 : node14755;
														assign node14755 = (inp[13]) ? node14763 : node14756;
															assign node14756 = (inp[2]) ? node14760 : node14757;
																assign node14757 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node14760 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node14763 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node14767 = (inp[1]) ? node14783 : node14768;
											assign node14768 = (inp[13]) ? node14776 : node14769;
												assign node14769 = (inp[2]) ? node14771 : 4'b0110;
													assign node14771 = (inp[10]) ? 4'b0111 : node14772;
														assign node14772 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node14776 = (inp[4]) ? node14780 : node14777;
													assign node14777 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node14780 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node14783 = (inp[9]) ? node14793 : node14784;
												assign node14784 = (inp[10]) ? node14786 : 4'b0110;
													assign node14786 = (inp[2]) ? node14788 : 4'b0111;
														assign node14788 = (inp[4]) ? node14790 : 4'b0011;
															assign node14790 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node14793 = (inp[10]) ? node14805 : node14794;
													assign node14794 = (inp[2]) ? node14800 : node14795;
														assign node14795 = (inp[13]) ? 4'b0011 : node14796;
															assign node14796 = (inp[4]) ? 4'b0011 : 4'b0110;
														assign node14800 = (inp[4]) ? 4'b0111 : node14801;
															assign node14801 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node14805 = (inp[4]) ? 4'b0010 : node14806;
														assign node14806 = (inp[2]) ? 4'b0110 : 4'b0111;
							assign node14810 = (inp[4]) ? node14962 : node14811;
								assign node14811 = (inp[15]) ? node14891 : node14812;
									assign node14812 = (inp[13]) ? node14848 : node14813;
										assign node14813 = (inp[0]) ? node14829 : node14814;
											assign node14814 = (inp[11]) ? node14822 : node14815;
												assign node14815 = (inp[1]) ? node14817 : 4'b0111;
													assign node14817 = (inp[9]) ? node14819 : 4'b0110;
														assign node14819 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node14822 = (inp[2]) ? node14824 : 4'b0110;
													assign node14824 = (inp[5]) ? 4'b0110 : node14825;
														assign node14825 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node14829 = (inp[2]) ? node14837 : node14830;
												assign node14830 = (inp[1]) ? 4'b0010 : node14831;
													assign node14831 = (inp[11]) ? node14833 : 4'b0111;
														assign node14833 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node14837 = (inp[11]) ? node14839 : 4'b0010;
													assign node14839 = (inp[5]) ? node14845 : node14840;
														assign node14840 = (inp[10]) ? 4'b0010 : node14841;
															assign node14841 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node14845 = (inp[1]) ? 4'b0111 : 4'b0011;
										assign node14848 = (inp[2]) ? node14874 : node14849;
											assign node14849 = (inp[1]) ? node14861 : node14850;
												assign node14850 = (inp[0]) ? node14856 : node14851;
													assign node14851 = (inp[11]) ? node14853 : 4'b0010;
														assign node14853 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node14856 = (inp[11]) ? 4'b0011 : node14857;
														assign node14857 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node14861 = (inp[5]) ? node14869 : node14862;
													assign node14862 = (inp[0]) ? 4'b0010 : node14863;
														assign node14863 = (inp[9]) ? 4'b0011 : node14864;
															assign node14864 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node14869 = (inp[0]) ? 4'b0111 : node14870;
														assign node14870 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node14874 = (inp[5]) ? node14886 : node14875;
												assign node14875 = (inp[1]) ? node14877 : 4'b0111;
													assign node14877 = (inp[9]) ? node14879 : 4'b0111;
														assign node14879 = (inp[10]) ? node14881 : 4'b0110;
															assign node14881 = (inp[11]) ? node14883 : 4'b0111;
																assign node14883 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node14886 = (inp[1]) ? 4'b0011 : node14887;
													assign node14887 = (inp[9]) ? 4'b0111 : 4'b0110;
									assign node14891 = (inp[11]) ? node14929 : node14892;
										assign node14892 = (inp[1]) ? node14908 : node14893;
											assign node14893 = (inp[2]) ? node14897 : node14894;
												assign node14894 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node14897 = (inp[0]) ? node14899 : 4'b0000;
													assign node14899 = (inp[9]) ? node14905 : node14900;
														assign node14900 = (inp[5]) ? node14902 : 4'b0000;
															assign node14902 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node14905 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node14908 = (inp[10]) ? node14918 : node14909;
												assign node14909 = (inp[2]) ? node14915 : node14910;
													assign node14910 = (inp[9]) ? 4'b0001 : node14911;
														assign node14911 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node14915 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node14918 = (inp[2]) ? node14924 : node14919;
													assign node14919 = (inp[13]) ? node14921 : 4'b0001;
														assign node14921 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node14924 = (inp[13]) ? 4'b0000 : node14925;
														assign node14925 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node14929 = (inp[9]) ? node14947 : node14930;
											assign node14930 = (inp[10]) ? node14938 : node14931;
												assign node14931 = (inp[13]) ? node14933 : 4'b0100;
													assign node14933 = (inp[0]) ? node14935 : 4'b0000;
														assign node14935 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node14938 = (inp[13]) ? node14944 : node14939;
													assign node14939 = (inp[0]) ? node14941 : 4'b0001;
														assign node14941 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node14944 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node14947 = (inp[10]) ? node14953 : node14948;
												assign node14948 = (inp[13]) ? node14950 : 4'b0000;
													assign node14950 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node14953 = (inp[2]) ? node14957 : node14954;
													assign node14954 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node14957 = (inp[1]) ? 4'b0100 : node14958;
														assign node14958 = (inp[13]) ? 4'b0100 : 4'b0001;
								assign node14962 = (inp[10]) ? node15048 : node14963;
									assign node14963 = (inp[15]) ? node15023 : node14964;
										assign node14964 = (inp[9]) ? node15004 : node14965;
											assign node14965 = (inp[0]) ? node14985 : node14966;
												assign node14966 = (inp[13]) ? node14976 : node14967;
													assign node14967 = (inp[1]) ? node14973 : node14968;
														assign node14968 = (inp[5]) ? node14970 : 4'b0000;
															assign node14970 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node14973 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node14976 = (inp[1]) ? node14980 : node14977;
														assign node14977 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node14980 = (inp[11]) ? node14982 : 4'b0001;
															assign node14982 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node14985 = (inp[5]) ? node14995 : node14986;
													assign node14986 = (inp[1]) ? node14992 : node14987;
														assign node14987 = (inp[13]) ? node14989 : 4'b0100;
															assign node14989 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node14992 = (inp[13]) ? 4'b0100 : 4'b0001;
													assign node14995 = (inp[2]) ? node14999 : node14996;
														assign node14996 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node14999 = (inp[13]) ? 4'b0000 : node15000;
															assign node15000 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node15004 = (inp[1]) ? node15018 : node15005;
												assign node15005 = (inp[13]) ? node15013 : node15006;
													assign node15006 = (inp[2]) ? node15008 : 4'b0000;
														assign node15008 = (inp[5]) ? 4'b0101 : node15009;
															assign node15009 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15013 = (inp[0]) ? node15015 : 4'b0100;
														assign node15015 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node15018 = (inp[13]) ? 4'b0001 : node15019;
													assign node15019 = (inp[11]) ? 4'b0100 : 4'b0001;
										assign node15023 = (inp[0]) ? node15031 : node15024;
											assign node15024 = (inp[9]) ? 4'b0000 : node15025;
												assign node15025 = (inp[1]) ? 4'b0000 : node15026;
													assign node15026 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node15031 = (inp[9]) ? node15043 : node15032;
												assign node15032 = (inp[5]) ? 4'b0100 : node15033;
													assign node15033 = (inp[1]) ? node15037 : node15034;
														assign node15034 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node15037 = (inp[13]) ? 4'b0000 : node15038;
															assign node15038 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node15043 = (inp[13]) ? 4'b0101 : node15044;
													assign node15044 = (inp[2]) ? 4'b0101 : 4'b0001;
									assign node15048 = (inp[15]) ? node15096 : node15049;
										assign node15049 = (inp[9]) ? node15065 : node15050;
											assign node15050 = (inp[11]) ? node15058 : node15051;
												assign node15051 = (inp[1]) ? 4'b0001 : node15052;
													assign node15052 = (inp[2]) ? 4'b0001 : node15053;
														assign node15053 = (inp[0]) ? 4'b0101 : 4'b0001;
												assign node15058 = (inp[5]) ? node15062 : node15059;
													assign node15059 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node15062 = (inp[0]) ? 4'b0001 : 4'b0101;
											assign node15065 = (inp[5]) ? node15081 : node15066;
												assign node15066 = (inp[11]) ? node15074 : node15067;
													assign node15067 = (inp[1]) ? node15069 : 4'b0101;
														assign node15069 = (inp[0]) ? 4'b0101 : node15070;
															assign node15070 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node15074 = (inp[2]) ? 4'b0101 : node15075;
														assign node15075 = (inp[0]) ? 4'b0001 : node15076;
															assign node15076 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node15081 = (inp[11]) ? node15089 : node15082;
													assign node15082 = (inp[0]) ? node15084 : 4'b0101;
														assign node15084 = (inp[1]) ? node15086 : 4'b0100;
															assign node15086 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node15089 = (inp[0]) ? 4'b0101 : node15090;
														assign node15090 = (inp[13]) ? node15092 : 4'b0000;
															assign node15092 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node15096 = (inp[13]) ? node15120 : node15097;
											assign node15097 = (inp[2]) ? node15109 : node15098;
												assign node15098 = (inp[11]) ? node15104 : node15099;
													assign node15099 = (inp[0]) ? node15101 : 4'b0001;
														assign node15101 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node15104 = (inp[1]) ? 4'b0001 : node15105;
														assign node15105 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node15109 = (inp[1]) ? node15115 : node15110;
													assign node15110 = (inp[5]) ? node15112 : 4'b0001;
														assign node15112 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node15115 = (inp[0]) ? node15117 : 4'b0100;
														assign node15117 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node15120 = (inp[1]) ? node15134 : node15121;
												assign node15121 = (inp[2]) ? node15127 : node15122;
													assign node15122 = (inp[9]) ? node15124 : 4'b0000;
														assign node15124 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node15127 = (inp[5]) ? 4'b0000 : node15128;
														assign node15128 = (inp[0]) ? node15130 : 4'b0100;
															assign node15130 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node15134 = (inp[2]) ? node15140 : node15135;
													assign node15135 = (inp[0]) ? node15137 : 4'b0101;
														assign node15137 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node15140 = (inp[0]) ? 4'b0000 : node15141;
														assign node15141 = (inp[9]) ? 4'b0001 : node15142;
															assign node15142 = (inp[5]) ? 4'b0000 : 4'b0001;
						assign node15147 = (inp[13]) ? node15373 : node15148;
							assign node15148 = (inp[4]) ? node15316 : node15149;
								assign node15149 = (inp[12]) ? node15231 : node15150;
									assign node15150 = (inp[15]) ? node15190 : node15151;
										assign node15151 = (inp[1]) ? node15169 : node15152;
											assign node15152 = (inp[5]) ? node15158 : node15153;
												assign node15153 = (inp[0]) ? 4'b0100 : node15154;
													assign node15154 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node15158 = (inp[0]) ? node15164 : node15159;
													assign node15159 = (inp[2]) ? 4'b0100 : node15160;
														assign node15160 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node15164 = (inp[2]) ? 4'b0101 : node15165;
														assign node15165 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node15169 = (inp[10]) ? node15183 : node15170;
												assign node15170 = (inp[9]) ? node15178 : node15171;
													assign node15171 = (inp[2]) ? node15173 : 4'b0000;
														assign node15173 = (inp[0]) ? node15175 : 4'b0001;
															assign node15175 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node15178 = (inp[11]) ? 4'b0001 : node15179;
														assign node15179 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node15183 = (inp[2]) ? node15185 : 4'b0000;
													assign node15185 = (inp[9]) ? 4'b0000 : node15186;
														assign node15186 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node15190 = (inp[5]) ? node15220 : node15191;
											assign node15191 = (inp[0]) ? node15207 : node15192;
												assign node15192 = (inp[10]) ? node15200 : node15193;
													assign node15193 = (inp[1]) ? node15195 : 4'b0000;
														assign node15195 = (inp[2]) ? node15197 : 4'b0001;
															assign node15197 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node15200 = (inp[1]) ? 4'b0000 : node15201;
														assign node15201 = (inp[2]) ? node15203 : 4'b0000;
															assign node15203 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node15207 = (inp[2]) ? node15215 : node15208;
													assign node15208 = (inp[10]) ? node15210 : 4'b0001;
														assign node15210 = (inp[9]) ? node15212 : 4'b0000;
															assign node15212 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node15215 = (inp[11]) ? 4'b0001 : node15216;
														assign node15216 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node15220 = (inp[9]) ? node15228 : node15221;
												assign node15221 = (inp[11]) ? node15223 : 4'b0000;
													assign node15223 = (inp[0]) ? node15225 : 4'b0000;
														assign node15225 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node15228 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node15231 = (inp[1]) ? node15267 : node15232;
										assign node15232 = (inp[15]) ? node15250 : node15233;
											assign node15233 = (inp[2]) ? node15239 : node15234;
												assign node15234 = (inp[9]) ? node15236 : 4'b0000;
													assign node15236 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node15239 = (inp[5]) ? node15247 : node15240;
													assign node15240 = (inp[10]) ? node15242 : 4'b0001;
														assign node15242 = (inp[9]) ? 4'b0001 : node15243;
															assign node15243 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15247 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node15250 = (inp[10]) ? node15262 : node15251;
												assign node15251 = (inp[5]) ? 4'b0101 : node15252;
													assign node15252 = (inp[11]) ? node15256 : node15253;
														assign node15253 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node15256 = (inp[9]) ? 4'b0101 : node15257;
															assign node15257 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node15262 = (inp[0]) ? 4'b0100 : node15263;
													assign node15263 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node15267 = (inp[5]) ? node15293 : node15268;
											assign node15268 = (inp[0]) ? node15284 : node15269;
												assign node15269 = (inp[11]) ? node15271 : 4'b0100;
													assign node15271 = (inp[2]) ? node15279 : node15272;
														assign node15272 = (inp[10]) ? node15274 : 4'b0101;
															assign node15274 = (inp[9]) ? node15276 : 4'b0100;
																assign node15276 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node15279 = (inp[15]) ? node15281 : 4'b0101;
															assign node15281 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node15284 = (inp[2]) ? node15286 : 4'b0101;
													assign node15286 = (inp[11]) ? 4'b0101 : node15287;
														assign node15287 = (inp[10]) ? node15289 : 4'b0100;
															assign node15289 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node15293 = (inp[0]) ? node15309 : node15294;
												assign node15294 = (inp[15]) ? node15304 : node15295;
													assign node15295 = (inp[11]) ? 4'b0100 : node15296;
														assign node15296 = (inp[10]) ? 4'b0101 : node15297;
															assign node15297 = (inp[9]) ? node15299 : 4'b0100;
																assign node15299 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node15304 = (inp[2]) ? node15306 : 4'b0101;
														assign node15306 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node15309 = (inp[10]) ? 4'b0100 : node15310;
													assign node15310 = (inp[15]) ? node15312 : 4'b0101;
														assign node15312 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node15316 = (inp[1]) ? node15352 : node15317;
									assign node15317 = (inp[11]) ? node15339 : node15318;
										assign node15318 = (inp[12]) ? node15330 : node15319;
											assign node15319 = (inp[9]) ? node15325 : node15320;
												assign node15320 = (inp[0]) ? node15322 : 4'b0100;
													assign node15322 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node15325 = (inp[0]) ? node15327 : 4'b0101;
													assign node15327 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node15330 = (inp[9]) ? node15334 : node15331;
												assign node15331 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node15334 = (inp[15]) ? 4'b0100 : node15335;
													assign node15335 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node15339 = (inp[12]) ? node15341 : 4'b0100;
											assign node15341 = (inp[9]) ? node15347 : node15342;
												assign node15342 = (inp[2]) ? node15344 : 4'b0101;
													assign node15344 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node15347 = (inp[0]) ? node15349 : 4'b0100;
													assign node15349 = (inp[15]) ? 4'b0100 : 4'b0101;
									assign node15352 = (inp[12]) ? node15360 : node15353;
										assign node15353 = (inp[15]) ? node15357 : node15354;
											assign node15354 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node15357 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node15360 = (inp[10]) ? node15368 : node15361;
											assign node15361 = (inp[5]) ? node15363 : 4'b0100;
												assign node15363 = (inp[9]) ? 4'b0101 : node15364;
													assign node15364 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node15368 = (inp[9]) ? 4'b0101 : node15369;
												assign node15369 = (inp[15]) ? 4'b0101 : 4'b0100;
							assign node15373 = (inp[4]) ? node15515 : node15374;
								assign node15374 = (inp[12]) ? node15452 : node15375;
									assign node15375 = (inp[1]) ? node15415 : node15376;
										assign node15376 = (inp[15]) ? node15398 : node15377;
											assign node15377 = (inp[10]) ? node15393 : node15378;
												assign node15378 = (inp[2]) ? node15388 : node15379;
													assign node15379 = (inp[9]) ? node15385 : node15380;
														assign node15380 = (inp[5]) ? 4'b0000 : node15381;
															assign node15381 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node15385 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15388 = (inp[5]) ? node15390 : 4'b0000;
														assign node15390 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node15393 = (inp[11]) ? 4'b0001 : node15394;
													assign node15394 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node15398 = (inp[11]) ? node15406 : node15399;
												assign node15399 = (inp[0]) ? node15401 : 4'b0100;
													assign node15401 = (inp[2]) ? 4'b0100 : node15402;
														assign node15402 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node15406 = (inp[9]) ? 4'b0101 : node15407;
													assign node15407 = (inp[0]) ? 4'b0100 : node15408;
														assign node15408 = (inp[5]) ? 4'b0101 : node15409;
															assign node15409 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node15415 = (inp[0]) ? node15437 : node15416;
											assign node15416 = (inp[5]) ? node15426 : node15417;
												assign node15417 = (inp[10]) ? node15419 : 4'b0101;
													assign node15419 = (inp[9]) ? node15423 : node15420;
														assign node15420 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node15423 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node15426 = (inp[11]) ? node15432 : node15427;
													assign node15427 = (inp[2]) ? 4'b0101 : node15428;
														assign node15428 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node15432 = (inp[15]) ? node15434 : 4'b0101;
														assign node15434 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node15437 = (inp[15]) ? node15447 : node15438;
												assign node15438 = (inp[11]) ? 4'b0101 : node15439;
													assign node15439 = (inp[9]) ? node15443 : node15440;
														assign node15440 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node15443 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node15447 = (inp[9]) ? 4'b0100 : node15448;
													assign node15448 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node15452 = (inp[1]) ? node15490 : node15453;
										assign node15453 = (inp[15]) ? node15473 : node15454;
											assign node15454 = (inp[10]) ? node15464 : node15455;
												assign node15455 = (inp[5]) ? 4'b0101 : node15456;
													assign node15456 = (inp[11]) ? node15458 : 4'b0101;
														assign node15458 = (inp[2]) ? 4'b0100 : node15459;
															assign node15459 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node15464 = (inp[2]) ? node15466 : 4'b0100;
													assign node15466 = (inp[9]) ? 4'b0101 : node15467;
														assign node15467 = (inp[5]) ? node15469 : 4'b0100;
															assign node15469 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node15473 = (inp[11]) ? node15483 : node15474;
												assign node15474 = (inp[2]) ? node15476 : 4'b0001;
													assign node15476 = (inp[9]) ? node15478 : 4'b0001;
														assign node15478 = (inp[5]) ? 4'b0000 : node15479;
															assign node15479 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node15483 = (inp[0]) ? 4'b0000 : node15484;
													assign node15484 = (inp[9]) ? node15486 : 4'b0000;
														assign node15486 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node15490 = (inp[5]) ? node15502 : node15491;
											assign node15491 = (inp[2]) ? node15493 : 4'b0001;
												assign node15493 = (inp[10]) ? 4'b0001 : node15494;
													assign node15494 = (inp[9]) ? node15498 : node15495;
														assign node15495 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node15498 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node15502 = (inp[11]) ? node15510 : node15503;
												assign node15503 = (inp[9]) ? node15507 : node15504;
													assign node15504 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node15507 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node15510 = (inp[2]) ? 4'b0000 : node15511;
													assign node15511 = (inp[9]) ? 4'b0001 : 4'b0000;
								assign node15515 = (inp[9]) ? node15529 : node15516;
									assign node15516 = (inp[1]) ? 4'b0001 : node15517;
										assign node15517 = (inp[12]) ? node15523 : node15518;
											assign node15518 = (inp[15]) ? 4'b0000 : node15519;
												assign node15519 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node15523 = (inp[15]) ? 4'b0001 : node15524;
												assign node15524 = (inp[0]) ? 4'b0001 : 4'b0000;
									assign node15529 = (inp[1]) ? 4'b0000 : node15530;
										assign node15530 = (inp[12]) ? node15536 : node15531;
											assign node15531 = (inp[15]) ? 4'b0001 : node15532;
												assign node15532 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node15536 = (inp[15]) ? 4'b0000 : node15537;
												assign node15537 = (inp[0]) ? 4'b0000 : 4'b0001;
			assign node15542 = (inp[12]) ? node17392 : node15543;
				assign node15543 = (inp[6]) ? node16699 : node15544;
					assign node15544 = (inp[14]) ? node16088 : node15545;
						assign node15545 = (inp[15]) ? node15853 : node15546;
							assign node15546 = (inp[4]) ? node15664 : node15547;
								assign node15547 = (inp[1]) ? node15597 : node15548;
									assign node15548 = (inp[2]) ? node15568 : node15549;
										assign node15549 = (inp[7]) ? node15557 : node15550;
											assign node15550 = (inp[10]) ? node15554 : node15551;
												assign node15551 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node15554 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node15557 = (inp[10]) ? node15563 : node15558;
												assign node15558 = (inp[11]) ? node15560 : 4'b0100;
													assign node15560 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node15563 = (inp[5]) ? node15565 : 4'b0101;
													assign node15565 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node15568 = (inp[7]) ? node15576 : node15569;
											assign node15569 = (inp[0]) ? 4'b0101 : node15570;
												assign node15570 = (inp[10]) ? 4'b0101 : node15571;
													assign node15571 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node15576 = (inp[11]) ? node15586 : node15577;
												assign node15577 = (inp[13]) ? node15579 : 4'b0001;
													assign node15579 = (inp[10]) ? node15583 : node15580;
														assign node15580 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node15583 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node15586 = (inp[9]) ? node15592 : node15587;
													assign node15587 = (inp[13]) ? node15589 : 4'b0000;
														assign node15589 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node15592 = (inp[10]) ? node15594 : 4'b0001;
														assign node15594 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node15597 = (inp[7]) ? node15631 : node15598;
										assign node15598 = (inp[2]) ? node15618 : node15599;
											assign node15599 = (inp[11]) ? node15613 : node15600;
												assign node15600 = (inp[9]) ? node15608 : node15601;
													assign node15601 = (inp[5]) ? 4'b0001 : node15602;
														assign node15602 = (inp[10]) ? node15604 : 4'b0000;
															assign node15604 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node15608 = (inp[13]) ? 4'b0000 : node15609;
														assign node15609 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node15613 = (inp[0]) ? 4'b0001 : node15614;
													assign node15614 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node15618 = (inp[13]) ? node15624 : node15619;
												assign node15619 = (inp[5]) ? node15621 : 4'b0101;
													assign node15621 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node15624 = (inp[11]) ? node15628 : node15625;
													assign node15625 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node15628 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node15631 = (inp[2]) ? node15649 : node15632;
											assign node15632 = (inp[10]) ? node15642 : node15633;
												assign node15633 = (inp[13]) ? 4'b0101 : node15634;
													assign node15634 = (inp[5]) ? node15638 : node15635;
														assign node15635 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node15638 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node15642 = (inp[5]) ? node15644 : 4'b0101;
													assign node15644 = (inp[13]) ? node15646 : 4'b0101;
														assign node15646 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node15649 = (inp[10]) ? node15657 : node15650;
												assign node15650 = (inp[5]) ? node15654 : node15651;
													assign node15651 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node15654 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node15657 = (inp[13]) ? node15661 : node15658;
													assign node15658 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15661 = (inp[5]) ? 4'b0000 : 4'b0001;
								assign node15664 = (inp[13]) ? node15750 : node15665;
									assign node15665 = (inp[9]) ? node15717 : node15666;
										assign node15666 = (inp[11]) ? node15692 : node15667;
											assign node15667 = (inp[1]) ? node15687 : node15668;
												assign node15668 = (inp[0]) ? node15680 : node15669;
													assign node15669 = (inp[5]) ? node15677 : node15670;
														assign node15670 = (inp[7]) ? node15674 : node15671;
															assign node15671 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node15674 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node15677 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node15680 = (inp[2]) ? node15682 : 4'b0101;
														assign node15682 = (inp[7]) ? 4'b0101 : node15683;
															assign node15683 = (inp[5]) ? 4'b0000 : 4'b0101;
												assign node15687 = (inp[10]) ? node15689 : 4'b0000;
													assign node15689 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node15692 = (inp[1]) ? node15706 : node15693;
												assign node15693 = (inp[10]) ? node15699 : node15694;
													assign node15694 = (inp[5]) ? node15696 : 4'b0000;
														assign node15696 = (inp[7]) ? 4'b0000 : 4'b0101;
													assign node15699 = (inp[2]) ? node15703 : node15700;
														assign node15700 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node15703 = (inp[5]) ? 4'b0001 : 4'b0100;
												assign node15706 = (inp[5]) ? node15712 : node15707;
													assign node15707 = (inp[7]) ? node15709 : 4'b0001;
														assign node15709 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node15712 = (inp[7]) ? node15714 : 4'b0101;
														assign node15714 = (inp[0]) ? 4'b0101 : 4'b0000;
										assign node15717 = (inp[0]) ? node15739 : node15718;
											assign node15718 = (inp[11]) ? node15728 : node15719;
												assign node15719 = (inp[2]) ? node15721 : 4'b0101;
													assign node15721 = (inp[10]) ? 4'b0001 : node15722;
														assign node15722 = (inp[5]) ? 4'b0101 : node15723;
															assign node15723 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node15728 = (inp[1]) ? node15730 : 4'b0100;
													assign node15730 = (inp[10]) ? node15732 : 4'b0001;
														assign node15732 = (inp[2]) ? node15734 : 4'b0100;
															assign node15734 = (inp[5]) ? 4'b0101 : node15735;
																assign node15735 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node15739 = (inp[11]) ? node15743 : node15740;
												assign node15740 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node15743 = (inp[7]) ? node15745 : 4'b0001;
													assign node15745 = (inp[2]) ? 4'b0100 : node15746;
														assign node15746 = (inp[5]) ? 4'b0001 : 4'b0101;
									assign node15750 = (inp[0]) ? node15806 : node15751;
										assign node15751 = (inp[1]) ? node15777 : node15752;
											assign node15752 = (inp[10]) ? node15764 : node15753;
												assign node15753 = (inp[11]) ? node15759 : node15754;
													assign node15754 = (inp[9]) ? 4'b0100 : node15755;
														assign node15755 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node15759 = (inp[9]) ? 4'b0001 : node15760;
														assign node15760 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node15764 = (inp[2]) ? node15772 : node15765;
													assign node15765 = (inp[9]) ? 4'b0000 : node15766;
														assign node15766 = (inp[7]) ? node15768 : 4'b0101;
															assign node15768 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node15772 = (inp[11]) ? 4'b0000 : node15773;
														assign node15773 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node15777 = (inp[7]) ? node15787 : node15778;
												assign node15778 = (inp[10]) ? node15784 : node15779;
													assign node15779 = (inp[11]) ? node15781 : 4'b0100;
														assign node15781 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node15784 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node15787 = (inp[9]) ? node15799 : node15788;
													assign node15788 = (inp[10]) ? node15794 : node15789;
														assign node15789 = (inp[5]) ? 4'b0100 : node15790;
															assign node15790 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node15794 = (inp[2]) ? node15796 : 4'b0001;
															assign node15796 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node15799 = (inp[10]) ? node15801 : 4'b0001;
														assign node15801 = (inp[5]) ? node15803 : 4'b0101;
															assign node15803 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node15806 = (inp[11]) ? node15834 : node15807;
											assign node15807 = (inp[9]) ? node15821 : node15808;
												assign node15808 = (inp[7]) ? node15816 : node15809;
													assign node15809 = (inp[2]) ? node15813 : node15810;
														assign node15810 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node15813 = (inp[5]) ? 4'b0000 : 4'b0101;
													assign node15816 = (inp[10]) ? node15818 : 4'b0100;
														assign node15818 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node15821 = (inp[10]) ? node15825 : node15822;
													assign node15822 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node15825 = (inp[7]) ? 4'b0100 : node15826;
														assign node15826 = (inp[5]) ? node15830 : node15827;
															assign node15827 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node15830 = (inp[2]) ? 4'b0000 : 4'b0101;
											assign node15834 = (inp[10]) ? node15848 : node15835;
												assign node15835 = (inp[5]) ? node15841 : node15836;
													assign node15836 = (inp[2]) ? 4'b0101 : node15837;
														assign node15837 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node15841 = (inp[1]) ? node15843 : 4'b0100;
														assign node15843 = (inp[7]) ? 4'b0000 : node15844;
															assign node15844 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node15848 = (inp[2]) ? 4'b0000 : node15849;
													assign node15849 = (inp[1]) ? 4'b0001 : 4'b0000;
							assign node15853 = (inp[7]) ? node15951 : node15854;
								assign node15854 = (inp[4]) ? node15894 : node15855;
									assign node15855 = (inp[2]) ? node15863 : node15856;
										assign node15856 = (inp[10]) ? node15860 : node15857;
											assign node15857 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node15860 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node15863 = (inp[9]) ? node15877 : node15864;
											assign node15864 = (inp[0]) ? node15870 : node15865;
												assign node15865 = (inp[10]) ? node15867 : 4'b0111;
													assign node15867 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node15870 = (inp[13]) ? 4'b0110 : node15871;
													assign node15871 = (inp[1]) ? 4'b0111 : node15872;
														assign node15872 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node15877 = (inp[11]) ? node15887 : node15878;
												assign node15878 = (inp[13]) ? 4'b0111 : node15879;
													assign node15879 = (inp[1]) ? node15883 : node15880;
														assign node15880 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node15883 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node15887 = (inp[5]) ? node15889 : 4'b0110;
													assign node15889 = (inp[10]) ? node15891 : 4'b0111;
														assign node15891 = (inp[1]) ? 4'b0110 : 4'b0111;
									assign node15894 = (inp[2]) ? node15928 : node15895;
										assign node15895 = (inp[9]) ? node15913 : node15896;
											assign node15896 = (inp[13]) ? node15908 : node15897;
												assign node15897 = (inp[5]) ? node15901 : node15898;
													assign node15898 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node15901 = (inp[1]) ? node15903 : 4'b0110;
														assign node15903 = (inp[11]) ? 4'b0110 : node15904;
															assign node15904 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node15908 = (inp[1]) ? node15910 : 4'b0110;
													assign node15910 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node15913 = (inp[13]) ? node15921 : node15914;
												assign node15914 = (inp[5]) ? node15916 : 4'b0111;
													assign node15916 = (inp[1]) ? 4'b0111 : node15917;
														assign node15917 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node15921 = (inp[0]) ? 4'b0110 : node15922;
													assign node15922 = (inp[10]) ? 4'b0111 : node15923;
														assign node15923 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node15928 = (inp[10]) ? node15940 : node15929;
											assign node15929 = (inp[1]) ? node15935 : node15930;
												assign node15930 = (inp[5]) ? 4'b0010 : node15931;
													assign node15931 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node15935 = (inp[11]) ? 4'b0011 : node15936;
													assign node15936 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node15940 = (inp[1]) ? node15946 : node15941;
												assign node15941 = (inp[5]) ? 4'b0011 : node15942;
													assign node15942 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node15946 = (inp[5]) ? 4'b0010 : node15947;
													assign node15947 = (inp[11]) ? 4'b0010 : 4'b0011;
								assign node15951 = (inp[1]) ? node16017 : node15952;
									assign node15952 = (inp[11]) ? node15982 : node15953;
										assign node15953 = (inp[9]) ? node15967 : node15954;
											assign node15954 = (inp[4]) ? node15962 : node15955;
												assign node15955 = (inp[2]) ? 4'b0111 : node15956;
													assign node15956 = (inp[0]) ? node15958 : 4'b0011;
														assign node15958 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node15962 = (inp[5]) ? 4'b0011 : node15963;
													assign node15963 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node15967 = (inp[0]) ? node15975 : node15968;
												assign node15968 = (inp[2]) ? node15972 : node15969;
													assign node15969 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node15972 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node15975 = (inp[13]) ? 4'b0111 : node15976;
													assign node15976 = (inp[4]) ? node15978 : 4'b0010;
														assign node15978 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node15982 = (inp[10]) ? node15998 : node15983;
											assign node15983 = (inp[5]) ? node15989 : node15984;
												assign node15984 = (inp[4]) ? node15986 : 4'b0111;
													assign node15986 = (inp[0]) ? 4'b0010 : 4'b0111;
												assign node15989 = (inp[9]) ? node15991 : 4'b0110;
													assign node15991 = (inp[0]) ? 4'b0010 : node15992;
														assign node15992 = (inp[13]) ? node15994 : 4'b0110;
															assign node15994 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node15998 = (inp[5]) ? node16006 : node15999;
												assign node15999 = (inp[9]) ? node16001 : 4'b0110;
													assign node16001 = (inp[2]) ? 4'b0011 : node16002;
														assign node16002 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node16006 = (inp[0]) ? node16010 : node16007;
													assign node16007 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node16010 = (inp[2]) ? node16014 : node16011;
														assign node16011 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16014 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node16017 = (inp[9]) ? node16065 : node16018;
										assign node16018 = (inp[10]) ? node16044 : node16019;
											assign node16019 = (inp[13]) ? node16037 : node16020;
												assign node16020 = (inp[0]) ? node16034 : node16021;
													assign node16021 = (inp[5]) ? node16029 : node16022;
														assign node16022 = (inp[2]) ? node16024 : 4'b0110;
															assign node16024 = (inp[4]) ? 4'b0011 : node16025;
																assign node16025 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node16029 = (inp[2]) ? 4'b0010 : node16030;
															assign node16030 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node16034 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node16037 = (inp[2]) ? node16041 : node16038;
													assign node16038 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node16041 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node16044 = (inp[13]) ? node16050 : node16045;
												assign node16045 = (inp[0]) ? 4'b0011 : node16046;
													assign node16046 = (inp[11]) ? 4'b0110 : 4'b0011;
												assign node16050 = (inp[11]) ? node16058 : node16051;
													assign node16051 = (inp[5]) ? node16055 : node16052;
														assign node16052 = (inp[0]) ? 4'b0010 : 4'b0110;
														assign node16055 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node16058 = (inp[5]) ? node16060 : 4'b0011;
														assign node16060 = (inp[0]) ? 4'b0010 : node16061;
															assign node16061 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node16065 = (inp[4]) ? node16079 : node16066;
											assign node16066 = (inp[2]) ? node16072 : node16067;
												assign node16067 = (inp[0]) ? 4'b0010 : node16068;
													assign node16068 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node16072 = (inp[11]) ? node16074 : 4'b0110;
													assign node16074 = (inp[10]) ? node16076 : 4'b0110;
														assign node16076 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node16079 = (inp[2]) ? 4'b0011 : node16080;
												assign node16080 = (inp[10]) ? node16082 : 4'b0111;
													assign node16082 = (inp[5]) ? 4'b0110 : node16083;
														assign node16083 = (inp[11]) ? 4'b0111 : 4'b0110;
						assign node16088 = (inp[11]) ? node16392 : node16089;
							assign node16089 = (inp[1]) ? node16237 : node16090;
								assign node16090 = (inp[10]) ? node16170 : node16091;
									assign node16091 = (inp[13]) ? node16139 : node16092;
										assign node16092 = (inp[7]) ? node16116 : node16093;
											assign node16093 = (inp[5]) ? node16103 : node16094;
												assign node16094 = (inp[2]) ? node16096 : 4'b0010;
													assign node16096 = (inp[15]) ? node16100 : node16097;
														assign node16097 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node16100 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node16103 = (inp[4]) ? node16107 : node16104;
													assign node16104 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node16107 = (inp[9]) ? node16111 : node16108;
														assign node16108 = (inp[15]) ? 4'b0011 : 4'b0110;
														assign node16111 = (inp[15]) ? node16113 : 4'b0011;
															assign node16113 = (inp[2]) ? 4'b0011 : 4'b0111;
											assign node16116 = (inp[5]) ? node16128 : node16117;
												assign node16117 = (inp[2]) ? node16123 : node16118;
													assign node16118 = (inp[4]) ? 4'b0110 : node16119;
														assign node16119 = (inp[15]) ? 4'b0010 : 4'b0110;
													assign node16123 = (inp[4]) ? 4'b0010 : node16124;
														assign node16124 = (inp[15]) ? 4'b0111 : 4'b0011;
												assign node16128 = (inp[9]) ? node16130 : 4'b0110;
													assign node16130 = (inp[0]) ? node16132 : 4'b0110;
														assign node16132 = (inp[15]) ? 4'b0010 : node16133;
															assign node16133 = (inp[2]) ? node16135 : 4'b0110;
																assign node16135 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node16139 = (inp[5]) ? node16153 : node16140;
											assign node16140 = (inp[2]) ? node16144 : node16141;
												assign node16141 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node16144 = (inp[4]) ? 4'b0010 : node16145;
													assign node16145 = (inp[15]) ? node16149 : node16146;
														assign node16146 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node16149 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node16153 = (inp[9]) ? node16161 : node16154;
												assign node16154 = (inp[0]) ? node16156 : 4'b0011;
													assign node16156 = (inp[4]) ? 4'b0111 : node16157;
														assign node16157 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node16161 = (inp[0]) ? node16163 : 4'b0111;
													assign node16163 = (inp[2]) ? node16165 : 4'b0111;
														assign node16165 = (inp[7]) ? node16167 : 4'b0111;
															assign node16167 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node16170 = (inp[15]) ? node16200 : node16171;
										assign node16171 = (inp[2]) ? node16187 : node16172;
											assign node16172 = (inp[13]) ? node16180 : node16173;
												assign node16173 = (inp[7]) ? node16177 : node16174;
													assign node16174 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node16177 = (inp[4]) ? 4'b0111 : 4'b0010;
												assign node16180 = (inp[5]) ? node16184 : node16181;
													assign node16181 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node16184 = (inp[7]) ? 4'b0011 : 4'b0110;
											assign node16187 = (inp[7]) ? node16193 : node16188;
												assign node16188 = (inp[9]) ? node16190 : 4'b0111;
													assign node16190 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node16193 = (inp[5]) ? node16197 : node16194;
													assign node16194 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node16197 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node16200 = (inp[7]) ? node16216 : node16201;
											assign node16201 = (inp[5]) ? node16209 : node16202;
												assign node16202 = (inp[2]) ? node16206 : node16203;
													assign node16203 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node16206 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node16209 = (inp[4]) ? node16213 : node16210;
													assign node16210 = (inp[2]) ? 4'b0110 : 4'b0011;
													assign node16213 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node16216 = (inp[9]) ? node16230 : node16217;
												assign node16217 = (inp[13]) ? node16221 : node16218;
													assign node16218 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node16221 = (inp[2]) ? node16225 : node16222;
														assign node16222 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node16225 = (inp[4]) ? 4'b0011 : node16226;
															assign node16226 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node16230 = (inp[4]) ? node16234 : node16231;
													assign node16231 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node16234 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node16237 = (inp[10]) ? node16313 : node16238;
									assign node16238 = (inp[2]) ? node16270 : node16239;
										assign node16239 = (inp[4]) ? node16253 : node16240;
											assign node16240 = (inp[15]) ? 4'b0011 : node16241;
												assign node16241 = (inp[13]) ? node16247 : node16242;
													assign node16242 = (inp[5]) ? 4'b0010 : node16243;
														assign node16243 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node16247 = (inp[9]) ? node16249 : 4'b0111;
														assign node16249 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node16253 = (inp[15]) ? node16265 : node16254;
												assign node16254 = (inp[7]) ? 4'b0111 : node16255;
													assign node16255 = (inp[0]) ? node16259 : node16256;
														assign node16256 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node16259 = (inp[5]) ? 4'b0010 : node16260;
															assign node16260 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node16265 = (inp[7]) ? 4'b0111 : node16266;
													assign node16266 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node16270 = (inp[4]) ? node16298 : node16271;
											assign node16271 = (inp[15]) ? node16285 : node16272;
												assign node16272 = (inp[13]) ? node16280 : node16273;
													assign node16273 = (inp[7]) ? node16277 : node16274;
														assign node16274 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node16277 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node16280 = (inp[5]) ? node16282 : 4'b0010;
														assign node16282 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node16285 = (inp[0]) ? node16291 : node16286;
													assign node16286 = (inp[5]) ? 4'b0111 : node16287;
														assign node16287 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node16291 = (inp[7]) ? node16295 : node16292;
														assign node16292 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node16295 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node16298 = (inp[7]) ? node16308 : node16299;
												assign node16299 = (inp[15]) ? node16305 : node16300;
													assign node16300 = (inp[13]) ? 4'b0110 : node16301;
														assign node16301 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node16305 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node16308 = (inp[13]) ? 4'b0011 : node16309;
													assign node16309 = (inp[15]) ? 4'b0011 : 4'b0010;
									assign node16313 = (inp[13]) ? node16349 : node16314;
										assign node16314 = (inp[7]) ? node16332 : node16315;
											assign node16315 = (inp[2]) ? node16325 : node16316;
												assign node16316 = (inp[0]) ? node16318 : 4'b0110;
													assign node16318 = (inp[9]) ? 4'b0111 : node16319;
														assign node16319 = (inp[15]) ? 4'b0010 : node16320;
															assign node16320 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node16325 = (inp[4]) ? node16329 : node16326;
													assign node16326 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node16329 = (inp[15]) ? 4'b0010 : 4'b0110;
											assign node16332 = (inp[15]) ? node16344 : node16333;
												assign node16333 = (inp[2]) ? node16339 : node16334;
													assign node16334 = (inp[9]) ? node16336 : 4'b0111;
														assign node16336 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node16339 = (inp[5]) ? 4'b0111 : node16340;
														assign node16340 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node16344 = (inp[5]) ? 4'b0110 : node16345;
													assign node16345 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node16349 = (inp[7]) ? node16365 : node16350;
											assign node16350 = (inp[5]) ? node16358 : node16351;
												assign node16351 = (inp[9]) ? node16355 : node16352;
													assign node16352 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node16355 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node16358 = (inp[15]) ? node16360 : 4'b0011;
													assign node16360 = (inp[2]) ? node16362 : 4'b0111;
														assign node16362 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node16365 = (inp[0]) ? node16383 : node16366;
												assign node16366 = (inp[9]) ? node16376 : node16367;
													assign node16367 = (inp[15]) ? node16371 : node16368;
														assign node16368 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node16371 = (inp[4]) ? node16373 : 4'b0010;
															assign node16373 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node16376 = (inp[15]) ? 4'b0010 : node16377;
														assign node16377 = (inp[2]) ? node16379 : 4'b0110;
															assign node16379 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node16383 = (inp[4]) ? 4'b0010 : node16384;
													assign node16384 = (inp[5]) ? 4'b0110 : node16385;
														assign node16385 = (inp[2]) ? node16387 : 4'b0110;
															assign node16387 = (inp[15]) ? 4'b0111 : 4'b0011;
							assign node16392 = (inp[7]) ? node16542 : node16393;
								assign node16393 = (inp[2]) ? node16467 : node16394;
									assign node16394 = (inp[15]) ? node16434 : node16395;
										assign node16395 = (inp[5]) ? node16419 : node16396;
											assign node16396 = (inp[4]) ? node16406 : node16397;
												assign node16397 = (inp[1]) ? node16403 : node16398;
													assign node16398 = (inp[10]) ? 4'b0011 : node16399;
														assign node16399 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node16403 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node16406 = (inp[10]) ? node16412 : node16407;
													assign node16407 = (inp[13]) ? 4'b0010 : node16408;
														assign node16408 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node16412 = (inp[0]) ? node16416 : node16413;
														assign node16413 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node16416 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node16419 = (inp[4]) ? node16421 : 4'b0110;
												assign node16421 = (inp[9]) ? node16427 : node16422;
													assign node16422 = (inp[10]) ? 4'b0011 : node16423;
														assign node16423 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node16427 = (inp[1]) ? node16429 : 4'b0010;
														assign node16429 = (inp[10]) ? node16431 : 4'b0010;
															assign node16431 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node16434 = (inp[4]) ? node16448 : node16435;
											assign node16435 = (inp[5]) ? node16443 : node16436;
												assign node16436 = (inp[1]) ? node16440 : node16437;
													assign node16437 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node16440 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node16443 = (inp[1]) ? node16445 : 4'b0011;
													assign node16445 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node16448 = (inp[5]) ? node16456 : node16449;
												assign node16449 = (inp[1]) ? node16453 : node16450;
													assign node16450 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node16453 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node16456 = (inp[9]) ? node16462 : node16457;
													assign node16457 = (inp[1]) ? node16459 : 4'b0110;
														assign node16459 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node16462 = (inp[1]) ? 4'b0110 : node16463;
														assign node16463 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node16467 = (inp[15]) ? node16501 : node16468;
										assign node16468 = (inp[5]) ? node16480 : node16469;
											assign node16469 = (inp[9]) ? node16471 : 4'b0110;
												assign node16471 = (inp[10]) ? 4'b0110 : node16472;
													assign node16472 = (inp[1]) ? 4'b0111 : node16473;
														assign node16473 = (inp[13]) ? node16475 : 4'b0110;
															assign node16475 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node16480 = (inp[4]) ? node16494 : node16481;
												assign node16481 = (inp[0]) ? node16487 : node16482;
													assign node16482 = (inp[10]) ? node16484 : 4'b0011;
														assign node16484 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node16487 = (inp[1]) ? node16489 : 4'b0010;
														assign node16489 = (inp[13]) ? 4'b0011 : node16490;
															assign node16490 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node16494 = (inp[1]) ? node16496 : 4'b0111;
													assign node16496 = (inp[13]) ? node16498 : 4'b0110;
														assign node16498 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node16501 = (inp[4]) ? node16517 : node16502;
											assign node16502 = (inp[5]) ? node16512 : node16503;
												assign node16503 = (inp[13]) ? node16505 : 4'b0111;
													assign node16505 = (inp[0]) ? node16507 : 4'b0110;
														assign node16507 = (inp[10]) ? 4'b0111 : node16508;
															assign node16508 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node16512 = (inp[9]) ? 4'b0110 : node16513;
													assign node16513 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node16517 = (inp[0]) ? node16533 : node16518;
												assign node16518 = (inp[5]) ? node16522 : node16519;
													assign node16519 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node16522 = (inp[13]) ? 4'b0010 : node16523;
														assign node16523 = (inp[9]) ? 4'b0010 : node16524;
															assign node16524 = (inp[1]) ? node16528 : node16525;
																assign node16525 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node16528 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node16533 = (inp[13]) ? node16535 : 4'b0011;
													assign node16535 = (inp[1]) ? 4'b0010 : node16536;
														assign node16536 = (inp[10]) ? node16538 : 4'b0011;
															assign node16538 = (inp[5]) ? 4'b0011 : 4'b0010;
								assign node16542 = (inp[2]) ? node16638 : node16543;
									assign node16543 = (inp[4]) ? node16589 : node16544;
										assign node16544 = (inp[15]) ? node16568 : node16545;
											assign node16545 = (inp[5]) ? node16565 : node16546;
												assign node16546 = (inp[1]) ? node16558 : node16547;
													assign node16547 = (inp[9]) ? node16549 : 4'b0111;
														assign node16549 = (inp[0]) ? node16553 : node16550;
															assign node16550 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node16553 = (inp[10]) ? node16555 : 4'b0111;
																assign node16555 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node16558 = (inp[10]) ? node16562 : node16559;
														assign node16559 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node16562 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node16565 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node16568 = (inp[1]) ? node16582 : node16569;
												assign node16569 = (inp[9]) ? node16571 : 4'b0010;
													assign node16571 = (inp[13]) ? node16573 : 4'b0010;
														assign node16573 = (inp[0]) ? 4'b0010 : node16574;
															assign node16574 = (inp[10]) ? node16578 : node16575;
																assign node16575 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node16578 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node16582 = (inp[9]) ? 4'b0011 : node16583;
													assign node16583 = (inp[10]) ? 4'b0010 : node16584;
														assign node16584 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node16589 = (inp[13]) ? node16615 : node16590;
											assign node16590 = (inp[9]) ? node16610 : node16591;
												assign node16591 = (inp[15]) ? node16597 : node16592;
													assign node16592 = (inp[0]) ? 4'b0110 : node16593;
														assign node16593 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node16597 = (inp[5]) ? node16605 : node16598;
														assign node16598 = (inp[0]) ? node16600 : 4'b0111;
															assign node16600 = (inp[1]) ? node16602 : 4'b0111;
																assign node16602 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node16605 = (inp[10]) ? 4'b0111 : node16606;
															assign node16606 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node16610 = (inp[0]) ? node16612 : 4'b0110;
													assign node16612 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node16615 = (inp[0]) ? node16627 : node16616;
												assign node16616 = (inp[9]) ? node16618 : 4'b0111;
													assign node16618 = (inp[15]) ? node16622 : node16619;
														assign node16619 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node16622 = (inp[1]) ? 4'b0111 : node16623;
															assign node16623 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node16627 = (inp[15]) ? node16633 : node16628;
													assign node16628 = (inp[1]) ? 4'b0110 : node16629;
														assign node16629 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node16633 = (inp[10]) ? 4'b0111 : node16634;
														assign node16634 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node16638 = (inp[4]) ? node16672 : node16639;
										assign node16639 = (inp[15]) ? node16665 : node16640;
											assign node16640 = (inp[5]) ? node16652 : node16641;
												assign node16641 = (inp[0]) ? node16647 : node16642;
													assign node16642 = (inp[1]) ? node16644 : 4'b0011;
														assign node16644 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node16647 = (inp[10]) ? 4'b0010 : node16648;
														assign node16648 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node16652 = (inp[1]) ? node16660 : node16653;
													assign node16653 = (inp[9]) ? node16657 : node16654;
														assign node16654 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node16657 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node16660 = (inp[0]) ? 4'b0110 : node16661;
														assign node16661 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node16665 = (inp[10]) ? node16669 : node16666;
												assign node16666 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node16669 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node16672 = (inp[15]) ? node16690 : node16673;
											assign node16673 = (inp[13]) ? node16685 : node16674;
												assign node16674 = (inp[5]) ? node16680 : node16675;
													assign node16675 = (inp[0]) ? 4'b0011 : node16676;
														assign node16676 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node16680 = (inp[1]) ? node16682 : 4'b0010;
														assign node16682 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node16685 = (inp[1]) ? node16687 : 4'b0011;
													assign node16687 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node16690 = (inp[5]) ? node16696 : node16691;
												assign node16691 = (inp[1]) ? 4'b0010 : node16692;
													assign node16692 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node16696 = (inp[1]) ? 4'b0011 : 4'b0010;
					assign node16699 = (inp[15]) ? node17139 : node16700;
						assign node16700 = (inp[14]) ? node16962 : node16701;
							assign node16701 = (inp[11]) ? node16813 : node16702;
								assign node16702 = (inp[13]) ? node16758 : node16703;
									assign node16703 = (inp[2]) ? node16717 : node16704;
										assign node16704 = (inp[5]) ? node16708 : node16705;
											assign node16705 = (inp[7]) ? 4'b0110 : 4'b0010;
											assign node16708 = (inp[7]) ? node16712 : node16709;
												assign node16709 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node16712 = (inp[4]) ? 4'b0010 : node16713;
													assign node16713 = (inp[10]) ? 4'b0010 : 4'b0011;
										assign node16717 = (inp[4]) ? node16743 : node16718;
											assign node16718 = (inp[1]) ? node16736 : node16719;
												assign node16719 = (inp[10]) ? node16725 : node16720;
													assign node16720 = (inp[7]) ? 4'b0110 : node16721;
														assign node16721 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node16725 = (inp[9]) ? 4'b0010 : node16726;
														assign node16726 = (inp[0]) ? node16728 : 4'b0010;
															assign node16728 = (inp[7]) ? node16732 : node16729;
																assign node16729 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node16732 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node16736 = (inp[5]) ? node16740 : node16737;
													assign node16737 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node16740 = (inp[7]) ? 4'b0010 : 4'b0111;
											assign node16743 = (inp[1]) ? node16751 : node16744;
												assign node16744 = (inp[7]) ? node16748 : node16745;
													assign node16745 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node16748 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node16751 = (inp[0]) ? node16753 : 4'b0010;
													assign node16753 = (inp[7]) ? node16755 : 4'b0110;
														assign node16755 = (inp[5]) ? 4'b0010 : 4'b0110;
									assign node16758 = (inp[1]) ? node16788 : node16759;
										assign node16759 = (inp[7]) ? node16767 : node16760;
											assign node16760 = (inp[5]) ? 4'b0111 : node16761;
												assign node16761 = (inp[2]) ? node16763 : 4'b0011;
													assign node16763 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node16767 = (inp[5]) ? node16773 : node16768;
												assign node16768 = (inp[4]) ? node16770 : 4'b0111;
													assign node16770 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node16773 = (inp[10]) ? node16783 : node16774;
													assign node16774 = (inp[0]) ? node16776 : 4'b0011;
														assign node16776 = (inp[4]) ? node16780 : node16777;
															assign node16777 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node16780 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node16783 = (inp[0]) ? 4'b0010 : node16784;
														assign node16784 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node16788 = (inp[0]) ? node16796 : node16789;
											assign node16789 = (inp[5]) ? node16793 : node16790;
												assign node16790 = (inp[4]) ? 4'b0011 : 4'b0110;
												assign node16793 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node16796 = (inp[2]) ? node16804 : node16797;
												assign node16797 = (inp[7]) ? node16801 : node16798;
													assign node16798 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node16801 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node16804 = (inp[7]) ? node16808 : node16805;
													assign node16805 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node16808 = (inp[5]) ? 4'b0011 : node16809;
														assign node16809 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node16813 = (inp[13]) ? node16883 : node16814;
									assign node16814 = (inp[10]) ? node16854 : node16815;
										assign node16815 = (inp[0]) ? node16839 : node16816;
											assign node16816 = (inp[2]) ? node16828 : node16817;
												assign node16817 = (inp[1]) ? node16823 : node16818;
													assign node16818 = (inp[9]) ? 4'b0011 : node16819;
														assign node16819 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node16823 = (inp[4]) ? node16825 : 4'b0011;
														assign node16825 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node16828 = (inp[1]) ? node16834 : node16829;
													assign node16829 = (inp[7]) ? 4'b0011 : node16830;
														assign node16830 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node16834 = (inp[7]) ? node16836 : 4'b0010;
														assign node16836 = (inp[4]) ? 4'b0111 : 4'b0110;
											assign node16839 = (inp[5]) ? node16847 : node16840;
												assign node16840 = (inp[7]) ? 4'b0111 : node16841;
													assign node16841 = (inp[4]) ? 4'b0011 : node16842;
														assign node16842 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node16847 = (inp[1]) ? node16849 : 4'b0111;
													assign node16849 = (inp[2]) ? node16851 : 4'b0110;
														assign node16851 = (inp[4]) ? 4'b0111 : 4'b0110;
										assign node16854 = (inp[5]) ? node16870 : node16855;
											assign node16855 = (inp[7]) ? node16857 : 4'b0011;
												assign node16857 = (inp[2]) ? node16859 : 4'b0111;
													assign node16859 = (inp[9]) ? node16865 : node16860;
														assign node16860 = (inp[1]) ? 4'b0110 : node16861;
															assign node16861 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node16865 = (inp[1]) ? node16867 : 4'b0110;
															assign node16867 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node16870 = (inp[7]) ? node16878 : node16871;
												assign node16871 = (inp[1]) ? node16873 : 4'b0111;
													assign node16873 = (inp[9]) ? 4'b0110 : node16874;
														assign node16874 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node16878 = (inp[4]) ? 4'b0011 : node16879;
													assign node16879 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node16883 = (inp[4]) ? node16929 : node16884;
										assign node16884 = (inp[9]) ? node16908 : node16885;
											assign node16885 = (inp[1]) ? node16897 : node16886;
												assign node16886 = (inp[0]) ? node16892 : node16887;
													assign node16887 = (inp[7]) ? 4'b0110 : node16888;
														assign node16888 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node16892 = (inp[7]) ? 4'b0010 : node16893;
														assign node16893 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node16897 = (inp[2]) ? node16905 : node16898;
													assign node16898 = (inp[10]) ? node16902 : node16899;
														assign node16899 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node16902 = (inp[0]) ? 4'b0010 : 4'b0110;
													assign node16905 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node16908 = (inp[10]) ? node16922 : node16909;
												assign node16909 = (inp[0]) ? node16915 : node16910;
													assign node16910 = (inp[2]) ? 4'b0010 : node16911;
														assign node16911 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node16915 = (inp[2]) ? node16919 : node16916;
														assign node16916 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node16919 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node16922 = (inp[2]) ? 4'b0111 : node16923;
													assign node16923 = (inp[5]) ? node16925 : 4'b0110;
														assign node16925 = (inp[1]) ? 4'b0110 : 4'b0011;
										assign node16929 = (inp[0]) ? node16939 : node16930;
											assign node16930 = (inp[7]) ? node16936 : node16931;
												assign node16931 = (inp[5]) ? node16933 : 4'b0010;
													assign node16933 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node16936 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node16939 = (inp[10]) ? node16949 : node16940;
												assign node16940 = (inp[1]) ? node16944 : node16941;
													assign node16941 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node16944 = (inp[2]) ? node16946 : 4'b0110;
														assign node16946 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node16949 = (inp[9]) ? node16955 : node16950;
													assign node16950 = (inp[2]) ? node16952 : 4'b0111;
														assign node16952 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node16955 = (inp[1]) ? node16957 : 4'b0110;
														assign node16957 = (inp[7]) ? 4'b0110 : node16958;
															assign node16958 = (inp[2]) ? 4'b0110 : 4'b0111;
							assign node16962 = (inp[9]) ? node17048 : node16963;
								assign node16963 = (inp[13]) ? node17011 : node16964;
									assign node16964 = (inp[1]) ? node16984 : node16965;
										assign node16965 = (inp[11]) ? node16971 : node16966;
											assign node16966 = (inp[2]) ? node16968 : 4'b0000;
												assign node16968 = (inp[7]) ? 4'b0100 : 4'b0001;
											assign node16971 = (inp[7]) ? node16977 : node16972;
												assign node16972 = (inp[5]) ? 4'b0101 : node16973;
													assign node16973 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node16977 = (inp[4]) ? 4'b0000 : node16978;
													assign node16978 = (inp[10]) ? 4'b0100 : node16979;
														assign node16979 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node16984 = (inp[5]) ? node17004 : node16985;
											assign node16985 = (inp[2]) ? node16997 : node16986;
												assign node16986 = (inp[10]) ? node16992 : node16987;
													assign node16987 = (inp[7]) ? node16989 : 4'b0100;
														assign node16989 = (inp[4]) ? 4'b0001 : 4'b0100;
													assign node16992 = (inp[4]) ? 4'b0100 : node16993;
														assign node16993 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node16997 = (inp[7]) ? node17001 : node16998;
													assign node16998 = (inp[4]) ? 4'b0100 : 4'b0001;
													assign node17001 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node17004 = (inp[4]) ? node17008 : node17005;
												assign node17005 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node17008 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node17011 = (inp[1]) ? node17031 : node17012;
										assign node17012 = (inp[7]) ? node17020 : node17013;
											assign node17013 = (inp[4]) ? node17017 : node17014;
												assign node17014 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node17017 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node17020 = (inp[4]) ? 4'b0001 : node17021;
												assign node17021 = (inp[11]) ? node17027 : node17022;
													assign node17022 = (inp[2]) ? node17024 : 4'b0101;
														assign node17024 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node17027 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node17031 = (inp[7]) ? node17043 : node17032;
											assign node17032 = (inp[4]) ? node17040 : node17033;
												assign node17033 = (inp[2]) ? node17037 : node17034;
													assign node17034 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node17037 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node17040 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node17043 = (inp[4]) ? 4'b0000 : node17044;
												assign node17044 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node17048 = (inp[4]) ? node17104 : node17049;
									assign node17049 = (inp[7]) ? node17073 : node17050;
										assign node17050 = (inp[5]) ? node17064 : node17051;
											assign node17051 = (inp[1]) ? node17055 : node17052;
												assign node17052 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node17055 = (inp[11]) ? 4'b0001 : node17056;
													assign node17056 = (inp[2]) ? node17060 : node17057;
														assign node17057 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node17060 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node17064 = (inp[2]) ? node17066 : 4'b0001;
												assign node17066 = (inp[13]) ? node17070 : node17067;
													assign node17067 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node17070 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node17073 = (inp[1]) ? node17091 : node17074;
											assign node17074 = (inp[5]) ? node17080 : node17075;
												assign node17075 = (inp[13]) ? 4'b0101 : node17076;
													assign node17076 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node17080 = (inp[0]) ? node17088 : node17081;
													assign node17081 = (inp[2]) ? node17085 : node17082;
														assign node17082 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node17085 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node17088 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node17091 = (inp[5]) ? node17099 : node17092;
												assign node17092 = (inp[13]) ? node17096 : node17093;
													assign node17093 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node17096 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node17099 = (inp[13]) ? 4'b0100 : node17100;
													assign node17100 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node17104 = (inp[7]) ? node17112 : node17105;
										assign node17105 = (inp[5]) ? node17109 : node17106;
											assign node17106 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node17109 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node17112 = (inp[11]) ? node17132 : node17113;
											assign node17113 = (inp[2]) ? node17119 : node17114;
												assign node17114 = (inp[0]) ? 4'b0000 : node17115;
													assign node17115 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node17119 = (inp[0]) ? node17125 : node17120;
													assign node17120 = (inp[10]) ? node17122 : 4'b0000;
														assign node17122 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node17125 = (inp[10]) ? node17127 : 4'b0001;
														assign node17127 = (inp[13]) ? node17129 : 4'b0000;
															assign node17129 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node17132 = (inp[1]) ? node17136 : node17133;
												assign node17133 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node17136 = (inp[13]) ? 4'b0000 : 4'b0001;
						assign node17139 = (inp[4]) ? node17257 : node17140;
							assign node17140 = (inp[5]) ? node17228 : node17141;
								assign node17141 = (inp[14]) ? node17201 : node17142;
									assign node17142 = (inp[7]) ? node17166 : node17143;
										assign node17143 = (inp[0]) ? node17151 : node17144;
											assign node17144 = (inp[1]) ? node17148 : node17145;
												assign node17145 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node17148 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node17151 = (inp[9]) ? node17159 : node17152;
												assign node17152 = (inp[11]) ? node17156 : node17153;
													assign node17153 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node17156 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node17159 = (inp[11]) ? node17163 : node17160;
													assign node17160 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node17163 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node17166 = (inp[13]) ? node17182 : node17167;
											assign node17167 = (inp[0]) ? 4'b0000 : node17168;
												assign node17168 = (inp[10]) ? node17174 : node17169;
													assign node17169 = (inp[11]) ? node17171 : 4'b0001;
														assign node17171 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node17174 = (inp[11]) ? 4'b0000 : node17175;
														assign node17175 = (inp[1]) ? 4'b0000 : node17176;
															assign node17176 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node17182 = (inp[10]) ? node17192 : node17183;
												assign node17183 = (inp[1]) ? 4'b0000 : node17184;
													assign node17184 = (inp[9]) ? 4'b0000 : node17185;
														assign node17185 = (inp[0]) ? 4'b0001 : node17186;
															assign node17186 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node17192 = (inp[9]) ? 4'b0001 : node17193;
													assign node17193 = (inp[11]) ? node17197 : node17194;
														assign node17194 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node17197 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node17201 = (inp[10]) ? node17209 : node17202;
										assign node17202 = (inp[2]) ? node17206 : node17203;
											assign node17203 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node17206 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node17209 = (inp[13]) ? node17223 : node17210;
											assign node17210 = (inp[7]) ? node17216 : node17211;
												assign node17211 = (inp[11]) ? node17213 : 4'b0101;
													assign node17213 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node17216 = (inp[2]) ? node17220 : node17217;
													assign node17217 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node17220 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node17223 = (inp[2]) ? 4'b0100 : node17224;
												assign node17224 = (inp[1]) ? 4'b0101 : 4'b0100;
								assign node17228 = (inp[2]) ? node17246 : node17229;
									assign node17229 = (inp[1]) ? node17239 : node17230;
										assign node17230 = (inp[14]) ? 4'b0100 : node17231;
											assign node17231 = (inp[7]) ? node17235 : node17232;
												assign node17232 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node17235 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node17239 = (inp[14]) ? 4'b0101 : node17240;
											assign node17240 = (inp[11]) ? 4'b0101 : node17241;
												assign node17241 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node17246 = (inp[1]) ? node17252 : node17247;
										assign node17247 = (inp[14]) ? 4'b0101 : node17248;
											assign node17248 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node17252 = (inp[11]) ? 4'b0100 : node17253;
											assign node17253 = (inp[14]) ? 4'b0100 : 4'b0101;
							assign node17257 = (inp[5]) ? node17365 : node17258;
								assign node17258 = (inp[14]) ? node17308 : node17259;
									assign node17259 = (inp[0]) ? node17281 : node17260;
										assign node17260 = (inp[9]) ? node17268 : node17261;
											assign node17261 = (inp[13]) ? node17263 : 4'b0101;
												assign node17263 = (inp[2]) ? 4'b0101 : node17264;
													assign node17264 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node17268 = (inp[7]) ? node17276 : node17269;
												assign node17269 = (inp[11]) ? 4'b0100 : node17270;
													assign node17270 = (inp[13]) ? node17272 : 4'b0100;
														assign node17272 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node17276 = (inp[1]) ? 4'b0101 : node17277;
													assign node17277 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node17281 = (inp[7]) ? node17303 : node17282;
											assign node17282 = (inp[10]) ? node17288 : node17283;
												assign node17283 = (inp[1]) ? 4'b0100 : node17284;
													assign node17284 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node17288 = (inp[2]) ? node17298 : node17289;
													assign node17289 = (inp[13]) ? node17293 : node17290;
														assign node17290 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node17293 = (inp[1]) ? 4'b0100 : node17294;
															assign node17294 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node17298 = (inp[11]) ? 4'b0101 : node17299;
														assign node17299 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node17303 = (inp[11]) ? node17305 : 4'b0100;
												assign node17305 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node17308 = (inp[0]) ? node17328 : node17309;
										assign node17309 = (inp[9]) ? node17317 : node17310;
											assign node17310 = (inp[1]) ? node17314 : node17311;
												assign node17311 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node17314 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node17317 = (inp[11]) ? node17323 : node17318;
												assign node17318 = (inp[1]) ? node17320 : 4'b0001;
													assign node17320 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node17323 = (inp[1]) ? 4'b0001 : node17324;
													assign node17324 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node17328 = (inp[9]) ? node17346 : node17329;
											assign node17329 = (inp[10]) ? 4'b0001 : node17330;
												assign node17330 = (inp[13]) ? node17340 : node17331;
													assign node17331 = (inp[11]) ? node17337 : node17332;
														assign node17332 = (inp[7]) ? 4'b0001 : node17333;
															assign node17333 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node17337 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node17340 = (inp[11]) ? 4'b0001 : node17341;
														assign node17341 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node17346 = (inp[13]) ? node17354 : node17347;
												assign node17347 = (inp[10]) ? 4'b0001 : node17348;
													assign node17348 = (inp[1]) ? node17350 : 4'b0000;
														assign node17350 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node17354 = (inp[10]) ? node17360 : node17355;
													assign node17355 = (inp[1]) ? node17357 : 4'b0001;
														assign node17357 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17360 = (inp[7]) ? node17362 : 4'b0000;
														assign node17362 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node17365 = (inp[1]) ? node17379 : node17366;
									assign node17366 = (inp[14]) ? 4'b0001 : node17367;
										assign node17367 = (inp[11]) ? node17373 : node17368;
											assign node17368 = (inp[7]) ? 4'b0000 : node17369;
												assign node17369 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node17373 = (inp[2]) ? 4'b0001 : node17374;
												assign node17374 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node17379 = (inp[14]) ? 4'b0000 : node17380;
										assign node17380 = (inp[11]) ? node17386 : node17381;
											assign node17381 = (inp[7]) ? 4'b0001 : node17382;
												assign node17382 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node17386 = (inp[2]) ? 4'b0000 : node17387;
												assign node17387 = (inp[7]) ? 4'b0000 : 4'b0001;
				assign node17392 = (inp[14]) ? node18234 : node17393;
					assign node17393 = (inp[15]) ? node18037 : node17394;
						assign node17394 = (inp[11]) ? node17754 : node17395;
							assign node17395 = (inp[13]) ? node17577 : node17396;
								assign node17396 = (inp[6]) ? node17504 : node17397;
									assign node17397 = (inp[5]) ? node17443 : node17398;
										assign node17398 = (inp[10]) ? node17416 : node17399;
											assign node17399 = (inp[7]) ? node17409 : node17400;
												assign node17400 = (inp[1]) ? node17404 : node17401;
													assign node17401 = (inp[4]) ? 4'b0011 : 4'b0110;
													assign node17404 = (inp[0]) ? node17406 : 4'b0111;
														assign node17406 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node17409 = (inp[2]) ? node17413 : node17410;
													assign node17410 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node17413 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node17416 = (inp[4]) ? node17428 : node17417;
												assign node17417 = (inp[7]) ? node17425 : node17418;
													assign node17418 = (inp[1]) ? node17422 : node17419;
														assign node17419 = (inp[0]) ? 4'b0111 : 4'b0011;
														assign node17422 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node17425 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node17428 = (inp[1]) ? node17436 : node17429;
													assign node17429 = (inp[2]) ? node17433 : node17430;
														assign node17430 = (inp[7]) ? 4'b0010 : 4'b0111;
														assign node17433 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node17436 = (inp[9]) ? 4'b0110 : node17437;
														assign node17437 = (inp[7]) ? 4'b0011 : node17438;
															assign node17438 = (inp[0]) ? 4'b0110 : 4'b0010;
										assign node17443 = (inp[0]) ? node17475 : node17444;
											assign node17444 = (inp[4]) ? node17456 : node17445;
												assign node17445 = (inp[1]) ? node17453 : node17446;
													assign node17446 = (inp[10]) ? 4'b0110 : node17447;
														assign node17447 = (inp[2]) ? node17449 : 4'b0010;
															assign node17449 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node17453 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node17456 = (inp[10]) ? node17468 : node17457;
													assign node17457 = (inp[9]) ? node17463 : node17458;
														assign node17458 = (inp[1]) ? node17460 : 4'b0110;
															assign node17460 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node17463 = (inp[1]) ? 4'b0110 : node17464;
															assign node17464 = (inp[2]) ? 4'b0110 : 4'b0011;
													assign node17468 = (inp[7]) ? node17470 : 4'b0010;
														assign node17470 = (inp[1]) ? 4'b0010 : node17471;
															assign node17471 = (inp[2]) ? 4'b0011 : 4'b0111;
											assign node17475 = (inp[4]) ? node17485 : node17476;
												assign node17476 = (inp[10]) ? node17480 : node17477;
													assign node17477 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node17480 = (inp[7]) ? node17482 : 4'b0011;
														assign node17482 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node17485 = (inp[10]) ? node17497 : node17486;
													assign node17486 = (inp[9]) ? 4'b0110 : node17487;
														assign node17487 = (inp[7]) ? node17493 : node17488;
															assign node17488 = (inp[2]) ? node17490 : 4'b0011;
																assign node17490 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node17493 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node17497 = (inp[2]) ? node17501 : node17498;
														assign node17498 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node17501 = (inp[1]) ? 4'b0110 : 4'b0111;
									assign node17504 = (inp[10]) ? node17552 : node17505;
										assign node17505 = (inp[2]) ? node17533 : node17506;
											assign node17506 = (inp[5]) ? node17512 : node17507;
												assign node17507 = (inp[7]) ? node17509 : 4'b0010;
													assign node17509 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node17512 = (inp[7]) ? node17524 : node17513;
													assign node17513 = (inp[9]) ? 4'b0111 : node17514;
														assign node17514 = (inp[0]) ? node17520 : node17515;
															assign node17515 = (inp[1]) ? 4'b0110 : node17516;
																assign node17516 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node17520 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node17524 = (inp[0]) ? 4'b0010 : node17525;
														assign node17525 = (inp[9]) ? node17527 : 4'b0011;
															assign node17527 = (inp[4]) ? 4'b0010 : node17528;
																assign node17528 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node17533 = (inp[1]) ? node17547 : node17534;
												assign node17534 = (inp[0]) ? node17540 : node17535;
													assign node17535 = (inp[5]) ? node17537 : 4'b0010;
														assign node17537 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node17540 = (inp[9]) ? node17544 : node17541;
														assign node17541 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node17544 = (inp[7]) ? 4'b0010 : 4'b0110;
												assign node17547 = (inp[4]) ? node17549 : 4'b0010;
													assign node17549 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node17552 = (inp[7]) ? node17564 : node17553;
											assign node17553 = (inp[5]) ? node17559 : node17554;
												assign node17554 = (inp[2]) ? node17556 : 4'b0010;
													assign node17556 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node17559 = (inp[1]) ? 4'b0110 : node17560;
													assign node17560 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node17564 = (inp[5]) ? node17574 : node17565;
												assign node17565 = (inp[1]) ? 4'b0110 : node17566;
													assign node17566 = (inp[2]) ? node17570 : node17567;
														assign node17567 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node17570 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node17574 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node17577 = (inp[0]) ? node17679 : node17578;
									assign node17578 = (inp[6]) ? node17642 : node17579;
										assign node17579 = (inp[7]) ? node17607 : node17580;
											assign node17580 = (inp[2]) ? node17596 : node17581;
												assign node17581 = (inp[5]) ? node17587 : node17582;
													assign node17582 = (inp[4]) ? node17584 : 4'b0010;
														assign node17584 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node17587 = (inp[1]) ? 4'b0011 : node17588;
														assign node17588 = (inp[4]) ? node17592 : node17589;
															assign node17589 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node17592 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node17596 = (inp[9]) ? node17598 : 4'b0110;
													assign node17598 = (inp[1]) ? node17602 : node17599;
														assign node17599 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node17602 = (inp[4]) ? node17604 : 4'b0111;
															assign node17604 = (inp[5]) ? 4'b0111 : 4'b0011;
											assign node17607 = (inp[2]) ? node17627 : node17608;
												assign node17608 = (inp[4]) ? node17616 : node17609;
													assign node17609 = (inp[1]) ? 4'b0110 : node17610;
														assign node17610 = (inp[9]) ? node17612 : 4'b0111;
															assign node17612 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node17616 = (inp[5]) ? node17624 : node17617;
														assign node17617 = (inp[9]) ? node17619 : 4'b0011;
															assign node17619 = (inp[1]) ? 4'b0010 : node17620;
																assign node17620 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node17624 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node17627 = (inp[5]) ? node17637 : node17628;
													assign node17628 = (inp[4]) ? node17632 : node17629;
														assign node17629 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node17632 = (inp[9]) ? 4'b0110 : node17633;
															assign node17633 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node17637 = (inp[10]) ? 4'b0010 : node17638;
														assign node17638 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node17642 = (inp[2]) ? node17666 : node17643;
											assign node17643 = (inp[5]) ? node17653 : node17644;
												assign node17644 = (inp[7]) ? node17648 : node17645;
													assign node17645 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node17648 = (inp[4]) ? node17650 : 4'b0111;
														assign node17650 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node17653 = (inp[7]) ? node17659 : node17654;
													assign node17654 = (inp[4]) ? node17656 : 4'b0110;
														assign node17656 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node17659 = (inp[1]) ? node17663 : node17660;
														assign node17660 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node17663 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node17666 = (inp[7]) ? node17674 : node17667;
												assign node17667 = (inp[5]) ? 4'b0111 : node17668;
													assign node17668 = (inp[1]) ? node17670 : 4'b0011;
														assign node17670 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node17674 = (inp[5]) ? 4'b0011 : node17675;
													assign node17675 = (inp[10]) ? 4'b0110 : 4'b0111;
									assign node17679 = (inp[5]) ? node17717 : node17680;
										assign node17680 = (inp[7]) ? node17696 : node17681;
											assign node17681 = (inp[6]) ? 4'b0011 : node17682;
												assign node17682 = (inp[1]) ? node17690 : node17683;
													assign node17683 = (inp[9]) ? node17687 : node17684;
														assign node17684 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node17687 = (inp[4]) ? 4'b0011 : 4'b0110;
													assign node17690 = (inp[2]) ? 4'b0011 : node17691;
														assign node17691 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node17696 = (inp[9]) ? node17702 : node17697;
												assign node17697 = (inp[6]) ? 4'b0111 : node17698;
													assign node17698 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node17702 = (inp[10]) ? node17708 : node17703;
													assign node17703 = (inp[1]) ? node17705 : 4'b0111;
														assign node17705 = (inp[6]) ? 4'b0111 : 4'b0110;
													assign node17708 = (inp[1]) ? 4'b0111 : node17709;
														assign node17709 = (inp[4]) ? node17713 : node17710;
															assign node17710 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node17713 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node17717 = (inp[2]) ? node17747 : node17718;
											assign node17718 = (inp[6]) ? node17732 : node17719;
												assign node17719 = (inp[7]) ? 4'b0110 : node17720;
													assign node17720 = (inp[4]) ? node17726 : node17721;
														assign node17721 = (inp[1]) ? node17723 : 4'b0011;
															assign node17723 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node17726 = (inp[1]) ? node17728 : 4'b0010;
															assign node17728 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node17732 = (inp[7]) ? node17740 : node17733;
													assign node17733 = (inp[4]) ? node17737 : node17734;
														assign node17734 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node17737 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node17740 = (inp[9]) ? node17742 : 4'b0011;
														assign node17742 = (inp[4]) ? 4'b0010 : node17743;
															assign node17743 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node17747 = (inp[7]) ? node17749 : 4'b0111;
												assign node17749 = (inp[4]) ? 4'b0011 : node17750;
													assign node17750 = (inp[6]) ? 4'b0011 : 4'b0010;
							assign node17754 = (inp[13]) ? node17878 : node17755;
								assign node17755 = (inp[6]) ? node17813 : node17756;
									assign node17756 = (inp[10]) ? node17784 : node17757;
										assign node17757 = (inp[2]) ? node17771 : node17758;
											assign node17758 = (inp[1]) ? node17762 : node17759;
												assign node17759 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node17762 = (inp[7]) ? node17766 : node17763;
													assign node17763 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node17766 = (inp[5]) ? node17768 : 4'b0011;
														assign node17768 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node17771 = (inp[9]) ? 4'b0110 : node17772;
												assign node17772 = (inp[5]) ? node17780 : node17773;
													assign node17773 = (inp[1]) ? 4'b0011 : node17774;
														assign node17774 = (inp[7]) ? node17776 : 4'b0110;
															assign node17776 = (inp[4]) ? 4'b0110 : 4'b0011;
													assign node17780 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node17784 = (inp[7]) ? node17796 : node17785;
											assign node17785 = (inp[2]) ? node17791 : node17786;
												assign node17786 = (inp[4]) ? node17788 : 4'b0011;
													assign node17788 = (inp[5]) ? 4'b0010 : 4'b0111;
												assign node17791 = (inp[4]) ? node17793 : 4'b0111;
													assign node17793 = (inp[5]) ? 4'b0111 : 4'b0011;
											assign node17796 = (inp[2]) ? node17808 : node17797;
												assign node17797 = (inp[1]) ? node17803 : node17798;
													assign node17798 = (inp[4]) ? node17800 : 4'b0110;
														assign node17800 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node17803 = (inp[4]) ? node17805 : 4'b0111;
														assign node17805 = (inp[5]) ? 4'b0111 : 4'b0010;
												assign node17808 = (inp[5]) ? 4'b0011 : node17809;
													assign node17809 = (inp[4]) ? 4'b0111 : 4'b0010;
									assign node17813 = (inp[1]) ? node17839 : node17814;
										assign node17814 = (inp[4]) ? node17828 : node17815;
											assign node17815 = (inp[2]) ? node17821 : node17816;
												assign node17816 = (inp[10]) ? node17818 : 4'b0111;
													assign node17818 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node17821 = (inp[10]) ? 4'b0111 : node17822;
													assign node17822 = (inp[5]) ? 4'b0011 : node17823;
														assign node17823 = (inp[7]) ? 4'b0110 : 4'b0011;
											assign node17828 = (inp[2]) ? node17830 : 4'b0010;
												assign node17830 = (inp[9]) ? node17832 : 4'b0011;
													assign node17832 = (inp[0]) ? 4'b0011 : node17833;
														assign node17833 = (inp[7]) ? node17835 : 4'b0111;
															assign node17835 = (inp[5]) ? 4'b0011 : 4'b0111;
										assign node17839 = (inp[4]) ? node17855 : node17840;
											assign node17840 = (inp[2]) ? node17848 : node17841;
												assign node17841 = (inp[7]) ? node17845 : node17842;
													assign node17842 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node17845 = (inp[5]) ? 4'b0010 : 4'b0111;
												assign node17848 = (inp[9]) ? 4'b0011 : node17849;
													assign node17849 = (inp[5]) ? 4'b0111 : node17850;
														assign node17850 = (inp[10]) ? 4'b0111 : 4'b0011;
											assign node17855 = (inp[2]) ? node17871 : node17856;
												assign node17856 = (inp[9]) ? node17866 : node17857;
													assign node17857 = (inp[0]) ? 4'b0011 : node17858;
														assign node17858 = (inp[10]) ? node17860 : 4'b0011;
															assign node17860 = (inp[7]) ? 4'b0111 : node17861;
																assign node17861 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node17866 = (inp[5]) ? node17868 : 4'b0111;
														assign node17868 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node17871 = (inp[5]) ? node17875 : node17872;
													assign node17872 = (inp[7]) ? 4'b0111 : 4'b0010;
													assign node17875 = (inp[7]) ? 4'b0011 : 4'b0111;
								assign node17878 = (inp[6]) ? node17954 : node17879;
									assign node17879 = (inp[10]) ? node17917 : node17880;
										assign node17880 = (inp[0]) ? node17896 : node17881;
											assign node17881 = (inp[7]) ? node17887 : node17882;
												assign node17882 = (inp[2]) ? 4'b0111 : node17883;
													assign node17883 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node17887 = (inp[2]) ? node17891 : node17888;
													assign node17888 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node17891 = (inp[4]) ? 4'b0111 : node17892;
														assign node17892 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node17896 = (inp[4]) ? node17908 : node17897;
												assign node17897 = (inp[9]) ? node17903 : node17898;
													assign node17898 = (inp[2]) ? 4'b0111 : node17899;
														assign node17899 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node17903 = (inp[2]) ? node17905 : 4'b0011;
														assign node17905 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node17908 = (inp[7]) ? 4'b0111 : node17909;
													assign node17909 = (inp[9]) ? 4'b0111 : node17910;
														assign node17910 = (inp[5]) ? 4'b0010 : node17911;
															assign node17911 = (inp[2]) ? 4'b0010 : 4'b0111;
										assign node17917 = (inp[5]) ? node17941 : node17918;
											assign node17918 = (inp[2]) ? node17930 : node17919;
												assign node17919 = (inp[1]) ? node17925 : node17920;
													assign node17920 = (inp[7]) ? 4'b0011 : node17921;
														assign node17921 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node17925 = (inp[7]) ? 4'b0110 : node17926;
														assign node17926 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node17930 = (inp[1]) ? node17936 : node17931;
													assign node17931 = (inp[4]) ? 4'b0110 : node17932;
														assign node17932 = (inp[0]) ? 4'b0011 : 4'b0110;
													assign node17936 = (inp[7]) ? node17938 : 4'b0011;
														assign node17938 = (inp[4]) ? 4'b0110 : 4'b0011;
											assign node17941 = (inp[2]) ? node17951 : node17942;
												assign node17942 = (inp[7]) ? node17946 : node17943;
													assign node17943 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node17946 = (inp[0]) ? 4'b0110 : node17947;
														assign node17947 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node17951 = (inp[7]) ? 4'b0010 : 4'b0110;
									assign node17954 = (inp[0]) ? node17998 : node17955;
										assign node17955 = (inp[4]) ? node17975 : node17956;
											assign node17956 = (inp[1]) ? node17962 : node17957;
												assign node17957 = (inp[7]) ? 4'b0010 : node17958;
													assign node17958 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node17962 = (inp[10]) ? node17964 : 4'b0110;
													assign node17964 = (inp[2]) ? node17966 : 4'b0110;
														assign node17966 = (inp[9]) ? node17972 : node17967;
															assign node17967 = (inp[7]) ? 4'b0110 : node17968;
																assign node17968 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node17972 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node17975 = (inp[1]) ? node17985 : node17976;
												assign node17976 = (inp[5]) ? node17982 : node17977;
													assign node17977 = (inp[7]) ? node17979 : 4'b0010;
														assign node17979 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node17982 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node17985 = (inp[10]) ? node17993 : node17986;
													assign node17986 = (inp[5]) ? node17990 : node17987;
														assign node17987 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node17990 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node17993 = (inp[9]) ? 4'b0110 : node17994;
														assign node17994 = (inp[7]) ? 4'b0110 : 4'b0011;
										assign node17998 = (inp[9]) ? node18018 : node17999;
											assign node17999 = (inp[5]) ? node18009 : node18000;
												assign node18000 = (inp[7]) ? 4'b0111 : node18001;
													assign node18001 = (inp[1]) ? node18003 : 4'b0010;
														assign node18003 = (inp[2]) ? 4'b0011 : node18004;
															assign node18004 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node18009 = (inp[7]) ? node18011 : 4'b0110;
													assign node18011 = (inp[1]) ? node18013 : 4'b0010;
														assign node18013 = (inp[10]) ? 4'b0010 : node18014;
															assign node18014 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node18018 = (inp[5]) ? node18032 : node18019;
												assign node18019 = (inp[7]) ? node18025 : node18020;
													assign node18020 = (inp[1]) ? node18022 : 4'b0010;
														assign node18022 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node18025 = (inp[10]) ? 4'b0110 : node18026;
														assign node18026 = (inp[4]) ? node18028 : 4'b0110;
															assign node18028 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node18032 = (inp[2]) ? node18034 : 4'b0011;
													assign node18034 = (inp[7]) ? 4'b0010 : 4'b0110;
						assign node18037 = (inp[5]) ? node18143 : node18038;
							assign node18038 = (inp[2]) ? node18086 : node18039;
								assign node18039 = (inp[6]) ? node18063 : node18040;
									assign node18040 = (inp[10]) ? node18052 : node18041;
										assign node18041 = (inp[7]) ? node18047 : node18042;
											assign node18042 = (inp[11]) ? node18044 : 4'b0000;
												assign node18044 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node18047 = (inp[11]) ? node18049 : 4'b0001;
												assign node18049 = (inp[4]) ? 4'b0000 : 4'b0001;
										assign node18052 = (inp[7]) ? node18058 : node18053;
											assign node18053 = (inp[13]) ? 4'b0001 : node18054;
												assign node18054 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node18058 = (inp[11]) ? node18060 : 4'b0000;
												assign node18060 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node18063 = (inp[1]) ? node18071 : node18064;
										assign node18064 = (inp[11]) ? node18068 : node18065;
											assign node18065 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node18068 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node18071 = (inp[10]) ? node18079 : node18072;
											assign node18072 = (inp[11]) ? node18076 : node18073;
												assign node18073 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node18076 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node18079 = (inp[7]) ? node18083 : node18080;
												assign node18080 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node18083 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node18086 = (inp[7]) ? node18112 : node18087;
									assign node18087 = (inp[10]) ? node18105 : node18088;
										assign node18088 = (inp[9]) ? node18098 : node18089;
											assign node18089 = (inp[6]) ? node18095 : node18090;
												assign node18090 = (inp[11]) ? 4'b0100 : node18091;
													assign node18091 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node18095 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node18098 = (inp[6]) ? 4'b0101 : node18099;
												assign node18099 = (inp[4]) ? node18101 : 4'b0100;
													assign node18101 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node18105 = (inp[11]) ? 4'b0101 : node18106;
											assign node18106 = (inp[4]) ? 4'b0100 : node18107;
												assign node18107 = (inp[6]) ? 4'b0100 : 4'b0101;
									assign node18112 = (inp[11]) ? node18138 : node18113;
										assign node18113 = (inp[6]) ? 4'b0101 : node18114;
											assign node18114 = (inp[13]) ? node18126 : node18115;
												assign node18115 = (inp[0]) ? node18117 : 4'b0101;
													assign node18117 = (inp[9]) ? node18119 : 4'b0100;
														assign node18119 = (inp[10]) ? node18123 : node18120;
															assign node18120 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node18123 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node18126 = (inp[9]) ? node18128 : 4'b0101;
													assign node18128 = (inp[1]) ? 4'b0101 : node18129;
														assign node18129 = (inp[4]) ? node18133 : node18130;
															assign node18130 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node18133 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node18138 = (inp[10]) ? 4'b0100 : node18139;
											assign node18139 = (inp[6]) ? 4'b0100 : 4'b0101;
							assign node18143 = (inp[2]) ? node18223 : node18144;
								assign node18144 = (inp[6]) ? node18160 : node18145;
									assign node18145 = (inp[0]) ? node18153 : node18146;
										assign node18146 = (inp[4]) ? node18150 : node18147;
											assign node18147 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node18150 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node18153 = (inp[10]) ? node18157 : node18154;
											assign node18154 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node18157 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node18160 = (inp[7]) ? node18192 : node18161;
										assign node18161 = (inp[0]) ? node18185 : node18162;
											assign node18162 = (inp[9]) ? node18168 : node18163;
												assign node18163 = (inp[1]) ? node18165 : 4'b0001;
													assign node18165 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node18168 = (inp[13]) ? node18178 : node18169;
													assign node18169 = (inp[10]) ? node18171 : 4'b0000;
														assign node18171 = (inp[1]) ? node18173 : 4'b0001;
															assign node18173 = (inp[11]) ? 4'b0000 : node18174;
																assign node18174 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node18178 = (inp[10]) ? 4'b0000 : node18179;
														assign node18179 = (inp[11]) ? 4'b0001 : node18180;
															assign node18180 = (inp[4]) ? 4'b0001 : 4'b0000;
											assign node18185 = (inp[4]) ? node18189 : node18186;
												assign node18186 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node18189 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node18192 = (inp[0]) ? node18210 : node18193;
											assign node18193 = (inp[9]) ? node18199 : node18194;
												assign node18194 = (inp[11]) ? node18196 : 4'b0001;
													assign node18196 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node18199 = (inp[1]) ? node18205 : node18200;
													assign node18200 = (inp[11]) ? node18202 : 4'b0000;
														assign node18202 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node18205 = (inp[4]) ? node18207 : 4'b0000;
														assign node18207 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node18210 = (inp[10]) ? node18216 : node18211;
												assign node18211 = (inp[11]) ? 4'b0000 : node18212;
													assign node18212 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node18216 = (inp[4]) ? node18220 : node18217;
													assign node18217 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node18220 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node18223 = (inp[11]) ? node18229 : node18224;
									assign node18224 = (inp[6]) ? 4'b0001 : node18225;
										assign node18225 = (inp[10]) ? 4'b0001 : 4'b0000;
									assign node18229 = (inp[6]) ? 4'b0000 : node18230;
										assign node18230 = (inp[10]) ? 4'b0000 : 4'b0001;
					assign node18234 = (inp[7]) ? node18480 : node18235;
						assign node18235 = (inp[15]) ? node18415 : node18236;
							assign node18236 = (inp[6]) ? node18376 : node18237;
								assign node18237 = (inp[2]) ? node18305 : node18238;
									assign node18238 = (inp[5]) ? node18254 : node18239;
										assign node18239 = (inp[4]) ? node18249 : node18240;
											assign node18240 = (inp[13]) ? node18244 : node18241;
												assign node18241 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node18244 = (inp[10]) ? 4'b0101 : node18245;
													assign node18245 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node18249 = (inp[1]) ? node18251 : 4'b0000;
												assign node18251 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node18254 = (inp[4]) ? node18278 : node18255;
											assign node18255 = (inp[9]) ? node18267 : node18256;
												assign node18256 = (inp[0]) ? node18258 : 4'b0001;
													assign node18258 = (inp[1]) ? 4'b0000 : node18259;
														assign node18259 = (inp[11]) ? node18263 : node18260;
															assign node18260 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node18263 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node18267 = (inp[0]) ? node18269 : 4'b0000;
													assign node18269 = (inp[11]) ? 4'b0000 : node18270;
														assign node18270 = (inp[1]) ? node18272 : 4'b0000;
															assign node18272 = (inp[10]) ? 4'b0001 : node18273;
																assign node18273 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node18278 = (inp[1]) ? node18286 : node18279;
												assign node18279 = (inp[13]) ? node18283 : node18280;
													assign node18280 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node18283 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node18286 = (inp[0]) ? node18296 : node18287;
													assign node18287 = (inp[11]) ? 4'b0000 : node18288;
														assign node18288 = (inp[9]) ? 4'b0001 : node18289;
															assign node18289 = (inp[13]) ? node18291 : 4'b0000;
																assign node18291 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node18296 = (inp[9]) ? node18298 : 4'b0001;
														assign node18298 = (inp[11]) ? node18302 : node18299;
															assign node18299 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node18302 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node18305 = (inp[5]) ? node18351 : node18306;
										assign node18306 = (inp[4]) ? node18330 : node18307;
											assign node18307 = (inp[9]) ? node18315 : node18308;
												assign node18308 = (inp[13]) ? 4'b0001 : node18309;
													assign node18309 = (inp[10]) ? 4'b0001 : node18310;
														assign node18310 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node18315 = (inp[13]) ? node18319 : node18316;
													assign node18316 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node18319 = (inp[0]) ? node18325 : node18320;
														assign node18320 = (inp[1]) ? node18322 : 4'b0000;
															assign node18322 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node18325 = (inp[1]) ? node18327 : 4'b0001;
															assign node18327 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node18330 = (inp[10]) ? node18338 : node18331;
												assign node18331 = (inp[13]) ? 4'b0100 : node18332;
													assign node18332 = (inp[11]) ? 4'b0101 : node18333;
														assign node18333 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node18338 = (inp[9]) ? node18340 : 4'b0101;
													assign node18340 = (inp[1]) ? 4'b0101 : node18341;
														assign node18341 = (inp[0]) ? node18347 : node18342;
															assign node18342 = (inp[11]) ? 4'b0101 : node18343;
																assign node18343 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node18347 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node18351 = (inp[13]) ? node18361 : node18352;
											assign node18352 = (inp[10]) ? node18358 : node18353;
												assign node18353 = (inp[11]) ? 4'b0100 : node18354;
													assign node18354 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node18358 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node18361 = (inp[4]) ? node18369 : node18362;
												assign node18362 = (inp[1]) ? 4'b0101 : node18363;
													assign node18363 = (inp[11]) ? 4'b0101 : node18364;
														assign node18364 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node18369 = (inp[9]) ? 4'b0101 : node18370;
													assign node18370 = (inp[10]) ? 4'b0100 : node18371;
														assign node18371 = (inp[0]) ? 4'b0101 : 4'b0100;
								assign node18376 = (inp[2]) ? node18400 : node18377;
									assign node18377 = (inp[13]) ? node18387 : node18378;
										assign node18378 = (inp[5]) ? node18384 : node18379;
											assign node18379 = (inp[4]) ? 4'b0100 : node18380;
												assign node18380 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node18384 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node18387 = (inp[1]) ? node18393 : node18388;
											assign node18388 = (inp[4]) ? node18390 : 4'b0101;
												assign node18390 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node18393 = (inp[5]) ? node18397 : node18394;
												assign node18394 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node18397 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node18400 = (inp[13]) ? node18408 : node18401;
										assign node18401 = (inp[5]) ? 4'b0101 : node18402;
											assign node18402 = (inp[1]) ? 4'b0100 : node18403;
												assign node18403 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node18408 = (inp[5]) ? 4'b0100 : node18409;
											assign node18409 = (inp[1]) ? 4'b0101 : node18410;
												assign node18410 = (inp[4]) ? 4'b0101 : 4'b0100;
							assign node18415 = (inp[6]) ? node18469 : node18416;
								assign node18416 = (inp[2]) ? node18454 : node18417;
									assign node18417 = (inp[10]) ? node18445 : node18418;
										assign node18418 = (inp[9]) ? node18432 : node18419;
											assign node18419 = (inp[13]) ? node18421 : 4'b0100;
												assign node18421 = (inp[1]) ? 4'b0100 : node18422;
													assign node18422 = (inp[0]) ? 4'b0100 : node18423;
														assign node18423 = (inp[11]) ? 4'b0101 : node18424;
															assign node18424 = (inp[4]) ? node18426 : 4'b0100;
																assign node18426 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node18432 = (inp[11]) ? node18438 : node18433;
												assign node18433 = (inp[4]) ? node18435 : 4'b0100;
													assign node18435 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node18438 = (inp[1]) ? node18440 : 4'b0101;
													assign node18440 = (inp[13]) ? 4'b0100 : node18441;
														assign node18441 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node18445 = (inp[5]) ? node18451 : node18446;
											assign node18446 = (inp[11]) ? node18448 : 4'b0101;
												assign node18448 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node18451 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node18454 = (inp[10]) ? node18462 : node18455;
										assign node18455 = (inp[5]) ? 4'b0001 : node18456;
											assign node18456 = (inp[11]) ? 4'b0000 : node18457;
												assign node18457 = (inp[4]) ? 4'b0000 : 4'b0001;
										assign node18462 = (inp[5]) ? 4'b0000 : node18463;
											assign node18463 = (inp[11]) ? 4'b0001 : node18464;
												assign node18464 = (inp[4]) ? 4'b0001 : 4'b0000;
								assign node18469 = (inp[5]) ? node18475 : node18470;
									assign node18470 = (inp[2]) ? 4'b0001 : node18471;
										assign node18471 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node18475 = (inp[2]) ? 4'b0000 : node18476;
										assign node18476 = (inp[4]) ? 4'b0000 : 4'b0001;
						assign node18480 = (inp[6]) ? node18664 : node18481;
							assign node18481 = (inp[2]) ? node18587 : node18482;
								assign node18482 = (inp[5]) ? node18532 : node18483;
									assign node18483 = (inp[4]) ? node18511 : node18484;
										assign node18484 = (inp[15]) ? node18504 : node18485;
											assign node18485 = (inp[11]) ? node18499 : node18486;
												assign node18486 = (inp[10]) ? node18494 : node18487;
													assign node18487 = (inp[0]) ? node18489 : 4'b0001;
														assign node18489 = (inp[13]) ? 4'b0000 : node18490;
															assign node18490 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node18494 = (inp[13]) ? 4'b0001 : node18495;
														assign node18495 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node18499 = (inp[10]) ? node18501 : 4'b0000;
													assign node18501 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node18504 = (inp[11]) ? node18508 : node18505;
												assign node18505 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node18508 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node18511 = (inp[10]) ? node18521 : node18512;
											assign node18512 = (inp[13]) ? 4'b0101 : node18513;
												assign node18513 = (inp[15]) ? 4'b0101 : node18514;
													assign node18514 = (inp[1]) ? 4'b0100 : node18515;
														assign node18515 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node18521 = (inp[15]) ? 4'b0100 : node18522;
												assign node18522 = (inp[9]) ? 4'b0101 : node18523;
													assign node18523 = (inp[0]) ? node18525 : 4'b0100;
														assign node18525 = (inp[1]) ? 4'b0101 : node18526;
															assign node18526 = (inp[13]) ? 4'b0101 : 4'b0100;
									assign node18532 = (inp[15]) ? node18564 : node18533;
										assign node18533 = (inp[4]) ? node18551 : node18534;
											assign node18534 = (inp[1]) ? node18536 : 4'b0100;
												assign node18536 = (inp[9]) ? node18542 : node18537;
													assign node18537 = (inp[11]) ? 4'b0100 : node18538;
														assign node18538 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node18542 = (inp[0]) ? node18548 : node18543;
														assign node18543 = (inp[13]) ? 4'b0100 : node18544;
															assign node18544 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node18548 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node18551 = (inp[13]) ? node18561 : node18552;
												assign node18552 = (inp[1]) ? 4'b0100 : node18553;
													assign node18553 = (inp[0]) ? 4'b0101 : node18554;
														assign node18554 = (inp[10]) ? 4'b0100 : node18555;
															assign node18555 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node18561 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node18564 = (inp[11]) ? node18572 : node18565;
											assign node18565 = (inp[10]) ? node18569 : node18566;
												assign node18566 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node18569 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node18572 = (inp[0]) ? node18580 : node18573;
												assign node18573 = (inp[10]) ? node18577 : node18574;
													assign node18574 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node18577 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node18580 = (inp[4]) ? node18584 : node18581;
													assign node18581 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node18584 = (inp[10]) ? 4'b0100 : 4'b0101;
								assign node18587 = (inp[10]) ? node18629 : node18588;
									assign node18588 = (inp[15]) ? node18622 : node18589;
										assign node18589 = (inp[4]) ? node18611 : node18590;
											assign node18590 = (inp[5]) ? node18604 : node18591;
												assign node18591 = (inp[9]) ? node18599 : node18592;
													assign node18592 = (inp[11]) ? node18594 : 4'b0101;
														assign node18594 = (inp[0]) ? node18596 : 4'b0100;
															assign node18596 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node18599 = (inp[13]) ? node18601 : 4'b0101;
														assign node18601 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node18604 = (inp[1]) ? node18608 : node18605;
													assign node18605 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node18608 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node18611 = (inp[13]) ? node18617 : node18612;
												assign node18612 = (inp[0]) ? node18614 : 4'b0000;
													assign node18614 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node18617 = (inp[11]) ? 4'b0001 : node18618;
													assign node18618 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node18622 = (inp[11]) ? 4'b0001 : node18623;
											assign node18623 = (inp[5]) ? 4'b0001 : node18624;
												assign node18624 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node18629 = (inp[15]) ? node18657 : node18630;
										assign node18630 = (inp[4]) ? node18646 : node18631;
											assign node18631 = (inp[5]) ? node18641 : node18632;
												assign node18632 = (inp[13]) ? node18636 : node18633;
													assign node18633 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node18636 = (inp[1]) ? node18638 : 4'b0101;
														assign node18638 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node18641 = (inp[9]) ? 4'b0000 : node18642;
													assign node18642 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node18646 = (inp[13]) ? node18652 : node18647;
												assign node18647 = (inp[1]) ? 4'b0001 : node18648;
													assign node18648 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node18652 = (inp[11]) ? 4'b0000 : node18653;
													assign node18653 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node18657 = (inp[11]) ? 4'b0000 : node18658;
											assign node18658 = (inp[5]) ? 4'b0000 : node18659;
												assign node18659 = (inp[4]) ? 4'b0000 : 4'b0001;
							assign node18664 = (inp[13]) ? node18684 : node18665;
								assign node18665 = (inp[15]) ? node18679 : node18666;
									assign node18666 = (inp[4]) ? 4'b0001 : node18667;
										assign node18667 = (inp[2]) ? node18673 : node18668;
											assign node18668 = (inp[1]) ? 4'b0000 : node18669;
												assign node18669 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node18673 = (inp[1]) ? 4'b0001 : node18674;
												assign node18674 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node18679 = (inp[4]) ? 4'b0000 : node18680;
										assign node18680 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node18684 = (inp[4]) ? 4'b0000 : node18685;
									assign node18685 = (inp[2]) ? node18695 : node18686;
										assign node18686 = (inp[10]) ? 4'b0001 : node18687;
											assign node18687 = (inp[1]) ? 4'b0001 : node18688;
												assign node18688 = (inp[15]) ? 4'b0001 : node18689;
													assign node18689 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node18695 = (inp[1]) ? 4'b0000 : node18696;
											assign node18696 = (inp[15]) ? 4'b0000 : node18697;
												assign node18697 = (inp[5]) ? 4'b0000 : 4'b0001;

endmodule