module dtc_split25_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node380;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node523;

	assign outp = (inp[3]) ? node386 : node1;
		assign node1 = (inp[9]) ? node165 : node2;
			assign node2 = (inp[1]) ? node68 : node3;
				assign node3 = (inp[4]) ? node27 : node4;
					assign node4 = (inp[6]) ? node14 : node5;
						assign node5 = (inp[0]) ? node11 : node6;
							assign node6 = (inp[5]) ? node8 : 3'b001;
								assign node8 = (inp[7]) ? 3'b001 : 3'b000;
							assign node11 = (inp[5]) ? 3'b001 : 3'b000;
						assign node14 = (inp[5]) ? node22 : node15;
							assign node15 = (inp[0]) ? node17 : 3'b000;
								assign node17 = (inp[7]) ? node19 : 3'b000;
									assign node19 = (inp[11]) ? 3'b000 : 3'b001;
							assign node22 = (inp[0]) ? 3'b000 : node23;
								assign node23 = (inp[8]) ? 3'b000 : 3'b001;
					assign node27 = (inp[0]) ? node43 : node28;
						assign node28 = (inp[6]) ? node30 : 3'b000;
							assign node30 = (inp[10]) ? node36 : node31;
								assign node31 = (inp[2]) ? node33 : 3'b000;
									assign node33 = (inp[5]) ? 3'b001 : 3'b000;
								assign node36 = (inp[7]) ? 3'b001 : node37;
									assign node37 = (inp[5]) ? node39 : 3'b001;
										assign node39 = (inp[8]) ? 3'b000 : 3'b000;
						assign node43 = (inp[2]) ? node63 : node44;
							assign node44 = (inp[7]) ? node56 : node45;
								assign node45 = (inp[8]) ? node51 : node46;
									assign node46 = (inp[6]) ? node48 : 3'b000;
										assign node48 = (inp[11]) ? 3'b001 : 3'b000;
									assign node51 = (inp[6]) ? node53 : 3'b001;
										assign node53 = (inp[5]) ? 3'b001 : 3'b000;
								assign node56 = (inp[10]) ? 3'b001 : node57;
									assign node57 = (inp[6]) ? node59 : 3'b001;
										assign node59 = (inp[5]) ? 3'b001 : 3'b000;
							assign node63 = (inp[5]) ? 3'b000 : node64;
								assign node64 = (inp[6]) ? 3'b000 : 3'b001;
				assign node68 = (inp[7]) ? node126 : node69;
					assign node69 = (inp[2]) ? node97 : node70;
						assign node70 = (inp[0]) ? node82 : node71;
							assign node71 = (inp[4]) ? 3'b000 : node72;
								assign node72 = (inp[6]) ? node76 : node73;
									assign node73 = (inp[5]) ? 3'b001 : 3'b000;
									assign node76 = (inp[5]) ? 3'b000 : node77;
										assign node77 = (inp[10]) ? 3'b000 : 3'b001;
							assign node82 = (inp[5]) ? node92 : node83;
								assign node83 = (inp[11]) ? node87 : node84;
									assign node84 = (inp[8]) ? 3'b001 : 3'b000;
									assign node87 = (inp[8]) ? 3'b000 : node88;
										assign node88 = (inp[4]) ? 3'b001 : 3'b000;
								assign node92 = (inp[4]) ? 3'b001 : node93;
									assign node93 = (inp[6]) ? 3'b000 : 3'b001;
						assign node97 = (inp[10]) ? node109 : node98;
							assign node98 = (inp[8]) ? 3'b001 : node99;
								assign node99 = (inp[5]) ? 3'b000 : node100;
									assign node100 = (inp[11]) ? node104 : node101;
										assign node101 = (inp[4]) ? 3'b000 : 3'b001;
										assign node104 = (inp[6]) ? 3'b001 : 3'b000;
							assign node109 = (inp[5]) ? node121 : node110;
								assign node110 = (inp[11]) ? node116 : node111;
									assign node111 = (inp[8]) ? 3'b000 : node112;
										assign node112 = (inp[6]) ? 3'b000 : 3'b000;
									assign node116 = (inp[0]) ? 3'b000 : node117;
										assign node117 = (inp[8]) ? 3'b000 : 3'b001;
								assign node121 = (inp[4]) ? node123 : 3'b001;
									assign node123 = (inp[0]) ? 3'b001 : 3'b000;
					assign node126 = (inp[6]) ? node150 : node127;
						assign node127 = (inp[4]) ? node139 : node128;
							assign node128 = (inp[8]) ? 3'b001 : node129;
								assign node129 = (inp[0]) ? 3'b000 : node130;
									assign node130 = (inp[11]) ? node134 : node131;
										assign node131 = (inp[5]) ? 3'b001 : 3'b000;
										assign node134 = (inp[2]) ? 3'b000 : 3'b001;
							assign node139 = (inp[0]) ? 3'b001 : node140;
								assign node140 = (inp[5]) ? node144 : node141;
									assign node141 = (inp[10]) ? 3'b001 : 3'b000;
									assign node144 = (inp[10]) ? node146 : 3'b001;
										assign node146 = (inp[11]) ? 3'b000 : 3'b001;
						assign node150 = (inp[0]) ? node160 : node151;
							assign node151 = (inp[2]) ? node153 : 3'b001;
								assign node153 = (inp[8]) ? 3'b000 : node154;
									assign node154 = (inp[10]) ? node156 : 3'b001;
										assign node156 = (inp[11]) ? 3'b000 : 3'b001;
							assign node160 = (inp[4]) ? 3'b000 : node161;
								assign node161 = (inp[8]) ? 3'b001 : 3'b000;
			assign node165 = (inp[4]) ? node271 : node166;
				assign node166 = (inp[6]) ? node220 : node167;
					assign node167 = (inp[0]) ? node193 : node168;
						assign node168 = (inp[5]) ? node180 : node169;
							assign node169 = (inp[1]) ? node173 : node170;
								assign node170 = (inp[7]) ? 3'b110 : 3'b010;
								assign node173 = (inp[7]) ? node177 : node174;
									assign node174 = (inp[10]) ? 3'b110 : 3'b101;
									assign node177 = (inp[2]) ? 3'b001 : 3'b010;
							assign node180 = (inp[1]) ? node184 : node181;
								assign node181 = (inp[7]) ? 3'b010 : 3'b100;
								assign node184 = (inp[11]) ? node190 : node185;
									assign node185 = (inp[10]) ? node187 : 3'b001;
										assign node187 = (inp[2]) ? 3'b101 : 3'b000;
									assign node190 = (inp[7]) ? 3'b110 : 3'b010;
						assign node193 = (inp[5]) ? node211 : node194;
							assign node194 = (inp[8]) ? node206 : node195;
								assign node195 = (inp[1]) ? node201 : node196;
									assign node196 = (inp[2]) ? 3'b001 : node197;
										assign node197 = (inp[11]) ? 3'b110 : 3'b010;
									assign node201 = (inp[7]) ? 3'b101 : node202;
										assign node202 = (inp[11]) ? 3'b001 : 3'b101;
								assign node206 = (inp[1]) ? node208 : 3'b001;
									assign node208 = (inp[7]) ? 3'b011 : 3'b000;
							assign node211 = (inp[1]) ? node213 : 3'b110;
								assign node213 = (inp[7]) ? node215 : 3'b111;
									assign node215 = (inp[2]) ? 3'b101 : node216;
										assign node216 = (inp[11]) ? 3'b001 : 3'b101;
					assign node220 = (inp[1]) ? node246 : node221;
						assign node221 = (inp[5]) ? node239 : node222;
							assign node222 = (inp[7]) ? node228 : node223;
								assign node223 = (inp[0]) ? 3'b101 : node224;
									assign node224 = (inp[10]) ? 3'b001 : 3'b101;
								assign node228 = (inp[10]) ? node234 : node229;
									assign node229 = (inp[0]) ? node231 : 3'b001;
										assign node231 = (inp[8]) ? 3'b101 : 3'b001;
									assign node234 = (inp[0]) ? node236 : 3'b101;
										assign node236 = (inp[8]) ? 3'b111 : 3'b011;
							assign node239 = (inp[0]) ? 3'b101 : node240;
								assign node240 = (inp[7]) ? node242 : 3'b110;
									assign node242 = (inp[10]) ? 3'b001 : 3'b010;
						assign node246 = (inp[0]) ? node260 : node247;
							assign node247 = (inp[2]) ? node251 : node248;
								assign node248 = (inp[7]) ? 3'b011 : 3'b001;
								assign node251 = (inp[5]) ? node257 : node252;
									assign node252 = (inp[7]) ? 3'b001 : node253;
										assign node253 = (inp[11]) ? 3'b101 : 3'b001;
									assign node257 = (inp[7]) ? 3'b101 : 3'b001;
							assign node260 = (inp[5]) ? node268 : node261;
								assign node261 = (inp[7]) ? 3'b111 : node262;
									assign node262 = (inp[8]) ? node264 : 3'b011;
										assign node264 = (inp[10]) ? 3'b111 : 3'b011;
								assign node268 = (inp[8]) ? 3'b011 : 3'b001;
				assign node271 = (inp[0]) ? node331 : node272;
					assign node272 = (inp[6]) ? node304 : node273;
						assign node273 = (inp[1]) ? node285 : node274;
							assign node274 = (inp[5]) ? node278 : node275;
								assign node275 = (inp[2]) ? 3'b100 : 3'b000;
								assign node278 = (inp[7]) ? 3'b000 : node279;
									assign node279 = (inp[2]) ? node281 : 3'b000;
										assign node281 = (inp[8]) ? 3'b000 : 3'b100;
							assign node285 = (inp[8]) ? node293 : node286;
								assign node286 = (inp[5]) ? 3'b000 : node287;
									assign node287 = (inp[11]) ? 3'b010 : node288;
										assign node288 = (inp[7]) ? 3'b000 : 3'b000;
								assign node293 = (inp[2]) ? node299 : node294;
									assign node294 = (inp[10]) ? node296 : 3'b000;
										assign node296 = (inp[11]) ? 3'b100 : 3'b100;
									assign node299 = (inp[5]) ? 3'b000 : node300;
										assign node300 = (inp[7]) ? 3'b010 : 3'b110;
						assign node304 = (inp[7]) ? node318 : node305;
							assign node305 = (inp[5]) ? node311 : node306;
								assign node306 = (inp[8]) ? 3'b010 : node307;
									assign node307 = (inp[1]) ? 3'b110 : 3'b100;
								assign node311 = (inp[1]) ? 3'b100 : node312;
									assign node312 = (inp[11]) ? 3'b100 : node313;
										assign node313 = (inp[8]) ? 3'b010 : 3'b100;
							assign node318 = (inp[1]) ? node324 : node319;
								assign node319 = (inp[10]) ? node321 : 3'b000;
									assign node321 = (inp[8]) ? 3'b110 : 3'b100;
								assign node324 = (inp[2]) ? node328 : node325;
									assign node325 = (inp[5]) ? 3'b010 : 3'b110;
									assign node328 = (inp[10]) ? 3'b101 : 3'b110;
					assign node331 = (inp[6]) ? node371 : node332;
						assign node332 = (inp[7]) ? node350 : node333;
							assign node333 = (inp[2]) ? node341 : node334;
								assign node334 = (inp[10]) ? node336 : 3'b100;
									assign node336 = (inp[11]) ? 3'b010 : node337;
										assign node337 = (inp[1]) ? 3'b100 : 3'b000;
								assign node341 = (inp[8]) ? node343 : 3'b010;
									assign node343 = (inp[10]) ? node347 : node344;
										assign node344 = (inp[11]) ? 3'b100 : 3'b000;
										assign node347 = (inp[5]) ? 3'b010 : 3'b000;
							assign node350 = (inp[10]) ? node364 : node351;
								assign node351 = (inp[8]) ? node357 : node352;
									assign node352 = (inp[5]) ? 3'b010 : node353;
										assign node353 = (inp[1]) ? 3'b110 : 3'b010;
									assign node357 = (inp[11]) ? node361 : node358;
										assign node358 = (inp[5]) ? 3'b100 : 3'b110;
										assign node361 = (inp[1]) ? 3'b010 : 3'b010;
								assign node364 = (inp[2]) ? node366 : 3'b010;
									assign node366 = (inp[11]) ? node368 : 3'b010;
										assign node368 = (inp[5]) ? 3'b100 : 3'b010;
						assign node371 = (inp[5]) ? node377 : node372;
							assign node372 = (inp[1]) ? node374 : 3'b001;
								assign node374 = (inp[7]) ? 3'b101 : 3'b001;
							assign node377 = (inp[1]) ? node383 : node378;
								assign node378 = (inp[10]) ? node380 : 3'b010;
									assign node380 = (inp[7]) ? 3'b110 : 3'b010;
								assign node383 = (inp[7]) ? 3'b001 : 3'b110;
		assign node386 = (inp[6]) ? node408 : node387;
			assign node387 = (inp[0]) ? node389 : 3'b000;
				assign node389 = (inp[1]) ? node391 : 3'b000;
					assign node391 = (inp[9]) ? node393 : 3'b000;
						assign node393 = (inp[4]) ? 3'b000 : node394;
							assign node394 = (inp[5]) ? node400 : node395;
								assign node395 = (inp[7]) ? 3'b100 : node396;
									assign node396 = (inp[8]) ? 3'b100 : 3'b000;
								assign node400 = (inp[7]) ? 3'b000 : node401;
									assign node401 = (inp[11]) ? 3'b000 : node402;
										assign node402 = (inp[8]) ? 3'b100 : 3'b000;
			assign node408 = (inp[9]) ? node478 : node409;
				assign node409 = (inp[4]) ? node425 : node410;
					assign node410 = (inp[0]) ? node418 : node411;
						assign node411 = (inp[7]) ? node413 : 3'b010;
							assign node413 = (inp[1]) ? node415 : 3'b010;
								assign node415 = (inp[2]) ? 3'b011 : 3'b010;
						assign node418 = (inp[5]) ? node420 : 3'b011;
							assign node420 = (inp[1]) ? node422 : 3'b010;
								assign node422 = (inp[7]) ? 3'b011 : 3'b010;
					assign node425 = (inp[0]) ? node445 : node426;
						assign node426 = (inp[5]) ? node432 : node427;
							assign node427 = (inp[10]) ? 3'b000 : node428;
								assign node428 = (inp[7]) ? 3'b010 : 3'b000;
							assign node432 = (inp[1]) ? node438 : node433;
								assign node433 = (inp[11]) ? node435 : 3'b000;
									assign node435 = (inp[8]) ? 3'b100 : 3'b000;
								assign node438 = (inp[11]) ? 3'b100 : node439;
									assign node439 = (inp[8]) ? 3'b100 : node440;
										assign node440 = (inp[7]) ? 3'b000 : 3'b000;
						assign node445 = (inp[7]) ? node455 : node446;
							assign node446 = (inp[10]) ? node450 : node447;
								assign node447 = (inp[11]) ? 3'b010 : 3'b110;
								assign node450 = (inp[1]) ? node452 : 3'b100;
									assign node452 = (inp[5]) ? 3'b100 : 3'b010;
							assign node455 = (inp[5]) ? node467 : node456;
								assign node456 = (inp[1]) ? node462 : node457;
									assign node457 = (inp[8]) ? node459 : 3'b010;
										assign node459 = (inp[10]) ? 3'b010 : 3'b110;
									assign node462 = (inp[10]) ? 3'b110 : node463;
										assign node463 = (inp[8]) ? 3'b101 : 3'b110;
								assign node467 = (inp[2]) ? node473 : node468;
									assign node468 = (inp[1]) ? 3'b010 : node469;
										assign node469 = (inp[11]) ? 3'b100 : 3'b010;
									assign node473 = (inp[10]) ? node475 : 3'b110;
										assign node475 = (inp[11]) ? 3'b010 : 3'b010;
				assign node478 = (inp[4]) ? node508 : node479;
					assign node479 = (inp[5]) ? node497 : node480;
						assign node480 = (inp[0]) ? node492 : node481;
							assign node481 = (inp[8]) ? node483 : 3'b000;
								assign node483 = (inp[7]) ? node487 : node484;
									assign node484 = (inp[2]) ? 3'b100 : 3'b000;
									assign node487 = (inp[1]) ? node489 : 3'b100;
										assign node489 = (inp[2]) ? 3'b010 : 3'b100;
							assign node492 = (inp[1]) ? node494 : 3'b010;
								assign node494 = (inp[7]) ? 3'b110 : 3'b010;
						assign node497 = (inp[0]) ? node503 : node498;
							assign node498 = (inp[11]) ? node500 : 3'b000;
								assign node500 = (inp[1]) ? 3'b110 : 3'b000;
							assign node503 = (inp[7]) ? node505 : 3'b100;
								assign node505 = (inp[1]) ? 3'b010 : 3'b100;
					assign node508 = (inp[0]) ? node510 : 3'b000;
						assign node510 = (inp[5]) ? 3'b000 : node511;
							assign node511 = (inp[2]) ? node521 : node512;
								assign node512 = (inp[1]) ? node514 : 3'b000;
									assign node514 = (inp[8]) ? node518 : node515;
										assign node515 = (inp[7]) ? 3'b100 : 3'b000;
										assign node518 = (inp[11]) ? 3'b000 : 3'b100;
								assign node521 = (inp[7]) ? node523 : 3'b000;
									assign node523 = (inp[10]) ? 3'b000 : 3'b100;

endmodule