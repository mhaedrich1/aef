module dtc_split66_bm9 (
	input  wire [8-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node9;
	wire [8-1:0] node12;
	wire [8-1:0] node15;
	wire [8-1:0] node16;
	wire [8-1:0] node17;
	wire [8-1:0] node20;
	wire [8-1:0] node23;
	wire [8-1:0] node24;
	wire [8-1:0] node27;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node32;
	wire [8-1:0] node33;
	wire [8-1:0] node36;
	wire [8-1:0] node39;
	wire [8-1:0] node41;
	wire [8-1:0] node44;
	wire [8-1:0] node45;
	wire [8-1:0] node47;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node54;
	wire [8-1:0] node57;
	wire [8-1:0] node58;
	wire [8-1:0] node59;
	wire [8-1:0] node60;
	wire [8-1:0] node61;
	wire [8-1:0] node64;
	wire [8-1:0] node67;
	wire [8-1:0] node68;
	wire [8-1:0] node71;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node76;
	wire [8-1:0] node79;
	wire [8-1:0] node82;
	wire [8-1:0] node84;
	wire [8-1:0] node87;
	wire [8-1:0] node88;
	wire [8-1:0] node89;
	wire [8-1:0] node90;
	wire [8-1:0] node93;
	wire [8-1:0] node96;
	wire [8-1:0] node97;
	wire [8-1:0] node101;
	wire [8-1:0] node102;
	wire [8-1:0] node103;
	wire [8-1:0] node106;
	wire [8-1:0] node109;
	wire [8-1:0] node110;
	wire [8-1:0] node113;
	wire [8-1:0] node116;
	wire [8-1:0] node117;
	wire [8-1:0] node118;
	wire [8-1:0] node119;
	wire [8-1:0] node120;
	wire [8-1:0] node121;
	wire [8-1:0] node125;
	wire [8-1:0] node127;
	wire [8-1:0] node130;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node135;
	wire [8-1:0] node138;
	wire [8-1:0] node139;
	wire [8-1:0] node142;
	wire [8-1:0] node145;
	wire [8-1:0] node146;
	wire [8-1:0] node147;
	wire [8-1:0] node149;
	wire [8-1:0] node152;
	wire [8-1:0] node153;
	wire [8-1:0] node156;
	wire [8-1:0] node159;
	wire [8-1:0] node160;
	wire [8-1:0] node161;
	wire [8-1:0] node164;
	wire [8-1:0] node167;
	wire [8-1:0] node168;
	wire [8-1:0] node171;
	wire [8-1:0] node174;
	wire [8-1:0] node175;
	wire [8-1:0] node176;
	wire [8-1:0] node177;
	wire [8-1:0] node179;
	wire [8-1:0] node182;
	wire [8-1:0] node183;
	wire [8-1:0] node186;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node191;
	wire [8-1:0] node194;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node206;
	wire [8-1:0] node207;
	wire [8-1:0] node210;
	wire [8-1:0] node213;
	wire [8-1:0] node214;
	wire [8-1:0] node217;
	wire [8-1:0] node220;
	wire [8-1:0] node221;
	wire [8-1:0] node222;
	wire [8-1:0] node225;
	wire [8-1:0] node228;
	wire [8-1:0] node229;
	wire [8-1:0] node232;

	assign outp = (inp[3]) ? node116 : node1;
		assign node1 = (inp[5]) ? node57 : node2;
			assign node2 = (inp[2]) ? node30 : node3;
				assign node3 = (inp[0]) ? node15 : node4;
					assign node4 = (inp[4]) ? node12 : node5;
						assign node5 = (inp[1]) ? node9 : node6;
							assign node6 = (inp[7]) ? 8'b00100000 : 8'b10000100;
							assign node9 = (inp[7]) ? 8'b00011110 : 8'b00100011;
						assign node12 = (inp[1]) ? 8'b01100011 : 8'b11101110;
					assign node15 = (inp[1]) ? node23 : node16;
						assign node16 = (inp[7]) ? node20 : node17;
							assign node17 = (inp[6]) ? 8'b11001000 : 8'b01000000;
							assign node20 = (inp[4]) ? 8'b01010011 : 8'b00000000;
						assign node23 = (inp[6]) ? node27 : node24;
							assign node24 = (inp[4]) ? 8'b01001101 : 8'b10000000;
							assign node27 = (inp[7]) ? 8'b00010100 : 8'b10010001;
				assign node30 = (inp[6]) ? node44 : node31;
					assign node31 = (inp[1]) ? node39 : node32;
						assign node32 = (inp[4]) ? node36 : node33;
							assign node33 = (inp[7]) ? 8'b00111001 : 8'b00100001;
							assign node36 = (inp[0]) ? 8'b01011011 : 8'b00010000;
						assign node39 = (inp[4]) ? node41 : 8'b01110110;
							assign node41 = (inp[7]) ? 8'b11111111 : 8'b10100001;
					assign node44 = (inp[4]) ? node50 : node45;
						assign node45 = (inp[1]) ? node47 : 8'b11100101;
							assign node47 = (inp[7]) ? 8'b00111000 : 8'b10101110;
						assign node50 = (inp[0]) ? node54 : node51;
							assign node51 = (inp[7]) ? 8'b11100111 : 8'b10100101;
							assign node54 = (inp[7]) ? 8'b10111111 : 8'b10110111;
			assign node57 = (inp[7]) ? node87 : node58;
				assign node58 = (inp[4]) ? node74 : node59;
					assign node59 = (inp[2]) ? node67 : node60;
						assign node60 = (inp[1]) ? node64 : node61;
							assign node61 = (inp[0]) ? 8'b11110101 : 8'b10010110;
							assign node64 = (inp[6]) ? 8'b11011010 : 8'b10010010;
						assign node67 = (inp[1]) ? node71 : node68;
							assign node68 = (inp[6]) ? 8'b10100111 : 8'b11111001;
							assign node71 = (inp[0]) ? 8'b01110001 : 8'b00010111;
					assign node74 = (inp[2]) ? node82 : node75;
						assign node75 = (inp[0]) ? node79 : node76;
							assign node76 = (inp[6]) ? 8'b01101010 : 8'b01010010;
							assign node79 = (inp[6]) ? 8'b00110100 : 8'b01100110;
						assign node82 = (inp[1]) ? node84 : 8'b10001010;
							assign node84 = (inp[6]) ? 8'b11000111 : 8'b01000000;
				assign node87 = (inp[2]) ? node101 : node88;
					assign node88 = (inp[1]) ? node96 : node89;
						assign node89 = (inp[6]) ? node93 : node90;
							assign node90 = (inp[0]) ? 8'b10111101 : 8'b00100000;
							assign node93 = (inp[4]) ? 8'b00001011 : 8'b10000011;
						assign node96 = (inp[4]) ? 8'b00010000 : node97;
							assign node97 = (inp[0]) ? 8'b01101110 : 8'b00000001;
					assign node101 = (inp[1]) ? node109 : node102;
						assign node102 = (inp[0]) ? node106 : node103;
							assign node103 = (inp[6]) ? 8'b00000100 : 8'b01011110;
							assign node106 = (inp[4]) ? 8'b00110110 : 8'b01100010;
						assign node109 = (inp[0]) ? node113 : node110;
							assign node110 = (inp[6]) ? 8'b01000001 : 8'b00101100;
							assign node113 = (inp[6]) ? 8'b00101100 : 8'b10000000;
		assign node116 = (inp[7]) ? node174 : node117;
			assign node117 = (inp[4]) ? node145 : node118;
				assign node118 = (inp[5]) ? node130 : node119;
					assign node119 = (inp[0]) ? node125 : node120;
						assign node120 = (inp[1]) ? 8'b00101101 : node121;
							assign node121 = (inp[2]) ? 8'b11111010 : 8'b10000010;
						assign node125 = (inp[1]) ? node127 : 8'b11001101;
							assign node127 = (inp[2]) ? 8'b11001111 : 8'b01011111;
					assign node130 = (inp[6]) ? node138 : node131;
						assign node131 = (inp[2]) ? node135 : node132;
							assign node132 = (inp[0]) ? 8'b10000000 : 8'b00110000;
							assign node135 = (inp[1]) ? 8'b01111001 : 8'b00110011;
						assign node138 = (inp[0]) ? node142 : node139;
							assign node139 = (inp[2]) ? 8'b01001000 : 8'b11000101;
							assign node142 = (inp[1]) ? 8'b00110010 : 8'b00100101;
				assign node145 = (inp[0]) ? node159 : node146;
					assign node146 = (inp[2]) ? node152 : node147;
						assign node147 = (inp[6]) ? node149 : 8'b10110010;
							assign node149 = (inp[5]) ? 8'b00000111 : 8'b00010100;
						assign node152 = (inp[1]) ? node156 : node153;
							assign node153 = (inp[6]) ? 8'b11100000 : 8'b10001100;
							assign node156 = (inp[5]) ? 8'b10001001 : 8'b01000110;
					assign node159 = (inp[1]) ? node167 : node160;
						assign node160 = (inp[6]) ? node164 : node161;
							assign node161 = (inp[2]) ? 8'b00100110 : 8'b00000000;
							assign node164 = (inp[2]) ? 8'b00010110 : 8'b00111101;
						assign node167 = (inp[2]) ? node171 : node168;
							assign node168 = (inp[5]) ? 8'b01001100 : 8'b01000011;
							assign node171 = (inp[6]) ? 8'b10010000 : 8'b00011100;
			assign node174 = (inp[5]) ? node204 : node175;
				assign node175 = (inp[2]) ? node189 : node176;
					assign node176 = (inp[0]) ? node182 : node177;
						assign node177 = (inp[6]) ? node179 : 8'b01111101;
							assign node179 = (inp[4]) ? 8'b01110101 : 8'b01000001;
						assign node182 = (inp[6]) ? node186 : node183;
							assign node183 = (inp[1]) ? 8'b11000000 : 8'b11001011;
							assign node186 = (inp[4]) ? 8'b01100101 : 8'b01000010;
					assign node189 = (inp[6]) ? node197 : node190;
						assign node190 = (inp[0]) ? node194 : node191;
							assign node191 = (inp[4]) ? 8'b00100011 : 8'b00100111;
							assign node194 = (inp[4]) ? 8'b00000001 : 8'b01101001;
						assign node197 = (inp[4]) ? node201 : node198;
							assign node198 = (inp[1]) ? 8'b00000001 : 8'b10100000;
							assign node201 = (inp[0]) ? 8'b00000000 : 8'b00010000;
				assign node204 = (inp[1]) ? node220 : node205;
					assign node205 = (inp[2]) ? node213 : node206;
						assign node206 = (inp[6]) ? node210 : node207;
							assign node207 = (inp[4]) ? 8'b11010101 : 8'b00011000;
							assign node210 = (inp[0]) ? 8'b00001001 : 8'b00010011;
						assign node213 = (inp[0]) ? node217 : node214;
							assign node214 = (inp[6]) ? 8'b10001101 : 8'b00001000;
							assign node217 = (inp[4]) ? 8'b01001110 : 8'b00101011;
					assign node220 = (inp[4]) ? node228 : node221;
						assign node221 = (inp[2]) ? node225 : node222;
							assign node222 = (inp[0]) ? 8'b00100001 : 8'b01000110;
							assign node225 = (inp[6]) ? 8'b11101001 : 8'b11000101;
						assign node228 = (inp[6]) ? node232 : node229;
							assign node229 = (inp[2]) ? 8'b10001000 : 8'b00101001;
							assign node232 = (inp[2]) ? 8'b01001000 : 8'b11100010;

endmodule