module dtc_split5_bm51 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node6;
	wire [2-1:0] node9;
	wire [2-1:0] node10;
	wire [2-1:0] node11;
	wire [2-1:0] node13;
	wire [2-1:0] node16;
	wire [2-1:0] node17;
	wire [2-1:0] node20;
	wire [2-1:0] node24;
	wire [2-1:0] node25;
	wire [2-1:0] node26;
	wire [2-1:0] node28;
	wire [2-1:0] node30;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node38;
	wire [2-1:0] node39;
	wire [2-1:0] node42;
	wire [2-1:0] node45;
	wire [2-1:0] node46;
	wire [2-1:0] node47;
	wire [2-1:0] node48;
	wire [2-1:0] node49;
	wire [2-1:0] node53;
	wire [2-1:0] node54;
	wire [2-1:0] node57;
	wire [2-1:0] node59;
	wire [2-1:0] node62;
	wire [2-1:0] node63;
	wire [2-1:0] node66;
	wire [2-1:0] node69;
	wire [2-1:0] node70;
	wire [2-1:0] node71;
	wire [2-1:0] node74;
	wire [2-1:0] node77;
	wire [2-1:0] node80;
	wire [2-1:0] node81;
	wire [2-1:0] node82;
	wire [2-1:0] node83;
	wire [2-1:0] node84;
	wire [2-1:0] node86;
	wire [2-1:0] node88;
	wire [2-1:0] node92;
	wire [2-1:0] node93;
	wire [2-1:0] node96;
	wire [2-1:0] node99;
	wire [2-1:0] node100;
	wire [2-1:0] node103;
	wire [2-1:0] node104;
	wire [2-1:0] node108;
	wire [2-1:0] node109;
	wire [2-1:0] node110;
	wire [2-1:0] node111;
	wire [2-1:0] node113;
	wire [2-1:0] node117;
	wire [2-1:0] node118;
	wire [2-1:0] node122;
	wire [2-1:0] node123;

	assign outp = (inp[7]) ? node80 : node1;
		assign node1 = (inp[0]) ? node45 : node2;
			assign node2 = (inp[6]) ? node24 : node3;
				assign node3 = (inp[2]) ? node9 : node4;
					assign node4 = (inp[4]) ? node6 : 2'b01;
						assign node6 = (inp[5]) ? 2'b00 : 2'b01;
					assign node9 = (inp[5]) ? 2'b10 : node10;
						assign node10 = (inp[3]) ? node16 : node11;
							assign node11 = (inp[4]) ? node13 : 2'b10;
								assign node13 = (inp[1]) ? 2'b10 : 2'b11;
							assign node16 = (inp[1]) ? node20 : node17;
								assign node17 = (inp[4]) ? 2'b11 : 2'b10;
								assign node20 = (inp[4]) ? 2'b10 : 2'b11;
				assign node24 = (inp[2]) ? node38 : node25;
					assign node25 = (inp[4]) ? node33 : node26;
						assign node26 = (inp[3]) ? node28 : 2'b10;
							assign node28 = (inp[5]) ? node30 : 2'b11;
								assign node30 = (inp[1]) ? 2'b11 : 2'b10;
						assign node33 = (inp[5]) ? 2'b10 : node34;
							assign node34 = (inp[3]) ? 2'b10 : 2'b11;
					assign node38 = (inp[1]) ? node42 : node39;
						assign node39 = (inp[4]) ? 2'b11 : 2'b10;
						assign node42 = (inp[5]) ? 2'b11 : 2'b10;
			assign node45 = (inp[2]) ? node69 : node46;
				assign node46 = (inp[6]) ? node62 : node47;
					assign node47 = (inp[1]) ? node53 : node48;
						assign node48 = (inp[4]) ? 2'b11 : node49;
							assign node49 = (inp[5]) ? 2'b11 : 2'b10;
						assign node53 = (inp[4]) ? node57 : node54;
							assign node54 = (inp[3]) ? 2'b10 : 2'b11;
							assign node57 = (inp[3]) ? node59 : 2'b10;
								assign node59 = (inp[5]) ? 2'b10 : 2'b11;
					assign node62 = (inp[5]) ? node66 : node63;
						assign node63 = (inp[1]) ? 2'b01 : 2'b00;
						assign node66 = (inp[1]) ? 2'b00 : 2'b01;
				assign node69 = (inp[6]) ? node77 : node70;
					assign node70 = (inp[1]) ? node74 : node71;
						assign node71 = (inp[3]) ? 2'b01 : 2'b00;
						assign node74 = (inp[3]) ? 2'b00 : 2'b01;
					assign node77 = (inp[1]) ? 2'b00 : 2'b01;
		assign node80 = (inp[6]) ? node108 : node81;
			assign node81 = (inp[2]) ? node99 : node82;
				assign node82 = (inp[0]) ? node92 : node83;
					assign node83 = (inp[5]) ? 2'b10 : node84;
						assign node84 = (inp[4]) ? node86 : 2'b10;
							assign node86 = (inp[1]) ? node88 : 2'b11;
								assign node88 = (inp[3]) ? 2'b11 : 2'b10;
					assign node92 = (inp[3]) ? node96 : node93;
						assign node93 = (inp[5]) ? 2'b11 : 2'b10;
						assign node96 = (inp[5]) ? 2'b10 : 2'b11;
				assign node99 = (inp[3]) ? node103 : node100;
					assign node100 = (inp[4]) ? 2'b01 : 2'b00;
					assign node103 = (inp[0]) ? 2'b00 : node104;
						assign node104 = (inp[4]) ? 2'b00 : 2'b01;
			assign node108 = (inp[2]) ? node122 : node109;
				assign node109 = (inp[5]) ? node117 : node110;
					assign node110 = (inp[0]) ? 2'b01 : node111;
						assign node111 = (inp[4]) ? node113 : 2'b01;
							assign node113 = (inp[1]) ? 2'b01 : 2'b00;
					assign node117 = (inp[0]) ? 2'b00 : node118;
						assign node118 = (inp[3]) ? 2'b01 : 2'b00;
				assign node122 = (inp[4]) ? 2'b00 : node123;
					assign node123 = (inp[0]) ? 2'b00 : 2'b01;

endmodule