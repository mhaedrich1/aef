module dtc_split875_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node25;
	wire [14-1:0] node26;
	wire [14-1:0] node29;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node34;
	wire [14-1:0] node37;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node44;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node54;
	wire [14-1:0] node57;
	wire [14-1:0] node58;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node64;
	wire [14-1:0] node68;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node73;
	wire [14-1:0] node74;
	wire [14-1:0] node77;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node84;
	wire [14-1:0] node87;
	wire [14-1:0] node88;
	wire [14-1:0] node89;
	wire [14-1:0] node92;
	wire [14-1:0] node95;
	wire [14-1:0] node96;
	wire [14-1:0] node99;
	wire [14-1:0] node102;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node105;
	wire [14-1:0] node107;
	wire [14-1:0] node109;
	wire [14-1:0] node112;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node117;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node127;
	wire [14-1:0] node128;
	wire [14-1:0] node131;
	wire [14-1:0] node134;
	wire [14-1:0] node135;
	wire [14-1:0] node138;
	wire [14-1:0] node141;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node146;
	wire [14-1:0] node149;
	wire [14-1:0] node151;
	wire [14-1:0] node154;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node158;
	wire [14-1:0] node161;
	wire [14-1:0] node164;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node173;
	wire [14-1:0] node176;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node183;
	wire [14-1:0] node186;
	wire [14-1:0] node187;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node192;
	wire [14-1:0] node196;
	wire [14-1:0] node198;
	wire [14-1:0] node199;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node209;
	wire [14-1:0] node212;
	wire [14-1:0] node213;
	wire [14-1:0] node214;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node222;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node231;
	wire [14-1:0] node234;
	wire [14-1:0] node235;
	wire [14-1:0] node239;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node244;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node251;
	wire [14-1:0] node254;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node264;
	wire [14-1:0] node267;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node272;
	wire [14-1:0] node275;
	wire [14-1:0] node276;
	wire [14-1:0] node280;
	wire [14-1:0] node282;
	wire [14-1:0] node283;
	wire [14-1:0] node285;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node292;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node299;
	wire [14-1:0] node300;
	wire [14-1:0] node302;
	wire [14-1:0] node305;
	wire [14-1:0] node306;
	wire [14-1:0] node309;
	wire [14-1:0] node312;
	wire [14-1:0] node313;
	wire [14-1:0] node314;
	wire [14-1:0] node315;
	wire [14-1:0] node318;
	wire [14-1:0] node321;
	wire [14-1:0] node322;
	wire [14-1:0] node325;
	wire [14-1:0] node330;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node335;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node341;
	wire [14-1:0] node344;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node349;
	wire [14-1:0] node352;
	wire [14-1:0] node353;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node360;
	wire [14-1:0] node363;
	wire [14-1:0] node366;
	wire [14-1:0] node367;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node374;
	wire [14-1:0] node377;
	wire [14-1:0] node378;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node389;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node396;
	wire [14-1:0] node399;
	wire [14-1:0] node400;
	wire [14-1:0] node401;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node416;
	wire [14-1:0] node419;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node425;
	wire [14-1:0] node426;
	wire [14-1:0] node427;
	wire [14-1:0] node429;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node436;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node444;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node452;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node458;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node472;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node484;
	wire [14-1:0] node487;
	wire [14-1:0] node488;
	wire [14-1:0] node491;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node499;
	wire [14-1:0] node502;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node509;
	wire [14-1:0] node512;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node520;
	wire [14-1:0] node521;
	wire [14-1:0] node522;
	wire [14-1:0] node525;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node532;
	wire [14-1:0] node535;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node540;
	wire [14-1:0] node544;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node550;
	wire [14-1:0] node553;
	wire [14-1:0] node554;
	wire [14-1:0] node557;
	wire [14-1:0] node560;
	wire [14-1:0] node561;
	wire [14-1:0] node562;
	wire [14-1:0] node565;
	wire [14-1:0] node570;
	wire [14-1:0] node572;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node575;
	wire [14-1:0] node577;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node584;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node589;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node597;
	wire [14-1:0] node600;
	wire [14-1:0] node601;
	wire [14-1:0] node602;
	wire [14-1:0] node604;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node611;
	wire [14-1:0] node614;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node619;
	wire [14-1:0] node623;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node631;
	wire [14-1:0] node634;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node639;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node646;
	wire [14-1:0] node649;
	wire [14-1:0] node650;
	wire [14-1:0] node651;
	wire [14-1:0] node653;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node660;
	wire [14-1:0] node663;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node668;
	wire [14-1:0] node671;
	wire [14-1:0] node672;
	wire [14-1:0] node675;
	wire [14-1:0] node678;
	wire [14-1:0] node679;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node683;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node690;
	wire [14-1:0] node693;
	wire [14-1:0] node694;
	wire [14-1:0] node697;
	wire [14-1:0] node698;
	wire [14-1:0] node701;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node710;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node720;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node725;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node728;
	wire [14-1:0] node731;
	wire [14-1:0] node734;
	wire [14-1:0] node736;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node741;
	wire [14-1:0] node744;
	wire [14-1:0] node747;
	wire [14-1:0] node748;
	wire [14-1:0] node752;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node758;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node765;
	wire [14-1:0] node768;
	wire [14-1:0] node770;
	wire [14-1:0] node773;
	wire [14-1:0] node774;
	wire [14-1:0] node775;
	wire [14-1:0] node777;
	wire [14-1:0] node778;
	wire [14-1:0] node781;
	wire [14-1:0] node784;
	wire [14-1:0] node785;
	wire [14-1:0] node787;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node799;
	wire [14-1:0] node802;
	wire [14-1:0] node803;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node812;
	wire [14-1:0] node815;
	wire [14-1:0] node816;
	wire [14-1:0] node819;
	wire [14-1:0] node822;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node826;
	wire [14-1:0] node829;
	wire [14-1:0] node830;
	wire [14-1:0] node833;
	wire [14-1:0] node836;
	wire [14-1:0] node837;
	wire [14-1:0] node840;
	wire [14-1:0] node843;
	wire [14-1:0] node844;
	wire [14-1:0] node845;
	wire [14-1:0] node846;
	wire [14-1:0] node847;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node856;
	wire [14-1:0] node857;
	wire [14-1:0] node858;
	wire [14-1:0] node861;
	wire [14-1:0] node864;
	wire [14-1:0] node866;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node871;
	wire [14-1:0] node873;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node882;
	wire [14-1:0] node884;
	wire [14-1:0] node885;
	wire [14-1:0] node886;
	wire [14-1:0] node887;
	wire [14-1:0] node888;
	wire [14-1:0] node891;
	wire [14-1:0] node894;
	wire [14-1:0] node895;
	wire [14-1:0] node899;
	wire [14-1:0] node900;
	wire [14-1:0] node901;
	wire [14-1:0] node904;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node911;
	wire [14-1:0] node914;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node919;
	wire [14-1:0] node921;
	wire [14-1:0] node924;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node929;
	wire [14-1:0] node933;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node937;
	wire [14-1:0] node938;
	wire [14-1:0] node939;
	wire [14-1:0] node940;
	wire [14-1:0] node941;
	wire [14-1:0] node944;
	wire [14-1:0] node947;
	wire [14-1:0] node948;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node955;
	wire [14-1:0] node958;
	wire [14-1:0] node961;
	wire [14-1:0] node962;
	wire [14-1:0] node963;
	wire [14-1:0] node964;
	wire [14-1:0] node967;
	wire [14-1:0] node970;
	wire [14-1:0] node971;
	wire [14-1:0] node975;
	wire [14-1:0] node976;
	wire [14-1:0] node977;
	wire [14-1:0] node980;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node988;
	wire [14-1:0] node989;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node996;
	wire [14-1:0] node999;
	wire [14-1:0] node1000;
	wire [14-1:0] node1003;
	wire [14-1:0] node1006;
	wire [14-1:0] node1007;
	wire [14-1:0] node1008;
	wire [14-1:0] node1011;
	wire [14-1:0] node1014;
	wire [14-1:0] node1015;
	wire [14-1:0] node1018;
	wire [14-1:0] node1021;
	wire [14-1:0] node1022;
	wire [14-1:0] node1023;
	wire [14-1:0] node1024;
	wire [14-1:0] node1027;
	wire [14-1:0] node1030;
	wire [14-1:0] node1031;
	wire [14-1:0] node1034;
	wire [14-1:0] node1037;
	wire [14-1:0] node1038;
	wire [14-1:0] node1039;
	wire [14-1:0] node1042;
	wire [14-1:0] node1048;
	wire [14-1:0] node1049;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1053;
	wire [14-1:0] node1054;
	wire [14-1:0] node1056;
	wire [14-1:0] node1057;
	wire [14-1:0] node1059;
	wire [14-1:0] node1062;
	wire [14-1:0] node1064;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1069;
	wire [14-1:0] node1070;
	wire [14-1:0] node1074;
	wire [14-1:0] node1075;
	wire [14-1:0] node1078;
	wire [14-1:0] node1081;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1086;
	wire [14-1:0] node1089;
	wire [14-1:0] node1090;
	wire [14-1:0] node1093;
	wire [14-1:0] node1096;
	wire [14-1:0] node1097;
	wire [14-1:0] node1098;
	wire [14-1:0] node1099;
	wire [14-1:0] node1100;
	wire [14-1:0] node1103;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1111;
	wire [14-1:0] node1112;
	wire [14-1:0] node1113;
	wire [14-1:0] node1116;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1123;
	wire [14-1:0] node1126;
	wire [14-1:0] node1127;
	wire [14-1:0] node1128;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1135;
	wire [14-1:0] node1138;
	wire [14-1:0] node1139;
	wire [14-1:0] node1140;
	wire [14-1:0] node1143;
	wire [14-1:0] node1146;
	wire [14-1:0] node1147;
	wire [14-1:0] node1150;
	wire [14-1:0] node1153;
	wire [14-1:0] node1154;
	wire [14-1:0] node1155;
	wire [14-1:0] node1156;
	wire [14-1:0] node1157;
	wire [14-1:0] node1158;
	wire [14-1:0] node1162;
	wire [14-1:0] node1163;
	wire [14-1:0] node1166;
	wire [14-1:0] node1169;
	wire [14-1:0] node1170;
	wire [14-1:0] node1171;
	wire [14-1:0] node1174;
	wire [14-1:0] node1177;
	wire [14-1:0] node1178;
	wire [14-1:0] node1182;
	wire [14-1:0] node1183;
	wire [14-1:0] node1184;
	wire [14-1:0] node1185;
	wire [14-1:0] node1188;
	wire [14-1:0] node1191;
	wire [14-1:0] node1192;
	wire [14-1:0] node1195;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1203;
	wire [14-1:0] node1206;
	wire [14-1:0] node1207;
	wire [14-1:0] node1210;
	wire [14-1:0] node1213;
	wire [14-1:0] node1214;
	wire [14-1:0] node1215;
	wire [14-1:0] node1216;
	wire [14-1:0] node1218;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1225;
	wire [14-1:0] node1229;
	wire [14-1:0] node1231;
	wire [14-1:0] node1232;
	wire [14-1:0] node1233;
	wire [14-1:0] node1236;
	wire [14-1:0] node1239;
	wire [14-1:0] node1240;
	wire [14-1:0] node1243;
	wire [14-1:0] node1246;
	wire [14-1:0] node1247;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1250;
	wire [14-1:0] node1251;
	wire [14-1:0] node1252;
	wire [14-1:0] node1255;
	wire [14-1:0] node1258;
	wire [14-1:0] node1259;
	wire [14-1:0] node1262;
	wire [14-1:0] node1265;
	wire [14-1:0] node1266;
	wire [14-1:0] node1267;
	wire [14-1:0] node1270;
	wire [14-1:0] node1273;
	wire [14-1:0] node1274;
	wire [14-1:0] node1277;
	wire [14-1:0] node1280;
	wire [14-1:0] node1281;
	wire [14-1:0] node1282;
	wire [14-1:0] node1284;
	wire [14-1:0] node1287;
	wire [14-1:0] node1288;
	wire [14-1:0] node1291;
	wire [14-1:0] node1294;
	wire [14-1:0] node1295;
	wire [14-1:0] node1296;
	wire [14-1:0] node1300;
	wire [14-1:0] node1302;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1307;
	wire [14-1:0] node1308;
	wire [14-1:0] node1309;
	wire [14-1:0] node1313;
	wire [14-1:0] node1314;
	wire [14-1:0] node1317;
	wire [14-1:0] node1320;
	wire [14-1:0] node1321;
	wire [14-1:0] node1323;
	wire [14-1:0] node1326;
	wire [14-1:0] node1327;
	wire [14-1:0] node1330;
	wire [14-1:0] node1333;
	wire [14-1:0] node1335;
	wire [14-1:0] node1336;
	wire [14-1:0] node1337;
	wire [14-1:0] node1340;
	wire [14-1:0] node1343;
	wire [14-1:0] node1344;
	wire [14-1:0] node1347;
	wire [14-1:0] node1350;
	wire [14-1:0] node1351;
	wire [14-1:0] node1352;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1356;
	wire [14-1:0] node1360;
	wire [14-1:0] node1361;
	wire [14-1:0] node1364;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1370;
	wire [14-1:0] node1373;
	wire [14-1:0] node1376;
	wire [14-1:0] node1377;
	wire [14-1:0] node1380;
	wire [14-1:0] node1385;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1389;
	wire [14-1:0] node1390;
	wire [14-1:0] node1391;
	wire [14-1:0] node1392;
	wire [14-1:0] node1394;
	wire [14-1:0] node1397;
	wire [14-1:0] node1398;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1404;
	wire [14-1:0] node1407;
	wire [14-1:0] node1410;
	wire [14-1:0] node1413;
	wire [14-1:0] node1414;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1419;
	wire [14-1:0] node1422;
	wire [14-1:0] node1425;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1431;
	wire [14-1:0] node1433;
	wire [14-1:0] node1436;
	wire [14-1:0] node1437;
	wire [14-1:0] node1438;
	wire [14-1:0] node1439;
	wire [14-1:0] node1441;
	wire [14-1:0] node1444;
	wire [14-1:0] node1445;
	wire [14-1:0] node1448;
	wire [14-1:0] node1451;
	wire [14-1:0] node1452;
	wire [14-1:0] node1453;
	wire [14-1:0] node1457;
	wire [14-1:0] node1459;
	wire [14-1:0] node1462;
	wire [14-1:0] node1463;
	wire [14-1:0] node1465;
	wire [14-1:0] node1466;
	wire [14-1:0] node1469;
	wire [14-1:0] node1475;
	wire [14-1:0] node1476;
	wire [14-1:0] node1477;
	wire [14-1:0] node1478;
	wire [14-1:0] node1479;
	wire [14-1:0] node1480;
	wire [14-1:0] node1481;
	wire [14-1:0] node1482;
	wire [14-1:0] node1484;
	wire [14-1:0] node1485;
	wire [14-1:0] node1486;
	wire [14-1:0] node1490;
	wire [14-1:0] node1491;
	wire [14-1:0] node1495;
	wire [14-1:0] node1496;
	wire [14-1:0] node1497;
	wire [14-1:0] node1498;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1506;
	wire [14-1:0] node1509;
	wire [14-1:0] node1510;
	wire [14-1:0] node1512;
	wire [14-1:0] node1515;
	wire [14-1:0] node1516;
	wire [14-1:0] node1519;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1524;
	wire [14-1:0] node1525;
	wire [14-1:0] node1526;
	wire [14-1:0] node1529;
	wire [14-1:0] node1532;
	wire [14-1:0] node1535;
	wire [14-1:0] node1536;
	wire [14-1:0] node1537;
	wire [14-1:0] node1540;
	wire [14-1:0] node1543;
	wire [14-1:0] node1544;
	wire [14-1:0] node1547;
	wire [14-1:0] node1550;
	wire [14-1:0] node1551;
	wire [14-1:0] node1552;
	wire [14-1:0] node1553;
	wire [14-1:0] node1556;
	wire [14-1:0] node1559;
	wire [14-1:0] node1560;
	wire [14-1:0] node1564;
	wire [14-1:0] node1565;
	wire [14-1:0] node1567;
	wire [14-1:0] node1570;
	wire [14-1:0] node1571;
	wire [14-1:0] node1574;
	wire [14-1:0] node1577;
	wire [14-1:0] node1578;
	wire [14-1:0] node1579;
	wire [14-1:0] node1580;
	wire [14-1:0] node1581;
	wire [14-1:0] node1582;
	wire [14-1:0] node1585;
	wire [14-1:0] node1588;
	wire [14-1:0] node1590;
	wire [14-1:0] node1593;
	wire [14-1:0] node1594;
	wire [14-1:0] node1595;
	wire [14-1:0] node1598;
	wire [14-1:0] node1601;
	wire [14-1:0] node1603;
	wire [14-1:0] node1606;
	wire [14-1:0] node1607;
	wire [14-1:0] node1608;
	wire [14-1:0] node1611;
	wire [14-1:0] node1612;
	wire [14-1:0] node1615;
	wire [14-1:0] node1618;
	wire [14-1:0] node1619;
	wire [14-1:0] node1622;
	wire [14-1:0] node1623;
	wire [14-1:0] node1626;
	wire [14-1:0] node1629;
	wire [14-1:0] node1630;
	wire [14-1:0] node1631;
	wire [14-1:0] node1632;
	wire [14-1:0] node1633;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1641;
	wire [14-1:0] node1645;
	wire [14-1:0] node1647;
	wire [14-1:0] node1648;
	wire [14-1:0] node1649;
	wire [14-1:0] node1652;
	wire [14-1:0] node1655;
	wire [14-1:0] node1658;
	wire [14-1:0] node1659;
	wire [14-1:0] node1660;
	wire [14-1:0] node1661;
	wire [14-1:0] node1662;
	wire [14-1:0] node1663;
	wire [14-1:0] node1664;
	wire [14-1:0] node1667;
	wire [14-1:0] node1670;
	wire [14-1:0] node1671;
	wire [14-1:0] node1675;
	wire [14-1:0] node1676;
	wire [14-1:0] node1677;
	wire [14-1:0] node1680;
	wire [14-1:0] node1683;
	wire [14-1:0] node1684;
	wire [14-1:0] node1687;
	wire [14-1:0] node1690;
	wire [14-1:0] node1691;
	wire [14-1:0] node1692;
	wire [14-1:0] node1693;
	wire [14-1:0] node1696;
	wire [14-1:0] node1699;
	wire [14-1:0] node1700;
	wire [14-1:0] node1704;
	wire [14-1:0] node1705;
	wire [14-1:0] node1706;
	wire [14-1:0] node1709;
	wire [14-1:0] node1712;
	wire [14-1:0] node1713;
	wire [14-1:0] node1717;
	wire [14-1:0] node1718;
	wire [14-1:0] node1719;
	wire [14-1:0] node1720;
	wire [14-1:0] node1723;
	wire [14-1:0] node1724;
	wire [14-1:0] node1727;
	wire [14-1:0] node1730;
	wire [14-1:0] node1731;
	wire [14-1:0] node1733;
	wire [14-1:0] node1736;
	wire [14-1:0] node1737;
	wire [14-1:0] node1740;
	wire [14-1:0] node1743;
	wire [14-1:0] node1745;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1751;
	wire [14-1:0] node1752;
	wire [14-1:0] node1755;
	wire [14-1:0] node1758;
	wire [14-1:0] node1759;
	wire [14-1:0] node1760;
	wire [14-1:0] node1762;
	wire [14-1:0] node1763;
	wire [14-1:0] node1764;
	wire [14-1:0] node1767;
	wire [14-1:0] node1770;
	wire [14-1:0] node1771;
	wire [14-1:0] node1774;
	wire [14-1:0] node1777;
	wire [14-1:0] node1778;
	wire [14-1:0] node1779;
	wire [14-1:0] node1780;
	wire [14-1:0] node1783;
	wire [14-1:0] node1786;
	wire [14-1:0] node1787;
	wire [14-1:0] node1790;
	wire [14-1:0] node1795;
	wire [14-1:0] node1796;
	wire [14-1:0] node1797;
	wire [14-1:0] node1798;
	wire [14-1:0] node1799;
	wire [14-1:0] node1800;
	wire [14-1:0] node1801;
	wire [14-1:0] node1802;
	wire [14-1:0] node1806;
	wire [14-1:0] node1808;
	wire [14-1:0] node1811;
	wire [14-1:0] node1812;
	wire [14-1:0] node1813;
	wire [14-1:0] node1817;
	wire [14-1:0] node1818;
	wire [14-1:0] node1821;
	wire [14-1:0] node1824;
	wire [14-1:0] node1825;
	wire [14-1:0] node1826;
	wire [14-1:0] node1829;
	wire [14-1:0] node1831;
	wire [14-1:0] node1834;
	wire [14-1:0] node1835;
	wire [14-1:0] node1836;
	wire [14-1:0] node1839;
	wire [14-1:0] node1842;
	wire [14-1:0] node1843;
	wire [14-1:0] node1846;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1851;
	wire [14-1:0] node1852;
	wire [14-1:0] node1853;
	wire [14-1:0] node1856;
	wire [14-1:0] node1859;
	wire [14-1:0] node1860;
	wire [14-1:0] node1863;
	wire [14-1:0] node1866;
	wire [14-1:0] node1867;
	wire [14-1:0] node1870;
	wire [14-1:0] node1871;
	wire [14-1:0] node1875;
	wire [14-1:0] node1876;
	wire [14-1:0] node1877;
	wire [14-1:0] node1878;
	wire [14-1:0] node1881;
	wire [14-1:0] node1884;
	wire [14-1:0] node1885;
	wire [14-1:0] node1888;
	wire [14-1:0] node1891;
	wire [14-1:0] node1892;
	wire [14-1:0] node1894;
	wire [14-1:0] node1897;
	wire [14-1:0] node1898;
	wire [14-1:0] node1901;
	wire [14-1:0] node1904;
	wire [14-1:0] node1905;
	wire [14-1:0] node1907;
	wire [14-1:0] node1908;
	wire [14-1:0] node1909;
	wire [14-1:0] node1910;
	wire [14-1:0] node1914;
	wire [14-1:0] node1915;
	wire [14-1:0] node1918;
	wire [14-1:0] node1921;
	wire [14-1:0] node1922;
	wire [14-1:0] node1925;
	wire [14-1:0] node1926;
	wire [14-1:0] node1929;
	wire [14-1:0] node1934;
	wire [14-1:0] node1935;
	wire [14-1:0] node1936;
	wire [14-1:0] node1937;
	wire [14-1:0] node1939;
	wire [14-1:0] node1940;
	wire [14-1:0] node1941;
	wire [14-1:0] node1942;
	wire [14-1:0] node1943;
	wire [14-1:0] node1946;
	wire [14-1:0] node1953;
	wire [14-1:0] node1954;
	wire [14-1:0] node1955;
	wire [14-1:0] node1956;
	wire [14-1:0] node1957;
	wire [14-1:0] node1959;
	wire [14-1:0] node1960;
	wire [14-1:0] node1963;
	wire [14-1:0] node1966;
	wire [14-1:0] node1967;
	wire [14-1:0] node1969;
	wire [14-1:0] node1972;
	wire [14-1:0] node1975;
	wire [14-1:0] node1976;
	wire [14-1:0] node1977;
	wire [14-1:0] node1978;
	wire [14-1:0] node1981;
	wire [14-1:0] node1984;
	wire [14-1:0] node1985;
	wire [14-1:0] node1988;
	wire [14-1:0] node1991;
	wire [14-1:0] node1992;
	wire [14-1:0] node1993;
	wire [14-1:0] node1996;
	wire [14-1:0] node1999;
	wire [14-1:0] node2000;
	wire [14-1:0] node2003;
	wire [14-1:0] node2006;
	wire [14-1:0] node2007;
	wire [14-1:0] node2008;
	wire [14-1:0] node2009;
	wire [14-1:0] node2010;
	wire [14-1:0] node2013;
	wire [14-1:0] node2016;
	wire [14-1:0] node2018;
	wire [14-1:0] node2021;
	wire [14-1:0] node2023;
	wire [14-1:0] node2024;
	wire [14-1:0] node2028;
	wire [14-1:0] node2029;
	wire [14-1:0] node2031;
	wire [14-1:0] node2032;
	wire [14-1:0] node2035;
	wire [14-1:0] node2039;
	wire [14-1:0] node2040;
	wire [14-1:0] node2041;
	wire [14-1:0] node2042;
	wire [14-1:0] node2043;
	wire [14-1:0] node2044;
	wire [14-1:0] node2047;
	wire [14-1:0] node2050;
	wire [14-1:0] node2051;
	wire [14-1:0] node2055;
	wire [14-1:0] node2057;
	wire [14-1:0] node2060;
	wire [14-1:0] node2061;
	wire [14-1:0] node2062;
	wire [14-1:0] node2063;
	wire [14-1:0] node2067;
	wire [14-1:0] node2069;
	wire [14-1:0] node2072;
	wire [14-1:0] node2073;
	wire [14-1:0] node2075;
	wire [14-1:0] node2080;
	wire [14-1:0] node2081;
	wire [14-1:0] node2083;
	wire [14-1:0] node2084;
	wire [14-1:0] node2086;
	wire [14-1:0] node2087;
	wire [14-1:0] node2089;
	wire [14-1:0] node2096;
	wire [14-1:0] node2097;
	wire [14-1:0] node2098;
	wire [14-1:0] node2099;
	wire [14-1:0] node2100;
	wire [14-1:0] node2101;
	wire [14-1:0] node2102;
	wire [14-1:0] node2103;
	wire [14-1:0] node2104;
	wire [14-1:0] node2105;
	wire [14-1:0] node2106;
	wire [14-1:0] node2111;
	wire [14-1:0] node2112;
	wire [14-1:0] node2113;
	wire [14-1:0] node2114;
	wire [14-1:0] node2117;
	wire [14-1:0] node2120;
	wire [14-1:0] node2121;
	wire [14-1:0] node2125;
	wire [14-1:0] node2126;
	wire [14-1:0] node2127;
	wire [14-1:0] node2132;
	wire [14-1:0] node2133;
	wire [14-1:0] node2134;
	wire [14-1:0] node2135;
	wire [14-1:0] node2136;
	wire [14-1:0] node2139;
	wire [14-1:0] node2142;
	wire [14-1:0] node2143;
	wire [14-1:0] node2146;
	wire [14-1:0] node2149;
	wire [14-1:0] node2150;
	wire [14-1:0] node2151;
	wire [14-1:0] node2154;
	wire [14-1:0] node2157;
	wire [14-1:0] node2158;
	wire [14-1:0] node2161;
	wire [14-1:0] node2164;
	wire [14-1:0] node2165;
	wire [14-1:0] node2166;
	wire [14-1:0] node2169;
	wire [14-1:0] node2172;
	wire [14-1:0] node2173;
	wire [14-1:0] node2176;
	wire [14-1:0] node2179;
	wire [14-1:0] node2180;
	wire [14-1:0] node2181;
	wire [14-1:0] node2183;
	wire [14-1:0] node2184;
	wire [14-1:0] node2185;
	wire [14-1:0] node2188;
	wire [14-1:0] node2191;
	wire [14-1:0] node2194;
	wire [14-1:0] node2195;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2200;
	wire [14-1:0] node2203;
	wire [14-1:0] node2206;
	wire [14-1:0] node2207;
	wire [14-1:0] node2208;
	wire [14-1:0] node2211;
	wire [14-1:0] node2214;
	wire [14-1:0] node2217;
	wire [14-1:0] node2218;
	wire [14-1:0] node2219;
	wire [14-1:0] node2220;
	wire [14-1:0] node2221;
	wire [14-1:0] node2224;
	wire [14-1:0] node2227;
	wire [14-1:0] node2230;
	wire [14-1:0] node2231;
	wire [14-1:0] node2232;
	wire [14-1:0] node2235;
	wire [14-1:0] node2238;
	wire [14-1:0] node2241;
	wire [14-1:0] node2242;
	wire [14-1:0] node2243;
	wire [14-1:0] node2244;
	wire [14-1:0] node2247;
	wire [14-1:0] node2250;
	wire [14-1:0] node2253;
	wire [14-1:0] node2254;
	wire [14-1:0] node2255;
	wire [14-1:0] node2258;
	wire [14-1:0] node2261;
	wire [14-1:0] node2264;
	wire [14-1:0] node2265;
	wire [14-1:0] node2266;
	wire [14-1:0] node2267;
	wire [14-1:0] node2269;
	wire [14-1:0] node2270;
	wire [14-1:0] node2271;
	wire [14-1:0] node2274;
	wire [14-1:0] node2277;
	wire [14-1:0] node2280;
	wire [14-1:0] node2281;
	wire [14-1:0] node2282;
	wire [14-1:0] node2283;
	wire [14-1:0] node2286;
	wire [14-1:0] node2289;
	wire [14-1:0] node2292;
	wire [14-1:0] node2293;
	wire [14-1:0] node2294;
	wire [14-1:0] node2297;
	wire [14-1:0] node2300;
	wire [14-1:0] node2303;
	wire [14-1:0] node2304;
	wire [14-1:0] node2305;
	wire [14-1:0] node2306;
	wire [14-1:0] node2307;
	wire [14-1:0] node2310;
	wire [14-1:0] node2313;
	wire [14-1:0] node2316;
	wire [14-1:0] node2317;
	wire [14-1:0] node2318;
	wire [14-1:0] node2321;
	wire [14-1:0] node2324;
	wire [14-1:0] node2327;
	wire [14-1:0] node2328;
	wire [14-1:0] node2329;
	wire [14-1:0] node2331;
	wire [14-1:0] node2334;
	wire [14-1:0] node2337;
	wire [14-1:0] node2338;
	wire [14-1:0] node2339;
	wire [14-1:0] node2342;
	wire [14-1:0] node2345;
	wire [14-1:0] node2348;
	wire [14-1:0] node2349;
	wire [14-1:0] node2350;
	wire [14-1:0] node2352;
	wire [14-1:0] node2353;
	wire [14-1:0] node2354;
	wire [14-1:0] node2357;
	wire [14-1:0] node2360;
	wire [14-1:0] node2363;
	wire [14-1:0] node2364;
	wire [14-1:0] node2365;
	wire [14-1:0] node2366;
	wire [14-1:0] node2369;
	wire [14-1:0] node2372;
	wire [14-1:0] node2375;
	wire [14-1:0] node2376;
	wire [14-1:0] node2377;
	wire [14-1:0] node2380;
	wire [14-1:0] node2383;
	wire [14-1:0] node2386;
	wire [14-1:0] node2387;
	wire [14-1:0] node2388;
	wire [14-1:0] node2389;
	wire [14-1:0] node2390;
	wire [14-1:0] node2393;
	wire [14-1:0] node2396;
	wire [14-1:0] node2397;
	wire [14-1:0] node2400;
	wire [14-1:0] node2403;
	wire [14-1:0] node2404;
	wire [14-1:0] node2405;
	wire [14-1:0] node2408;
	wire [14-1:0] node2411;
	wire [14-1:0] node2412;
	wire [14-1:0] node2415;
	wire [14-1:0] node2418;
	wire [14-1:0] node2419;
	wire [14-1:0] node2420;
	wire [14-1:0] node2423;
	wire [14-1:0] node2426;
	wire [14-1:0] node2427;
	wire [14-1:0] node2430;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2437;
	wire [14-1:0] node2438;
	wire [14-1:0] node2439;
	wire [14-1:0] node2440;
	wire [14-1:0] node2443;
	wire [14-1:0] node2446;
	wire [14-1:0] node2447;
	wire [14-1:0] node2450;
	wire [14-1:0] node2453;
	wire [14-1:0] node2454;
	wire [14-1:0] node2456;
	wire [14-1:0] node2459;
	wire [14-1:0] node2460;
	wire [14-1:0] node2463;
	wire [14-1:0] node2466;
	wire [14-1:0] node2467;
	wire [14-1:0] node2468;
	wire [14-1:0] node2469;
	wire [14-1:0] node2472;
	wire [14-1:0] node2475;
	wire [14-1:0] node2476;
	wire [14-1:0] node2479;
	wire [14-1:0] node2482;
	wire [14-1:0] node2483;
	wire [14-1:0] node2484;
	wire [14-1:0] node2487;
	wire [14-1:0] node2490;
	wire [14-1:0] node2491;
	wire [14-1:0] node2494;
	wire [14-1:0] node2497;
	wire [14-1:0] node2498;
	wire [14-1:0] node2499;
	wire [14-1:0] node2501;
	wire [14-1:0] node2502;
	wire [14-1:0] node2505;
	wire [14-1:0] node2508;
	wire [14-1:0] node2509;
	wire [14-1:0] node2510;
	wire [14-1:0] node2513;
	wire [14-1:0] node2516;
	wire [14-1:0] node2517;
	wire [14-1:0] node2520;
	wire [14-1:0] node2523;
	wire [14-1:0] node2524;
	wire [14-1:0] node2525;
	wire [14-1:0] node2526;
	wire [14-1:0] node2529;
	wire [14-1:0] node2532;
	wire [14-1:0] node2533;
	wire [14-1:0] node2536;
	wire [14-1:0] node2539;
	wire [14-1:0] node2540;
	wire [14-1:0] node2541;
	wire [14-1:0] node2544;
	wire [14-1:0] node2547;
	wire [14-1:0] node2548;
	wire [14-1:0] node2551;
	wire [14-1:0] node2554;
	wire [14-1:0] node2556;
	wire [14-1:0] node2557;
	wire [14-1:0] node2558;
	wire [14-1:0] node2559;
	wire [14-1:0] node2561;
	wire [14-1:0] node2564;
	wire [14-1:0] node2565;
	wire [14-1:0] node2568;
	wire [14-1:0] node2571;
	wire [14-1:0] node2572;
	wire [14-1:0] node2573;
	wire [14-1:0] node2576;
	wire [14-1:0] node2579;
	wire [14-1:0] node2580;
	wire [14-1:0] node2583;
	wire [14-1:0] node2586;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2589;
	wire [14-1:0] node2592;
	wire [14-1:0] node2595;
	wire [14-1:0] node2596;
	wire [14-1:0] node2599;
	wire [14-1:0] node2602;
	wire [14-1:0] node2603;
	wire [14-1:0] node2604;
	wire [14-1:0] node2607;
	wire [14-1:0] node2610;
	wire [14-1:0] node2611;
	wire [14-1:0] node2614;
	wire [14-1:0] node2617;
	wire [14-1:0] node2618;
	wire [14-1:0] node2619;
	wire [14-1:0] node2620;
	wire [14-1:0] node2622;
	wire [14-1:0] node2623;
	wire [14-1:0] node2624;
	wire [14-1:0] node2627;
	wire [14-1:0] node2630;
	wire [14-1:0] node2631;
	wire [14-1:0] node2634;
	wire [14-1:0] node2637;
	wire [14-1:0] node2638;
	wire [14-1:0] node2639;
	wire [14-1:0] node2640;
	wire [14-1:0] node2643;
	wire [14-1:0] node2646;
	wire [14-1:0] node2647;
	wire [14-1:0] node2650;
	wire [14-1:0] node2653;
	wire [14-1:0] node2654;
	wire [14-1:0] node2655;
	wire [14-1:0] node2658;
	wire [14-1:0] node2661;
	wire [14-1:0] node2662;
	wire [14-1:0] node2665;
	wire [14-1:0] node2670;
	wire [14-1:0] node2671;
	wire [14-1:0] node2672;
	wire [14-1:0] node2673;
	wire [14-1:0] node2674;
	wire [14-1:0] node2675;
	wire [14-1:0] node2676;
	wire [14-1:0] node2678;
	wire [14-1:0] node2679;
	wire [14-1:0] node2682;
	wire [14-1:0] node2686;
	wire [14-1:0] node2687;
	wire [14-1:0] node2688;
	wire [14-1:0] node2689;
	wire [14-1:0] node2692;
	wire [14-1:0] node2695;
	wire [14-1:0] node2696;
	wire [14-1:0] node2699;
	wire [14-1:0] node2702;
	wire [14-1:0] node2703;
	wire [14-1:0] node2706;
	wire [14-1:0] node2709;
	wire [14-1:0] node2710;
	wire [14-1:0] node2711;
	wire [14-1:0] node2712;
	wire [14-1:0] node2713;
	wire [14-1:0] node2716;
	wire [14-1:0] node2719;
	wire [14-1:0] node2720;
	wire [14-1:0] node2723;
	wire [14-1:0] node2726;
	wire [14-1:0] node2727;
	wire [14-1:0] node2730;
	wire [14-1:0] node2733;
	wire [14-1:0] node2734;
	wire [14-1:0] node2735;
	wire [14-1:0] node2736;
	wire [14-1:0] node2739;
	wire [14-1:0] node2742;
	wire [14-1:0] node2745;
	wire [14-1:0] node2746;
	wire [14-1:0] node2747;
	wire [14-1:0] node2750;
	wire [14-1:0] node2753;
	wire [14-1:0] node2756;
	wire [14-1:0] node2757;
	wire [14-1:0] node2758;
	wire [14-1:0] node2759;
	wire [14-1:0] node2760;
	wire [14-1:0] node2761;
	wire [14-1:0] node2764;
	wire [14-1:0] node2767;
	wire [14-1:0] node2770;
	wire [14-1:0] node2771;
	wire [14-1:0] node2772;
	wire [14-1:0] node2775;
	wire [14-1:0] node2778;
	wire [14-1:0] node2781;
	wire [14-1:0] node2782;
	wire [14-1:0] node2783;
	wire [14-1:0] node2784;
	wire [14-1:0] node2787;
	wire [14-1:0] node2790;
	wire [14-1:0] node2793;
	wire [14-1:0] node2794;
	wire [14-1:0] node2795;
	wire [14-1:0] node2798;
	wire [14-1:0] node2801;
	wire [14-1:0] node2804;
	wire [14-1:0] node2805;
	wire [14-1:0] node2806;
	wire [14-1:0] node2807;
	wire [14-1:0] node2808;
	wire [14-1:0] node2811;
	wire [14-1:0] node2814;
	wire [14-1:0] node2817;
	wire [14-1:0] node2818;
	wire [14-1:0] node2819;
	wire [14-1:0] node2822;
	wire [14-1:0] node2825;
	wire [14-1:0] node2828;
	wire [14-1:0] node2829;
	wire [14-1:0] node2830;
	wire [14-1:0] node2831;
	wire [14-1:0] node2834;
	wire [14-1:0] node2837;
	wire [14-1:0] node2840;
	wire [14-1:0] node2841;
	wire [14-1:0] node2842;
	wire [14-1:0] node2845;
	wire [14-1:0] node2848;
	wire [14-1:0] node2851;
	wire [14-1:0] node2852;
	wire [14-1:0] node2853;
	wire [14-1:0] node2854;
	wire [14-1:0] node2855;
	wire [14-1:0] node2856;
	wire [14-1:0] node2857;
	wire [14-1:0] node2860;
	wire [14-1:0] node2863;
	wire [14-1:0] node2864;
	wire [14-1:0] node2867;
	wire [14-1:0] node2870;
	wire [14-1:0] node2871;
	wire [14-1:0] node2872;
	wire [14-1:0] node2875;
	wire [14-1:0] node2878;
	wire [14-1:0] node2879;
	wire [14-1:0] node2882;
	wire [14-1:0] node2885;
	wire [14-1:0] node2886;
	wire [14-1:0] node2887;
	wire [14-1:0] node2888;
	wire [14-1:0] node2891;
	wire [14-1:0] node2894;
	wire [14-1:0] node2895;
	wire [14-1:0] node2898;
	wire [14-1:0] node2901;
	wire [14-1:0] node2902;
	wire [14-1:0] node2903;
	wire [14-1:0] node2906;
	wire [14-1:0] node2909;
	wire [14-1:0] node2910;
	wire [14-1:0] node2913;
	wire [14-1:0] node2916;
	wire [14-1:0] node2918;
	wire [14-1:0] node2919;
	wire [14-1:0] node2920;
	wire [14-1:0] node2921;
	wire [14-1:0] node2924;
	wire [14-1:0] node2927;
	wire [14-1:0] node2928;
	wire [14-1:0] node2931;
	wire [14-1:0] node2934;
	wire [14-1:0] node2935;
	wire [14-1:0] node2936;
	wire [14-1:0] node2939;
	wire [14-1:0] node2942;
	wire [14-1:0] node2943;
	wire [14-1:0] node2946;
	wire [14-1:0] node2949;
	wire [14-1:0] node2950;
	wire [14-1:0] node2951;
	wire [14-1:0] node2952;
	wire [14-1:0] node2954;
	wire [14-1:0] node2956;
	wire [14-1:0] node2959;
	wire [14-1:0] node2960;
	wire [14-1:0] node2961;
	wire [14-1:0] node2964;
	wire [14-1:0] node2967;
	wire [14-1:0] node2968;
	wire [14-1:0] node2971;
	wire [14-1:0] node2976;
	wire [14-1:0] node2978;
	wire [14-1:0] node2979;
	wire [14-1:0] node2980;
	wire [14-1:0] node2981;
	wire [14-1:0] node2982;
	wire [14-1:0] node2983;
	wire [14-1:0] node2984;
	wire [14-1:0] node2990;
	wire [14-1:0] node2991;
	wire [14-1:0] node2992;
	wire [14-1:0] node2994;
	wire [14-1:0] node2998;
	wire [14-1:0] node3000;
	wire [14-1:0] node3001;
	wire [14-1:0] node3007;
	wire [14-1:0] node3008;
	wire [14-1:0] node3009;
	wire [14-1:0] node3010;
	wire [14-1:0] node3011;
	wire [14-1:0] node3012;
	wire [14-1:0] node3013;
	wire [14-1:0] node3014;
	wire [14-1:0] node3015;
	wire [14-1:0] node3017;
	wire [14-1:0] node3020;
	wire [14-1:0] node3021;
	wire [14-1:0] node3024;
	wire [14-1:0] node3027;
	wire [14-1:0] node3028;
	wire [14-1:0] node3029;
	wire [14-1:0] node3032;
	wire [14-1:0] node3035;
	wire [14-1:0] node3036;
	wire [14-1:0] node3039;
	wire [14-1:0] node3042;
	wire [14-1:0] node3043;
	wire [14-1:0] node3044;
	wire [14-1:0] node3046;
	wire [14-1:0] node3049;
	wire [14-1:0] node3050;
	wire [14-1:0] node3053;
	wire [14-1:0] node3056;
	wire [14-1:0] node3057;
	wire [14-1:0] node3058;
	wire [14-1:0] node3061;
	wire [14-1:0] node3064;
	wire [14-1:0] node3065;
	wire [14-1:0] node3068;
	wire [14-1:0] node3071;
	wire [14-1:0] node3072;
	wire [14-1:0] node3073;
	wire [14-1:0] node3074;
	wire [14-1:0] node3075;
	wire [14-1:0] node3078;
	wire [14-1:0] node3081;
	wire [14-1:0] node3082;
	wire [14-1:0] node3085;
	wire [14-1:0] node3088;
	wire [14-1:0] node3089;
	wire [14-1:0] node3090;
	wire [14-1:0] node3093;
	wire [14-1:0] node3096;
	wire [14-1:0] node3097;
	wire [14-1:0] node3100;
	wire [14-1:0] node3105;
	wire [14-1:0] node3106;
	wire [14-1:0] node3107;
	wire [14-1:0] node3108;
	wire [14-1:0] node3109;
	wire [14-1:0] node3111;
	wire [14-1:0] node3114;
	wire [14-1:0] node3115;
	wire [14-1:0] node3118;
	wire [14-1:0] node3121;
	wire [14-1:0] node3122;
	wire [14-1:0] node3123;
	wire [14-1:0] node3126;
	wire [14-1:0] node3129;
	wire [14-1:0] node3130;
	wire [14-1:0] node3133;
	wire [14-1:0] node3136;
	wire [14-1:0] node3137;
	wire [14-1:0] node3138;
	wire [14-1:0] node3140;
	wire [14-1:0] node3143;
	wire [14-1:0] node3144;
	wire [14-1:0] node3147;
	wire [14-1:0] node3150;
	wire [14-1:0] node3151;
	wire [14-1:0] node3152;
	wire [14-1:0] node3155;
	wire [14-1:0] node3158;
	wire [14-1:0] node3159;
	wire [14-1:0] node3162;
	wire [14-1:0] node3165;
	wire [14-1:0] node3166;
	wire [14-1:0] node3167;
	wire [14-1:0] node3168;
	wire [14-1:0] node3169;
	wire [14-1:0] node3172;
	wire [14-1:0] node3175;
	wire [14-1:0] node3176;
	wire [14-1:0] node3179;
	wire [14-1:0] node3182;
	wire [14-1:0] node3183;
	wire [14-1:0] node3184;
	wire [14-1:0] node3187;
	wire [14-1:0] node3190;
	wire [14-1:0] node3191;
	wire [14-1:0] node3194;
	wire [14-1:0] node3198;
	wire [14-1:0] node3199;
	wire [14-1:0] node3200;
	wire [14-1:0] node3201;
	wire [14-1:0] node3202;
	wire [14-1:0] node3203;
	wire [14-1:0] node3204;
	wire [14-1:0] node3206;
	wire [14-1:0] node3209;
	wire [14-1:0] node3210;
	wire [14-1:0] node3213;
	wire [14-1:0] node3216;
	wire [14-1:0] node3217;
	wire [14-1:0] node3218;
	wire [14-1:0] node3221;
	wire [14-1:0] node3224;
	wire [14-1:0] node3225;
	wire [14-1:0] node3228;
	wire [14-1:0] node3231;
	wire [14-1:0] node3232;
	wire [14-1:0] node3233;
	wire [14-1:0] node3234;
	wire [14-1:0] node3237;
	wire [14-1:0] node3240;
	wire [14-1:0] node3241;
	wire [14-1:0] node3244;
	wire [14-1:0] node3248;
	wire [14-1:0] node3249;
	wire [14-1:0] node3251;
	wire [14-1:0] node3253;
	wire [14-1:0] node3254;
	wire [14-1:0] node3258;
	wire [14-1:0] node3259;
	wire [14-1:0] node3260;
	wire [14-1:0] node3261;
	wire [14-1:0] node3264;
	wire [14-1:0] node3267;
	wire [14-1:0] node3268;
	wire [14-1:0] node3271;
	wire [14-1:0] node3274;
	wire [14-1:0] node3275;
	wire [14-1:0] node3276;
	wire [14-1:0] node3279;
	wire [14-1:0] node3283;
	wire [14-1:0] node3285;
	wire [14-1:0] node3286;
	wire [14-1:0] node3288;
	wire [14-1:0] node3289;
	wire [14-1:0] node3291;
	wire [14-1:0] node3295;
	wire [14-1:0] node3296;
	wire [14-1:0] node3297;
	wire [14-1:0] node3298;
	wire [14-1:0] node3301;
	wire [14-1:0] node3304;
	wire [14-1:0] node3305;
	wire [14-1:0] node3308;
	wire [14-1:0] node3311;
	wire [14-1:0] node3312;
	wire [14-1:0] node3313;
	wire [14-1:0] node3316;
	wire [14-1:0] node3321;
	wire [14-1:0] node3322;
	wire [14-1:0] node3323;
	wire [14-1:0] node3324;
	wire [14-1:0] node3325;
	wire [14-1:0] node3326;
	wire [14-1:0] node3327;
	wire [14-1:0] node3328;
	wire [14-1:0] node3329;
	wire [14-1:0] node3332;
	wire [14-1:0] node3335;
	wire [14-1:0] node3336;
	wire [14-1:0] node3339;
	wire [14-1:0] node3342;
	wire [14-1:0] node3343;
	wire [14-1:0] node3344;
	wire [14-1:0] node3347;
	wire [14-1:0] node3350;
	wire [14-1:0] node3351;
	wire [14-1:0] node3354;
	wire [14-1:0] node3357;
	wire [14-1:0] node3358;
	wire [14-1:0] node3359;
	wire [14-1:0] node3360;
	wire [14-1:0] node3363;
	wire [14-1:0] node3366;
	wire [14-1:0] node3367;
	wire [14-1:0] node3370;
	wire [14-1:0] node3374;
	wire [14-1:0] node3376;
	wire [14-1:0] node3377;
	wire [14-1:0] node3378;
	wire [14-1:0] node3379;
	wire [14-1:0] node3382;
	wire [14-1:0] node3385;
	wire [14-1:0] node3386;
	wire [14-1:0] node3389;
	wire [14-1:0] node3392;
	wire [14-1:0] node3393;
	wire [14-1:0] node3394;
	wire [14-1:0] node3397;
	wire [14-1:0] node3401;
	wire [14-1:0] node3402;
	wire [14-1:0] node3404;
	wire [14-1:0] node3405;
	wire [14-1:0] node3406;
	wire [14-1:0] node3407;
	wire [14-1:0] node3410;
	wire [14-1:0] node3413;
	wire [14-1:0] node3414;
	wire [14-1:0] node3417;
	wire [14-1:0] node3420;
	wire [14-1:0] node3421;
	wire [14-1:0] node3422;
	wire [14-1:0] node3425;
	wire [14-1:0] node3430;
	wire [14-1:0] node3431;
	wire [14-1:0] node3432;
	wire [14-1:0] node3433;
	wire [14-1:0] node3435;
	wire [14-1:0] node3436;
	wire [14-1:0] node3438;
	wire [14-1:0] node3442;
	wire [14-1:0] node3443;
	wire [14-1:0] node3444;
	wire [14-1:0] node3445;
	wire [14-1:0] node3453;
	wire [14-1:0] node3454;
	wire [14-1:0] node3456;
	wire [14-1:0] node3457;
	wire [14-1:0] node3458;
	wire [14-1:0] node3459;
	wire [14-1:0] node3461;
	wire [14-1:0] node3462;
	wire [14-1:0] node3466;
	wire [14-1:0] node3467;
	wire [14-1:0] node3468;
	wire [14-1:0] node3473;
	wire [14-1:0] node3475;
	wire [14-1:0] node3476;
	wire [14-1:0] node3477;
	wire [14-1:0] node3484;
	wire [14-1:0] node3485;
	wire [14-1:0] node3486;
	wire [14-1:0] node3487;
	wire [14-1:0] node3488;
	wire [14-1:0] node3489;
	wire [14-1:0] node3490;
	wire [14-1:0] node3491;
	wire [14-1:0] node3492;
	wire [14-1:0] node3494;
	wire [14-1:0] node3495;
	wire [14-1:0] node3498;
	wire [14-1:0] node3502;
	wire [14-1:0] node3503;
	wire [14-1:0] node3504;
	wire [14-1:0] node3505;
	wire [14-1:0] node3508;
	wire [14-1:0] node3511;
	wire [14-1:0] node3512;
	wire [14-1:0] node3516;
	wire [14-1:0] node3517;
	wire [14-1:0] node3520;
	wire [14-1:0] node3523;
	wire [14-1:0] node3524;
	wire [14-1:0] node3525;
	wire [14-1:0] node3526;
	wire [14-1:0] node3527;
	wire [14-1:0] node3530;
	wire [14-1:0] node3533;
	wire [14-1:0] node3536;
	wire [14-1:0] node3537;
	wire [14-1:0] node3538;
	wire [14-1:0] node3541;
	wire [14-1:0] node3544;
	wire [14-1:0] node3547;
	wire [14-1:0] node3548;
	wire [14-1:0] node3549;
	wire [14-1:0] node3550;
	wire [14-1:0] node3553;
	wire [14-1:0] node3556;
	wire [14-1:0] node3559;
	wire [14-1:0] node3560;
	wire [14-1:0] node3561;
	wire [14-1:0] node3564;
	wire [14-1:0] node3567;
	wire [14-1:0] node3570;
	wire [14-1:0] node3571;
	wire [14-1:0] node3572;
	wire [14-1:0] node3573;
	wire [14-1:0] node3574;
	wire [14-1:0] node3575;
	wire [14-1:0] node3578;
	wire [14-1:0] node3581;
	wire [14-1:0] node3584;
	wire [14-1:0] node3585;
	wire [14-1:0] node3586;
	wire [14-1:0] node3589;
	wire [14-1:0] node3592;
	wire [14-1:0] node3595;
	wire [14-1:0] node3596;
	wire [14-1:0] node3597;
	wire [14-1:0] node3598;
	wire [14-1:0] node3601;
	wire [14-1:0] node3604;
	wire [14-1:0] node3607;
	wire [14-1:0] node3608;
	wire [14-1:0] node3609;
	wire [14-1:0] node3612;
	wire [14-1:0] node3615;
	wire [14-1:0] node3618;
	wire [14-1:0] node3619;
	wire [14-1:0] node3620;
	wire [14-1:0] node3621;
	wire [14-1:0] node3622;
	wire [14-1:0] node3625;
	wire [14-1:0] node3628;
	wire [14-1:0] node3631;
	wire [14-1:0] node3632;
	wire [14-1:0] node3633;
	wire [14-1:0] node3637;
	wire [14-1:0] node3640;
	wire [14-1:0] node3641;
	wire [14-1:0] node3642;
	wire [14-1:0] node3643;
	wire [14-1:0] node3646;
	wire [14-1:0] node3649;
	wire [14-1:0] node3652;
	wire [14-1:0] node3653;
	wire [14-1:0] node3654;
	wire [14-1:0] node3657;
	wire [14-1:0] node3660;
	wire [14-1:0] node3663;
	wire [14-1:0] node3664;
	wire [14-1:0] node3665;
	wire [14-1:0] node3666;
	wire [14-1:0] node3667;
	wire [14-1:0] node3668;
	wire [14-1:0] node3669;
	wire [14-1:0] node3672;
	wire [14-1:0] node3675;
	wire [14-1:0] node3676;
	wire [14-1:0] node3679;
	wire [14-1:0] node3682;
	wire [14-1:0] node3683;
	wire [14-1:0] node3684;
	wire [14-1:0] node3687;
	wire [14-1:0] node3690;
	wire [14-1:0] node3691;
	wire [14-1:0] node3694;
	wire [14-1:0] node3697;
	wire [14-1:0] node3698;
	wire [14-1:0] node3699;
	wire [14-1:0] node3700;
	wire [14-1:0] node3703;
	wire [14-1:0] node3706;
	wire [14-1:0] node3707;
	wire [14-1:0] node3710;
	wire [14-1:0] node3713;
	wire [14-1:0] node3714;
	wire [14-1:0] node3715;
	wire [14-1:0] node3718;
	wire [14-1:0] node3721;
	wire [14-1:0] node3722;
	wire [14-1:0] node3725;
	wire [14-1:0] node3728;
	wire [14-1:0] node3730;
	wire [14-1:0] node3731;
	wire [14-1:0] node3732;
	wire [14-1:0] node3734;
	wire [14-1:0] node3737;
	wire [14-1:0] node3738;
	wire [14-1:0] node3741;
	wire [14-1:0] node3744;
	wire [14-1:0] node3745;
	wire [14-1:0] node3746;
	wire [14-1:0] node3749;
	wire [14-1:0] node3752;
	wire [14-1:0] node3753;
	wire [14-1:0] node3757;
	wire [14-1:0] node3758;
	wire [14-1:0] node3759;
	wire [14-1:0] node3760;
	wire [14-1:0] node3762;
	wire [14-1:0] node3763;
	wire [14-1:0] node3766;
	wire [14-1:0] node3769;
	wire [14-1:0] node3770;
	wire [14-1:0] node3771;
	wire [14-1:0] node3774;
	wire [14-1:0] node3777;
	wire [14-1:0] node3778;
	wire [14-1:0] node3781;
	wire [14-1:0] node3786;
	wire [14-1:0] node3787;
	wire [14-1:0] node3788;
	wire [14-1:0] node3789;
	wire [14-1:0] node3790;
	wire [14-1:0] node3791;
	wire [14-1:0] node3792;
	wire [14-1:0] node3793;
	wire [14-1:0] node3796;
	wire [14-1:0] node3799;
	wire [14-1:0] node3800;
	wire [14-1:0] node3803;
	wire [14-1:0] node3806;
	wire [14-1:0] node3807;
	wire [14-1:0] node3808;
	wire [14-1:0] node3811;
	wire [14-1:0] node3814;
	wire [14-1:0] node3815;
	wire [14-1:0] node3818;
	wire [14-1:0] node3822;
	wire [14-1:0] node3823;
	wire [14-1:0] node3824;
	wire [14-1:0] node3825;
	wire [14-1:0] node3828;
	wire [14-1:0] node3831;
	wire [14-1:0] node3832;
	wire [14-1:0] node3835;
	wire [14-1:0] node3838;
	wire [14-1:0] node3839;
	wire [14-1:0] node3840;
	wire [14-1:0] node3843;
	wire [14-1:0] node3846;
	wire [14-1:0] node3847;
	wire [14-1:0] node3850;
	wire [14-1:0] node3853;
	wire [14-1:0] node3854;
	wire [14-1:0] node3855;
	wire [14-1:0] node3856;
	wire [14-1:0] node3857;
	wire [14-1:0] node3858;
	wire [14-1:0] node3862;
	wire [14-1:0] node3863;
	wire [14-1:0] node3866;
	wire [14-1:0] node3869;
	wire [14-1:0] node3871;
	wire [14-1:0] node3872;
	wire [14-1:0] node3875;
	wire [14-1:0] node3878;
	wire [14-1:0] node3880;
	wire [14-1:0] node3882;
	wire [14-1:0] node3883;
	wire [14-1:0] node3886;
	wire [14-1:0] node3890;
	wire [14-1:0] node3891;
	wire [14-1:0] node3892;
	wire [14-1:0] node3893;
	wire [14-1:0] node3894;
	wire [14-1:0] node3895;
	wire [14-1:0] node3896;
	wire [14-1:0] node3899;
	wire [14-1:0] node3902;
	wire [14-1:0] node3903;
	wire [14-1:0] node3907;
	wire [14-1:0] node3909;
	wire [14-1:0] node3910;
	wire [14-1:0] node3913;
	wire [14-1:0] node3916;
	wire [14-1:0] node3917;
	wire [14-1:0] node3919;
	wire [14-1:0] node3920;
	wire [14-1:0] node3923;
	wire [14-1:0] node3929;
	wire [14-1:0] node3930;
	wire [14-1:0] node3931;
	wire [14-1:0] node3932;
	wire [14-1:0] node3933;
	wire [14-1:0] node3934;
	wire [14-1:0] node3936;
	wire [14-1:0] node3937;
	wire [14-1:0] node3939;
	wire [14-1:0] node3942;
	wire [14-1:0] node3948;
	wire [14-1:0] node3949;
	wire [14-1:0] node3950;
	wire [14-1:0] node3951;
	wire [14-1:0] node3952;
	wire [14-1:0] node3953;
	wire [14-1:0] node3954;
	wire [14-1:0] node3957;
	wire [14-1:0] node3960;
	wire [14-1:0] node3963;
	wire [14-1:0] node3964;
	wire [14-1:0] node3965;
	wire [14-1:0] node3968;
	wire [14-1:0] node3971;
	wire [14-1:0] node3974;
	wire [14-1:0] node3975;
	wire [14-1:0] node3976;
	wire [14-1:0] node3977;
	wire [14-1:0] node3980;
	wire [14-1:0] node3983;
	wire [14-1:0] node3986;
	wire [14-1:0] node3987;
	wire [14-1:0] node3988;
	wire [14-1:0] node3991;
	wire [14-1:0] node3994;
	wire [14-1:0] node3997;
	wire [14-1:0] node3998;
	wire [14-1:0] node3999;
	wire [14-1:0] node4000;
	wire [14-1:0] node4001;
	wire [14-1:0] node4004;
	wire [14-1:0] node4007;
	wire [14-1:0] node4008;
	wire [14-1:0] node4011;
	wire [14-1:0] node4014;
	wire [14-1:0] node4016;
	wire [14-1:0] node4017;
	wire [14-1:0] node4020;
	wire [14-1:0] node4023;
	wire [14-1:0] node4024;
	wire [14-1:0] node4025;
	wire [14-1:0] node4026;
	wire [14-1:0] node4029;
	wire [14-1:0] node4034;
	wire [14-1:0] node4035;
	wire [14-1:0] node4036;
	wire [14-1:0] node4037;
	wire [14-1:0] node4038;
	wire [14-1:0] node4039;
	wire [14-1:0] node4042;
	wire [14-1:0] node4046;
	wire [14-1:0] node4047;
	wire [14-1:0] node4050;
	wire [14-1:0] node4053;
	wire [14-1:0] node4054;
	wire [14-1:0] node4055;
	wire [14-1:0] node4056;
	wire [14-1:0] node4059;
	wire [14-1:0] node4062;
	wire [14-1:0] node4064;
	wire [14-1:0] node4068;
	wire [14-1:0] node4069;
	wire [14-1:0] node4070;
	wire [14-1:0] node4071;
	wire [14-1:0] node4072;
	wire [14-1:0] node4075;
	wire [14-1:0] node4078;
	wire [14-1:0] node4080;
	wire [14-1:0] node4086;
	wire [14-1:0] node4087;
	wire [14-1:0] node4088;
	wire [14-1:0] node4089;
	wire [14-1:0] node4090;
	wire [14-1:0] node4091;
	wire [14-1:0] node4092;
	wire [14-1:0] node4094;
	wire [14-1:0] node4095;
	wire [14-1:0] node4096;
	wire [14-1:0] node4101;
	wire [14-1:0] node4102;
	wire [14-1:0] node4103;
	wire [14-1:0] node4104;
	wire [14-1:0] node4107;
	wire [14-1:0] node4116;
	wire [14-1:0] node4117;
	wire [14-1:0] node4118;
	wire [14-1:0] node4119;
	wire [14-1:0] node4120;
	wire [14-1:0] node4121;
	wire [14-1:0] node4123;
	wire [14-1:0] node4125;
	wire [14-1:0] node4128;
	wire [14-1:0] node4129;
	wire [14-1:0] node4130;
	wire [14-1:0] node4138;
	wire [14-1:0] node4139;
	wire [14-1:0] node4140;
	wire [14-1:0] node4141;
	wire [14-1:0] node4142;
	wire [14-1:0] node4143;
	wire [14-1:0] node4145;
	wire [14-1:0] node4152;
	wire [14-1:0] node4153;
	wire [14-1:0] node4154;
	wire [14-1:0] node4155;
	wire [14-1:0] node4156;
	wire [14-1:0] node4157;
	wire [14-1:0] node4164;
	wire [14-1:0] node4166;
	wire [14-1:0] node4168;
	wire [14-1:0] node4170;
	wire [14-1:0] node4171;
	wire [14-1:0] node4174;

	assign outp = (inp[13]) ? node2096 : node1;
		assign node1 = (inp[8]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[11]) ? node1475 : node4;
				assign node4 = (inp[7]) ? node1048 : node5;
					assign node5 = (inp[12]) ? node623 : node6;
						assign node6 = (inp[2]) ? node330 : node7;
							assign node7 = (inp[6]) ? node203 : node8;
								assign node8 = (inp[5]) ? node102 : node9;
									assign node9 = (inp[4]) ? node47 : node10;
										assign node10 = (inp[10]) ? node18 : node11;
											assign node11 = (inp[3]) ? 14'b00000000000001 : node12;
												assign node12 = (inp[0]) ? 14'b00000000000001 : node13;
													assign node13 = (inp[9]) ? 14'b00000000000001 : 14'b10000000001000;
											assign node18 = (inp[9]) ? node32 : node19;
												assign node19 = (inp[3]) ? node25 : node20;
													assign node20 = (inp[0]) ? 14'b01111110100010 : node21;
														assign node21 = (inp[1]) ? 14'b01111010000010 : 14'b00000000000001;
													assign node25 = (inp[0]) ? node29 : node26;
														assign node26 = (inp[1]) ? 14'b01111010110010 : 14'b01111110110010;
														assign node29 = (inp[1]) ? 14'b01101010100010 : 14'b01101110100010;
												assign node32 = (inp[0]) ? node40 : node33;
													assign node33 = (inp[3]) ? node37 : node34;
														assign node34 = (inp[1]) ? 14'b01101000000010 : 14'b01101100000010;
														assign node37 = (inp[1]) ? 14'b01111010010010 : 14'b01111110010010;
													assign node40 = (inp[3]) ? node44 : node41;
														assign node41 = (inp[1]) ? 14'b00000000000001 : 14'b01111110000010;
														assign node44 = (inp[1]) ? 14'b01101010000010 : 14'b00000000000001;
										assign node47 = (inp[10]) ? node71 : node48;
											assign node48 = (inp[3]) ? node62 : node49;
												assign node49 = (inp[9]) ? node57 : node50;
													assign node50 = (inp[0]) ? node54 : node51;
														assign node51 = (inp[1]) ? 14'b01111010000110 : 14'b00000000000001;
														assign node54 = (inp[1]) ? 14'b01111010100110 : 14'b01111110100110;
													assign node57 = (inp[1]) ? 14'b00000000000001 : node58;
														assign node58 = (inp[0]) ? 14'b01111110000110 : 14'b01101100000110;
												assign node62 = (inp[0]) ? node68 : node63;
													assign node63 = (inp[9]) ? 14'b01111110010110 : node64;
														assign node64 = (inp[1]) ? 14'b01111010110110 : 14'b01111110110110;
													assign node68 = (inp[9]) ? 14'b01101010000110 : 14'b01101110100110;
											assign node71 = (inp[9]) ? node87 : node72;
												assign node72 = (inp[3]) ? node80 : node73;
													assign node73 = (inp[0]) ? node77 : node74;
														assign node74 = (inp[1]) ? 14'b01111010000000 : 14'b00000000000001;
														assign node77 = (inp[1]) ? 14'b01111010100000 : 14'b01111110100000;
													assign node80 = (inp[0]) ? node84 : node81;
														assign node81 = (inp[1]) ? 14'b01111010110000 : 14'b01111110110000;
														assign node84 = (inp[1]) ? 14'b01101010100000 : 14'b01101110100000;
												assign node87 = (inp[0]) ? node95 : node88;
													assign node88 = (inp[3]) ? node92 : node89;
														assign node89 = (inp[1]) ? 14'b01101000000000 : 14'b01101100000000;
														assign node92 = (inp[1]) ? 14'b01111010010000 : 14'b01111110010000;
													assign node95 = (inp[1]) ? node99 : node96;
														assign node96 = (inp[3]) ? 14'b00000000000001 : 14'b01111110000000;
														assign node99 = (inp[3]) ? 14'b01101010000000 : 14'b00000000000001;
									assign node102 = (inp[9]) ? node154 : node103;
										assign node103 = (inp[1]) ? node125 : node104;
											assign node104 = (inp[0]) ? node112 : node105;
												assign node105 = (inp[3]) ? node107 : 14'b00000000000001;
													assign node107 = (inp[10]) ? node109 : 14'b01110110110110;
														assign node109 = (inp[4]) ? 14'b01110110110000 : 14'b01110110110010;
												assign node112 = (inp[3]) ? node120 : node113;
													assign node113 = (inp[4]) ? node117 : node114;
														assign node114 = (inp[10]) ? 14'b01110110100010 : 14'b00110110100010;
														assign node117 = (inp[10]) ? 14'b01110110100000 : 14'b01110110100110;
													assign node120 = (inp[10]) ? 14'b01100110100000 : node121;
														assign node121 = (inp[4]) ? 14'b01100110100110 : 14'b00100110100010;
											assign node125 = (inp[3]) ? node141 : node126;
												assign node126 = (inp[0]) ? node134 : node127;
													assign node127 = (inp[4]) ? node131 : node128;
														assign node128 = (inp[10]) ? 14'b01110010000010 : 14'b00110010000010;
														assign node131 = (inp[10]) ? 14'b01110010000000 : 14'b01110010000110;
													assign node134 = (inp[4]) ? node138 : node135;
														assign node135 = (inp[10]) ? 14'b01110010100010 : 14'b00110010100010;
														assign node138 = (inp[10]) ? 14'b01110010100000 : 14'b01110010100110;
												assign node141 = (inp[0]) ? node149 : node142;
													assign node142 = (inp[10]) ? node146 : node143;
														assign node143 = (inp[4]) ? 14'b01110010110110 : 14'b00110010110010;
														assign node146 = (inp[4]) ? 14'b01110010110000 : 14'b01110010110010;
													assign node149 = (inp[10]) ? node151 : 14'b01100010100110;
														assign node151 = (inp[4]) ? 14'b01100010100000 : 14'b01100010100010;
										assign node154 = (inp[0]) ? node186 : node155;
											assign node155 = (inp[3]) ? node171 : node156;
												assign node156 = (inp[1]) ? node164 : node157;
													assign node157 = (inp[10]) ? node161 : node158;
														assign node158 = (inp[4]) ? 14'b01100100000110 : 14'b00100100000010;
														assign node161 = (inp[4]) ? 14'b01100100000000 : 14'b01100100000010;
													assign node164 = (inp[10]) ? node168 : node165;
														assign node165 = (inp[4]) ? 14'b01100000000110 : 14'b00100000000010;
														assign node168 = (inp[4]) ? 14'b01100000000000 : 14'b01100000000010;
												assign node171 = (inp[1]) ? node179 : node172;
													assign node172 = (inp[4]) ? node176 : node173;
														assign node173 = (inp[10]) ? 14'b01110110010010 : 14'b00110110010010;
														assign node176 = (inp[10]) ? 14'b01110110010000 : 14'b01110110010110;
													assign node179 = (inp[10]) ? node183 : node180;
														assign node180 = (inp[4]) ? 14'b01110010010110 : 14'b00110010010010;
														assign node183 = (inp[4]) ? 14'b01110010010000 : 14'b01110010010010;
											assign node186 = (inp[1]) ? node196 : node187;
												assign node187 = (inp[3]) ? 14'b00000000000001 : node188;
													assign node188 = (inp[4]) ? node192 : node189;
														assign node189 = (inp[10]) ? 14'b01110110000010 : 14'b00110110000010;
														assign node192 = (inp[10]) ? 14'b01110110000000 : 14'b01110110000110;
												assign node196 = (inp[3]) ? node198 : 14'b00000000000001;
													assign node198 = (inp[4]) ? 14'b01100010000110 : node199;
														assign node199 = (inp[10]) ? 14'b01100010000010 : 14'b00100010000010;
								assign node203 = (inp[3]) ? node295 : node204;
									assign node204 = (inp[1]) ? node254 : node205;
										assign node205 = (inp[5]) ? node225 : node206;
											assign node206 = (inp[10]) ? node212 : node207;
												assign node207 = (inp[4]) ? node209 : 14'b00000000000001;
													assign node209 = (inp[9]) ? 14'b01111100010110 : 14'b01111100110110;
												assign node212 = (inp[9]) ? node218 : node213;
													assign node213 = (inp[4]) ? 14'b01111100110000 : node214;
														assign node214 = (inp[0]) ? 14'b01111100100010 : 14'b01111100110010;
													assign node218 = (inp[4]) ? node222 : node219;
														assign node219 = (inp[0]) ? 14'b01111100000010 : 14'b01111100010010;
														assign node222 = (inp[0]) ? 14'b01111100000000 : 14'b01111100010000;
											assign node225 = (inp[0]) ? node239 : node226;
												assign node226 = (inp[9]) ? node234 : node227;
													assign node227 = (inp[10]) ? node231 : node228;
														assign node228 = (inp[4]) ? 14'b01110100110110 : 14'b00110100110010;
														assign node231 = (inp[4]) ? 14'b01110100110000 : 14'b01110100110010;
													assign node234 = (inp[4]) ? 14'b01110100010110 : node235;
														assign node235 = (inp[10]) ? 14'b01110100010010 : 14'b00110100010010;
												assign node239 = (inp[9]) ? node247 : node240;
													assign node240 = (inp[4]) ? node244 : node241;
														assign node241 = (inp[10]) ? 14'b01110100100010 : 14'b00110100100010;
														assign node244 = (inp[10]) ? 14'b01110100100000 : 14'b01110100100110;
													assign node247 = (inp[10]) ? node251 : node248;
														assign node248 = (inp[4]) ? 14'b01110100000110 : 14'b00110100000010;
														assign node251 = (inp[4]) ? 14'b01110100000000 : 14'b01110100000010;
										assign node254 = (inp[0]) ? node280 : node255;
											assign node255 = (inp[10]) ? node267 : node256;
												assign node256 = (inp[4]) ? node260 : node257;
													assign node257 = (inp[5]) ? 14'b00110000110010 : 14'b00000000000001;
													assign node260 = (inp[5]) ? node264 : node261;
														assign node261 = (inp[9]) ? 14'b01111000010110 : 14'b01111000110110;
														assign node264 = (inp[9]) ? 14'b01110000010110 : 14'b01110000110110;
												assign node267 = (inp[5]) ? node275 : node268;
													assign node268 = (inp[9]) ? node272 : node269;
														assign node269 = (inp[4]) ? 14'b01111000110000 : 14'b01111000110010;
														assign node272 = (inp[4]) ? 14'b01111000010000 : 14'b01111000010010;
													assign node275 = (inp[9]) ? 14'b01110000010000 : node276;
														assign node276 = (inp[4]) ? 14'b01110000110000 : 14'b01110000110010;
											assign node280 = (inp[9]) ? node282 : 14'b00000000000001;
												assign node282 = (inp[10]) ? node288 : node283;
													assign node283 = (inp[5]) ? node285 : 14'b00000000000001;
														assign node285 = (inp[4]) ? 14'b01110000000110 : 14'b00110000000010;
													assign node288 = (inp[4]) ? node292 : node289;
														assign node289 = (inp[5]) ? 14'b01110000000010 : 14'b01111000000010;
														assign node292 = (inp[5]) ? 14'b01110000000000 : 14'b01111000000000;
									assign node295 = (inp[9]) ? 14'b00000000000001 : node296;
										assign node296 = (inp[0]) ? node312 : node297;
											assign node297 = (inp[1]) ? node299 : 14'b00000000000001;
												assign node299 = (inp[5]) ? node305 : node300;
													assign node300 = (inp[10]) ? node302 : 14'b01111000100110;
														assign node302 = (inp[4]) ? 14'b01111000100000 : 14'b01111000100010;
													assign node305 = (inp[10]) ? node309 : node306;
														assign node306 = (inp[4]) ? 14'b01110000100110 : 14'b00110000100010;
														assign node309 = (inp[4]) ? 14'b01110000100000 : 14'b01110000100010;
											assign node312 = (inp[1]) ? 14'b00000000000001 : node313;
												assign node313 = (inp[4]) ? node321 : node314;
													assign node314 = (inp[10]) ? node318 : node315;
														assign node315 = (inp[5]) ? 14'b00100110000010 : 14'b00000000000001;
														assign node318 = (inp[5]) ? 14'b01100110000010 : 14'b01101110000010;
													assign node321 = (inp[10]) ? node325 : node322;
														assign node322 = (inp[5]) ? 14'b01100110000110 : 14'b01101110000110;
														assign node325 = (inp[5]) ? 14'b01100110000000 : 14'b01101110000000;
							assign node330 = (inp[10]) ? node516 : node331;
								assign node331 = (inp[4]) ? node423 : node332;
									assign node332 = (inp[9]) ? node382 : node333;
										assign node333 = (inp[6]) ? node357 : node334;
											assign node334 = (inp[0]) ? node344 : node335;
												assign node335 = (inp[3]) ? node337 : 14'b00000000000001;
													assign node337 = (inp[5]) ? node341 : node338;
														assign node338 = (inp[1]) ? 14'b00011010110000 : 14'b00011110110000;
														assign node341 = (inp[1]) ? 14'b00010010110000 : 14'b00010110110000;
												assign node344 = (inp[3]) ? node352 : node345;
													assign node345 = (inp[1]) ? node349 : node346;
														assign node346 = (inp[5]) ? 14'b00010110100000 : 14'b00011110100000;
														assign node349 = (inp[5]) ? 14'b00010010100000 : 14'b00011010100000;
													assign node352 = (inp[1]) ? 14'b00000010100000 : node353;
														assign node353 = (inp[5]) ? 14'b00000110100000 : 14'b00001110100000;
											assign node357 = (inp[3]) ? node371 : node358;
												assign node358 = (inp[0]) ? node366 : node359;
													assign node359 = (inp[5]) ? node363 : node360;
														assign node360 = (inp[1]) ? 14'b00011000110000 : 14'b00011100110000;
														assign node363 = (inp[1]) ? 14'b00010000110000 : 14'b00010100110000;
													assign node366 = (inp[1]) ? 14'b00000000000001 : node367;
														assign node367 = (inp[5]) ? 14'b00010100100000 : 14'b00011100100000;
												assign node371 = (inp[0]) ? node377 : node372;
													assign node372 = (inp[1]) ? node374 : 14'b00000000000001;
														assign node374 = (inp[5]) ? 14'b00010000100000 : 14'b00011000100000;
													assign node377 = (inp[1]) ? 14'b00000000000001 : node378;
														assign node378 = (inp[5]) ? 14'b00000110000000 : 14'b00001110000000;
										assign node382 = (inp[3]) ? node410 : node383;
											assign node383 = (inp[1]) ? node399 : node384;
												assign node384 = (inp[5]) ? node392 : node385;
													assign node385 = (inp[6]) ? node389 : node386;
														assign node386 = (inp[0]) ? 14'b00011110000000 : 14'b00001100000000;
														assign node389 = (inp[0]) ? 14'b00011100000000 : 14'b00011100010000;
													assign node392 = (inp[0]) ? node396 : node393;
														assign node393 = (inp[6]) ? 14'b00010100010000 : 14'b00000100000000;
														assign node396 = (inp[6]) ? 14'b00010100000000 : 14'b00010110000000;
												assign node399 = (inp[6]) ? node405 : node400;
													assign node400 = (inp[0]) ? 14'b00000000000001 : node401;
														assign node401 = (inp[5]) ? 14'b00000000000000 : 14'b00001000000000;
													assign node405 = (inp[0]) ? 14'b00011000000000 : node406;
														assign node406 = (inp[5]) ? 14'b00010000010000 : 14'b00011000010000;
											assign node410 = (inp[6]) ? 14'b00000000000001 : node411;
												assign node411 = (inp[0]) ? node419 : node412;
													assign node412 = (inp[1]) ? node416 : node413;
														assign node413 = (inp[5]) ? 14'b00010110010000 : 14'b00011110010000;
														assign node416 = (inp[5]) ? 14'b00010010010000 : 14'b00011010010000;
													assign node419 = (inp[1]) ? 14'b00000010000000 : 14'b00000000000001;
									assign node423 = (inp[6]) ? node477 : node424;
										assign node424 = (inp[9]) ? node452 : node425;
											assign node425 = (inp[3]) ? node439 : node426;
												assign node426 = (inp[0]) ? node432 : node427;
													assign node427 = (inp[1]) ? node429 : 14'b00000000000001;
														assign node429 = (inp[5]) ? 14'b00110010000110 : 14'b00111010000110;
													assign node432 = (inp[1]) ? node436 : node433;
														assign node433 = (inp[5]) ? 14'b00110110100110 : 14'b00111110100110;
														assign node436 = (inp[5]) ? 14'b00110010100110 : 14'b00111010100110;
												assign node439 = (inp[0]) ? node447 : node440;
													assign node440 = (inp[5]) ? node444 : node441;
														assign node441 = (inp[1]) ? 14'b00111010110110 : 14'b00111110110110;
														assign node444 = (inp[1]) ? 14'b00110010110110 : 14'b00110110110110;
													assign node447 = (inp[1]) ? 14'b00101010100110 : node448;
														assign node448 = (inp[5]) ? 14'b00100110100110 : 14'b00101110100110;
											assign node452 = (inp[0]) ? node468 : node453;
												assign node453 = (inp[3]) ? node461 : node454;
													assign node454 = (inp[5]) ? node458 : node455;
														assign node455 = (inp[1]) ? 14'b00101000000110 : 14'b00101100000110;
														assign node458 = (inp[1]) ? 14'b00100000000110 : 14'b00100100000110;
													assign node461 = (inp[1]) ? node465 : node462;
														assign node462 = (inp[5]) ? 14'b00110110010110 : 14'b00111110010110;
														assign node465 = (inp[5]) ? 14'b00110010010110 : 14'b00111010010110;
												assign node468 = (inp[3]) ? node472 : node469;
													assign node469 = (inp[1]) ? 14'b00000000000001 : 14'b00110110000110;
													assign node472 = (inp[1]) ? node474 : 14'b00000000000001;
														assign node474 = (inp[5]) ? 14'b00100010000110 : 14'b00101010000110;
										assign node477 = (inp[3]) ? node505 : node478;
											assign node478 = (inp[1]) ? node494 : node479;
												assign node479 = (inp[0]) ? node487 : node480;
													assign node480 = (inp[9]) ? node484 : node481;
														assign node481 = (inp[5]) ? 14'b00110100110110 : 14'b00111100110110;
														assign node484 = (inp[5]) ? 14'b00110100010110 : 14'b00111100010110;
													assign node487 = (inp[5]) ? node491 : node488;
														assign node488 = (inp[9]) ? 14'b00111100000110 : 14'b00111100100110;
														assign node491 = (inp[9]) ? 14'b00110100000110 : 14'b00110100100110;
												assign node494 = (inp[0]) ? node502 : node495;
													assign node495 = (inp[5]) ? node499 : node496;
														assign node496 = (inp[9]) ? 14'b00111000010110 : 14'b00111000110110;
														assign node499 = (inp[9]) ? 14'b00110000010110 : 14'b00110000110110;
													assign node502 = (inp[9]) ? 14'b00110000000110 : 14'b00000000000001;
											assign node505 = (inp[9]) ? 14'b00000000000001 : node506;
												assign node506 = (inp[1]) ? node512 : node507;
													assign node507 = (inp[0]) ? node509 : 14'b00000000000001;
														assign node509 = (inp[5]) ? 14'b00100110000110 : 14'b00101110000110;
													assign node512 = (inp[0]) ? 14'b00000000000001 : 14'b00110000100110;
								assign node516 = (inp[4]) ? node570 : node517;
									assign node517 = (inp[5]) ? 14'b00000000000001 : node518;
										assign node518 = (inp[1]) ? node544 : node519;
											assign node519 = (inp[3]) ? node535 : node520;
												assign node520 = (inp[6]) ? node528 : node521;
													assign node521 = (inp[0]) ? node525 : node522;
														assign node522 = (inp[9]) ? 14'b00101100000010 : 14'b00000000000001;
														assign node525 = (inp[9]) ? 14'b00111110000010 : 14'b00111110100010;
													assign node528 = (inp[0]) ? node532 : node529;
														assign node529 = (inp[9]) ? 14'b00111100010010 : 14'b00111100110010;
														assign node532 = (inp[9]) ? 14'b00111100000010 : 14'b00111100100010;
												assign node535 = (inp[9]) ? 14'b00000000000001 : node536;
													assign node536 = (inp[6]) ? node540 : node537;
														assign node537 = (inp[0]) ? 14'b00101110100010 : 14'b00111110110010;
														assign node540 = (inp[0]) ? 14'b00101110000010 : 14'b00000000000001;
											assign node544 = (inp[6]) ? node560 : node545;
												assign node545 = (inp[9]) ? node553 : node546;
													assign node546 = (inp[0]) ? node550 : node547;
														assign node547 = (inp[3]) ? 14'b00111010110010 : 14'b00111010000010;
														assign node550 = (inp[3]) ? 14'b00101010100010 : 14'b00111010100010;
													assign node553 = (inp[3]) ? node557 : node554;
														assign node554 = (inp[0]) ? 14'b00000000000001 : 14'b00101000000010;
														assign node557 = (inp[0]) ? 14'b00101010000010 : 14'b00111010010010;
												assign node560 = (inp[3]) ? 14'b00000000000001 : node561;
													assign node561 = (inp[0]) ? node565 : node562;
														assign node562 = (inp[9]) ? 14'b00111000010010 : 14'b00111000110010;
														assign node565 = (inp[9]) ? 14'b00111000000010 : 14'b00000000000001;
									assign node570 = (inp[5]) ? node572 : 14'b00000000000001;
										assign node572 = (inp[6]) ? node600 : node573;
											assign node573 = (inp[1]) ? node587 : node574;
												assign node574 = (inp[0]) ? node580 : node575;
													assign node575 = (inp[9]) ? node577 : 14'b00000000000001;
														assign node577 = (inp[3]) ? 14'b00110110010000 : 14'b00100100000000;
													assign node580 = (inp[9]) ? node584 : node581;
														assign node581 = (inp[3]) ? 14'b00100110100000 : 14'b00110110100000;
														assign node584 = (inp[3]) ? 14'b00000000000001 : 14'b00110110000000;
												assign node587 = (inp[3]) ? node593 : node588;
													assign node588 = (inp[0]) ? 14'b00000000000001 : node589;
														assign node589 = (inp[9]) ? 14'b00100000000000 : 14'b00110010000000;
													assign node593 = (inp[0]) ? node597 : node594;
														assign node594 = (inp[9]) ? 14'b00110010010000 : 14'b00110010110000;
														assign node597 = (inp[9]) ? 14'b00100010000000 : 14'b00100010100000;
											assign node600 = (inp[3]) ? node614 : node601;
												assign node601 = (inp[0]) ? node607 : node602;
													assign node602 = (inp[1]) ? node604 : 14'b00110100110000;
														assign node604 = (inp[9]) ? 14'b00110000010000 : 14'b00110000110000;
													assign node607 = (inp[1]) ? node611 : node608;
														assign node608 = (inp[9]) ? 14'b00110100000000 : 14'b00110100100000;
														assign node611 = (inp[9]) ? 14'b00110000000000 : 14'b00000000000001;
												assign node614 = (inp[9]) ? 14'b00000000000001 : node615;
													assign node615 = (inp[1]) ? node619 : node616;
														assign node616 = (inp[0]) ? 14'b00100110000000 : 14'b00000000000001;
														assign node619 = (inp[0]) ? 14'b00000000000001 : 14'b00110000100000;
						assign node623 = (inp[4]) ? node933 : node624;
							assign node624 = (inp[10]) ? node792 : node625;
								assign node625 = (inp[6]) ? node723 : node626;
									assign node626 = (inp[9]) ? node678 : node627;
										assign node627 = (inp[3]) ? node649 : node628;
											assign node628 = (inp[1]) ? node634 : node629;
												assign node629 = (inp[0]) ? node631 : 14'b00000000000001;
													assign node631 = (inp[2]) ? 14'b00010110100110 : 14'b01010110100110;
												assign node634 = (inp[2]) ? node642 : node635;
													assign node635 = (inp[5]) ? node639 : node636;
														assign node636 = (inp[0]) ? 14'b01011010100110 : 14'b01011010000110;
														assign node639 = (inp[0]) ? 14'b01010010100110 : 14'b01010010000110;
													assign node642 = (inp[0]) ? node646 : node643;
														assign node643 = (inp[5]) ? 14'b00010010000110 : 14'b00011010000110;
														assign node646 = (inp[5]) ? 14'b00010010100110 : 14'b00011010100110;
											assign node649 = (inp[0]) ? node663 : node650;
												assign node650 = (inp[5]) ? node656 : node651;
													assign node651 = (inp[1]) ? node653 : 14'b01011110110110;
														assign node653 = (inp[2]) ? 14'b00011010110110 : 14'b01011010110110;
													assign node656 = (inp[1]) ? node660 : node657;
														assign node657 = (inp[2]) ? 14'b00010110110110 : 14'b01010110110110;
														assign node660 = (inp[2]) ? 14'b00010010110110 : 14'b01010010110110;
												assign node663 = (inp[2]) ? node671 : node664;
													assign node664 = (inp[1]) ? node668 : node665;
														assign node665 = (inp[5]) ? 14'b01000110100110 : 14'b01001110100110;
														assign node668 = (inp[5]) ? 14'b01000010100110 : 14'b01001010100110;
													assign node671 = (inp[1]) ? node675 : node672;
														assign node672 = (inp[5]) ? 14'b00000110100110 : 14'b00001110100110;
														assign node675 = (inp[5]) ? 14'b00000010100110 : 14'b00001010100110;
										assign node678 = (inp[0]) ? node704 : node679;
											assign node679 = (inp[3]) ? node693 : node680;
												assign node680 = (inp[5]) ? node686 : node681;
													assign node681 = (inp[2]) ? node683 : 14'b01001000000110;
														assign node683 = (inp[1]) ? 14'b00001000000110 : 14'b00001100000110;
													assign node686 = (inp[2]) ? node690 : node687;
														assign node687 = (inp[1]) ? 14'b01000000000110 : 14'b01000100000110;
														assign node690 = (inp[1]) ? 14'b00000000000110 : 14'b00000100000110;
												assign node693 = (inp[1]) ? node697 : node694;
													assign node694 = (inp[2]) ? 14'b00010110010110 : 14'b01010110010110;
													assign node697 = (inp[2]) ? node701 : node698;
														assign node698 = (inp[5]) ? 14'b01010010010110 : 14'b01011010010110;
														assign node701 = (inp[5]) ? 14'b00010010010110 : 14'b00011010010110;
											assign node704 = (inp[1]) ? node714 : node705;
												assign node705 = (inp[3]) ? 14'b00000000000001 : node706;
													assign node706 = (inp[5]) ? node710 : node707;
														assign node707 = (inp[2]) ? 14'b00011110000110 : 14'b01011110000110;
														assign node710 = (inp[2]) ? 14'b00010110000110 : 14'b01010110000110;
												assign node714 = (inp[3]) ? node716 : 14'b00000000000001;
													assign node716 = (inp[2]) ? node720 : node717;
														assign node717 = (inp[5]) ? 14'b01000010000110 : 14'b01001010000110;
														assign node720 = (inp[5]) ? 14'b00000010000110 : 14'b00001010000110;
									assign node723 = (inp[3]) ? node773 : node724;
										assign node724 = (inp[0]) ? node752 : node725;
											assign node725 = (inp[1]) ? node739 : node726;
												assign node726 = (inp[9]) ? node734 : node727;
													assign node727 = (inp[5]) ? node731 : node728;
														assign node728 = (inp[2]) ? 14'b00011100110110 : 14'b01011100110110;
														assign node731 = (inp[2]) ? 14'b00010100110110 : 14'b01010100110110;
													assign node734 = (inp[5]) ? node736 : 14'b01011100010110;
														assign node736 = (inp[2]) ? 14'b00010100010110 : 14'b01010100010110;
												assign node739 = (inp[5]) ? node747 : node740;
													assign node740 = (inp[2]) ? node744 : node741;
														assign node741 = (inp[9]) ? 14'b01011000010110 : 14'b01011000110110;
														assign node744 = (inp[9]) ? 14'b00011000010110 : 14'b00011000110110;
													assign node747 = (inp[2]) ? 14'b00010000110110 : node748;
														assign node748 = (inp[9]) ? 14'b01010000010110 : 14'b01010000110110;
											assign node752 = (inp[1]) ? node768 : node753;
												assign node753 = (inp[9]) ? node761 : node754;
													assign node754 = (inp[5]) ? node758 : node755;
														assign node755 = (inp[2]) ? 14'b00011100100110 : 14'b01011100100110;
														assign node758 = (inp[2]) ? 14'b00010100100110 : 14'b01010100100110;
													assign node761 = (inp[5]) ? node765 : node762;
														assign node762 = (inp[2]) ? 14'b00011100000110 : 14'b01011100000110;
														assign node765 = (inp[2]) ? 14'b00010100000110 : 14'b01010100000110;
												assign node768 = (inp[9]) ? node770 : 14'b00000000000001;
													assign node770 = (inp[5]) ? 14'b00010000000110 : 14'b00011000000110;
										assign node773 = (inp[9]) ? 14'b00000000000001 : node774;
											assign node774 = (inp[0]) ? node784 : node775;
												assign node775 = (inp[1]) ? node777 : 14'b00000000000001;
													assign node777 = (inp[2]) ? node781 : node778;
														assign node778 = (inp[5]) ? 14'b01010000100110 : 14'b01011000100110;
														assign node781 = (inp[5]) ? 14'b00010000100110 : 14'b00011000100110;
												assign node784 = (inp[1]) ? 14'b00000000000001 : node785;
													assign node785 = (inp[2]) ? node787 : 14'b01001110000110;
														assign node787 = (inp[5]) ? 14'b00000110000110 : 14'b00001110000110;
								assign node792 = (inp[5]) ? node882 : node793;
									assign node793 = (inp[6]) ? node843 : node794;
										assign node794 = (inp[9]) ? node822 : node795;
											assign node795 = (inp[1]) ? node807 : node796;
												assign node796 = (inp[3]) ? node802 : node797;
													assign node797 = (inp[0]) ? node799 : 14'b00000000000001;
														assign node799 = (inp[2]) ? 14'b00011110100010 : 14'b01011110100010;
													assign node802 = (inp[0]) ? 14'b00001110100010 : node803;
														assign node803 = (inp[2]) ? 14'b00011110110010 : 14'b01011110110010;
												assign node807 = (inp[2]) ? node815 : node808;
													assign node808 = (inp[0]) ? node812 : node809;
														assign node809 = (inp[3]) ? 14'b01011010110010 : 14'b01011010000010;
														assign node812 = (inp[3]) ? 14'b01001010100010 : 14'b01011010100010;
													assign node815 = (inp[3]) ? node819 : node816;
														assign node816 = (inp[0]) ? 14'b00011010100010 : 14'b00011010000010;
														assign node819 = (inp[0]) ? 14'b00001010100010 : 14'b00011010110010;
											assign node822 = (inp[0]) ? node836 : node823;
												assign node823 = (inp[3]) ? node829 : node824;
													assign node824 = (inp[1]) ? node826 : 14'b01001100000010;
														assign node826 = (inp[2]) ? 14'b00001000000010 : 14'b01001000000010;
													assign node829 = (inp[2]) ? node833 : node830;
														assign node830 = (inp[1]) ? 14'b01011010010010 : 14'b01011110010010;
														assign node833 = (inp[1]) ? 14'b00011010010010 : 14'b00011110010010;
												assign node836 = (inp[3]) ? node840 : node837;
													assign node837 = (inp[1]) ? 14'b00000000000001 : 14'b01011110000010;
													assign node840 = (inp[1]) ? 14'b00001010000010 : 14'b00000000000001;
										assign node843 = (inp[3]) ? node869 : node844;
											assign node844 = (inp[0]) ? node856 : node845;
												assign node845 = (inp[2]) ? node853 : node846;
													assign node846 = (inp[9]) ? node850 : node847;
														assign node847 = (inp[1]) ? 14'b01011000110010 : 14'b01011100110010;
														assign node850 = (inp[1]) ? 14'b01011000010010 : 14'b01011100010010;
													assign node853 = (inp[1]) ? 14'b00011000110010 : 14'b00011100110010;
												assign node856 = (inp[1]) ? node864 : node857;
													assign node857 = (inp[9]) ? node861 : node858;
														assign node858 = (inp[2]) ? 14'b00011100100010 : 14'b01011100100010;
														assign node861 = (inp[2]) ? 14'b00011100000010 : 14'b01011100000010;
													assign node864 = (inp[9]) ? node866 : 14'b00000000000001;
														assign node866 = (inp[2]) ? 14'b00011000000010 : 14'b01011000000010;
											assign node869 = (inp[9]) ? 14'b00000000000001 : node870;
												assign node870 = (inp[0]) ? node876 : node871;
													assign node871 = (inp[1]) ? node873 : 14'b00000000000001;
														assign node873 = (inp[2]) ? 14'b00011000100010 : 14'b01011000100010;
													assign node876 = (inp[1]) ? 14'b00000000000001 : node877;
														assign node877 = (inp[2]) ? 14'b00001110000010 : 14'b01001110000010;
									assign node882 = (inp[2]) ? node884 : 14'b00000000000001;
										assign node884 = (inp[9]) ? node914 : node885;
											assign node885 = (inp[6]) ? node899 : node886;
												assign node886 = (inp[3]) ? node894 : node887;
													assign node887 = (inp[0]) ? node891 : node888;
														assign node888 = (inp[1]) ? 14'b00010010000010 : 14'b00000000000001;
														assign node891 = (inp[1]) ? 14'b00010010100010 : 14'b00010110100010;
													assign node894 = (inp[0]) ? 14'b00000010100010 : node895;
														assign node895 = (inp[1]) ? 14'b00010010110010 : 14'b00010110110010;
												assign node899 = (inp[3]) ? node907 : node900;
													assign node900 = (inp[1]) ? node904 : node901;
														assign node901 = (inp[0]) ? 14'b00010100100010 : 14'b00010100110010;
														assign node904 = (inp[0]) ? 14'b00000000000001 : 14'b00010000110010;
													assign node907 = (inp[1]) ? node911 : node908;
														assign node908 = (inp[0]) ? 14'b00000110000010 : 14'b00000000000001;
														assign node911 = (inp[0]) ? 14'b00000000000001 : 14'b00010000100010;
											assign node914 = (inp[3]) ? node924 : node915;
												assign node915 = (inp[6]) ? node919 : node916;
													assign node916 = (inp[0]) ? 14'b00000000000001 : 14'b00000000000010;
													assign node919 = (inp[0]) ? node921 : 14'b00010000010010;
														assign node921 = (inp[1]) ? 14'b00010000000010 : 14'b00010100000010;
												assign node924 = (inp[6]) ? 14'b00000000000001 : node925;
													assign node925 = (inp[0]) ? node929 : node926;
														assign node926 = (inp[1]) ? 14'b00010010010010 : 14'b00010110010010;
														assign node929 = (inp[1]) ? 14'b00000010000010 : 14'b00000000000001;
							assign node933 = (inp[2]) ? 14'b00000000000001 : node934;
								assign node934 = (inp[5]) ? node988 : node935;
									assign node935 = (inp[10]) ? node937 : 14'b00000000000001;
										assign node937 = (inp[1]) ? node961 : node938;
											assign node938 = (inp[0]) ? node952 : node939;
												assign node939 = (inp[6]) ? node947 : node940;
													assign node940 = (inp[3]) ? node944 : node941;
														assign node941 = (inp[9]) ? 14'b00101100000000 : 14'b00000000000001;
														assign node944 = (inp[9]) ? 14'b00111110010000 : 14'b00111110110000;
													assign node947 = (inp[3]) ? 14'b00000000000001 : node948;
														assign node948 = (inp[9]) ? 14'b00111100010000 : 14'b00111100110000;
												assign node952 = (inp[3]) ? node958 : node953;
													assign node953 = (inp[6]) ? node955 : 14'b00111110000000;
														assign node955 = (inp[9]) ? 14'b00111100000000 : 14'b00111100100000;
													assign node958 = (inp[6]) ? 14'b00101110000000 : 14'b00101110100000;
											assign node961 = (inp[9]) ? node975 : node962;
												assign node962 = (inp[6]) ? node970 : node963;
													assign node963 = (inp[3]) ? node967 : node964;
														assign node964 = (inp[0]) ? 14'b00111010100000 : 14'b00111010000000;
														assign node967 = (inp[0]) ? 14'b00101010100000 : 14'b00111010110000;
													assign node970 = (inp[0]) ? 14'b00000000000001 : node971;
														assign node971 = (inp[3]) ? 14'b00111000100000 : 14'b00111000110000;
												assign node975 = (inp[6]) ? node983 : node976;
													assign node976 = (inp[3]) ? node980 : node977;
														assign node977 = (inp[0]) ? 14'b00000000000001 : 14'b00101000000000;
														assign node980 = (inp[0]) ? 14'b00101010000000 : 14'b00111010010000;
													assign node983 = (inp[3]) ? 14'b00000000000001 : node984;
														assign node984 = (inp[0]) ? 14'b00111000000000 : 14'b00111000010000;
									assign node988 = (inp[10]) ? 14'b00000000000001 : node989;
										assign node989 = (inp[6]) ? node1021 : node990;
											assign node990 = (inp[9]) ? node1006 : node991;
												assign node991 = (inp[3]) ? node999 : node992;
													assign node992 = (inp[0]) ? node996 : node993;
														assign node993 = (inp[1]) ? 14'b01010010000010 : 14'b00000000000001;
														assign node996 = (inp[1]) ? 14'b01010010100010 : 14'b01010110100010;
													assign node999 = (inp[0]) ? node1003 : node1000;
														assign node1000 = (inp[1]) ? 14'b01010010110010 : 14'b01010110110010;
														assign node1003 = (inp[1]) ? 14'b01000010100010 : 14'b01000110100010;
												assign node1006 = (inp[0]) ? node1014 : node1007;
													assign node1007 = (inp[3]) ? node1011 : node1008;
														assign node1008 = (inp[1]) ? 14'b01000000000010 : 14'b01000100000010;
														assign node1011 = (inp[1]) ? 14'b01010010010010 : 14'b01010110010010;
													assign node1014 = (inp[3]) ? node1018 : node1015;
														assign node1015 = (inp[1]) ? 14'b00000000000001 : 14'b01010110000010;
														assign node1018 = (inp[1]) ? 14'b01000010000010 : 14'b00000000000001;
											assign node1021 = (inp[3]) ? node1037 : node1022;
												assign node1022 = (inp[1]) ? node1030 : node1023;
													assign node1023 = (inp[9]) ? node1027 : node1024;
														assign node1024 = (inp[0]) ? 14'b01010100100010 : 14'b01010100110010;
														assign node1027 = (inp[0]) ? 14'b01010100000010 : 14'b01010100010010;
													assign node1030 = (inp[0]) ? node1034 : node1031;
														assign node1031 = (inp[9]) ? 14'b01010000010010 : 14'b01010000110010;
														assign node1034 = (inp[9]) ? 14'b01010000000010 : 14'b00000000000001;
												assign node1037 = (inp[9]) ? 14'b00000000000001 : node1038;
													assign node1038 = (inp[1]) ? node1042 : node1039;
														assign node1039 = (inp[0]) ? 14'b01000110000010 : 14'b00000000000001;
														assign node1042 = (inp[0]) ? 14'b00000000000001 : 14'b01010000100010;
					assign node1048 = (inp[0]) ? 14'b00000000000001 : node1049;
						assign node1049 = (inp[3]) ? node1385 : node1050;
							assign node1050 = (inp[12]) ? node1246 : node1051;
								assign node1051 = (inp[2]) ? node1153 : node1052;
									assign node1052 = (inp[10]) ? node1096 : node1053;
										assign node1053 = (inp[4]) ? node1067 : node1054;
											assign node1054 = (inp[5]) ? node1056 : 14'b00000000000001;
												assign node1056 = (inp[9]) ? node1062 : node1057;
													assign node1057 = (inp[1]) ? node1059 : 14'b00100100110010;
														assign node1059 = (inp[6]) ? 14'b00100000110010 : 14'b00100010110010;
													assign node1062 = (inp[1]) ? node1064 : 14'b00100110010010;
														assign node1064 = (inp[6]) ? 14'b00100000010010 : 14'b00100010010010;
											assign node1067 = (inp[5]) ? node1081 : node1068;
												assign node1068 = (inp[1]) ? node1074 : node1069;
													assign node1069 = (inp[9]) ? 14'b01101100010110 : node1070;
														assign node1070 = (inp[6]) ? 14'b01101100110110 : 14'b01101110110110;
													assign node1074 = (inp[6]) ? node1078 : node1075;
														assign node1075 = (inp[9]) ? 14'b01101010010110 : 14'b01101010110110;
														assign node1078 = (inp[9]) ? 14'b01101000010110 : 14'b01101000110110;
												assign node1081 = (inp[6]) ? node1089 : node1082;
													assign node1082 = (inp[1]) ? node1086 : node1083;
														assign node1083 = (inp[9]) ? 14'b01100110010110 : 14'b01100110110110;
														assign node1086 = (inp[9]) ? 14'b01100010010110 : 14'b01100010110110;
													assign node1089 = (inp[9]) ? node1093 : node1090;
														assign node1090 = (inp[1]) ? 14'b01100000110110 : 14'b01100100110110;
														assign node1093 = (inp[1]) ? 14'b01100000010110 : 14'b01100100010110;
										assign node1096 = (inp[1]) ? node1126 : node1097;
											assign node1097 = (inp[9]) ? node1111 : node1098;
												assign node1098 = (inp[4]) ? node1106 : node1099;
													assign node1099 = (inp[6]) ? node1103 : node1100;
														assign node1100 = (inp[5]) ? 14'b01100110110010 : 14'b01101110110010;
														assign node1103 = (inp[5]) ? 14'b01100100110010 : 14'b01101100110010;
													assign node1106 = (inp[6]) ? 14'b01101100110000 : node1107;
														assign node1107 = (inp[5]) ? 14'b01100110110000 : 14'b01101110110000;
												assign node1111 = (inp[4]) ? node1119 : node1112;
													assign node1112 = (inp[5]) ? node1116 : node1113;
														assign node1113 = (inp[6]) ? 14'b01101100010010 : 14'b01101110010010;
														assign node1116 = (inp[6]) ? 14'b01100100010010 : 14'b01100110010010;
													assign node1119 = (inp[6]) ? node1123 : node1120;
														assign node1120 = (inp[5]) ? 14'b01100110010000 : 14'b01101110010000;
														assign node1123 = (inp[5]) ? 14'b01100100010000 : 14'b01101100010000;
											assign node1126 = (inp[6]) ? node1138 : node1127;
												assign node1127 = (inp[9]) ? node1131 : node1128;
													assign node1128 = (inp[4]) ? 14'b01101010110000 : 14'b01101010110010;
													assign node1131 = (inp[5]) ? node1135 : node1132;
														assign node1132 = (inp[4]) ? 14'b01101010010000 : 14'b01101010010010;
														assign node1135 = (inp[4]) ? 14'b01100010010000 : 14'b01100010010010;
												assign node1138 = (inp[9]) ? node1146 : node1139;
													assign node1139 = (inp[5]) ? node1143 : node1140;
														assign node1140 = (inp[4]) ? 14'b01101000110000 : 14'b01101000110010;
														assign node1143 = (inp[4]) ? 14'b01100000110000 : 14'b01100000110010;
													assign node1146 = (inp[4]) ? node1150 : node1147;
														assign node1147 = (inp[5]) ? 14'b01100000010010 : 14'b01101000010010;
														assign node1150 = (inp[5]) ? 14'b01100000010000 : 14'b01101000010000;
									assign node1153 = (inp[10]) ? node1213 : node1154;
										assign node1154 = (inp[4]) ? node1182 : node1155;
											assign node1155 = (inp[9]) ? node1169 : node1156;
												assign node1156 = (inp[1]) ? node1162 : node1157;
													assign node1157 = (inp[6]) ? 14'b00001100110000 : node1158;
														assign node1158 = (inp[5]) ? 14'b00000110110000 : 14'b00001110110000;
													assign node1162 = (inp[5]) ? node1166 : node1163;
														assign node1163 = (inp[6]) ? 14'b00001000110000 : 14'b00001010110000;
														assign node1166 = (inp[6]) ? 14'b00000000110000 : 14'b00000010110000;
												assign node1169 = (inp[1]) ? node1177 : node1170;
													assign node1170 = (inp[5]) ? node1174 : node1171;
														assign node1171 = (inp[6]) ? 14'b00001100010000 : 14'b00001110010000;
														assign node1174 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
													assign node1177 = (inp[6]) ? 14'b00001000010000 : node1178;
														assign node1178 = (inp[5]) ? 14'b00000010010000 : 14'b00001010010000;
											assign node1182 = (inp[9]) ? node1198 : node1183;
												assign node1183 = (inp[5]) ? node1191 : node1184;
													assign node1184 = (inp[6]) ? node1188 : node1185;
														assign node1185 = (inp[1]) ? 14'b00101010110110 : 14'b00101110110110;
														assign node1188 = (inp[1]) ? 14'b00101000110110 : 14'b00101100110110;
													assign node1191 = (inp[6]) ? node1195 : node1192;
														assign node1192 = (inp[1]) ? 14'b00100010110110 : 14'b00100110110110;
														assign node1195 = (inp[1]) ? 14'b00100000110110 : 14'b00100100110110;
												assign node1198 = (inp[6]) ? node1206 : node1199;
													assign node1199 = (inp[5]) ? node1203 : node1200;
														assign node1200 = (inp[1]) ? 14'b00101010010110 : 14'b00101110010110;
														assign node1203 = (inp[1]) ? 14'b00100010010110 : 14'b00100110010110;
													assign node1206 = (inp[5]) ? node1210 : node1207;
														assign node1207 = (inp[1]) ? 14'b00101000010110 : 14'b00101100010110;
														assign node1210 = (inp[1]) ? 14'b00100000010110 : 14'b00100100010110;
										assign node1213 = (inp[5]) ? node1229 : node1214;
											assign node1214 = (inp[4]) ? 14'b00000000000001 : node1215;
												assign node1215 = (inp[1]) ? node1221 : node1216;
													assign node1216 = (inp[9]) ? node1218 : 14'b00101100110010;
														assign node1218 = (inp[6]) ? 14'b00101100010010 : 14'b00101110010010;
													assign node1221 = (inp[9]) ? node1225 : node1222;
														assign node1222 = (inp[6]) ? 14'b00101000110010 : 14'b00101010110010;
														assign node1225 = (inp[6]) ? 14'b00101000010010 : 14'b00101010010010;
											assign node1229 = (inp[4]) ? node1231 : 14'b00000000000001;
												assign node1231 = (inp[9]) ? node1239 : node1232;
													assign node1232 = (inp[6]) ? node1236 : node1233;
														assign node1233 = (inp[1]) ? 14'b00100010110000 : 14'b00100110110000;
														assign node1236 = (inp[1]) ? 14'b00100000110000 : 14'b00100100110000;
													assign node1239 = (inp[1]) ? node1243 : node1240;
														assign node1240 = (inp[6]) ? 14'b00100100010000 : 14'b00100110010000;
														assign node1243 = (inp[6]) ? 14'b00100000010000 : 14'b00100010010000;
								assign node1246 = (inp[4]) ? node1350 : node1247;
									assign node1247 = (inp[10]) ? node1305 : node1248;
										assign node1248 = (inp[9]) ? node1280 : node1249;
											assign node1249 = (inp[2]) ? node1265 : node1250;
												assign node1250 = (inp[5]) ? node1258 : node1251;
													assign node1251 = (inp[6]) ? node1255 : node1252;
														assign node1252 = (inp[1]) ? 14'b01001010110110 : 14'b01001110110110;
														assign node1255 = (inp[1]) ? 14'b01001000110110 : 14'b01001100110110;
													assign node1258 = (inp[1]) ? node1262 : node1259;
														assign node1259 = (inp[6]) ? 14'b01000100110110 : 14'b01000110110110;
														assign node1262 = (inp[6]) ? 14'b01000000110110 : 14'b01000010110110;
												assign node1265 = (inp[1]) ? node1273 : node1266;
													assign node1266 = (inp[6]) ? node1270 : node1267;
														assign node1267 = (inp[5]) ? 14'b00000110110110 : 14'b00001110110110;
														assign node1270 = (inp[5]) ? 14'b00000100110110 : 14'b00001100110110;
													assign node1273 = (inp[5]) ? node1277 : node1274;
														assign node1274 = (inp[6]) ? 14'b00001000110110 : 14'b00001010110110;
														assign node1277 = (inp[6]) ? 14'b00000000110110 : 14'b00000010110110;
											assign node1280 = (inp[5]) ? node1294 : node1281;
												assign node1281 = (inp[6]) ? node1287 : node1282;
													assign node1282 = (inp[2]) ? node1284 : 14'b01001010010110;
														assign node1284 = (inp[1]) ? 14'b00001010010110 : 14'b00001110010110;
													assign node1287 = (inp[1]) ? node1291 : node1288;
														assign node1288 = (inp[2]) ? 14'b00001100010110 : 14'b01001100010110;
														assign node1291 = (inp[2]) ? 14'b00001000010110 : 14'b01001000010110;
												assign node1294 = (inp[6]) ? node1300 : node1295;
													assign node1295 = (inp[2]) ? 14'b00000010010110 : node1296;
														assign node1296 = (inp[1]) ? 14'b01000010010110 : 14'b01000110010110;
													assign node1300 = (inp[2]) ? node1302 : 14'b01000000010110;
														assign node1302 = (inp[1]) ? 14'b00000000010110 : 14'b00000100010110;
										assign node1305 = (inp[5]) ? node1333 : node1306;
											assign node1306 = (inp[6]) ? node1320 : node1307;
												assign node1307 = (inp[2]) ? node1313 : node1308;
													assign node1308 = (inp[9]) ? 14'b01001010010010 : node1309;
														assign node1309 = (inp[1]) ? 14'b01001010110010 : 14'b01001110110010;
													assign node1313 = (inp[1]) ? node1317 : node1314;
														assign node1314 = (inp[9]) ? 14'b00001110010010 : 14'b00001110110010;
														assign node1317 = (inp[9]) ? 14'b00001010010010 : 14'b00001010110010;
												assign node1320 = (inp[9]) ? node1326 : node1321;
													assign node1321 = (inp[2]) ? node1323 : 14'b01001000110010;
														assign node1323 = (inp[1]) ? 14'b00001000110010 : 14'b00001100110010;
													assign node1326 = (inp[1]) ? node1330 : node1327;
														assign node1327 = (inp[2]) ? 14'b00001100010010 : 14'b01001100010010;
														assign node1330 = (inp[2]) ? 14'b00001000010010 : 14'b01001000010010;
											assign node1333 = (inp[2]) ? node1335 : 14'b00000000000001;
												assign node1335 = (inp[6]) ? node1343 : node1336;
													assign node1336 = (inp[9]) ? node1340 : node1337;
														assign node1337 = (inp[1]) ? 14'b00000010110010 : 14'b00000110110010;
														assign node1340 = (inp[1]) ? 14'b00000010010010 : 14'b00000110010010;
													assign node1343 = (inp[9]) ? node1347 : node1344;
														assign node1344 = (inp[1]) ? 14'b00000000110010 : 14'b00000100110010;
														assign node1347 = (inp[1]) ? 14'b00000000010010 : 14'b00000100010010;
									assign node1350 = (inp[2]) ? 14'b00000000000001 : node1351;
										assign node1351 = (inp[10]) ? node1367 : node1352;
											assign node1352 = (inp[5]) ? node1354 : 14'b00000000000001;
												assign node1354 = (inp[9]) ? node1360 : node1355;
													assign node1355 = (inp[1]) ? 14'b01000000110010 : node1356;
														assign node1356 = (inp[6]) ? 14'b01000100110010 : 14'b01000110110010;
													assign node1360 = (inp[1]) ? node1364 : node1361;
														assign node1361 = (inp[6]) ? 14'b01000100010010 : 14'b01000110010010;
														assign node1364 = (inp[6]) ? 14'b01000000010010 : 14'b01000010010010;
											assign node1367 = (inp[5]) ? 14'b00000000000001 : node1368;
												assign node1368 = (inp[6]) ? node1376 : node1369;
													assign node1369 = (inp[9]) ? node1373 : node1370;
														assign node1370 = (inp[1]) ? 14'b00101010110000 : 14'b00101110110000;
														assign node1373 = (inp[1]) ? 14'b00101010010000 : 14'b00101110010000;
													assign node1376 = (inp[9]) ? node1380 : node1377;
														assign node1377 = (inp[1]) ? 14'b00101000110000 : 14'b00101100110000;
														assign node1380 = (inp[1]) ? 14'b00101000010000 : 14'b00101100010000;
							assign node1385 = (inp[6]) ? node1387 : 14'b00000000000001;
								assign node1387 = (inp[9]) ? 14'b00000000000001 : node1388;
									assign node1388 = (inp[12]) ? node1436 : node1389;
										assign node1389 = (inp[2]) ? node1413 : node1390;
											assign node1390 = (inp[5]) ? node1402 : node1391;
												assign node1391 = (inp[4]) ? node1397 : node1392;
													assign node1392 = (inp[10]) ? node1394 : 14'b00000000000001;
														assign node1394 = (inp[1]) ? 14'b01101000100010 : 14'b01101100100010;
													assign node1397 = (inp[10]) ? 14'b01101000100000 : node1398;
														assign node1398 = (inp[1]) ? 14'b01101000100110 : 14'b01101100100110;
												assign node1402 = (inp[1]) ? node1410 : node1403;
													assign node1403 = (inp[10]) ? node1407 : node1404;
														assign node1404 = (inp[4]) ? 14'b01100100100110 : 14'b00100100100010;
														assign node1407 = (inp[4]) ? 14'b01100100100000 : 14'b01100100100010;
													assign node1410 = (inp[4]) ? 14'b01100000100000 : 14'b01100000100010;
											assign node1413 = (inp[10]) ? node1425 : node1414;
												assign node1414 = (inp[4]) ? node1422 : node1415;
													assign node1415 = (inp[1]) ? node1419 : node1416;
														assign node1416 = (inp[5]) ? 14'b00000100100000 : 14'b00001100100000;
														assign node1419 = (inp[5]) ? 14'b00000000100000 : 14'b00001000100000;
													assign node1422 = (inp[1]) ? 14'b00101000100110 : 14'b00100100100110;
												assign node1425 = (inp[5]) ? node1431 : node1426;
													assign node1426 = (inp[4]) ? 14'b00000000000001 : node1427;
														assign node1427 = (inp[1]) ? 14'b00101000100010 : 14'b00101100100010;
													assign node1431 = (inp[4]) ? node1433 : 14'b00000000000001;
														assign node1433 = (inp[1]) ? 14'b00100000100000 : 14'b00100100100000;
										assign node1436 = (inp[4]) ? node1462 : node1437;
											assign node1437 = (inp[10]) ? node1451 : node1438;
												assign node1438 = (inp[5]) ? node1444 : node1439;
													assign node1439 = (inp[1]) ? node1441 : 14'b01001100100110;
														assign node1441 = (inp[2]) ? 14'b00001000100110 : 14'b01001000100110;
													assign node1444 = (inp[1]) ? node1448 : node1445;
														assign node1445 = (inp[2]) ? 14'b00000100100110 : 14'b01000100100110;
														assign node1448 = (inp[2]) ? 14'b00000000100110 : 14'b01000000100110;
												assign node1451 = (inp[5]) ? node1457 : node1452;
													assign node1452 = (inp[2]) ? 14'b00001000100010 : node1453;
														assign node1453 = (inp[1]) ? 14'b01001000100010 : 14'b01001100100010;
													assign node1457 = (inp[2]) ? node1459 : 14'b00000000000001;
														assign node1459 = (inp[1]) ? 14'b00000000100010 : 14'b00000100100010;
											assign node1462 = (inp[2]) ? 14'b00000000000001 : node1463;
												assign node1463 = (inp[1]) ? node1465 : 14'b00000000000001;
													assign node1465 = (inp[10]) ? node1469 : node1466;
														assign node1466 = (inp[5]) ? 14'b01000000100010 : 14'b00000000000001;
														assign node1469 = (inp[5]) ? 14'b00000000000001 : 14'b00101000100000;
				assign node1475 = (inp[10]) ? 14'b00000000000001 : node1476;
					assign node1476 = (inp[4]) ? node1934 : node1477;
						assign node1477 = (inp[7]) ? node1795 : node1478;
							assign node1478 = (inp[6]) ? node1658 : node1479;
								assign node1479 = (inp[9]) ? node1577 : node1480;
									assign node1480 = (inp[1]) ? node1522 : node1481;
										assign node1481 = (inp[0]) ? node1495 : node1482;
											assign node1482 = (inp[3]) ? node1484 : 14'b00000000000001;
												assign node1484 = (inp[12]) ? node1490 : node1485;
													assign node1485 = (inp[2]) ? 14'b00111110110100 : node1486;
														assign node1486 = (inp[5]) ? 14'b01110110110100 : 14'b01111110110100;
													assign node1490 = (inp[2]) ? 14'b00010110110100 : node1491;
														assign node1491 = (inp[5]) ? 14'b01010110110100 : 14'b01011110110100;
											assign node1495 = (inp[3]) ? node1509 : node1496;
												assign node1496 = (inp[12]) ? node1502 : node1497;
													assign node1497 = (inp[2]) ? 14'b00111110100100 : node1498;
														assign node1498 = (inp[5]) ? 14'b01110110100100 : 14'b01111110100100;
													assign node1502 = (inp[2]) ? node1506 : node1503;
														assign node1503 = (inp[5]) ? 14'b01010110100100 : 14'b01011110100100;
														assign node1506 = (inp[5]) ? 14'b00010110100100 : 14'b00011110100100;
												assign node1509 = (inp[5]) ? node1515 : node1510;
													assign node1510 = (inp[2]) ? node1512 : 14'b01101110100100;
														assign node1512 = (inp[12]) ? 14'b00001110100100 : 14'b00101110100100;
													assign node1515 = (inp[2]) ? node1519 : node1516;
														assign node1516 = (inp[12]) ? 14'b01000110100100 : 14'b01100110100100;
														assign node1519 = (inp[12]) ? 14'b00000110100100 : 14'b00100110100100;
										assign node1522 = (inp[2]) ? node1550 : node1523;
											assign node1523 = (inp[12]) ? node1535 : node1524;
												assign node1524 = (inp[3]) ? node1532 : node1525;
													assign node1525 = (inp[5]) ? node1529 : node1526;
														assign node1526 = (inp[0]) ? 14'b01111010100100 : 14'b01111010000100;
														assign node1529 = (inp[0]) ? 14'b01110010100100 : 14'b01110010000100;
													assign node1532 = (inp[5]) ? 14'b01110010110100 : 14'b01111010110100;
												assign node1535 = (inp[5]) ? node1543 : node1536;
													assign node1536 = (inp[0]) ? node1540 : node1537;
														assign node1537 = (inp[3]) ? 14'b01011010110100 : 14'b01011010000100;
														assign node1540 = (inp[3]) ? 14'b01001010100100 : 14'b01011010100100;
													assign node1543 = (inp[3]) ? node1547 : node1544;
														assign node1544 = (inp[0]) ? 14'b01010010100100 : 14'b01010010000100;
														assign node1547 = (inp[0]) ? 14'b01000010100100 : 14'b01010010110100;
											assign node1550 = (inp[5]) ? node1564 : node1551;
												assign node1551 = (inp[12]) ? node1559 : node1552;
													assign node1552 = (inp[0]) ? node1556 : node1553;
														assign node1553 = (inp[3]) ? 14'b00111010110100 : 14'b00111010000100;
														assign node1556 = (inp[3]) ? 14'b00101010100100 : 14'b00111010100100;
													assign node1559 = (inp[0]) ? 14'b00001010100100 : node1560;
														assign node1560 = (inp[3]) ? 14'b00011010110100 : 14'b00011010000100;
												assign node1564 = (inp[12]) ? node1570 : node1565;
													assign node1565 = (inp[0]) ? node1567 : 14'b00110010110100;
														assign node1567 = (inp[3]) ? 14'b00100010100100 : 14'b00110010100100;
													assign node1570 = (inp[3]) ? node1574 : node1571;
														assign node1571 = (inp[0]) ? 14'b00010010100100 : 14'b00010010000100;
														assign node1574 = (inp[0]) ? 14'b00000010100100 : 14'b00010010110100;
									assign node1577 = (inp[0]) ? node1629 : node1578;
										assign node1578 = (inp[3]) ? node1606 : node1579;
											assign node1579 = (inp[1]) ? node1593 : node1580;
												assign node1580 = (inp[5]) ? node1588 : node1581;
													assign node1581 = (inp[12]) ? node1585 : node1582;
														assign node1582 = (inp[2]) ? 14'b00101100000100 : 14'b01101100000100;
														assign node1585 = (inp[2]) ? 14'b00001100000100 : 14'b01001100000100;
													assign node1588 = (inp[12]) ? node1590 : 14'b01100100000100;
														assign node1590 = (inp[2]) ? 14'b00000100000100 : 14'b01000100000100;
												assign node1593 = (inp[5]) ? node1601 : node1594;
													assign node1594 = (inp[2]) ? node1598 : node1595;
														assign node1595 = (inp[12]) ? 14'b01001000000100 : 14'b01101000000100;
														assign node1598 = (inp[12]) ? 14'b00001000000100 : 14'b00101000000100;
													assign node1601 = (inp[2]) ? node1603 : 14'b01100000000100;
														assign node1603 = (inp[12]) ? 14'b00000000000100 : 14'b00100000000100;
											assign node1606 = (inp[5]) ? node1618 : node1607;
												assign node1607 = (inp[12]) ? node1611 : node1608;
													assign node1608 = (inp[1]) ? 14'b01111010010100 : 14'b01111110010100;
													assign node1611 = (inp[2]) ? node1615 : node1612;
														assign node1612 = (inp[1]) ? 14'b01011010010100 : 14'b01011110010100;
														assign node1615 = (inp[1]) ? 14'b00011010010100 : 14'b00011110010100;
												assign node1618 = (inp[2]) ? node1622 : node1619;
													assign node1619 = (inp[1]) ? 14'b01010010010100 : 14'b01010110010100;
													assign node1622 = (inp[1]) ? node1626 : node1623;
														assign node1623 = (inp[12]) ? 14'b00010110010100 : 14'b00110110010100;
														assign node1626 = (inp[12]) ? 14'b00010010010100 : 14'b00110010010100;
										assign node1629 = (inp[1]) ? node1645 : node1630;
											assign node1630 = (inp[3]) ? 14'b00000000000001 : node1631;
												assign node1631 = (inp[2]) ? node1637 : node1632;
													assign node1632 = (inp[12]) ? 14'b01010110000100 : node1633;
														assign node1633 = (inp[5]) ? 14'b01110110000100 : 14'b01111110000100;
													assign node1637 = (inp[12]) ? node1641 : node1638;
														assign node1638 = (inp[5]) ? 14'b00110110000100 : 14'b00111110000100;
														assign node1641 = (inp[5]) ? 14'b00010110000100 : 14'b00011110000100;
											assign node1645 = (inp[3]) ? node1647 : 14'b00000000000001;
												assign node1647 = (inp[2]) ? node1655 : node1648;
													assign node1648 = (inp[12]) ? node1652 : node1649;
														assign node1649 = (inp[5]) ? 14'b01100010000100 : 14'b01101010000100;
														assign node1652 = (inp[5]) ? 14'b01000010000100 : 14'b01001010000100;
													assign node1655 = (inp[12]) ? 14'b00001010000100 : 14'b00101010000100;
								assign node1658 = (inp[3]) ? node1758 : node1659;
									assign node1659 = (inp[1]) ? node1717 : node1660;
										assign node1660 = (inp[9]) ? node1690 : node1661;
											assign node1661 = (inp[12]) ? node1675 : node1662;
												assign node1662 = (inp[5]) ? node1670 : node1663;
													assign node1663 = (inp[2]) ? node1667 : node1664;
														assign node1664 = (inp[0]) ? 14'b01111100100100 : 14'b01111100110100;
														assign node1667 = (inp[0]) ? 14'b00111100100100 : 14'b00111100110100;
													assign node1670 = (inp[2]) ? 14'b00110100110100 : node1671;
														assign node1671 = (inp[0]) ? 14'b01110100100100 : 14'b01110100110100;
												assign node1675 = (inp[5]) ? node1683 : node1676;
													assign node1676 = (inp[2]) ? node1680 : node1677;
														assign node1677 = (inp[0]) ? 14'b01011100100100 : 14'b01011100110100;
														assign node1680 = (inp[0]) ? 14'b00011100100100 : 14'b00011100110100;
													assign node1683 = (inp[0]) ? node1687 : node1684;
														assign node1684 = (inp[2]) ? 14'b00010100110100 : 14'b01010100110100;
														assign node1687 = (inp[2]) ? 14'b00010100100100 : 14'b01010100100100;
											assign node1690 = (inp[5]) ? node1704 : node1691;
												assign node1691 = (inp[12]) ? node1699 : node1692;
													assign node1692 = (inp[0]) ? node1696 : node1693;
														assign node1693 = (inp[2]) ? 14'b00111100010100 : 14'b01111100010100;
														assign node1696 = (inp[2]) ? 14'b00111100000100 : 14'b01111100000100;
													assign node1699 = (inp[2]) ? 14'b00011100010100 : node1700;
														assign node1700 = (inp[0]) ? 14'b01011100000100 : 14'b01011100010100;
												assign node1704 = (inp[12]) ? node1712 : node1705;
													assign node1705 = (inp[0]) ? node1709 : node1706;
														assign node1706 = (inp[2]) ? 14'b00110100010100 : 14'b01110100010100;
														assign node1709 = (inp[2]) ? 14'b00110100000100 : 14'b01110100000100;
													assign node1712 = (inp[0]) ? 14'b00010100000100 : node1713;
														assign node1713 = (inp[2]) ? 14'b00010100010100 : 14'b01010100010100;
										assign node1717 = (inp[0]) ? node1743 : node1718;
											assign node1718 = (inp[9]) ? node1730 : node1719;
												assign node1719 = (inp[2]) ? node1723 : node1720;
													assign node1720 = (inp[12]) ? 14'b01011000110100 : 14'b01111000110100;
													assign node1723 = (inp[12]) ? node1727 : node1724;
														assign node1724 = (inp[5]) ? 14'b00110000110100 : 14'b00111000110100;
														assign node1727 = (inp[5]) ? 14'b00010000110100 : 14'b00011000110100;
												assign node1730 = (inp[5]) ? node1736 : node1731;
													assign node1731 = (inp[2]) ? node1733 : 14'b01011000010100;
														assign node1733 = (inp[12]) ? 14'b00011000010100 : 14'b00111000010100;
													assign node1736 = (inp[2]) ? node1740 : node1737;
														assign node1737 = (inp[12]) ? 14'b01010000010100 : 14'b01110000010100;
														assign node1740 = (inp[12]) ? 14'b00010000010100 : 14'b00110000010100;
											assign node1743 = (inp[9]) ? node1745 : 14'b00000000000001;
												assign node1745 = (inp[12]) ? node1751 : node1746;
													assign node1746 = (inp[5]) ? 14'b01110000000100 : node1747;
														assign node1747 = (inp[2]) ? 14'b00111000000100 : 14'b01111000000100;
													assign node1751 = (inp[2]) ? node1755 : node1752;
														assign node1752 = (inp[5]) ? 14'b01010000000100 : 14'b01011000000100;
														assign node1755 = (inp[5]) ? 14'b00010000000100 : 14'b00011000000100;
									assign node1758 = (inp[9]) ? 14'b00000000000001 : node1759;
										assign node1759 = (inp[1]) ? node1777 : node1760;
											assign node1760 = (inp[0]) ? node1762 : 14'b00000000000001;
												assign node1762 = (inp[12]) ? node1770 : node1763;
													assign node1763 = (inp[5]) ? node1767 : node1764;
														assign node1764 = (inp[2]) ? 14'b00101110000100 : 14'b01101110000100;
														assign node1767 = (inp[2]) ? 14'b00100110000100 : 14'b01100110000100;
													assign node1770 = (inp[2]) ? node1774 : node1771;
														assign node1771 = (inp[5]) ? 14'b01000110000100 : 14'b01001110000100;
														assign node1774 = (inp[5]) ? 14'b00000110000100 : 14'b00001110000100;
											assign node1777 = (inp[0]) ? 14'b00000000000001 : node1778;
												assign node1778 = (inp[2]) ? node1786 : node1779;
													assign node1779 = (inp[5]) ? node1783 : node1780;
														assign node1780 = (inp[12]) ? 14'b01011000100100 : 14'b01111000100100;
														assign node1783 = (inp[12]) ? 14'b01010000100100 : 14'b01110000100100;
													assign node1786 = (inp[5]) ? node1790 : node1787;
														assign node1787 = (inp[12]) ? 14'b00011000100100 : 14'b00111000100100;
														assign node1790 = (inp[12]) ? 14'b00010000100100 : 14'b00110000100100;
							assign node1795 = (inp[0]) ? 14'b00000000000001 : node1796;
								assign node1796 = (inp[3]) ? node1904 : node1797;
									assign node1797 = (inp[5]) ? node1849 : node1798;
										assign node1798 = (inp[2]) ? node1824 : node1799;
											assign node1799 = (inp[12]) ? node1811 : node1800;
												assign node1800 = (inp[6]) ? node1806 : node1801;
													assign node1801 = (inp[9]) ? 14'b01101010010100 : node1802;
														assign node1802 = (inp[1]) ? 14'b01101010110100 : 14'b01101110110100;
													assign node1806 = (inp[9]) ? node1808 : 14'b01101000110100;
														assign node1808 = (inp[1]) ? 14'b01101000010100 : 14'b01101100010100;
												assign node1811 = (inp[9]) ? node1817 : node1812;
													assign node1812 = (inp[1]) ? 14'b01001000110100 : node1813;
														assign node1813 = (inp[6]) ? 14'b01001100110100 : 14'b01001110110100;
													assign node1817 = (inp[6]) ? node1821 : node1818;
														assign node1818 = (inp[1]) ? 14'b01001010010100 : 14'b01001110010100;
														assign node1821 = (inp[1]) ? 14'b01001000010100 : 14'b01001100010100;
											assign node1824 = (inp[9]) ? node1834 : node1825;
												assign node1825 = (inp[1]) ? node1829 : node1826;
													assign node1826 = (inp[12]) ? 14'b00001100110100 : 14'b00101100110100;
													assign node1829 = (inp[12]) ? node1831 : 14'b00101000110100;
														assign node1831 = (inp[6]) ? 14'b00001000110100 : 14'b00001010110100;
												assign node1834 = (inp[12]) ? node1842 : node1835;
													assign node1835 = (inp[1]) ? node1839 : node1836;
														assign node1836 = (inp[6]) ? 14'b00101100010100 : 14'b00101110010100;
														assign node1839 = (inp[6]) ? 14'b00101000010100 : 14'b00101010010100;
													assign node1842 = (inp[1]) ? node1846 : node1843;
														assign node1843 = (inp[6]) ? 14'b00001100010100 : 14'b00001110010100;
														assign node1846 = (inp[6]) ? 14'b00001000010100 : 14'b00001010010100;
										assign node1849 = (inp[6]) ? node1875 : node1850;
											assign node1850 = (inp[1]) ? node1866 : node1851;
												assign node1851 = (inp[12]) ? node1859 : node1852;
													assign node1852 = (inp[2]) ? node1856 : node1853;
														assign node1853 = (inp[9]) ? 14'b01100110010100 : 14'b01100110110100;
														assign node1856 = (inp[9]) ? 14'b00100110010100 : 14'b00100110110100;
													assign node1859 = (inp[2]) ? node1863 : node1860;
														assign node1860 = (inp[9]) ? 14'b01000110010100 : 14'b01000110110100;
														assign node1863 = (inp[9]) ? 14'b00000110010100 : 14'b00000110110100;
												assign node1866 = (inp[9]) ? node1870 : node1867;
													assign node1867 = (inp[2]) ? 14'b00000010110100 : 14'b01000010110100;
													assign node1870 = (inp[2]) ? 14'b00000010010100 : node1871;
														assign node1871 = (inp[12]) ? 14'b01000010010100 : 14'b01100010010100;
											assign node1875 = (inp[2]) ? node1891 : node1876;
												assign node1876 = (inp[1]) ? node1884 : node1877;
													assign node1877 = (inp[12]) ? node1881 : node1878;
														assign node1878 = (inp[9]) ? 14'b01100100010100 : 14'b01100100110100;
														assign node1881 = (inp[9]) ? 14'b01000100010100 : 14'b01000100110100;
													assign node1884 = (inp[9]) ? node1888 : node1885;
														assign node1885 = (inp[12]) ? 14'b01000000110100 : 14'b01100000110100;
														assign node1888 = (inp[12]) ? 14'b01000000010100 : 14'b01100000010100;
												assign node1891 = (inp[12]) ? node1897 : node1892;
													assign node1892 = (inp[1]) ? node1894 : 14'b00100100110100;
														assign node1894 = (inp[9]) ? 14'b00100000010100 : 14'b00100000110100;
													assign node1897 = (inp[9]) ? node1901 : node1898;
														assign node1898 = (inp[1]) ? 14'b00000000110100 : 14'b00000100110100;
														assign node1901 = (inp[1]) ? 14'b00000000010100 : 14'b00000100010100;
									assign node1904 = (inp[9]) ? 14'b00000000000001 : node1905;
										assign node1905 = (inp[6]) ? node1907 : 14'b00000000000001;
											assign node1907 = (inp[1]) ? node1921 : node1908;
												assign node1908 = (inp[12]) ? node1914 : node1909;
													assign node1909 = (inp[2]) ? 14'b00101100100100 : node1910;
														assign node1910 = (inp[5]) ? 14'b01100100100100 : 14'b01101100100100;
													assign node1914 = (inp[2]) ? node1918 : node1915;
														assign node1915 = (inp[5]) ? 14'b01000100100100 : 14'b01001100100100;
														assign node1918 = (inp[5]) ? 14'b00000100100100 : 14'b00001100100100;
												assign node1921 = (inp[2]) ? node1925 : node1922;
													assign node1922 = (inp[12]) ? 14'b01000000100100 : 14'b01100000100100;
													assign node1925 = (inp[5]) ? node1929 : node1926;
														assign node1926 = (inp[12]) ? 14'b00001000100100 : 14'b00101000100100;
														assign node1929 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
						assign node1934 = (inp[2]) ? node2080 : node1935;
							assign node1935 = (inp[12]) ? node1953 : node1936;
								assign node1936 = (inp[1]) ? 14'b00000000000001 : node1937;
									assign node1937 = (inp[3]) ? node1939 : 14'b00000000000001;
										assign node1939 = (inp[9]) ? 14'b00000000000001 : node1940;
											assign node1940 = (inp[0]) ? 14'b00000000000001 : node1941;
												assign node1941 = (inp[5]) ? 14'b00000000000001 : node1942;
													assign node1942 = (inp[7]) ? node1946 : node1943;
														assign node1943 = (inp[6]) ? 14'b10000001001000 : 14'b00000000000001;
														assign node1946 = (inp[6]) ? 14'b00000000000001 : 14'b10000001000000;
								assign node1953 = (inp[0]) ? node2039 : node1954;
									assign node1954 = (inp[3]) ? node2006 : node1955;
										assign node1955 = (inp[7]) ? node1975 : node1956;
											assign node1956 = (inp[6]) ? node1966 : node1957;
												assign node1957 = (inp[1]) ? node1959 : 14'b00000000000001;
													assign node1959 = (inp[9]) ? node1963 : node1960;
														assign node1960 = (inp[5]) ? 14'b01010010000000 : 14'b01011010000000;
														assign node1963 = (inp[5]) ? 14'b01000000000000 : 14'b01001000000000;
												assign node1966 = (inp[5]) ? node1972 : node1967;
													assign node1967 = (inp[1]) ? node1969 : 14'b01011100010000;
														assign node1969 = (inp[9]) ? 14'b01011000010000 : 14'b01011000110000;
													assign node1972 = (inp[1]) ? 14'b01010000110000 : 14'b01010100110000;
											assign node1975 = (inp[5]) ? node1991 : node1976;
												assign node1976 = (inp[1]) ? node1984 : node1977;
													assign node1977 = (inp[6]) ? node1981 : node1978;
														assign node1978 = (inp[9]) ? 14'b01001110010000 : 14'b01001110110000;
														assign node1981 = (inp[9]) ? 14'b01001100010000 : 14'b01001100110000;
													assign node1984 = (inp[9]) ? node1988 : node1985;
														assign node1985 = (inp[6]) ? 14'b01001000110000 : 14'b01001010110000;
														assign node1988 = (inp[6]) ? 14'b01001000010000 : 14'b01001010010000;
												assign node1991 = (inp[6]) ? node1999 : node1992;
													assign node1992 = (inp[9]) ? node1996 : node1993;
														assign node1993 = (inp[1]) ? 14'b01000010110000 : 14'b01000110110000;
														assign node1996 = (inp[1]) ? 14'b01000010010000 : 14'b01000110010000;
													assign node1999 = (inp[1]) ? node2003 : node2000;
														assign node2000 = (inp[9]) ? 14'b01000100010000 : 14'b01000100110000;
														assign node2003 = (inp[9]) ? 14'b01000000010000 : 14'b01000000110000;
										assign node2006 = (inp[7]) ? node2028 : node2007;
											assign node2007 = (inp[6]) ? node2021 : node2008;
												assign node2008 = (inp[9]) ? node2016 : node2009;
													assign node2009 = (inp[1]) ? node2013 : node2010;
														assign node2010 = (inp[5]) ? 14'b01010110110000 : 14'b01011110110000;
														assign node2013 = (inp[5]) ? 14'b01010010110000 : 14'b01011010110000;
													assign node2016 = (inp[5]) ? node2018 : 14'b01011010010000;
														assign node2018 = (inp[1]) ? 14'b01010010010000 : 14'b01010110010000;
												assign node2021 = (inp[1]) ? node2023 : 14'b00000000000001;
													assign node2023 = (inp[9]) ? 14'b00000000000001 : node2024;
														assign node2024 = (inp[5]) ? 14'b01010000100000 : 14'b01011000100000;
											assign node2028 = (inp[9]) ? 14'b00000000000001 : node2029;
												assign node2029 = (inp[6]) ? node2031 : 14'b00000000000001;
													assign node2031 = (inp[5]) ? node2035 : node2032;
														assign node2032 = (inp[1]) ? 14'b01001000100000 : 14'b01001100100000;
														assign node2035 = (inp[1]) ? 14'b01000000100000 : 14'b01000100100000;
									assign node2039 = (inp[7]) ? 14'b00000000000001 : node2040;
										assign node2040 = (inp[1]) ? node2060 : node2041;
											assign node2041 = (inp[9]) ? node2055 : node2042;
												assign node2042 = (inp[3]) ? node2050 : node2043;
													assign node2043 = (inp[5]) ? node2047 : node2044;
														assign node2044 = (inp[6]) ? 14'b01011100100000 : 14'b01011110100000;
														assign node2047 = (inp[6]) ? 14'b01010100100000 : 14'b01010110100000;
													assign node2050 = (inp[5]) ? 14'b01000110100000 : node2051;
														assign node2051 = (inp[6]) ? 14'b01001110000000 : 14'b01001110100000;
												assign node2055 = (inp[6]) ? node2057 : 14'b00000000000001;
													assign node2057 = (inp[5]) ? 14'b01010100000000 : 14'b01011100000000;
											assign node2060 = (inp[6]) ? node2072 : node2061;
												assign node2061 = (inp[9]) ? node2067 : node2062;
													assign node2062 = (inp[3]) ? 14'b01001010100000 : node2063;
														assign node2063 = (inp[5]) ? 14'b01010010100000 : 14'b01011010100000;
													assign node2067 = (inp[3]) ? node2069 : 14'b00000000000001;
														assign node2069 = (inp[5]) ? 14'b01000010000000 : 14'b01001010000000;
												assign node2072 = (inp[3]) ? 14'b00000000000001 : node2073;
													assign node2073 = (inp[9]) ? node2075 : 14'b00000000000001;
														assign node2075 = (inp[5]) ? 14'b01010000000000 : 14'b01011000000000;
							assign node2080 = (inp[3]) ? 14'b00000000000001 : node2081;
								assign node2081 = (inp[1]) ? node2083 : 14'b00000000000001;
									assign node2083 = (inp[9]) ? 14'b00000000000001 : node2084;
										assign node2084 = (inp[6]) ? node2086 : 14'b00000000000001;
											assign node2086 = (inp[7]) ? 14'b00000000000001 : node2087;
												assign node2087 = (inp[12]) ? node2089 : 14'b00000000000001;
													assign node2089 = (inp[5]) ? 14'b00000000000001 : 14'b10000000000000;
		assign node2096 = (inp[0]) ? node3484 : node2097;
			assign node2097 = (inp[5]) ? node3007 : node2098;
				assign node2098 = (inp[6]) ? node2670 : node2099;
					assign node2099 = (inp[2]) ? node2433 : node2100;
						assign node2100 = (inp[4]) ? node2264 : node2101;
							assign node2101 = (inp[12]) ? node2179 : node2102;
								assign node2102 = (inp[7]) ? node2132 : node2103;
									assign node2103 = (inp[10]) ? node2111 : node2104;
										assign node2104 = (inp[3]) ? 14'b00000000000001 : node2105;
											assign node2105 = (inp[1]) ? 14'b00000000000001 : node2106;
												assign node2106 = (inp[9]) ? 14'b00000000000001 : 14'b10000000001000;
										assign node2111 = (inp[8]) ? node2125 : node2112;
											assign node2112 = (inp[3]) ? node2120 : node2113;
												assign node2113 = (inp[1]) ? node2117 : node2114;
													assign node2114 = (inp[9]) ? 14'b01100100000010 : 14'b00000000000001;
													assign node2117 = (inp[9]) ? 14'b01110110000010 : 14'b01110110100010;
												assign node2120 = (inp[1]) ? 14'b01100110100010 : node2121;
													assign node2121 = (inp[9]) ? 14'b01110110010010 : 14'b01110110110010;
											assign node2125 = (inp[3]) ? 14'b00000000000001 : node2126;
												assign node2126 = (inp[1]) ? 14'b00000000000001 : node2127;
													assign node2127 = (inp[9]) ? 14'b00000000000001 : 14'b10000000001000;
									assign node2132 = (inp[8]) ? node2164 : node2133;
										assign node2133 = (inp[10]) ? node2149 : node2134;
											assign node2134 = (inp[3]) ? node2142 : node2135;
												assign node2135 = (inp[1]) ? node2139 : node2136;
													assign node2136 = (inp[9]) ? 14'b00000000000010 : 14'b00000000000001;
													assign node2139 = (inp[9]) ? 14'b00010010000010 : 14'b00010010100010;
												assign node2142 = (inp[1]) ? node2146 : node2143;
													assign node2143 = (inp[9]) ? 14'b00010010010010 : 14'b00010010110010;
													assign node2146 = (inp[9]) ? 14'b00000010000010 : 14'b00000010100010;
											assign node2149 = (inp[3]) ? node2157 : node2150;
												assign node2150 = (inp[1]) ? node2154 : node2151;
													assign node2151 = (inp[9]) ? 14'b01100000000010 : 14'b00000000000001;
													assign node2154 = (inp[9]) ? 14'b01110010000010 : 14'b01110010100010;
												assign node2157 = (inp[1]) ? node2161 : node2158;
													assign node2158 = (inp[9]) ? 14'b01110010010010 : 14'b01110010110010;
													assign node2161 = (inp[9]) ? 14'b01100010000010 : 14'b01100010100010;
										assign node2164 = (inp[1]) ? node2172 : node2165;
											assign node2165 = (inp[3]) ? node2169 : node2166;
												assign node2166 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000001;
												assign node2169 = (inp[9]) ? 14'b00010010010000 : 14'b00010010110000;
											assign node2172 = (inp[9]) ? node2176 : node2173;
												assign node2173 = (inp[3]) ? 14'b00000010100000 : 14'b00010010100000;
												assign node2176 = (inp[3]) ? 14'b00000010000000 : 14'b00010010000000;
								assign node2179 = (inp[3]) ? node2217 : node2180;
									assign node2180 = (inp[1]) ? node2194 : node2181;
										assign node2181 = (inp[9]) ? node2183 : 14'b00000000000001;
											assign node2183 = (inp[8]) ? node2191 : node2184;
												assign node2184 = (inp[10]) ? node2188 : node2185;
													assign node2185 = (inp[7]) ? 14'b00000000000000 : 14'b01000000000100;
													assign node2188 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
												assign node2191 = (inp[7]) ? 14'b01000000000100 : 14'b01000100000100;
										assign node2194 = (inp[9]) ? node2206 : node2195;
											assign node2195 = (inp[8]) ? node2203 : node2196;
												assign node2196 = (inp[10]) ? node2200 : node2197;
													assign node2197 = (inp[7]) ? 14'b00010010100000 : 14'b01010010100100;
													assign node2200 = (inp[7]) ? 14'b01110010100000 : 14'b01110110100000;
												assign node2203 = (inp[7]) ? 14'b01010010100100 : 14'b01010110100100;
											assign node2206 = (inp[8]) ? node2214 : node2207;
												assign node2207 = (inp[10]) ? node2211 : node2208;
													assign node2208 = (inp[7]) ? 14'b00010010000000 : 14'b01010010000100;
													assign node2211 = (inp[7]) ? 14'b01110010000000 : 14'b01110110000000;
												assign node2214 = (inp[7]) ? 14'b01010010000100 : 14'b01010110000100;
									assign node2217 = (inp[1]) ? node2241 : node2218;
										assign node2218 = (inp[9]) ? node2230 : node2219;
											assign node2219 = (inp[8]) ? node2227 : node2220;
												assign node2220 = (inp[10]) ? node2224 : node2221;
													assign node2221 = (inp[7]) ? 14'b00010010110000 : 14'b01010010110100;
													assign node2224 = (inp[7]) ? 14'b01110010110000 : 14'b01110110110000;
												assign node2227 = (inp[7]) ? 14'b01010010110100 : 14'b01010110110100;
											assign node2230 = (inp[8]) ? node2238 : node2231;
												assign node2231 = (inp[10]) ? node2235 : node2232;
													assign node2232 = (inp[7]) ? 14'b00010010010000 : 14'b01010010010100;
													assign node2235 = (inp[7]) ? 14'b01110010010000 : 14'b01110110010000;
												assign node2238 = (inp[7]) ? 14'b01010010010100 : 14'b01010110010100;
										assign node2241 = (inp[9]) ? node2253 : node2242;
											assign node2242 = (inp[8]) ? node2250 : node2243;
												assign node2243 = (inp[10]) ? node2247 : node2244;
													assign node2244 = (inp[7]) ? 14'b00000010100000 : 14'b01000010100100;
													assign node2247 = (inp[7]) ? 14'b01100010100000 : 14'b01100110100000;
												assign node2250 = (inp[7]) ? 14'b01000010100100 : 14'b01000110100100;
											assign node2253 = (inp[8]) ? node2261 : node2254;
												assign node2254 = (inp[10]) ? node2258 : node2255;
													assign node2255 = (inp[7]) ? 14'b00000010000000 : 14'b01000010000100;
													assign node2258 = (inp[7]) ? 14'b01100010000000 : 14'b01100110000000;
												assign node2261 = (inp[7]) ? 14'b01000010000100 : 14'b01000110000100;
							assign node2264 = (inp[7]) ? node2348 : node2265;
								assign node2265 = (inp[1]) ? node2303 : node2266;
									assign node2266 = (inp[3]) ? node2280 : node2267;
										assign node2267 = (inp[9]) ? node2269 : 14'b00000000000001;
											assign node2269 = (inp[8]) ? node2277 : node2270;
												assign node2270 = (inp[10]) ? node2274 : node2271;
													assign node2271 = (inp[12]) ? 14'b00100100000100 : 14'b00100100000110;
													assign node2274 = (inp[12]) ? 14'b00100100000000 : 14'b00100100000010;
												assign node2277 = (inp[12]) ? 14'b00000100000100 : 14'b00100100000100;
										assign node2280 = (inp[9]) ? node2292 : node2281;
											assign node2281 = (inp[8]) ? node2289 : node2282;
												assign node2282 = (inp[12]) ? node2286 : node2283;
													assign node2283 = (inp[10]) ? 14'b00110110110010 : 14'b00110110110110;
													assign node2286 = (inp[10]) ? 14'b00110110110000 : 14'b00110110110100;
												assign node2289 = (inp[12]) ? 14'b00010110110100 : 14'b00110110110100;
											assign node2292 = (inp[8]) ? node2300 : node2293;
												assign node2293 = (inp[10]) ? node2297 : node2294;
													assign node2294 = (inp[12]) ? 14'b00110110010100 : 14'b00110110010110;
													assign node2297 = (inp[12]) ? 14'b00110110010000 : 14'b00110110010010;
												assign node2300 = (inp[12]) ? 14'b00010110010100 : 14'b00110110010100;
									assign node2303 = (inp[9]) ? node2327 : node2304;
										assign node2304 = (inp[3]) ? node2316 : node2305;
											assign node2305 = (inp[8]) ? node2313 : node2306;
												assign node2306 = (inp[12]) ? node2310 : node2307;
													assign node2307 = (inp[10]) ? 14'b00110110100010 : 14'b00110110100110;
													assign node2310 = (inp[10]) ? 14'b00110110100000 : 14'b00110110100100;
												assign node2313 = (inp[12]) ? 14'b00010110100100 : 14'b00110110100100;
											assign node2316 = (inp[8]) ? node2324 : node2317;
												assign node2317 = (inp[12]) ? node2321 : node2318;
													assign node2318 = (inp[10]) ? 14'b00100110100010 : 14'b00100110100110;
													assign node2321 = (inp[10]) ? 14'b00100110100000 : 14'b00100110100100;
												assign node2324 = (inp[12]) ? 14'b00000110100100 : 14'b00100110100100;
										assign node2327 = (inp[3]) ? node2337 : node2328;
											assign node2328 = (inp[8]) ? node2334 : node2329;
												assign node2329 = (inp[10]) ? node2331 : 14'b00110110000110;
													assign node2331 = (inp[12]) ? 14'b00110110000000 : 14'b00110110000010;
												assign node2334 = (inp[12]) ? 14'b00010110000100 : 14'b00110110000100;
											assign node2337 = (inp[8]) ? node2345 : node2338;
												assign node2338 = (inp[10]) ? node2342 : node2339;
													assign node2339 = (inp[12]) ? 14'b00100110000100 : 14'b00100110000110;
													assign node2342 = (inp[12]) ? 14'b00100110000000 : 14'b00100110000010;
												assign node2345 = (inp[12]) ? 14'b00000110000100 : 14'b00100110000100;
								assign node2348 = (inp[9]) ? node2386 : node2349;
									assign node2349 = (inp[3]) ? node2363 : node2350;
										assign node2350 = (inp[1]) ? node2352 : 14'b00000000000001;
											assign node2352 = (inp[8]) ? node2360 : node2353;
												assign node2353 = (inp[10]) ? node2357 : node2354;
													assign node2354 = (inp[12]) ? 14'b00110010100100 : 14'b00110010100110;
													assign node2357 = (inp[12]) ? 14'b00110010100000 : 14'b00110010100010;
												assign node2360 = (inp[12]) ? 14'b00010010100100 : 14'b00110010100100;
										assign node2363 = (inp[1]) ? node2375 : node2364;
											assign node2364 = (inp[8]) ? node2372 : node2365;
												assign node2365 = (inp[12]) ? node2369 : node2366;
													assign node2366 = (inp[10]) ? 14'b00110010110010 : 14'b00110010110110;
													assign node2369 = (inp[10]) ? 14'b00110010110000 : 14'b00110010110100;
												assign node2372 = (inp[12]) ? 14'b00010010110100 : 14'b00110010110100;
											assign node2375 = (inp[8]) ? node2383 : node2376;
												assign node2376 = (inp[12]) ? node2380 : node2377;
													assign node2377 = (inp[10]) ? 14'b00100010100010 : 14'b00100010100110;
													assign node2380 = (inp[10]) ? 14'b00100010100000 : 14'b00100010100100;
												assign node2383 = (inp[12]) ? 14'b00000010100100 : 14'b00100010100100;
									assign node2386 = (inp[8]) ? node2418 : node2387;
										assign node2387 = (inp[12]) ? node2403 : node2388;
											assign node2388 = (inp[10]) ? node2396 : node2389;
												assign node2389 = (inp[3]) ? node2393 : node2390;
													assign node2390 = (inp[1]) ? 14'b00110010000110 : 14'b00100000000110;
													assign node2393 = (inp[1]) ? 14'b00100010000110 : 14'b00110010010110;
												assign node2396 = (inp[1]) ? node2400 : node2397;
													assign node2397 = (inp[3]) ? 14'b00110010010010 : 14'b00100000000010;
													assign node2400 = (inp[3]) ? 14'b00100010000010 : 14'b00110010000010;
											assign node2403 = (inp[10]) ? node2411 : node2404;
												assign node2404 = (inp[3]) ? node2408 : node2405;
													assign node2405 = (inp[1]) ? 14'b00110010000100 : 14'b00100000000100;
													assign node2408 = (inp[1]) ? 14'b00100010000100 : 14'b00110010010100;
												assign node2411 = (inp[1]) ? node2415 : node2412;
													assign node2412 = (inp[3]) ? 14'b00110010010000 : 14'b00100000000000;
													assign node2415 = (inp[3]) ? 14'b00100010000000 : 14'b00110010000000;
										assign node2418 = (inp[12]) ? node2426 : node2419;
											assign node2419 = (inp[1]) ? node2423 : node2420;
												assign node2420 = (inp[3]) ? 14'b00110010010100 : 14'b00100000000100;
												assign node2423 = (inp[3]) ? 14'b00100010000100 : 14'b00110010000100;
											assign node2426 = (inp[1]) ? node2430 : node2427;
												assign node2427 = (inp[3]) ? 14'b00010010010100 : 14'b00000000000100;
												assign node2430 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
						assign node2433 = (inp[4]) ? node2617 : node2434;
							assign node2434 = (inp[10]) ? node2554 : node2435;
								assign node2435 = (inp[7]) ? node2497 : node2436;
									assign node2436 = (inp[12]) ? node2466 : node2437;
										assign node2437 = (inp[8]) ? node2453 : node2438;
											assign node2438 = (inp[9]) ? node2446 : node2439;
												assign node2439 = (inp[1]) ? node2443 : node2440;
													assign node2440 = (inp[3]) ? 14'b01110110110110 : 14'b00000000000001;
													assign node2443 = (inp[3]) ? 14'b01100110100110 : 14'b01110110100110;
												assign node2446 = (inp[3]) ? node2450 : node2447;
													assign node2447 = (inp[1]) ? 14'b01110110000110 : 14'b01100100000110;
													assign node2450 = (inp[1]) ? 14'b01100110000110 : 14'b01110110010110;
											assign node2453 = (inp[3]) ? node2459 : node2454;
												assign node2454 = (inp[9]) ? node2456 : 14'b00000000000001;
													assign node2456 = (inp[1]) ? 14'b01110110000100 : 14'b01100100000100;
												assign node2459 = (inp[1]) ? node2463 : node2460;
													assign node2460 = (inp[9]) ? 14'b01110110010100 : 14'b01110110110100;
													assign node2463 = (inp[9]) ? 14'b01100110000100 : 14'b01100110100100;
										assign node2466 = (inp[8]) ? node2482 : node2467;
											assign node2467 = (inp[1]) ? node2475 : node2468;
												assign node2468 = (inp[3]) ? node2472 : node2469;
													assign node2469 = (inp[9]) ? 14'b01100100000100 : 14'b00000000000001;
													assign node2472 = (inp[9]) ? 14'b01110110010100 : 14'b01110110110100;
												assign node2475 = (inp[3]) ? node2479 : node2476;
													assign node2476 = (inp[9]) ? 14'b01110110000100 : 14'b01110110100100;
													assign node2479 = (inp[9]) ? 14'b01100110000100 : 14'b01100110100100;
											assign node2482 = (inp[1]) ? node2490 : node2483;
												assign node2483 = (inp[3]) ? node2487 : node2484;
													assign node2484 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
													assign node2487 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
												assign node2490 = (inp[3]) ? node2494 : node2491;
													assign node2491 = (inp[9]) ? 14'b01010110000000 : 14'b01010110100000;
													assign node2494 = (inp[9]) ? 14'b01000110000000 : 14'b01000110100000;
									assign node2497 = (inp[1]) ? node2523 : node2498;
										assign node2498 = (inp[3]) ? node2508 : node2499;
											assign node2499 = (inp[9]) ? node2501 : 14'b00000000000001;
												assign node2501 = (inp[8]) ? node2505 : node2502;
													assign node2502 = (inp[12]) ? 14'b01100000000100 : 14'b01100000000110;
													assign node2505 = (inp[12]) ? 14'b01000000000000 : 14'b01100000000100;
											assign node2508 = (inp[9]) ? node2516 : node2509;
												assign node2509 = (inp[12]) ? node2513 : node2510;
													assign node2510 = (inp[8]) ? 14'b01110010110100 : 14'b01110010110110;
													assign node2513 = (inp[8]) ? 14'b01010010110000 : 14'b01110010110100;
												assign node2516 = (inp[12]) ? node2520 : node2517;
													assign node2517 = (inp[8]) ? 14'b01110010010100 : 14'b01110010010110;
													assign node2520 = (inp[8]) ? 14'b01010010010000 : 14'b01110010010100;
										assign node2523 = (inp[9]) ? node2539 : node2524;
											assign node2524 = (inp[3]) ? node2532 : node2525;
												assign node2525 = (inp[8]) ? node2529 : node2526;
													assign node2526 = (inp[12]) ? 14'b01110010100100 : 14'b01110010100110;
													assign node2529 = (inp[12]) ? 14'b01010010100000 : 14'b01110010100100;
												assign node2532 = (inp[12]) ? node2536 : node2533;
													assign node2533 = (inp[8]) ? 14'b01100010100100 : 14'b01100010100110;
													assign node2536 = (inp[8]) ? 14'b01000010100000 : 14'b01100010100100;
											assign node2539 = (inp[12]) ? node2547 : node2540;
												assign node2540 = (inp[3]) ? node2544 : node2541;
													assign node2541 = (inp[8]) ? 14'b01110010000100 : 14'b01110010000110;
													assign node2544 = (inp[8]) ? 14'b01100010000100 : 14'b01100010000110;
												assign node2547 = (inp[8]) ? node2551 : node2548;
													assign node2548 = (inp[11]) ? 14'b01100010000100 : 14'b01110010000100;
													assign node2551 = (inp[3]) ? 14'b01000010000000 : 14'b01010010000000;
								assign node2554 = (inp[8]) ? node2556 : 14'b00000000000001;
									assign node2556 = (inp[12]) ? node2586 : node2557;
										assign node2557 = (inp[9]) ? node2571 : node2558;
											assign node2558 = (inp[1]) ? node2564 : node2559;
												assign node2559 = (inp[3]) ? node2561 : 14'b00000000000001;
													assign node2561 = (inp[7]) ? 14'b01110010110100 : 14'b01110110110100;
												assign node2564 = (inp[7]) ? node2568 : node2565;
													assign node2565 = (inp[3]) ? 14'b01100110100100 : 14'b01110110100100;
													assign node2568 = (inp[3]) ? 14'b01100010100100 : 14'b01110010100100;
											assign node2571 = (inp[7]) ? node2579 : node2572;
												assign node2572 = (inp[3]) ? node2576 : node2573;
													assign node2573 = (inp[1]) ? 14'b01110110000100 : 14'b01100100000100;
													assign node2576 = (inp[1]) ? 14'b01100110000100 : 14'b01110110010100;
												assign node2579 = (inp[1]) ? node2583 : node2580;
													assign node2580 = (inp[3]) ? 14'b01110010010100 : 14'b01100000000100;
													assign node2583 = (inp[3]) ? 14'b01100010000100 : 14'b01110010000100;
										assign node2586 = (inp[7]) ? node2602 : node2587;
											assign node2587 = (inp[1]) ? node2595 : node2588;
												assign node2588 = (inp[3]) ? node2592 : node2589;
													assign node2589 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
													assign node2592 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
												assign node2595 = (inp[9]) ? node2599 : node2596;
													assign node2596 = (inp[3]) ? 14'b01000110100000 : 14'b01010110100000;
													assign node2599 = (inp[3]) ? 14'b01000110000000 : 14'b01010110000000;
											assign node2602 = (inp[9]) ? node2610 : node2603;
												assign node2603 = (inp[1]) ? node2607 : node2604;
													assign node2604 = (inp[3]) ? 14'b01010010110000 : 14'b00000000000001;
													assign node2607 = (inp[3]) ? 14'b01000010100000 : 14'b01010010100000;
												assign node2610 = (inp[1]) ? node2614 : node2611;
													assign node2611 = (inp[3]) ? 14'b01010010010000 : 14'b01000000000000;
													assign node2614 = (inp[3]) ? 14'b01000010000000 : 14'b01010010000000;
							assign node2617 = (inp[7]) ? 14'b00000000000001 : node2618;
								assign node2618 = (inp[8]) ? 14'b00000000000001 : node2619;
									assign node2619 = (inp[10]) ? node2637 : node2620;
										assign node2620 = (inp[12]) ? node2622 : 14'b00000000000001;
											assign node2622 = (inp[9]) ? node2630 : node2623;
												assign node2623 = (inp[3]) ? node2627 : node2624;
													assign node2624 = (inp[1]) ? 14'b00010110100100 : 14'b00000000000001;
													assign node2627 = (inp[1]) ? 14'b00000110100100 : 14'b00010110110100;
												assign node2630 = (inp[3]) ? node2634 : node2631;
													assign node2631 = (inp[1]) ? 14'b00010110000100 : 14'b00000100000100;
													assign node2634 = (inp[1]) ? 14'b00000110000100 : 14'b00010110010100;
										assign node2637 = (inp[12]) ? node2653 : node2638;
											assign node2638 = (inp[3]) ? node2646 : node2639;
												assign node2639 = (inp[1]) ? node2643 : node2640;
													assign node2640 = (inp[9]) ? 14'b00000100000010 : 14'b00000000000001;
													assign node2643 = (inp[9]) ? 14'b00010110000010 : 14'b00010110100010;
												assign node2646 = (inp[1]) ? node2650 : node2647;
													assign node2647 = (inp[9]) ? 14'b00010110010010 : 14'b00010110110010;
													assign node2650 = (inp[9]) ? 14'b00000110000010 : 14'b00000110100010;
											assign node2653 = (inp[1]) ? node2661 : node2654;
												assign node2654 = (inp[3]) ? node2658 : node2655;
													assign node2655 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
													assign node2658 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
												assign node2661 = (inp[9]) ? node2665 : node2662;
													assign node2662 = (inp[3]) ? 14'b00000110100000 : 14'b00010110100000;
													assign node2665 = (inp[3]) ? 14'b00000110000000 : 14'b00010110000000;
					assign node2670 = (inp[3]) ? node2976 : node2671;
						assign node2671 = (inp[2]) ? node2851 : node2672;
							assign node2672 = (inp[4]) ? node2756 : node2673;
								assign node2673 = (inp[12]) ? node2709 : node2674;
									assign node2674 = (inp[7]) ? node2686 : node2675;
										assign node2675 = (inp[8]) ? 14'b00000000000001 : node2676;
											assign node2676 = (inp[10]) ? node2678 : 14'b00000000000001;
												assign node2678 = (inp[9]) ? node2682 : node2679;
													assign node2679 = (inp[1]) ? 14'b01110100100010 : 14'b01110100110010;
													assign node2682 = (inp[1]) ? 14'b01110100000010 : 14'b01110100010010;
										assign node2686 = (inp[8]) ? node2702 : node2687;
											assign node2687 = (inp[10]) ? node2695 : node2688;
												assign node2688 = (inp[1]) ? node2692 : node2689;
													assign node2689 = (inp[9]) ? 14'b00010000010010 : 14'b00010000110010;
													assign node2692 = (inp[9]) ? 14'b00010000000010 : 14'b00010000100010;
												assign node2695 = (inp[9]) ? node2699 : node2696;
													assign node2696 = (inp[1]) ? 14'b01110000100010 : 14'b01110000110010;
													assign node2699 = (inp[1]) ? 14'b01110000000010 : 14'b01110000010010;
											assign node2702 = (inp[9]) ? node2706 : node2703;
												assign node2703 = (inp[1]) ? 14'b00010000100000 : 14'b00010000110000;
												assign node2706 = (inp[1]) ? 14'b00010000000000 : 14'b00010000010000;
									assign node2709 = (inp[1]) ? node2733 : node2710;
										assign node2710 = (inp[8]) ? node2726 : node2711;
											assign node2711 = (inp[10]) ? node2719 : node2712;
												assign node2712 = (inp[7]) ? node2716 : node2713;
													assign node2713 = (inp[9]) ? 14'b01010000010100 : 14'b01010000110100;
													assign node2716 = (inp[9]) ? 14'b00010000010000 : 14'b00010000110000;
												assign node2719 = (inp[7]) ? node2723 : node2720;
													assign node2720 = (inp[9]) ? 14'b01110100010000 : 14'b01110100110000;
													assign node2723 = (inp[9]) ? 14'b01110000010000 : 14'b01110000110000;
											assign node2726 = (inp[9]) ? node2730 : node2727;
												assign node2727 = (inp[7]) ? 14'b01010000110100 : 14'b01010100110100;
												assign node2730 = (inp[7]) ? 14'b01010000010100 : 14'b01010100010100;
										assign node2733 = (inp[9]) ? node2745 : node2734;
											assign node2734 = (inp[8]) ? node2742 : node2735;
												assign node2735 = (inp[10]) ? node2739 : node2736;
													assign node2736 = (inp[7]) ? 14'b00010000100000 : 14'b01010000100100;
													assign node2739 = (inp[7]) ? 14'b01110000100000 : 14'b01110100100000;
												assign node2742 = (inp[7]) ? 14'b01010000100100 : 14'b01010100100100;
											assign node2745 = (inp[8]) ? node2753 : node2746;
												assign node2746 = (inp[10]) ? node2750 : node2747;
													assign node2747 = (inp[7]) ? 14'b00010000000000 : 14'b01010000000100;
													assign node2750 = (inp[11]) ? 14'b01110000000000 : 14'b01110100000000;
												assign node2753 = (inp[7]) ? 14'b01010000000100 : 14'b01010100000100;
								assign node2756 = (inp[9]) ? node2804 : node2757;
									assign node2757 = (inp[7]) ? node2781 : node2758;
										assign node2758 = (inp[1]) ? node2770 : node2759;
											assign node2759 = (inp[8]) ? node2767 : node2760;
												assign node2760 = (inp[10]) ? node2764 : node2761;
													assign node2761 = (inp[12]) ? 14'b00110100110100 : 14'b00110100110110;
													assign node2764 = (inp[12]) ? 14'b00110100110000 : 14'b00110100110010;
												assign node2767 = (inp[12]) ? 14'b00010100110100 : 14'b00110100110100;
											assign node2770 = (inp[8]) ? node2778 : node2771;
												assign node2771 = (inp[12]) ? node2775 : node2772;
													assign node2772 = (inp[10]) ? 14'b00110100100010 : 14'b00110100100110;
													assign node2775 = (inp[10]) ? 14'b00110100100000 : 14'b00110100100100;
												assign node2778 = (inp[12]) ? 14'b00010100100100 : 14'b00110100100100;
										assign node2781 = (inp[1]) ? node2793 : node2782;
											assign node2782 = (inp[8]) ? node2790 : node2783;
												assign node2783 = (inp[10]) ? node2787 : node2784;
													assign node2784 = (inp[12]) ? 14'b00110000110100 : 14'b00110000110110;
													assign node2787 = (inp[12]) ? 14'b00110000110000 : 14'b00110000110010;
												assign node2790 = (inp[12]) ? 14'b00010000110100 : 14'b00110000110100;
											assign node2793 = (inp[8]) ? node2801 : node2794;
												assign node2794 = (inp[10]) ? node2798 : node2795;
													assign node2795 = (inp[12]) ? 14'b00110000100100 : 14'b00110000100110;
													assign node2798 = (inp[12]) ? 14'b00110000100000 : 14'b00110000100010;
												assign node2801 = (inp[12]) ? 14'b00010000100100 : 14'b00110000100100;
									assign node2804 = (inp[7]) ? node2828 : node2805;
										assign node2805 = (inp[1]) ? node2817 : node2806;
											assign node2806 = (inp[8]) ? node2814 : node2807;
												assign node2807 = (inp[10]) ? node2811 : node2808;
													assign node2808 = (inp[12]) ? 14'b00110100010100 : 14'b00110100010110;
													assign node2811 = (inp[12]) ? 14'b00110100010000 : 14'b00110100010010;
												assign node2814 = (inp[12]) ? 14'b00010100010100 : 14'b00110100010100;
											assign node2817 = (inp[8]) ? node2825 : node2818;
												assign node2818 = (inp[10]) ? node2822 : node2819;
													assign node2819 = (inp[12]) ? 14'b00110100000100 : 14'b00110100000110;
													assign node2822 = (inp[12]) ? 14'b00110100000000 : 14'b00110100000010;
												assign node2825 = (inp[12]) ? 14'b00010100000100 : 14'b00110100000100;
										assign node2828 = (inp[1]) ? node2840 : node2829;
											assign node2829 = (inp[8]) ? node2837 : node2830;
												assign node2830 = (inp[12]) ? node2834 : node2831;
													assign node2831 = (inp[10]) ? 14'b00110000010010 : 14'b00110000010110;
													assign node2834 = (inp[10]) ? 14'b00110000010000 : 14'b00110000010100;
												assign node2837 = (inp[12]) ? 14'b00010000010100 : 14'b00110000010100;
											assign node2840 = (inp[8]) ? node2848 : node2841;
												assign node2841 = (inp[10]) ? node2845 : node2842;
													assign node2842 = (inp[12]) ? 14'b00110000000100 : 14'b00110000000110;
													assign node2845 = (inp[12]) ? 14'b00110000000000 : 14'b00110000000010;
												assign node2848 = (inp[12]) ? 14'b00010000000100 : 14'b00110000000100;
							assign node2851 = (inp[4]) ? node2949 : node2852;
								assign node2852 = (inp[10]) ? node2916 : node2853;
									assign node2853 = (inp[9]) ? node2885 : node2854;
										assign node2854 = (inp[7]) ? node2870 : node2855;
											assign node2855 = (inp[1]) ? node2863 : node2856;
												assign node2856 = (inp[8]) ? node2860 : node2857;
													assign node2857 = (inp[12]) ? 14'b01110100110100 : 14'b01110100110110;
													assign node2860 = (inp[12]) ? 14'b01010100110000 : 14'b01110100110100;
												assign node2863 = (inp[8]) ? node2867 : node2864;
													assign node2864 = (inp[12]) ? 14'b01110100100100 : 14'b01110100100110;
													assign node2867 = (inp[12]) ? 14'b01010100100000 : 14'b01110100100100;
											assign node2870 = (inp[1]) ? node2878 : node2871;
												assign node2871 = (inp[8]) ? node2875 : node2872;
													assign node2872 = (inp[12]) ? 14'b01110000110100 : 14'b01110000110110;
													assign node2875 = (inp[12]) ? 14'b01010000110000 : 14'b01110000110100;
												assign node2878 = (inp[12]) ? node2882 : node2879;
													assign node2879 = (inp[8]) ? 14'b01110000100100 : 14'b01110000100110;
													assign node2882 = (inp[8]) ? 14'b01010000100000 : 14'b01110000100100;
										assign node2885 = (inp[7]) ? node2901 : node2886;
											assign node2886 = (inp[1]) ? node2894 : node2887;
												assign node2887 = (inp[8]) ? node2891 : node2888;
													assign node2888 = (inp[12]) ? 14'b01110100010100 : 14'b01110100010110;
													assign node2891 = (inp[12]) ? 14'b01010100010000 : 14'b01110100010100;
												assign node2894 = (inp[12]) ? node2898 : node2895;
													assign node2895 = (inp[8]) ? 14'b01110100000100 : 14'b01110100000110;
													assign node2898 = (inp[8]) ? 14'b01010100000000 : 14'b01110100000100;
											assign node2901 = (inp[8]) ? node2909 : node2902;
												assign node2902 = (inp[12]) ? node2906 : node2903;
													assign node2903 = (inp[1]) ? 14'b01110000000110 : 14'b01110000010110;
													assign node2906 = (inp[1]) ? 14'b01110000000100 : 14'b01110000010100;
												assign node2909 = (inp[12]) ? node2913 : node2910;
													assign node2910 = (inp[1]) ? 14'b01110000000100 : 14'b01110000010100;
													assign node2913 = (inp[1]) ? 14'b01010000000000 : 14'b01010000010000;
									assign node2916 = (inp[8]) ? node2918 : 14'b00000000000001;
										assign node2918 = (inp[12]) ? node2934 : node2919;
											assign node2919 = (inp[9]) ? node2927 : node2920;
												assign node2920 = (inp[1]) ? node2924 : node2921;
													assign node2921 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
													assign node2924 = (inp[7]) ? 14'b01110000100100 : 14'b01110100100100;
												assign node2927 = (inp[1]) ? node2931 : node2928;
													assign node2928 = (inp[7]) ? 14'b01110000010100 : 14'b01110100010100;
													assign node2931 = (inp[7]) ? 14'b01110000000100 : 14'b01110100000100;
											assign node2934 = (inp[9]) ? node2942 : node2935;
												assign node2935 = (inp[1]) ? node2939 : node2936;
													assign node2936 = (inp[7]) ? 14'b01010000110000 : 14'b01010100110000;
													assign node2939 = (inp[7]) ? 14'b01010000100000 : 14'b01010100100000;
												assign node2942 = (inp[1]) ? node2946 : node2943;
													assign node2943 = (inp[7]) ? 14'b01010000010000 : 14'b01010100010000;
													assign node2946 = (inp[7]) ? 14'b01010000000000 : 14'b01010100000000;
								assign node2949 = (inp[7]) ? 14'b00000000000001 : node2950;
									assign node2950 = (inp[8]) ? 14'b00000000000001 : node2951;
										assign node2951 = (inp[10]) ? node2959 : node2952;
											assign node2952 = (inp[12]) ? node2954 : 14'b00000000000001;
												assign node2954 = (inp[9]) ? node2956 : 14'b00010100100100;
													assign node2956 = (inp[1]) ? 14'b00010100000100 : 14'b00010100010100;
											assign node2959 = (inp[12]) ? node2967 : node2960;
												assign node2960 = (inp[9]) ? node2964 : node2961;
													assign node2961 = (inp[1]) ? 14'b00010100100010 : 14'b00010100110010;
													assign node2964 = (inp[1]) ? 14'b00010100000010 : 14'b00010100010010;
												assign node2967 = (inp[9]) ? node2971 : node2968;
													assign node2968 = (inp[1]) ? 14'b00010100100000 : 14'b00010100110000;
													assign node2971 = (inp[1]) ? 14'b00010100000000 : 14'b00010100010000;
						assign node2976 = (inp[2]) ? node2978 : 14'b00000000000001;
							assign node2978 = (inp[9]) ? 14'b00000000000001 : node2979;
								assign node2979 = (inp[12]) ? 14'b00000000000001 : node2980;
									assign node2980 = (inp[4]) ? node2990 : node2981;
										assign node2981 = (inp[8]) ? 14'b00000000000001 : node2982;
											assign node2982 = (inp[7]) ? 14'b00000000000001 : node2983;
												assign node2983 = (inp[1]) ? 14'b00000000000001 : node2984;
													assign node2984 = (inp[10]) ? 14'b10000001001000 : 14'b00000000000001;
										assign node2990 = (inp[7]) ? node2998 : node2991;
											assign node2991 = (inp[1]) ? 14'b00000000000001 : node2992;
												assign node2992 = (inp[10]) ? node2994 : 14'b10000001001010;
													assign node2994 = (inp[8]) ? 14'b10000001001010 : 14'b00000000000001;
											assign node2998 = (inp[1]) ? node3000 : 14'b00000000000001;
												assign node3000 = (inp[10]) ? 14'b10000000000000 : node3001;
													assign node3001 = (inp[8]) ? 14'b10000000000000 : 14'b00000000000001;
				assign node3007 = (inp[12]) ? node3321 : node3008;
					assign node3008 = (inp[2]) ? node3198 : node3009;
						assign node3009 = (inp[8]) ? node3105 : node3010;
							assign node3010 = (inp[10]) ? 14'b00000000000001 : node3011;
								assign node3011 = (inp[6]) ? node3071 : node3012;
									assign node3012 = (inp[4]) ? node3042 : node3013;
										assign node3013 = (inp[9]) ? node3027 : node3014;
											assign node3014 = (inp[3]) ? node3020 : node3015;
												assign node3015 = (inp[1]) ? node3017 : 14'b00000000000001;
													assign node3017 = (inp[7]) ? 14'b01010010100110 : 14'b01010110100110;
												assign node3020 = (inp[1]) ? node3024 : node3021;
													assign node3021 = (inp[7]) ? 14'b01010010110110 : 14'b01010110110110;
													assign node3024 = (inp[7]) ? 14'b01000010100110 : 14'b01000110100110;
											assign node3027 = (inp[7]) ? node3035 : node3028;
												assign node3028 = (inp[1]) ? node3032 : node3029;
													assign node3029 = (inp[3]) ? 14'b01010110010110 : 14'b01000100000110;
													assign node3032 = (inp[3]) ? 14'b01000110000110 : 14'b01010110000110;
												assign node3035 = (inp[1]) ? node3039 : node3036;
													assign node3036 = (inp[3]) ? 14'b01010010010110 : 14'b01000000000110;
													assign node3039 = (inp[3]) ? 14'b01000010000110 : 14'b01010010000110;
										assign node3042 = (inp[3]) ? node3056 : node3043;
											assign node3043 = (inp[1]) ? node3049 : node3044;
												assign node3044 = (inp[9]) ? node3046 : 14'b00000000000001;
													assign node3046 = (inp[7]) ? 14'b00000000000110 : 14'b00000100000110;
												assign node3049 = (inp[9]) ? node3053 : node3050;
													assign node3050 = (inp[7]) ? 14'b00010010100110 : 14'b00010110100110;
													assign node3053 = (inp[7]) ? 14'b00010010000110 : 14'b00010110000110;
											assign node3056 = (inp[1]) ? node3064 : node3057;
												assign node3057 = (inp[9]) ? node3061 : node3058;
													assign node3058 = (inp[7]) ? 14'b00010010110110 : 14'b00010110110110;
													assign node3061 = (inp[7]) ? 14'b00010010010110 : 14'b00010110010110;
												assign node3064 = (inp[9]) ? node3068 : node3065;
													assign node3065 = (inp[7]) ? 14'b00000010100110 : 14'b00000110100110;
													assign node3068 = (inp[7]) ? 14'b00000010000110 : 14'b00000110000110;
									assign node3071 = (inp[3]) ? 14'b00000000000001 : node3072;
										assign node3072 = (inp[1]) ? node3088 : node3073;
											assign node3073 = (inp[7]) ? node3081 : node3074;
												assign node3074 = (inp[4]) ? node3078 : node3075;
													assign node3075 = (inp[9]) ? 14'b01010100010110 : 14'b01010100110110;
													assign node3078 = (inp[9]) ? 14'b00010100010110 : 14'b00010100110110;
												assign node3081 = (inp[9]) ? node3085 : node3082;
													assign node3082 = (inp[4]) ? 14'b00010000110110 : 14'b01010000110110;
													assign node3085 = (inp[4]) ? 14'b00010000010110 : 14'b01010000010110;
											assign node3088 = (inp[9]) ? node3096 : node3089;
												assign node3089 = (inp[7]) ? node3093 : node3090;
													assign node3090 = (inp[4]) ? 14'b00010100100110 : 14'b01010100100110;
													assign node3093 = (inp[4]) ? 14'b00010000100110 : 14'b01010000100110;
												assign node3096 = (inp[7]) ? node3100 : node3097;
													assign node3097 = (inp[4]) ? 14'b00010100000110 : 14'b01010100000110;
													assign node3100 = (inp[4]) ? 14'b00010000000110 : 14'b01010000000110;
							assign node3105 = (inp[6]) ? node3165 : node3106;
								assign node3106 = (inp[7]) ? node3136 : node3107;
									assign node3107 = (inp[3]) ? node3121 : node3108;
										assign node3108 = (inp[1]) ? node3114 : node3109;
											assign node3109 = (inp[9]) ? node3111 : 14'b00000000000001;
												assign node3111 = (inp[4]) ? 14'b00100100000000 : 14'b01100100000000;
											assign node3114 = (inp[9]) ? node3118 : node3115;
												assign node3115 = (inp[4]) ? 14'b00110110100000 : 14'b01110110100000;
												assign node3118 = (inp[4]) ? 14'b00110110000000 : 14'b01110110000000;
										assign node3121 = (inp[1]) ? node3129 : node3122;
											assign node3122 = (inp[9]) ? node3126 : node3123;
												assign node3123 = (inp[4]) ? 14'b00110110110000 : 14'b01110110110000;
												assign node3126 = (inp[4]) ? 14'b00110110010000 : 14'b01110110010000;
											assign node3129 = (inp[4]) ? node3133 : node3130;
												assign node3130 = (inp[9]) ? 14'b01100110000000 : 14'b01100110100000;
												assign node3133 = (inp[9]) ? 14'b00100110000000 : 14'b00100110100000;
									assign node3136 = (inp[3]) ? node3150 : node3137;
										assign node3137 = (inp[1]) ? node3143 : node3138;
											assign node3138 = (inp[9]) ? node3140 : 14'b00000000000001;
												assign node3140 = (inp[4]) ? 14'b00100000000000 : 14'b01100000000000;
											assign node3143 = (inp[9]) ? node3147 : node3144;
												assign node3144 = (inp[4]) ? 14'b00110010100000 : 14'b01110010100000;
												assign node3147 = (inp[4]) ? 14'b00110010000000 : 14'b01110010000000;
										assign node3150 = (inp[1]) ? node3158 : node3151;
											assign node3151 = (inp[9]) ? node3155 : node3152;
												assign node3152 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110000;
												assign node3155 = (inp[4]) ? 14'b00110010010000 : 14'b01110010010000;
											assign node3158 = (inp[9]) ? node3162 : node3159;
												assign node3159 = (inp[4]) ? 14'b00100010100000 : 14'b01100010100000;
												assign node3162 = (inp[4]) ? 14'b00100010000000 : 14'b01100010000000;
								assign node3165 = (inp[3]) ? 14'b00000000000001 : node3166;
									assign node3166 = (inp[1]) ? node3182 : node3167;
										assign node3167 = (inp[9]) ? node3175 : node3168;
											assign node3168 = (inp[7]) ? node3172 : node3169;
												assign node3169 = (inp[4]) ? 14'b00110100110000 : 14'b01110100110000;
												assign node3172 = (inp[4]) ? 14'b00110000110000 : 14'b01110000110000;
											assign node3175 = (inp[4]) ? node3179 : node3176;
												assign node3176 = (inp[7]) ? 14'b01110000010000 : 14'b01110100010000;
												assign node3179 = (inp[7]) ? 14'b00110000010000 : 14'b00110100010000;
										assign node3182 = (inp[4]) ? node3190 : node3183;
											assign node3183 = (inp[7]) ? node3187 : node3184;
												assign node3184 = (inp[9]) ? 14'b01110100000000 : 14'b01110100100000;
												assign node3187 = (inp[9]) ? 14'b01110000000000 : 14'b01110000100000;
											assign node3190 = (inp[9]) ? node3194 : node3191;
												assign node3191 = (inp[7]) ? 14'b00110000100000 : 14'b00110100100000;
												assign node3194 = (inp[7]) ? 14'b00110000000000 : 14'b00110100000000;
						assign node3198 = (inp[7]) ? 14'b00000000000001 : node3199;
							assign node3199 = (inp[10]) ? node3283 : node3200;
								assign node3200 = (inp[8]) ? node3248 : node3201;
									assign node3201 = (inp[6]) ? node3231 : node3202;
										assign node3202 = (inp[1]) ? node3216 : node3203;
											assign node3203 = (inp[3]) ? node3209 : node3204;
												assign node3204 = (inp[9]) ? node3206 : 14'b00000000000001;
													assign node3206 = (inp[4]) ? 14'b01000000000010 : 14'b01000100000010;
												assign node3209 = (inp[9]) ? node3213 : node3210;
													assign node3210 = (inp[4]) ? 14'b01010010110010 : 14'b01010110110010;
													assign node3213 = (inp[4]) ? 14'b01010010010010 : 14'b01010110010010;
											assign node3216 = (inp[4]) ? node3224 : node3217;
												assign node3217 = (inp[9]) ? node3221 : node3218;
													assign node3218 = (inp[3]) ? 14'b01000110100010 : 14'b01010110100010;
													assign node3221 = (inp[3]) ? 14'b01000110000010 : 14'b01010110000010;
												assign node3224 = (inp[3]) ? node3228 : node3225;
													assign node3225 = (inp[9]) ? 14'b01010010000010 : 14'b01010010100010;
													assign node3228 = (inp[9]) ? 14'b01000010000010 : 14'b01000010100010;
										assign node3231 = (inp[3]) ? 14'b00000000000001 : node3232;
											assign node3232 = (inp[1]) ? node3240 : node3233;
												assign node3233 = (inp[9]) ? node3237 : node3234;
													assign node3234 = (inp[4]) ? 14'b01010000110010 : 14'b01010100110010;
													assign node3237 = (inp[4]) ? 14'b01010000010010 : 14'b01010100010010;
												assign node3240 = (inp[4]) ? node3244 : node3241;
													assign node3241 = (inp[9]) ? 14'b01010100000010 : 14'b01010100100010;
													assign node3244 = (inp[9]) ? 14'b01010000000010 : 14'b01010000100010;
									assign node3248 = (inp[4]) ? node3258 : node3249;
										assign node3249 = (inp[3]) ? node3251 : 14'b00000000000001;
											assign node3251 = (inp[6]) ? node3253 : 14'b00000000000001;
												assign node3253 = (inp[1]) ? 14'b00000000000001 : node3254;
													assign node3254 = (inp[9]) ? 14'b00000000000001 : 14'b10000001001000;
										assign node3258 = (inp[3]) ? node3274 : node3259;
											assign node3259 = (inp[1]) ? node3267 : node3260;
												assign node3260 = (inp[6]) ? node3264 : node3261;
													assign node3261 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
													assign node3264 = (inp[9]) ? 14'b00010100010000 : 14'b00010100110000;
												assign node3267 = (inp[6]) ? node3271 : node3268;
													assign node3268 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
													assign node3271 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
											assign node3274 = (inp[6]) ? 14'b00000000000001 : node3275;
												assign node3275 = (inp[1]) ? node3279 : node3276;
													assign node3276 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
													assign node3279 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
								assign node3283 = (inp[8]) ? node3285 : 14'b00000000000001;
									assign node3285 = (inp[4]) ? node3295 : node3286;
										assign node3286 = (inp[3]) ? node3288 : 14'b00000000000001;
											assign node3288 = (inp[9]) ? 14'b00000000000001 : node3289;
												assign node3289 = (inp[6]) ? node3291 : 14'b00000000000001;
													assign node3291 = (inp[1]) ? 14'b00000000000001 : 14'b10000001001000;
										assign node3295 = (inp[6]) ? node3311 : node3296;
											assign node3296 = (inp[9]) ? node3304 : node3297;
												assign node3297 = (inp[3]) ? node3301 : node3298;
													assign node3298 = (inp[1]) ? 14'b00010110100000 : 14'b00000000000001;
													assign node3301 = (inp[1]) ? 14'b00000110100000 : 14'b00010110110000;
												assign node3304 = (inp[3]) ? node3308 : node3305;
													assign node3305 = (inp[1]) ? 14'b00010110000000 : 14'b00000100000000;
													assign node3308 = (inp[1]) ? 14'b00000110000000 : 14'b00010110010000;
											assign node3311 = (inp[3]) ? 14'b00000000000001 : node3312;
												assign node3312 = (inp[1]) ? node3316 : node3313;
													assign node3313 = (inp[9]) ? 14'b00010100010000 : 14'b00010100110000;
													assign node3316 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
					assign node3321 = (inp[10]) ? node3453 : node3322;
						assign node3322 = (inp[8]) ? node3430 : node3323;
							assign node3323 = (inp[4]) ? node3401 : node3324;
								assign node3324 = (inp[7]) ? node3374 : node3325;
									assign node3325 = (inp[6]) ? node3357 : node3326;
										assign node3326 = (inp[2]) ? node3342 : node3327;
											assign node3327 = (inp[3]) ? node3335 : node3328;
												assign node3328 = (inp[1]) ? node3332 : node3329;
													assign node3329 = (inp[9]) ? 14'b01000100000100 : 14'b00000000000001;
													assign node3332 = (inp[9]) ? 14'b01010110000100 : 14'b01010110100100;
												assign node3335 = (inp[1]) ? node3339 : node3336;
													assign node3336 = (inp[9]) ? 14'b01010110010100 : 14'b01010110110100;
													assign node3339 = (inp[9]) ? 14'b01000110000100 : 14'b01000110100100;
											assign node3342 = (inp[1]) ? node3350 : node3343;
												assign node3343 = (inp[3]) ? node3347 : node3344;
													assign node3344 = (inp[9]) ? 14'b01000100000000 : 14'b00000000000001;
													assign node3347 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
												assign node3350 = (inp[3]) ? node3354 : node3351;
													assign node3351 = (inp[9]) ? 14'b01010110000000 : 14'b01010110100000;
													assign node3354 = (inp[9]) ? 14'b01000110000000 : 14'b01000110100000;
										assign node3357 = (inp[3]) ? 14'b00000000000001 : node3358;
											assign node3358 = (inp[1]) ? node3366 : node3359;
												assign node3359 = (inp[2]) ? node3363 : node3360;
													assign node3360 = (inp[9]) ? 14'b01010100010100 : 14'b01010100110100;
													assign node3363 = (inp[9]) ? 14'b01010100010000 : 14'b01010100110000;
												assign node3366 = (inp[2]) ? node3370 : node3367;
													assign node3367 = (inp[9]) ? 14'b01010100000100 : 14'b01010100100100;
													assign node3370 = (inp[9]) ? 14'b01010100000000 : 14'b01010100100000;
									assign node3374 = (inp[2]) ? node3376 : 14'b00000000000001;
										assign node3376 = (inp[6]) ? node3392 : node3377;
											assign node3377 = (inp[3]) ? node3385 : node3378;
												assign node3378 = (inp[1]) ? node3382 : node3379;
													assign node3379 = (inp[9]) ? 14'b01000000000000 : 14'b00000000000001;
													assign node3382 = (inp[9]) ? 14'b01010010000000 : 14'b01010010100000;
												assign node3385 = (inp[1]) ? node3389 : node3386;
													assign node3386 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
													assign node3389 = (inp[9]) ? 14'b01000010000000 : 14'b01000010100000;
											assign node3392 = (inp[3]) ? 14'b00000000000001 : node3393;
												assign node3393 = (inp[9]) ? node3397 : node3394;
													assign node3394 = (inp[1]) ? 14'b01010000100000 : 14'b01010000110000;
													assign node3397 = (inp[1]) ? 14'b01010000000000 : 14'b01010000010000;
								assign node3401 = (inp[2]) ? 14'b00000000000001 : node3402;
									assign node3402 = (inp[7]) ? node3404 : 14'b00000000000001;
										assign node3404 = (inp[6]) ? node3420 : node3405;
											assign node3405 = (inp[1]) ? node3413 : node3406;
												assign node3406 = (inp[3]) ? node3410 : node3407;
													assign node3407 = (inp[9]) ? 14'b00000000000100 : 14'b00000000000001;
													assign node3410 = (inp[9]) ? 14'b00010010010100 : 14'b00010010110100;
												assign node3413 = (inp[9]) ? node3417 : node3414;
													assign node3414 = (inp[3]) ? 14'b00000010100100 : 14'b00010010100100;
													assign node3417 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
											assign node3420 = (inp[3]) ? 14'b00000000000001 : node3421;
												assign node3421 = (inp[9]) ? node3425 : node3422;
													assign node3422 = (inp[1]) ? 14'b00010000100100 : 14'b00010000110100;
													assign node3425 = (inp[1]) ? 14'b00010000000100 : 14'b00010000010100;
							assign node3430 = (inp[1]) ? 14'b00000000000001 : node3431;
								assign node3431 = (inp[9]) ? 14'b00000000000001 : node3432;
									assign node3432 = (inp[3]) ? node3442 : node3433;
										assign node3433 = (inp[2]) ? node3435 : 14'b00000000000001;
											assign node3435 = (inp[6]) ? 14'b00000000000001 : node3436;
												assign node3436 = (inp[7]) ? node3438 : 14'b00000000000001;
													assign node3438 = (inp[4]) ? 14'b10001001000010 : 14'b10001000001000;
										assign node3442 = (inp[7]) ? 14'b00000000000001 : node3443;
											assign node3443 = (inp[2]) ? 14'b00000000000001 : node3444;
												assign node3444 = (inp[4]) ? 14'b00000000000001 : node3445;
													assign node3445 = (inp[6]) ? 14'b10001000000010 : 14'b00000000000001;
						assign node3453 = (inp[9]) ? 14'b00000000000001 : node3454;
							assign node3454 = (inp[8]) ? node3456 : 14'b00000000000001;
								assign node3456 = (inp[1]) ? 14'b00000000000001 : node3457;
									assign node3457 = (inp[4]) ? node3473 : node3458;
										assign node3458 = (inp[3]) ? node3466 : node3459;
											assign node3459 = (inp[7]) ? node3461 : 14'b00000000000001;
												assign node3461 = (inp[6]) ? 14'b00000000000001 : node3462;
													assign node3462 = (inp[2]) ? 14'b10001000001000 : 14'b00000000000001;
											assign node3466 = (inp[2]) ? 14'b00000000000001 : node3467;
												assign node3467 = (inp[7]) ? 14'b00000000000001 : node3468;
													assign node3468 = (inp[6]) ? 14'b10001000000010 : 14'b00000000000001;
										assign node3473 = (inp[2]) ? node3475 : 14'b00000000000001;
											assign node3475 = (inp[6]) ? 14'b00000000000001 : node3476;
												assign node3476 = (inp[3]) ? 14'b00000000000001 : node3477;
													assign node3477 = (inp[7]) ? 14'b10001001000010 : 14'b00000000000001;
			assign node3484 = (inp[1]) ? node4086 : node3485;
				assign node3485 = (inp[3]) ? node3929 : node3486;
					assign node3486 = (inp[5]) ? node3786 : node3487;
						assign node3487 = (inp[2]) ? node3663 : node3488;
							assign node3488 = (inp[4]) ? node3570 : node3489;
								assign node3489 = (inp[12]) ? node3523 : node3490;
									assign node3490 = (inp[7]) ? node3502 : node3491;
										assign node3491 = (inp[8]) ? 14'b00000000000001 : node3492;
											assign node3492 = (inp[10]) ? node3494 : 14'b00000000000001;
												assign node3494 = (inp[9]) ? node3498 : node3495;
													assign node3495 = (inp[6]) ? 14'b01100100110010 : 14'b01100110110010;
													assign node3498 = (inp[6]) ? 14'b01100100010010 : 14'b01100110010010;
										assign node3502 = (inp[8]) ? node3516 : node3503;
											assign node3503 = (inp[10]) ? node3511 : node3504;
												assign node3504 = (inp[9]) ? node3508 : node3505;
													assign node3505 = (inp[6]) ? 14'b00000000110010 : 14'b00000010110010;
													assign node3508 = (inp[6]) ? 14'b00000000010010 : 14'b00000010010010;
												assign node3511 = (inp[6]) ? 14'b01100000010010 : node3512;
													assign node3512 = (inp[9]) ? 14'b01100010010010 : 14'b01100010110010;
											assign node3516 = (inp[9]) ? node3520 : node3517;
												assign node3517 = (inp[6]) ? 14'b00000000110000 : 14'b00000010110000;
												assign node3520 = (inp[6]) ? 14'b00000000010000 : 14'b00000010010000;
									assign node3523 = (inp[6]) ? node3547 : node3524;
										assign node3524 = (inp[9]) ? node3536 : node3525;
											assign node3525 = (inp[8]) ? node3533 : node3526;
												assign node3526 = (inp[10]) ? node3530 : node3527;
													assign node3527 = (inp[7]) ? 14'b00000010110000 : 14'b01000010110100;
													assign node3530 = (inp[7]) ? 14'b01100010110000 : 14'b01100110110000;
												assign node3533 = (inp[7]) ? 14'b01000010110100 : 14'b01000110110100;
											assign node3536 = (inp[8]) ? node3544 : node3537;
												assign node3537 = (inp[10]) ? node3541 : node3538;
													assign node3538 = (inp[7]) ? 14'b00000010010000 : 14'b01000010010100;
													assign node3541 = (inp[7]) ? 14'b01100010010000 : 14'b01100110010000;
												assign node3544 = (inp[7]) ? 14'b01000010010100 : 14'b01000110010100;
										assign node3547 = (inp[9]) ? node3559 : node3548;
											assign node3548 = (inp[8]) ? node3556 : node3549;
												assign node3549 = (inp[10]) ? node3553 : node3550;
													assign node3550 = (inp[7]) ? 14'b00000000110000 : 14'b01000000110100;
													assign node3553 = (inp[7]) ? 14'b01100000110000 : 14'b01100100110000;
												assign node3556 = (inp[7]) ? 14'b01000000110100 : 14'b01000100110100;
											assign node3559 = (inp[8]) ? node3567 : node3560;
												assign node3560 = (inp[10]) ? node3564 : node3561;
													assign node3561 = (inp[7]) ? 14'b00000000010000 : 14'b01000000010100;
													assign node3564 = (inp[7]) ? 14'b01100000010000 : 14'b01100100010000;
												assign node3567 = (inp[7]) ? 14'b01000000010100 : 14'b01000100010100;
								assign node3570 = (inp[6]) ? node3618 : node3571;
									assign node3571 = (inp[9]) ? node3595 : node3572;
										assign node3572 = (inp[7]) ? node3584 : node3573;
											assign node3573 = (inp[8]) ? node3581 : node3574;
												assign node3574 = (inp[10]) ? node3578 : node3575;
													assign node3575 = (inp[12]) ? 14'b00100110110100 : 14'b00100110110110;
													assign node3578 = (inp[12]) ? 14'b00100110110000 : 14'b00100110110010;
												assign node3581 = (inp[12]) ? 14'b00000110110100 : 14'b00100110110100;
											assign node3584 = (inp[8]) ? node3592 : node3585;
												assign node3585 = (inp[12]) ? node3589 : node3586;
													assign node3586 = (inp[10]) ? 14'b00100010110010 : 14'b00100010110110;
													assign node3589 = (inp[10]) ? 14'b00100010110000 : 14'b00100010110100;
												assign node3592 = (inp[12]) ? 14'b00000010110100 : 14'b00100010110100;
										assign node3595 = (inp[7]) ? node3607 : node3596;
											assign node3596 = (inp[8]) ? node3604 : node3597;
												assign node3597 = (inp[10]) ? node3601 : node3598;
													assign node3598 = (inp[12]) ? 14'b00100110010100 : 14'b00100110010110;
													assign node3601 = (inp[12]) ? 14'b00100110010000 : 14'b00100110010010;
												assign node3604 = (inp[12]) ? 14'b00000110010100 : 14'b00100110010100;
											assign node3607 = (inp[8]) ? node3615 : node3608;
												assign node3608 = (inp[10]) ? node3612 : node3609;
													assign node3609 = (inp[12]) ? 14'b00100010010100 : 14'b00100010010110;
													assign node3612 = (inp[12]) ? 14'b00100010010000 : 14'b00100010010010;
												assign node3615 = (inp[12]) ? 14'b00000010010100 : 14'b00100010010100;
									assign node3618 = (inp[7]) ? node3640 : node3619;
										assign node3619 = (inp[9]) ? node3631 : node3620;
											assign node3620 = (inp[8]) ? node3628 : node3621;
												assign node3621 = (inp[10]) ? node3625 : node3622;
													assign node3622 = (inp[12]) ? 14'b00100100110100 : 14'b00100100110110;
													assign node3625 = (inp[12]) ? 14'b00100100110000 : 14'b00100100110010;
												assign node3628 = (inp[12]) ? 14'b00000100110100 : 14'b00100100110100;
											assign node3631 = (inp[8]) ? node3637 : node3632;
												assign node3632 = (inp[12]) ? 14'b00100100010100 : node3633;
													assign node3633 = (inp[10]) ? 14'b00100100010010 : 14'b00100100010110;
												assign node3637 = (inp[12]) ? 14'b00000100010100 : 14'b00100100010100;
										assign node3640 = (inp[9]) ? node3652 : node3641;
											assign node3641 = (inp[8]) ? node3649 : node3642;
												assign node3642 = (inp[12]) ? node3646 : node3643;
													assign node3643 = (inp[10]) ? 14'b00100000110010 : 14'b00100000110110;
													assign node3646 = (inp[10]) ? 14'b00100000110000 : 14'b00100000110100;
												assign node3649 = (inp[12]) ? 14'b00000000110100 : 14'b00100000110100;
											assign node3652 = (inp[8]) ? node3660 : node3653;
												assign node3653 = (inp[12]) ? node3657 : node3654;
													assign node3654 = (inp[10]) ? 14'b00100000010010 : 14'b00100000010110;
													assign node3657 = (inp[10]) ? 14'b00100000010000 : 14'b00100000010100;
												assign node3660 = (inp[12]) ? 14'b00000000010100 : 14'b00100000010100;
							assign node3663 = (inp[4]) ? node3757 : node3664;
								assign node3664 = (inp[10]) ? node3728 : node3665;
									assign node3665 = (inp[6]) ? node3697 : node3666;
										assign node3666 = (inp[9]) ? node3682 : node3667;
											assign node3667 = (inp[7]) ? node3675 : node3668;
												assign node3668 = (inp[12]) ? node3672 : node3669;
													assign node3669 = (inp[8]) ? 14'b01100110110100 : 14'b01100110110110;
													assign node3672 = (inp[8]) ? 14'b01000110110000 : 14'b01100110110100;
												assign node3675 = (inp[12]) ? node3679 : node3676;
													assign node3676 = (inp[8]) ? 14'b01100010110100 : 14'b01100010110110;
													assign node3679 = (inp[8]) ? 14'b01000010110000 : 14'b01100010110100;
											assign node3682 = (inp[7]) ? node3690 : node3683;
												assign node3683 = (inp[8]) ? node3687 : node3684;
													assign node3684 = (inp[12]) ? 14'b01100110010100 : 14'b01100110010110;
													assign node3687 = (inp[12]) ? 14'b01000110010000 : 14'b01100110010100;
												assign node3690 = (inp[8]) ? node3694 : node3691;
													assign node3691 = (inp[12]) ? 14'b01100010010100 : 14'b01100010010110;
													assign node3694 = (inp[12]) ? 14'b01000010010000 : 14'b01100010010100;
										assign node3697 = (inp[9]) ? node3713 : node3698;
											assign node3698 = (inp[7]) ? node3706 : node3699;
												assign node3699 = (inp[12]) ? node3703 : node3700;
													assign node3700 = (inp[8]) ? 14'b01100100110100 : 14'b01100100110110;
													assign node3703 = (inp[8]) ? 14'b01000100110000 : 14'b01100100110100;
												assign node3706 = (inp[12]) ? node3710 : node3707;
													assign node3707 = (inp[8]) ? 14'b01100000110100 : 14'b01100000110110;
													assign node3710 = (inp[8]) ? 14'b01000000110000 : 14'b01100000110100;
											assign node3713 = (inp[7]) ? node3721 : node3714;
												assign node3714 = (inp[12]) ? node3718 : node3715;
													assign node3715 = (inp[8]) ? 14'b01100100010100 : 14'b01100100010110;
													assign node3718 = (inp[8]) ? 14'b01000100010000 : 14'b01100100010100;
												assign node3721 = (inp[12]) ? node3725 : node3722;
													assign node3722 = (inp[8]) ? 14'b01100000010100 : 14'b01100000010110;
													assign node3725 = (inp[8]) ? 14'b01000000010000 : 14'b01100000010100;
									assign node3728 = (inp[8]) ? node3730 : 14'b00000000000001;
										assign node3730 = (inp[12]) ? node3744 : node3731;
											assign node3731 = (inp[6]) ? node3737 : node3732;
												assign node3732 = (inp[9]) ? node3734 : 14'b01100110110100;
													assign node3734 = (inp[7]) ? 14'b01100010010100 : 14'b01100110010100;
												assign node3737 = (inp[9]) ? node3741 : node3738;
													assign node3738 = (inp[7]) ? 14'b01100000110100 : 14'b01100100110100;
													assign node3741 = (inp[7]) ? 14'b01100000010100 : 14'b01100100010100;
											assign node3744 = (inp[7]) ? node3752 : node3745;
												assign node3745 = (inp[9]) ? node3749 : node3746;
													assign node3746 = (inp[6]) ? 14'b01000100110000 : 14'b01000110110000;
													assign node3749 = (inp[11]) ? 14'b01000110010000 : 14'b01000100010000;
												assign node3752 = (inp[9]) ? 14'b01000010010000 : node3753;
													assign node3753 = (inp[6]) ? 14'b01000000110000 : 14'b01000010110000;
								assign node3757 = (inp[8]) ? 14'b00000000000001 : node3758;
									assign node3758 = (inp[7]) ? 14'b00000000000001 : node3759;
										assign node3759 = (inp[12]) ? node3769 : node3760;
											assign node3760 = (inp[10]) ? node3762 : 14'b00000000000001;
												assign node3762 = (inp[6]) ? node3766 : node3763;
													assign node3763 = (inp[9]) ? 14'b00000110010010 : 14'b00000110110010;
													assign node3766 = (inp[9]) ? 14'b00000100010010 : 14'b00000100110010;
											assign node3769 = (inp[6]) ? node3777 : node3770;
												assign node3770 = (inp[9]) ? node3774 : node3771;
													assign node3771 = (inp[10]) ? 14'b00000110110000 : 14'b00000110110100;
													assign node3774 = (inp[10]) ? 14'b00000110010000 : 14'b00000110010100;
												assign node3777 = (inp[9]) ? node3781 : node3778;
													assign node3778 = (inp[10]) ? 14'b00000100110000 : 14'b00000100110100;
													assign node3781 = (inp[10]) ? 14'b00000100010000 : 14'b00000100010100;
						assign node3786 = (inp[12]) ? node3890 : node3787;
							assign node3787 = (inp[2]) ? node3853 : node3788;
								assign node3788 = (inp[8]) ? node3822 : node3789;
									assign node3789 = (inp[10]) ? 14'b00000000000001 : node3790;
										assign node3790 = (inp[4]) ? node3806 : node3791;
											assign node3791 = (inp[7]) ? node3799 : node3792;
												assign node3792 = (inp[9]) ? node3796 : node3793;
													assign node3793 = (inp[6]) ? 14'b01000100110110 : 14'b01000110110110;
													assign node3796 = (inp[6]) ? 14'b01000100010110 : 14'b01000110010110;
												assign node3799 = (inp[6]) ? node3803 : node3800;
													assign node3800 = (inp[9]) ? 14'b01000010010110 : 14'b01000010110110;
													assign node3803 = (inp[9]) ? 14'b01000000010110 : 14'b01000000110110;
											assign node3806 = (inp[7]) ? node3814 : node3807;
												assign node3807 = (inp[6]) ? node3811 : node3808;
													assign node3808 = (inp[9]) ? 14'b00000110010110 : 14'b00000110110110;
													assign node3811 = (inp[9]) ? 14'b00000100010110 : 14'b00000100110110;
												assign node3814 = (inp[9]) ? node3818 : node3815;
													assign node3815 = (inp[6]) ? 14'b00000000110110 : 14'b00000010110110;
													assign node3818 = (inp[6]) ? 14'b00000000010110 : 14'b00000010010110;
									assign node3822 = (inp[4]) ? node3838 : node3823;
										assign node3823 = (inp[9]) ? node3831 : node3824;
											assign node3824 = (inp[7]) ? node3828 : node3825;
												assign node3825 = (inp[6]) ? 14'b01100100110000 : 14'b01100110110000;
												assign node3828 = (inp[6]) ? 14'b01100000110000 : 14'b01100010110000;
											assign node3831 = (inp[7]) ? node3835 : node3832;
												assign node3832 = (inp[6]) ? 14'b01100100010000 : 14'b01100110010000;
												assign node3835 = (inp[6]) ? 14'b01100000010000 : 14'b01100010010000;
										assign node3838 = (inp[7]) ? node3846 : node3839;
											assign node3839 = (inp[6]) ? node3843 : node3840;
												assign node3840 = (inp[9]) ? 14'b00100110010000 : 14'b00100110110000;
												assign node3843 = (inp[9]) ? 14'b00100100010000 : 14'b00100100110000;
											assign node3846 = (inp[6]) ? node3850 : node3847;
												assign node3847 = (inp[9]) ? 14'b00100010010000 : 14'b00100010110000;
												assign node3850 = (inp[9]) ? 14'b00100000010000 : 14'b00100000110000;
								assign node3853 = (inp[7]) ? 14'b00000000000001 : node3854;
									assign node3854 = (inp[10]) ? node3878 : node3855;
										assign node3855 = (inp[8]) ? node3869 : node3856;
											assign node3856 = (inp[4]) ? node3862 : node3857;
												assign node3857 = (inp[6]) ? 14'b01000100010010 : node3858;
													assign node3858 = (inp[9]) ? 14'b01000110010010 : 14'b01000110110010;
												assign node3862 = (inp[9]) ? node3866 : node3863;
													assign node3863 = (inp[6]) ? 14'b01000000110010 : 14'b01000010110010;
													assign node3866 = (inp[6]) ? 14'b01000000010010 : 14'b01000010010010;
											assign node3869 = (inp[4]) ? node3871 : 14'b00000000000001;
												assign node3871 = (inp[6]) ? node3875 : node3872;
													assign node3872 = (inp[9]) ? 14'b00000110010000 : 14'b00000110110000;
													assign node3875 = (inp[9]) ? 14'b00000100010000 : 14'b00000100110000;
										assign node3878 = (inp[4]) ? node3880 : 14'b00000000000001;
											assign node3880 = (inp[8]) ? node3882 : 14'b00000000000001;
												assign node3882 = (inp[9]) ? node3886 : node3883;
													assign node3883 = (inp[6]) ? 14'b00000100110000 : 14'b00000110110000;
													assign node3886 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
							assign node3890 = (inp[8]) ? 14'b00000000000001 : node3891;
								assign node3891 = (inp[10]) ? 14'b00000000000001 : node3892;
									assign node3892 = (inp[4]) ? node3916 : node3893;
										assign node3893 = (inp[7]) ? node3907 : node3894;
											assign node3894 = (inp[6]) ? node3902 : node3895;
												assign node3895 = (inp[2]) ? node3899 : node3896;
													assign node3896 = (inp[9]) ? 14'b01000110010100 : 14'b01000110110100;
													assign node3899 = (inp[9]) ? 14'b01000110010000 : 14'b01000110110000;
												assign node3902 = (inp[9]) ? 14'b01000100010000 : node3903;
													assign node3903 = (inp[2]) ? 14'b01000100110000 : 14'b01000100110100;
											assign node3907 = (inp[2]) ? node3909 : 14'b00000000000001;
												assign node3909 = (inp[9]) ? node3913 : node3910;
													assign node3910 = (inp[6]) ? 14'b01000000110000 : 14'b01000010110000;
													assign node3913 = (inp[6]) ? 14'b01000000010000 : 14'b01000010010000;
										assign node3916 = (inp[2]) ? 14'b00000000000001 : node3917;
											assign node3917 = (inp[7]) ? node3919 : 14'b00000000000001;
												assign node3919 = (inp[9]) ? node3923 : node3920;
													assign node3920 = (inp[6]) ? 14'b00000000110100 : 14'b00000010110100;
													assign node3923 = (inp[6]) ? 14'b00000000010100 : 14'b00000010010100;
					assign node3929 = (inp[9]) ? 14'b00000000000001 : node3930;
						assign node3930 = (inp[6]) ? node3948 : node3931;
							assign node3931 = (inp[7]) ? 14'b00000000000001 : node3932;
								assign node3932 = (inp[4]) ? 14'b00000000000001 : node3933;
									assign node3933 = (inp[12]) ? 14'b00000000000001 : node3934;
										assign node3934 = (inp[2]) ? node3936 : 14'b00000000000001;
											assign node3936 = (inp[8]) ? node3942 : node3937;
												assign node3937 = (inp[10]) ? node3939 : 14'b00000000000001;
													assign node3939 = (inp[5]) ? 14'b00000000000001 : 14'b10000001000000;
												assign node3942 = (inp[5]) ? 14'b10000001000000 : 14'b00000000000001;
							assign node3948 = (inp[5]) ? node4034 : node3949;
								assign node3949 = (inp[2]) ? node3997 : node3950;
									assign node3950 = (inp[4]) ? node3974 : node3951;
										assign node3951 = (inp[12]) ? node3963 : node3952;
											assign node3952 = (inp[8]) ? node3960 : node3953;
												assign node3953 = (inp[10]) ? node3957 : node3954;
													assign node3954 = (inp[7]) ? 14'b00000000100010 : 14'b00000000000001;
													assign node3957 = (inp[7]) ? 14'b01100000100010 : 14'b01100100100010;
												assign node3960 = (inp[7]) ? 14'b00000000100000 : 14'b00000000000001;
											assign node3963 = (inp[8]) ? node3971 : node3964;
												assign node3964 = (inp[10]) ? node3968 : node3965;
													assign node3965 = (inp[7]) ? 14'b00000000100000 : 14'b01000000100100;
													assign node3968 = (inp[7]) ? 14'b01100000100000 : 14'b01100100100000;
												assign node3971 = (inp[7]) ? 14'b01000000100100 : 14'b01000100100100;
										assign node3974 = (inp[7]) ? node3986 : node3975;
											assign node3975 = (inp[8]) ? node3983 : node3976;
												assign node3976 = (inp[10]) ? node3980 : node3977;
													assign node3977 = (inp[12]) ? 14'b00100100100100 : 14'b00100100100110;
													assign node3980 = (inp[12]) ? 14'b00100100100000 : 14'b00100100100010;
												assign node3983 = (inp[12]) ? 14'b00000100100100 : 14'b00100100100100;
											assign node3986 = (inp[8]) ? node3994 : node3987;
												assign node3987 = (inp[10]) ? node3991 : node3988;
													assign node3988 = (inp[12]) ? 14'b00100000100100 : 14'b00100000100110;
													assign node3991 = (inp[12]) ? 14'b00100000100000 : 14'b00100000100010;
												assign node3994 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
									assign node3997 = (inp[4]) ? node4023 : node3998;
										assign node3998 = (inp[10]) ? node4014 : node3999;
											assign node3999 = (inp[7]) ? node4007 : node4000;
												assign node4000 = (inp[8]) ? node4004 : node4001;
													assign node4001 = (inp[12]) ? 14'b01100100100100 : 14'b01100100100110;
													assign node4004 = (inp[12]) ? 14'b01000100100000 : 14'b01100100100100;
												assign node4007 = (inp[8]) ? node4011 : node4008;
													assign node4008 = (inp[12]) ? 14'b01100000100100 : 14'b01100000100110;
													assign node4011 = (inp[12]) ? 14'b01000000100000 : 14'b01100000100100;
											assign node4014 = (inp[8]) ? node4016 : 14'b00000000000001;
												assign node4016 = (inp[12]) ? node4020 : node4017;
													assign node4017 = (inp[7]) ? 14'b01100000100100 : 14'b01100100100100;
													assign node4020 = (inp[7]) ? 14'b01000000100000 : 14'b01000100100000;
										assign node4023 = (inp[8]) ? 14'b00000000000001 : node4024;
											assign node4024 = (inp[7]) ? 14'b00000000000001 : node4025;
												assign node4025 = (inp[12]) ? node4029 : node4026;
													assign node4026 = (inp[10]) ? 14'b00000100100010 : 14'b00000000000001;
													assign node4029 = (inp[10]) ? 14'b00000100100000 : 14'b00000100100100;
								assign node4034 = (inp[12]) ? node4068 : node4035;
									assign node4035 = (inp[2]) ? node4053 : node4036;
										assign node4036 = (inp[8]) ? node4046 : node4037;
											assign node4037 = (inp[10]) ? 14'b00000000000001 : node4038;
												assign node4038 = (inp[4]) ? node4042 : node4039;
													assign node4039 = (inp[7]) ? 14'b01000000100110 : 14'b01000100100110;
													assign node4042 = (inp[7]) ? 14'b00000000100110 : 14'b00000100100110;
											assign node4046 = (inp[4]) ? node4050 : node4047;
												assign node4047 = (inp[7]) ? 14'b01100000100000 : 14'b01100100100000;
												assign node4050 = (inp[7]) ? 14'b00100000100000 : 14'b00100100100000;
										assign node4053 = (inp[7]) ? 14'b00000000000001 : node4054;
											assign node4054 = (inp[10]) ? node4062 : node4055;
												assign node4055 = (inp[8]) ? node4059 : node4056;
													assign node4056 = (inp[4]) ? 14'b01000000100010 : 14'b01000100100010;
													assign node4059 = (inp[4]) ? 14'b00000100100000 : 14'b00000000000001;
												assign node4062 = (inp[8]) ? node4064 : 14'b00000000000001;
													assign node4064 = (inp[4]) ? 14'b00000100100000 : 14'b00000000000001;
									assign node4068 = (inp[8]) ? 14'b00000000000001 : node4069;
										assign node4069 = (inp[10]) ? 14'b00000000000001 : node4070;
											assign node4070 = (inp[4]) ? node4078 : node4071;
												assign node4071 = (inp[7]) ? node4075 : node4072;
													assign node4072 = (inp[2]) ? 14'b01000100100000 : 14'b01000100100100;
													assign node4075 = (inp[2]) ? 14'b01000000100000 : 14'b00000000000001;
												assign node4078 = (inp[7]) ? node4080 : 14'b00000000000001;
													assign node4080 = (inp[2]) ? 14'b00000000000001 : 14'b00000000100100;
				assign node4086 = (inp[8]) ? node4116 : node4087;
					assign node4087 = (inp[12]) ? 14'b00000000000001 : node4088;
						assign node4088 = (inp[7]) ? 14'b00000000000001 : node4089;
							assign node4089 = (inp[5]) ? 14'b00000000000001 : node4090;
								assign node4090 = (inp[6]) ? 14'b00000000000001 : node4091;
									assign node4091 = (inp[2]) ? node4101 : node4092;
										assign node4092 = (inp[9]) ? node4094 : 14'b00000000000001;
											assign node4094 = (inp[10]) ? 14'b00000000000001 : node4095;
												assign node4095 = (inp[4]) ? 14'b00000000000001 : node4096;
													assign node4096 = (inp[3]) ? 14'b10000000000010 : 14'b00000000000001;
										assign node4101 = (inp[9]) ? 14'b00000000000001 : node4102;
											assign node4102 = (inp[3]) ? 14'b00000000000001 : node4103;
												assign node4103 = (inp[10]) ? node4107 : node4104;
													assign node4104 = (inp[4]) ? 14'b10000001000010 : 14'b00000000000001;
													assign node4107 = (inp[4]) ? 14'b00000000000001 : 14'b10000000001010;
					assign node4116 = (inp[5]) ? node4138 : node4117;
						assign node4117 = (inp[7]) ? 14'b00000000000001 : node4118;
							assign node4118 = (inp[6]) ? 14'b00000000000001 : node4119;
								assign node4119 = (inp[12]) ? 14'b00000000000001 : node4120;
									assign node4120 = (inp[9]) ? node4128 : node4121;
										assign node4121 = (inp[2]) ? node4123 : 14'b00000000000001;
											assign node4123 = (inp[4]) ? node4125 : 14'b00000000000001;
												assign node4125 = (inp[3]) ? 14'b00000000000001 : 14'b10000001000010;
										assign node4128 = (inp[2]) ? 14'b00000000000001 : node4129;
											assign node4129 = (inp[4]) ? 14'b00000000000001 : node4130;
												assign node4130 = (inp[3]) ? 14'b10000000000010 : 14'b00000000000001;
						assign node4138 = (inp[2]) ? node4152 : node4139;
							assign node4139 = (inp[6]) ? 14'b00000000000001 : node4140;
								assign node4140 = (inp[3]) ? 14'b00000000000001 : node4141;
									assign node4141 = (inp[9]) ? 14'b00000000000001 : node4142;
										assign node4142 = (inp[4]) ? 14'b00000000000001 : node4143;
											assign node4143 = (inp[12]) ? node4145 : 14'b00000000000001;
												assign node4145 = (inp[7]) ? 14'b00000000000001 : 14'b10001001001000;
							assign node4152 = (inp[7]) ? node4164 : node4153;
								assign node4153 = (inp[9]) ? 14'b00000000000001 : node4154;
									assign node4154 = (inp[3]) ? 14'b00000000000001 : node4155;
										assign node4155 = (inp[4]) ? 14'b00000000000001 : node4156;
											assign node4156 = (inp[12]) ? 14'b00000000000001 : node4157;
												assign node4157 = (inp[6]) ? 14'b00000000000001 : 14'b10000000001010;
								assign node4164 = (inp[3]) ? node4166 : 14'b00000000000001;
									assign node4166 = (inp[9]) ? node4168 : 14'b00000000000001;
										assign node4168 = (inp[12]) ? node4170 : 14'b00000000000001;
											assign node4170 = (inp[4]) ? node4174 : node4171;
												assign node4171 = (inp[6]) ? 14'b10001001000000 : 14'b10001000000000;
												assign node4174 = (inp[6]) ? 14'b10001001001010 : 14'b10001000001010;

endmodule