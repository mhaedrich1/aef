module dtc_split25_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node868;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node988;

	assign outp = (inp[3]) ? node576 : node1;
		assign node1 = (inp[4]) ? node271 : node2;
			assign node2 = (inp[9]) ? node126 : node3;
				assign node3 = (inp[7]) ? node79 : node4;
					assign node4 = (inp[11]) ? node42 : node5;
						assign node5 = (inp[1]) ? node27 : node6;
							assign node6 = (inp[6]) ? node14 : node7;
								assign node7 = (inp[2]) ? 3'b001 : node8;
									assign node8 = (inp[0]) ? node10 : 3'b001;
										assign node10 = (inp[5]) ? 3'b001 : 3'b111;
								assign node14 = (inp[2]) ? node20 : node15;
									assign node15 = (inp[8]) ? 3'b111 : node16;
										assign node16 = (inp[0]) ? 3'b001 : 3'b011;
									assign node20 = (inp[8]) ? node24 : node21;
										assign node21 = (inp[0]) ? 3'b101 : 3'b101;
										assign node24 = (inp[0]) ? 3'b011 : 3'b001;
							assign node27 = (inp[5]) ? node35 : node28;
								assign node28 = (inp[10]) ? node30 : 3'b001;
									assign node30 = (inp[0]) ? node32 : 3'b011;
										assign node32 = (inp[2]) ? 3'b011 : 3'b111;
								assign node35 = (inp[10]) ? 3'b011 : node36;
									assign node36 = (inp[6]) ? 3'b111 : node37;
										assign node37 = (inp[0]) ? 3'b011 : 3'b111;
						assign node42 = (inp[2]) ? node60 : node43;
							assign node43 = (inp[10]) ? node53 : node44;
								assign node44 = (inp[5]) ? node50 : node45;
									assign node45 = (inp[8]) ? 3'b111 : node46;
										assign node46 = (inp[0]) ? 3'b011 : 3'b111;
									assign node50 = (inp[0]) ? 3'b111 : 3'b011;
								assign node53 = (inp[5]) ? node55 : 3'b011;
									assign node55 = (inp[1]) ? 3'b011 : node56;
										assign node56 = (inp[8]) ? 3'b101 : 3'b001;
							assign node60 = (inp[0]) ? node74 : node61;
								assign node61 = (inp[10]) ? node69 : node62;
									assign node62 = (inp[5]) ? node66 : node63;
										assign node63 = (inp[8]) ? 3'b101 : 3'b111;
										assign node66 = (inp[1]) ? 3'b011 : 3'b111;
									assign node69 = (inp[8]) ? 3'b101 : node70;
										assign node70 = (inp[6]) ? 3'b011 : 3'b001;
								assign node74 = (inp[5]) ? node76 : 3'b111;
									assign node76 = (inp[8]) ? 3'b111 : 3'b101;
					assign node79 = (inp[5]) ? node105 : node80;
						assign node80 = (inp[1]) ? node90 : node81;
							assign node81 = (inp[2]) ? node83 : 3'b111;
								assign node83 = (inp[10]) ? node85 : 3'b111;
									assign node85 = (inp[6]) ? node87 : 3'b111;
										assign node87 = (inp[11]) ? 3'b111 : 3'b101;
							assign node90 = (inp[6]) ? node98 : node91;
								assign node91 = (inp[10]) ? node93 : 3'b011;
									assign node93 = (inp[2]) ? node95 : 3'b111;
										assign node95 = (inp[8]) ? 3'b001 : 3'b111;
								assign node98 = (inp[2]) ? node100 : 3'b111;
									assign node100 = (inp[0]) ? 3'b111 : node101;
										assign node101 = (inp[8]) ? 3'b101 : 3'b111;
						assign node105 = (inp[0]) ? node117 : node106;
							assign node106 = (inp[6]) ? node114 : node107;
								assign node107 = (inp[1]) ? node109 : 3'b111;
									assign node109 = (inp[2]) ? 3'b011 : node110;
										assign node110 = (inp[10]) ? 3'b011 : 3'b101;
								assign node114 = (inp[11]) ? 3'b101 : 3'b111;
							assign node117 = (inp[1]) ? node119 : 3'b011;
								assign node119 = (inp[6]) ? 3'b111 : node120;
									assign node120 = (inp[2]) ? node122 : 3'b011;
										assign node122 = (inp[8]) ? 3'b111 : 3'b011;
				assign node126 = (inp[6]) ? node200 : node127;
					assign node127 = (inp[0]) ? node167 : node128;
						assign node128 = (inp[10]) ? node146 : node129;
							assign node129 = (inp[7]) ? node137 : node130;
								assign node130 = (inp[1]) ? node132 : 3'b110;
									assign node132 = (inp[11]) ? 3'b110 : node133;
										assign node133 = (inp[5]) ? 3'b001 : 3'b101;
								assign node137 = (inp[1]) ? 3'b110 : node138;
									assign node138 = (inp[8]) ? node142 : node139;
										assign node139 = (inp[11]) ? 3'b000 : 3'b001;
										assign node142 = (inp[2]) ? 3'b001 : 3'b101;
							assign node146 = (inp[5]) ? node154 : node147;
								assign node147 = (inp[7]) ? node149 : 3'b110;
									assign node149 = (inp[11]) ? node151 : 3'b001;
										assign node151 = (inp[1]) ? 3'b001 : 3'b110;
								assign node154 = (inp[8]) ? node162 : node155;
									assign node155 = (inp[1]) ? node159 : node156;
										assign node156 = (inp[7]) ? 3'b010 : 3'b100;
										assign node159 = (inp[7]) ? 3'b110 : 3'b010;
									assign node162 = (inp[7]) ? node164 : 3'b010;
										assign node164 = (inp[11]) ? 3'b010 : 3'b110;
						assign node167 = (inp[1]) ? node187 : node168;
							assign node168 = (inp[7]) ? node180 : node169;
								assign node169 = (inp[10]) ? node175 : node170;
									assign node170 = (inp[2]) ? node172 : 3'b101;
										assign node172 = (inp[8]) ? 3'b010 : 3'b001;
									assign node175 = (inp[8]) ? 3'b110 : node176;
										assign node176 = (inp[5]) ? 3'b010 : 3'b110;
								assign node180 = (inp[8]) ? 3'b001 : node181;
									assign node181 = (inp[10]) ? node183 : 3'b101;
										assign node183 = (inp[5]) ? 3'b110 : 3'b101;
							assign node187 = (inp[8]) ? node195 : node188;
								assign node188 = (inp[2]) ? 3'b101 : node189;
									assign node189 = (inp[11]) ? node191 : 3'b101;
										assign node191 = (inp[10]) ? 3'b001 : 3'b001;
								assign node195 = (inp[10]) ? 3'b101 : node196;
									assign node196 = (inp[11]) ? 3'b101 : 3'b111;
					assign node200 = (inp[0]) ? node244 : node201;
						assign node201 = (inp[7]) ? node225 : node202;
							assign node202 = (inp[5]) ? node214 : node203;
								assign node203 = (inp[2]) ? node209 : node204;
									assign node204 = (inp[8]) ? 3'b101 : node205;
										assign node205 = (inp[1]) ? 3'b101 : 3'b001;
									assign node209 = (inp[10]) ? node211 : 3'b011;
										assign node211 = (inp[1]) ? 3'b101 : 3'b001;
								assign node214 = (inp[10]) ? node218 : node215;
									assign node215 = (inp[8]) ? 3'b101 : 3'b001;
									assign node218 = (inp[1]) ? node222 : node219;
										assign node219 = (inp[11]) ? 3'b110 : 3'b010;
										assign node222 = (inp[8]) ? 3'b001 : 3'b110;
							assign node225 = (inp[11]) ? node231 : node226;
								assign node226 = (inp[8]) ? 3'b011 : node227;
									assign node227 = (inp[2]) ? 3'b011 : 3'b101;
								assign node231 = (inp[1]) ? node239 : node232;
									assign node232 = (inp[8]) ? node236 : node233;
										assign node233 = (inp[5]) ? 3'b001 : 3'b101;
										assign node236 = (inp[5]) ? 3'b101 : 3'b001;
									assign node239 = (inp[8]) ? 3'b011 : node240;
										assign node240 = (inp[2]) ? 3'b011 : 3'b101;
						assign node244 = (inp[1]) ? node262 : node245;
							assign node245 = (inp[10]) ? node253 : node246;
								assign node246 = (inp[7]) ? 3'b111 : node247;
									assign node247 = (inp[11]) ? 3'b101 : node248;
										assign node248 = (inp[5]) ? 3'b011 : 3'b111;
								assign node253 = (inp[5]) ? node259 : node254;
									assign node254 = (inp[11]) ? node256 : 3'b011;
										assign node256 = (inp[7]) ? 3'b011 : 3'b001;
									assign node259 = (inp[11]) ? 3'b001 : 3'b101;
							assign node262 = (inp[11]) ? node264 : 3'b111;
								assign node264 = (inp[5]) ? node266 : 3'b111;
									assign node266 = (inp[10]) ? 3'b011 : node267;
										assign node267 = (inp[7]) ? 3'b111 : 3'b011;
			assign node271 = (inp[0]) ? node419 : node272;
				assign node272 = (inp[9]) ? node356 : node273;
					assign node273 = (inp[11]) ? node315 : node274;
						assign node274 = (inp[1]) ? node294 : node275;
							assign node275 = (inp[8]) ? node283 : node276;
								assign node276 = (inp[5]) ? node280 : node277;
									assign node277 = (inp[10]) ? 3'b010 : 3'b011;
									assign node280 = (inp[10]) ? 3'b001 : 3'b101;
								assign node283 = (inp[2]) ? node289 : node284;
									assign node284 = (inp[6]) ? 3'b001 : node285;
										assign node285 = (inp[5]) ? 3'b001 : 3'b101;
									assign node289 = (inp[6]) ? 3'b101 : node290;
										assign node290 = (inp[7]) ? 3'b001 : 3'b001;
							assign node294 = (inp[10]) ? node306 : node295;
								assign node295 = (inp[6]) ? node301 : node296;
									assign node296 = (inp[5]) ? node298 : 3'b101;
										assign node298 = (inp[7]) ? 3'b001 : 3'b010;
									assign node301 = (inp[8]) ? 3'b110 : node302;
										assign node302 = (inp[7]) ? 3'b000 : 3'b010;
								assign node306 = (inp[5]) ? node310 : node307;
									assign node307 = (inp[7]) ? 3'b111 : 3'b001;
									assign node310 = (inp[6]) ? 3'b101 : node311;
										assign node311 = (inp[8]) ? 3'b000 : 3'b010;
						assign node315 = (inp[8]) ? node335 : node316;
							assign node316 = (inp[2]) ? node330 : node317;
								assign node317 = (inp[10]) ? node323 : node318;
									assign node318 = (inp[1]) ? node320 : 3'b101;
										assign node320 = (inp[6]) ? 3'b000 : 3'b000;
									assign node323 = (inp[7]) ? node327 : node324;
										assign node324 = (inp[1]) ? 3'b010 : 3'b000;
										assign node327 = (inp[6]) ? 3'b101 : 3'b110;
								assign node330 = (inp[5]) ? 3'b110 : node331;
									assign node331 = (inp[10]) ? 3'b001 : 3'b010;
							assign node335 = (inp[1]) ? node345 : node336;
								assign node336 = (inp[7]) ? node340 : node337;
									assign node337 = (inp[2]) ? 3'b011 : 3'b010;
									assign node340 = (inp[2]) ? node342 : 3'b010;
										assign node342 = (inp[6]) ? 3'b110 : 3'b010;
								assign node345 = (inp[7]) ? node349 : node346;
									assign node346 = (inp[10]) ? 3'b110 : 3'b010;
									assign node349 = (inp[6]) ? node353 : node350;
										assign node350 = (inp[5]) ? 3'b000 : 3'b001;
										assign node353 = (inp[5]) ? 3'b111 : 3'b110;
					assign node356 = (inp[6]) ? node384 : node357;
						assign node357 = (inp[1]) ? node365 : node358;
							assign node358 = (inp[5]) ? node360 : 3'b100;
								assign node360 = (inp[10]) ? 3'b000 : node361;
									assign node361 = (inp[7]) ? 3'b100 : 3'b000;
							assign node365 = (inp[10]) ? node375 : node366;
								assign node366 = (inp[5]) ? node370 : node367;
									assign node367 = (inp[7]) ? 3'b110 : 3'b010;
									assign node370 = (inp[7]) ? node372 : 3'b100;
										assign node372 = (inp[2]) ? 3'b000 : 3'b010;
								assign node375 = (inp[5]) ? node379 : node376;
									assign node376 = (inp[7]) ? 3'b010 : 3'b100;
									assign node379 = (inp[7]) ? 3'b100 : node380;
										assign node380 = (inp[11]) ? 3'b000 : 3'b100;
						assign node384 = (inp[10]) ? node400 : node385;
							assign node385 = (inp[8]) ? node397 : node386;
								assign node386 = (inp[7]) ? node394 : node387;
									assign node387 = (inp[5]) ? node391 : node388;
										assign node388 = (inp[1]) ? 3'b111 : 3'b110;
										assign node391 = (inp[1]) ? 3'b110 : 3'b010;
									assign node394 = (inp[11]) ? 3'b010 : 3'b001;
								assign node397 = (inp[5]) ? 3'b000 : 3'b001;
							assign node400 = (inp[11]) ? node408 : node401;
								assign node401 = (inp[2]) ? node403 : 3'b010;
									assign node403 = (inp[7]) ? 3'b110 : node404;
										assign node404 = (inp[1]) ? 3'b010 : 3'b000;
								assign node408 = (inp[2]) ? node414 : node409;
									assign node409 = (inp[7]) ? node411 : 3'b100;
										assign node411 = (inp[5]) ? 3'b100 : 3'b110;
									assign node414 = (inp[5]) ? 3'b110 : node415;
										assign node415 = (inp[1]) ? 3'b000 : 3'b110;
				assign node419 = (inp[9]) ? node491 : node420;
					assign node420 = (inp[8]) ? node460 : node421;
						assign node421 = (inp[6]) ? node443 : node422;
							assign node422 = (inp[7]) ? node430 : node423;
								assign node423 = (inp[2]) ? node427 : node424;
									assign node424 = (inp[1]) ? 3'b000 : 3'b001;
									assign node427 = (inp[10]) ? 3'b110 : 3'b011;
								assign node430 = (inp[5]) ? node438 : node431;
									assign node431 = (inp[11]) ? node435 : node432;
										assign node432 = (inp[2]) ? 3'b111 : 3'b011;
										assign node435 = (inp[10]) ? 3'b111 : 3'b100;
									assign node438 = (inp[10]) ? 3'b001 : node439;
										assign node439 = (inp[1]) ? 3'b001 : 3'b101;
							assign node443 = (inp[1]) ? node453 : node444;
								assign node444 = (inp[2]) ? node450 : node445;
									assign node445 = (inp[10]) ? node447 : 3'b100;
										assign node447 = (inp[11]) ? 3'b111 : 3'b001;
									assign node450 = (inp[11]) ? 3'b001 : 3'b000;
								assign node453 = (inp[5]) ? 3'b101 : node454;
									assign node454 = (inp[2]) ? node456 : 3'b101;
										assign node456 = (inp[7]) ? 3'b001 : 3'b011;
						assign node460 = (inp[11]) ? node478 : node461;
							assign node461 = (inp[2]) ? node471 : node462;
								assign node462 = (inp[10]) ? node466 : node463;
									assign node463 = (inp[1]) ? 3'b101 : 3'b011;
									assign node466 = (inp[1]) ? node468 : 3'b111;
										assign node468 = (inp[5]) ? 3'b111 : 3'b011;
								assign node471 = (inp[5]) ? 3'b011 : node472;
									assign node472 = (inp[1]) ? node474 : 3'b001;
										assign node474 = (inp[6]) ? 3'b001 : 3'b011;
							assign node478 = (inp[6]) ? node488 : node479;
								assign node479 = (inp[1]) ? node485 : node480;
									assign node480 = (inp[10]) ? node482 : 3'b101;
										assign node482 = (inp[5]) ? 3'b000 : 3'b111;
									assign node485 = (inp[5]) ? 3'b001 : 3'b101;
								assign node488 = (inp[1]) ? 3'b111 : 3'b101;
					assign node491 = (inp[6]) ? node531 : node492;
						assign node492 = (inp[7]) ? node510 : node493;
							assign node493 = (inp[5]) ? node501 : node494;
								assign node494 = (inp[2]) ? 3'b110 : node495;
									assign node495 = (inp[11]) ? 3'b010 : node496;
										assign node496 = (inp[8]) ? 3'b010 : 3'b110;
								assign node501 = (inp[10]) ? node507 : node502;
									assign node502 = (inp[1]) ? node504 : 3'b010;
										assign node504 = (inp[8]) ? 3'b110 : 3'b010;
									assign node507 = (inp[11]) ? 3'b100 : 3'b010;
							assign node510 = (inp[1]) ? node518 : node511;
								assign node511 = (inp[10]) ? node515 : node512;
									assign node512 = (inp[8]) ? 3'b110 : 3'b010;
									assign node515 = (inp[5]) ? 3'b100 : 3'b010;
								assign node518 = (inp[10]) ? node524 : node519;
									assign node519 = (inp[5]) ? node521 : 3'b101;
										assign node521 = (inp[8]) ? 3'b001 : 3'b101;
									assign node524 = (inp[5]) ? node528 : node525;
										assign node525 = (inp[2]) ? 3'b001 : 3'b000;
										assign node528 = (inp[2]) ? 3'b110 : 3'b010;
						assign node531 = (inp[1]) ? node553 : node532;
							assign node532 = (inp[2]) ? node542 : node533;
								assign node533 = (inp[10]) ? node537 : node534;
									assign node534 = (inp[5]) ? 3'b111 : 3'b011;
									assign node537 = (inp[5]) ? node539 : 3'b110;
										assign node539 = (inp[8]) ? 3'b110 : 3'b010;
								assign node542 = (inp[8]) ? node550 : node543;
									assign node543 = (inp[10]) ? node547 : node544;
										assign node544 = (inp[5]) ? 3'b001 : 3'b101;
										assign node547 = (inp[5]) ? 3'b000 : 3'b001;
									assign node550 = (inp[10]) ? 3'b001 : 3'b011;
							assign node553 = (inp[5]) ? node565 : node554;
								assign node554 = (inp[10]) ? node560 : node555;
									assign node555 = (inp[7]) ? 3'b011 : node556;
										assign node556 = (inp[8]) ? 3'b011 : 3'b001;
									assign node560 = (inp[7]) ? 3'b101 : node561;
										assign node561 = (inp[8]) ? 3'b100 : 3'b101;
								assign node565 = (inp[10]) ? node571 : node566;
									assign node566 = (inp[7]) ? 3'b101 : node567;
										assign node567 = (inp[8]) ? 3'b101 : 3'b001;
									assign node571 = (inp[8]) ? 3'b001 : node572;
										assign node572 = (inp[11]) ? 3'b110 : 3'b001;
		assign node576 = (inp[4]) ? node846 : node577;
			assign node577 = (inp[9]) ? node729 : node578;
				assign node578 = (inp[0]) ? node662 : node579;
					assign node579 = (inp[6]) ? node625 : node580;
						assign node580 = (inp[11]) ? node604 : node581;
							assign node581 = (inp[7]) ? node595 : node582;
								assign node582 = (inp[8]) ? node588 : node583;
									assign node583 = (inp[1]) ? 3'b100 : node584;
										assign node584 = (inp[2]) ? 3'b000 : 3'b000;
									assign node588 = (inp[1]) ? node592 : node589;
										assign node589 = (inp[10]) ? 3'b000 : 3'b000;
										assign node592 = (inp[10]) ? 3'b000 : 3'b010;
								assign node595 = (inp[1]) ? node601 : node596;
									assign node596 = (inp[2]) ? node598 : 3'b000;
										assign node598 = (inp[10]) ? 3'b010 : 3'b000;
									assign node601 = (inp[10]) ? 3'b110 : 3'b011;
							assign node604 = (inp[1]) ? node614 : node605;
								assign node605 = (inp[8]) ? node609 : node606;
									assign node606 = (inp[2]) ? 3'b100 : 3'b000;
									assign node609 = (inp[5]) ? 3'b100 : node610;
										assign node610 = (inp[10]) ? 3'b100 : 3'b100;
								assign node614 = (inp[5]) ? node620 : node615;
									assign node615 = (inp[10]) ? 3'b100 : node616;
										assign node616 = (inp[2]) ? 3'b000 : 3'b010;
									assign node620 = (inp[10]) ? 3'b000 : node621;
										assign node621 = (inp[7]) ? 3'b000 : 3'b100;
						assign node625 = (inp[7]) ? node641 : node626;
							assign node626 = (inp[1]) ? node634 : node627;
								assign node627 = (inp[10]) ? node629 : 3'b100;
									assign node629 = (inp[5]) ? node631 : 3'b000;
										assign node631 = (inp[11]) ? 3'b100 : 3'b000;
								assign node634 = (inp[5]) ? node638 : node635;
									assign node635 = (inp[2]) ? 3'b000 : 3'b110;
									assign node638 = (inp[10]) ? 3'b010 : 3'b110;
							assign node641 = (inp[8]) ? node651 : node642;
								assign node642 = (inp[1]) ? node648 : node643;
									assign node643 = (inp[11]) ? node645 : 3'b110;
										assign node645 = (inp[10]) ? 3'b110 : 3'b100;
									assign node648 = (inp[5]) ? 3'b010 : 3'b110;
								assign node651 = (inp[5]) ? node657 : node652;
									assign node652 = (inp[1]) ? node654 : 3'b010;
										assign node654 = (inp[2]) ? 3'b011 : 3'b010;
									assign node657 = (inp[10]) ? 3'b110 : node658;
										assign node658 = (inp[11]) ? 3'b101 : 3'b111;
					assign node662 = (inp[6]) ? node692 : node663;
						assign node663 = (inp[10]) ? node681 : node664;
							assign node664 = (inp[7]) ? node674 : node665;
								assign node665 = (inp[2]) ? node671 : node666;
									assign node666 = (inp[1]) ? 3'b110 : node667;
										assign node667 = (inp[5]) ? 3'b010 : 3'b110;
									assign node671 = (inp[11]) ? 3'b110 : 3'b100;
								assign node674 = (inp[11]) ? node678 : node675;
									assign node675 = (inp[5]) ? 3'b110 : 3'b011;
									assign node678 = (inp[1]) ? 3'b101 : 3'b100;
							assign node681 = (inp[5]) ? node689 : node682;
								assign node682 = (inp[11]) ? node684 : 3'b110;
									assign node684 = (inp[8]) ? node686 : 3'b010;
										assign node686 = (inp[2]) ? 3'b010 : 3'b010;
								assign node689 = (inp[7]) ? 3'b010 : 3'b100;
						assign node692 = (inp[7]) ? node712 : node693;
							assign node693 = (inp[10]) ? node705 : node694;
								assign node694 = (inp[5]) ? node700 : node695;
									assign node695 = (inp[2]) ? node697 : 3'b111;
										assign node697 = (inp[1]) ? 3'b011 : 3'b000;
									assign node700 = (inp[2]) ? node702 : 3'b001;
										assign node702 = (inp[1]) ? 3'b101 : 3'b001;
								assign node705 = (inp[11]) ? 3'b110 : node706;
									assign node706 = (inp[5]) ? 3'b110 : node707;
										assign node707 = (inp[8]) ? 3'b001 : 3'b000;
							assign node712 = (inp[5]) ? node724 : node713;
								assign node713 = (inp[10]) ? node717 : node714;
									assign node714 = (inp[1]) ? 3'b011 : 3'b010;
									assign node717 = (inp[1]) ? node721 : node718;
										assign node718 = (inp[11]) ? 3'b001 : 3'b101;
										assign node721 = (inp[11]) ? 3'b101 : 3'b011;
								assign node724 = (inp[10]) ? 3'b001 : node725;
									assign node725 = (inp[1]) ? 3'b101 : 3'b001;
				assign node729 = (inp[0]) ? node777 : node730;
					assign node730 = (inp[10]) ? node766 : node731;
						assign node731 = (inp[6]) ? node741 : node732;
							assign node732 = (inp[8]) ? node734 : 3'b000;
								assign node734 = (inp[5]) ? 3'b000 : node735;
									assign node735 = (inp[1]) ? node737 : 3'b000;
										assign node737 = (inp[11]) ? 3'b100 : 3'b000;
							assign node741 = (inp[1]) ? node753 : node742;
								assign node742 = (inp[8]) ? node750 : node743;
									assign node743 = (inp[5]) ? node747 : node744;
										assign node744 = (inp[7]) ? 3'b010 : 3'b000;
										assign node747 = (inp[7]) ? 3'b100 : 3'b000;
									assign node750 = (inp[7]) ? 3'b010 : 3'b000;
								assign node753 = (inp[2]) ? node761 : node754;
									assign node754 = (inp[11]) ? node758 : node755;
										assign node755 = (inp[8]) ? 3'b010 : 3'b000;
										assign node758 = (inp[7]) ? 3'b100 : 3'b000;
									assign node761 = (inp[8]) ? node763 : 3'b010;
										assign node763 = (inp[5]) ? 3'b100 : 3'b110;
						assign node766 = (inp[7]) ? node768 : 3'b000;
							assign node768 = (inp[8]) ? node770 : 3'b000;
								assign node770 = (inp[6]) ? node772 : 3'b000;
									assign node772 = (inp[1]) ? 3'b100 : node773;
										assign node773 = (inp[5]) ? 3'b000 : 3'b100;
					assign node777 = (inp[6]) ? node815 : node778;
						assign node778 = (inp[5]) ? node802 : node779;
							assign node779 = (inp[11]) ? node793 : node780;
								assign node780 = (inp[8]) ? node788 : node781;
									assign node781 = (inp[10]) ? node785 : node782;
										assign node782 = (inp[1]) ? 3'b000 : 3'b100;
										assign node785 = (inp[2]) ? 3'b100 : 3'b000;
									assign node788 = (inp[1]) ? 3'b010 : node789;
										assign node789 = (inp[10]) ? 3'b100 : 3'b010;
								assign node793 = (inp[8]) ? node797 : node794;
									assign node794 = (inp[10]) ? 3'b000 : 3'b100;
									assign node797 = (inp[10]) ? 3'b100 : node798;
										assign node798 = (inp[2]) ? 3'b110 : 3'b100;
							assign node802 = (inp[1]) ? node804 : 3'b000;
								assign node804 = (inp[8]) ? node810 : node805;
									assign node805 = (inp[11]) ? 3'b100 : node806;
										assign node806 = (inp[7]) ? 3'b010 : 3'b000;
									assign node810 = (inp[7]) ? 3'b100 : node811;
										assign node811 = (inp[2]) ? 3'b100 : 3'b000;
						assign node815 = (inp[5]) ? node831 : node816;
							assign node816 = (inp[10]) ? node826 : node817;
								assign node817 = (inp[11]) ? node823 : node818;
									assign node818 = (inp[1]) ? 3'b001 : node819;
										assign node819 = (inp[7]) ? 3'b001 : 3'b110;
									assign node823 = (inp[1]) ? 3'b110 : 3'b010;
								assign node826 = (inp[7]) ? node828 : 3'b010;
									assign node828 = (inp[8]) ? 3'b110 : 3'b010;
							assign node831 = (inp[10]) ? node839 : node832;
								assign node832 = (inp[11]) ? node834 : 3'b110;
									assign node834 = (inp[7]) ? node836 : 3'b010;
										assign node836 = (inp[1]) ? 3'b110 : 3'b010;
								assign node839 = (inp[1]) ? 3'b100 : node840;
									assign node840 = (inp[2]) ? 3'b100 : node841;
										assign node841 = (inp[7]) ? 3'b100 : 3'b000;
			assign node846 = (inp[6]) ? node886 : node847;
				assign node847 = (inp[0]) ? node849 : 3'b000;
					assign node849 = (inp[7]) ? node859 : node850;
						assign node850 = (inp[8]) ? node852 : 3'b000;
							assign node852 = (inp[1]) ? node854 : 3'b000;
								assign node854 = (inp[5]) ? 3'b000 : node855;
									assign node855 = (inp[9]) ? 3'b000 : 3'b001;
						assign node859 = (inp[9]) ? node877 : node860;
							assign node860 = (inp[11]) ? node868 : node861;
								assign node861 = (inp[8]) ? 3'b000 : node862;
									assign node862 = (inp[5]) ? 3'b100 : node863;
										assign node863 = (inp[1]) ? 3'b100 : 3'b100;
								assign node868 = (inp[8]) ? node870 : 3'b000;
									assign node870 = (inp[2]) ? node874 : node871;
										assign node871 = (inp[10]) ? 3'b000 : 3'b110;
										assign node874 = (inp[5]) ? 3'b010 : 3'b000;
							assign node877 = (inp[11]) ? 3'b000 : node878;
								assign node878 = (inp[10]) ? 3'b000 : node879;
									assign node879 = (inp[1]) ? node881 : 3'b010;
										assign node881 = (inp[5]) ? 3'b000 : 3'b100;
				assign node886 = (inp[9]) ? node962 : node887;
					assign node887 = (inp[0]) ? node923 : node888;
						assign node888 = (inp[10]) ? node910 : node889;
							assign node889 = (inp[7]) ? node901 : node890;
								assign node890 = (inp[5]) ? node896 : node891;
									assign node891 = (inp[1]) ? 3'b000 : node892;
										assign node892 = (inp[11]) ? 3'b100 : 3'b000;
									assign node896 = (inp[1]) ? 3'b100 : node897;
										assign node897 = (inp[8]) ? 3'b000 : 3'b000;
								assign node901 = (inp[8]) ? node905 : node902;
									assign node902 = (inp[2]) ? 3'b110 : 3'b100;
									assign node905 = (inp[11]) ? node907 : 3'b010;
										assign node907 = (inp[5]) ? 3'b100 : 3'b110;
							assign node910 = (inp[11]) ? 3'b000 : node911;
								assign node911 = (inp[8]) ? node919 : node912;
									assign node912 = (inp[5]) ? node916 : node913;
										assign node913 = (inp[7]) ? 3'b000 : 3'b000;
										assign node916 = (inp[1]) ? 3'b100 : 3'b000;
									assign node919 = (inp[5]) ? 3'b000 : 3'b100;
						assign node923 = (inp[5]) ? node941 : node924;
							assign node924 = (inp[10]) ? node932 : node925;
								assign node925 = (inp[7]) ? 3'b001 : node926;
									assign node926 = (inp[11]) ? 3'b110 : node927;
										assign node927 = (inp[1]) ? 3'b001 : 3'b000;
								assign node932 = (inp[8]) ? node936 : node933;
									assign node933 = (inp[7]) ? 3'b110 : 3'b100;
									assign node936 = (inp[11]) ? 3'b010 : node937;
										assign node937 = (inp[7]) ? 3'b001 : 3'b110;
							assign node941 = (inp[10]) ? node953 : node942;
								assign node942 = (inp[11]) ? node948 : node943;
									assign node943 = (inp[7]) ? 3'b001 : node944;
										assign node944 = (inp[8]) ? 3'b010 : 3'b000;
									assign node948 = (inp[7]) ? 3'b110 : node949;
										assign node949 = (inp[1]) ? 3'b010 : 3'b100;
								assign node953 = (inp[11]) ? node957 : node954;
									assign node954 = (inp[7]) ? 3'b010 : 3'b100;
									assign node957 = (inp[7]) ? 3'b100 : node958;
										assign node958 = (inp[1]) ? 3'b100 : 3'b000;
					assign node962 = (inp[1]) ? node970 : node963;
						assign node963 = (inp[5]) ? 3'b000 : node964;
							assign node964 = (inp[11]) ? 3'b000 : node965;
								assign node965 = (inp[10]) ? 3'b000 : 3'b010;
						assign node970 = (inp[10]) ? node984 : node971;
							assign node971 = (inp[8]) ? node977 : node972;
								assign node972 = (inp[0]) ? node974 : 3'b000;
									assign node974 = (inp[5]) ? 3'b000 : 3'b100;
								assign node977 = (inp[0]) ? node981 : node978;
									assign node978 = (inp[7]) ? 3'b100 : 3'b000;
									assign node981 = (inp[7]) ? 3'b010 : 3'b100;
							assign node984 = (inp[0]) ? node986 : 3'b000;
								assign node986 = (inp[2]) ? node988 : 3'b000;
									assign node988 = (inp[7]) ? 3'b100 : 3'b000;

endmodule