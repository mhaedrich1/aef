module dtc_split125_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node13;
	wire [1-1:0] node14;
	wire [1-1:0] node16;
	wire [1-1:0] node18;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node26;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node31;
	wire [1-1:0] node32;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node76;
	wire [1-1:0] node77;
	wire [1-1:0] node78;
	wire [1-1:0] node80;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node118;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node129;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node152;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node159;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node172;
	wire [1-1:0] node173;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node198;
	wire [1-1:0] node200;
	wire [1-1:0] node202;
	wire [1-1:0] node203;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node210;
	wire [1-1:0] node211;
	wire [1-1:0] node216;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node224;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node230;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node250;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node264;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node268;
	wire [1-1:0] node270;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node276;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node282;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node316;
	wire [1-1:0] node317;
	wire [1-1:0] node318;
	wire [1-1:0] node323;
	wire [1-1:0] node324;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node328;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node348;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node363;
	wire [1-1:0] node364;
	wire [1-1:0] node365;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node372;
	wire [1-1:0] node373;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node384;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node394;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node402;
	wire [1-1:0] node403;
	wire [1-1:0] node405;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node410;
	wire [1-1:0] node411;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node421;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node430;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node446;
	wire [1-1:0] node447;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node454;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node462;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node482;
	wire [1-1:0] node486;
	wire [1-1:0] node487;
	wire [1-1:0] node488;

	assign outp = (inp[10]) ? node262 : node1;
		assign node1 = (inp[4]) ? node109 : node2;
			assign node2 = (inp[6]) ? node42 : node3;
				assign node3 = (inp[2]) ? node5 : 1'b1;
					assign node5 = (inp[12]) ? node13 : node6;
						assign node6 = (inp[8]) ? node8 : 1'b1;
							assign node8 = (inp[3]) ? node10 : 1'b1;
								assign node10 = (inp[0]) ? 1'b0 : 1'b1;
						assign node13 = (inp[7]) ? node21 : node14;
							assign node14 = (inp[11]) ? node16 : 1'b1;
								assign node16 = (inp[5]) ? node18 : 1'b1;
									assign node18 = (inp[0]) ? 1'b0 : 1'b1;
							assign node21 = (inp[9]) ? node29 : node22;
								assign node22 = (inp[0]) ? node24 : 1'b1;
									assign node24 = (inp[11]) ? node26 : 1'b1;
										assign node26 = (inp[8]) ? 1'b0 : 1'b1;
								assign node29 = (inp[0]) ? 1'b0 : node30;
									assign node30 = (inp[8]) ? node36 : node31;
										assign node31 = (inp[5]) ? 1'b1 : node32;
											assign node32 = (inp[1]) ? 1'b0 : 1'b1;
										assign node36 = (inp[1]) ? 1'b0 : node37;
											assign node37 = (inp[11]) ? 1'b0 : 1'b1;
				assign node42 = (inp[12]) ? node76 : node43;
					assign node43 = (inp[0]) ? node53 : node44;
						assign node44 = (inp[2]) ? node46 : 1'b1;
							assign node46 = (inp[1]) ? node48 : 1'b1;
								assign node48 = (inp[11]) ? node50 : 1'b1;
									assign node50 = (inp[9]) ? 1'b0 : 1'b1;
						assign node53 = (inp[9]) ? node65 : node54;
							assign node54 = (inp[8]) ? node56 : 1'b1;
								assign node56 = (inp[5]) ? node58 : 1'b1;
									assign node58 = (inp[11]) ? 1'b0 : node59;
										assign node59 = (inp[3]) ? node61 : 1'b1;
											assign node61 = (inp[1]) ? 1'b0 : 1'b1;
							assign node65 = (inp[7]) ? node71 : node66;
								assign node66 = (inp[3]) ? 1'b1 : node67;
									assign node67 = (inp[11]) ? 1'b0 : 1'b1;
								assign node71 = (inp[1]) ? 1'b0 : node72;
									assign node72 = (inp[5]) ? 1'b0 : 1'b1;
					assign node76 = (inp[3]) ? node100 : node77;
						assign node77 = (inp[7]) ? node85 : node78;
							assign node78 = (inp[5]) ? node80 : 1'b1;
								assign node80 = (inp[1]) ? node82 : 1'b1;
									assign node82 = (inp[2]) ? 1'b0 : 1'b1;
							assign node85 = (inp[1]) ? node95 : node86;
								assign node86 = (inp[5]) ? node88 : 1'b1;
									assign node88 = (inp[0]) ? 1'b0 : node89;
										assign node89 = (inp[11]) ? node91 : 1'b1;
											assign node91 = (inp[8]) ? 1'b0 : 1'b1;
								assign node95 = (inp[2]) ? 1'b0 : node96;
									assign node96 = (inp[0]) ? 1'b0 : 1'b1;
						assign node100 = (inp[1]) ? 1'b0 : node101;
							assign node101 = (inp[0]) ? node103 : 1'b1;
								assign node103 = (inp[8]) ? 1'b0 : node104;
									assign node104 = (inp[5]) ? 1'b0 : 1'b1;
			assign node109 = (inp[5]) ? node193 : node110;
				assign node110 = (inp[6]) ? node148 : node111;
					assign node111 = (inp[2]) ? node121 : node112;
						assign node112 = (inp[1]) ? node114 : 1'b1;
							assign node114 = (inp[0]) ? node116 : 1'b1;
								assign node116 = (inp[3]) ? node118 : 1'b1;
									assign node118 = (inp[11]) ? 1'b0 : 1'b1;
						assign node121 = (inp[9]) ? node133 : node122;
							assign node122 = (inp[8]) ? node124 : 1'b1;
								assign node124 = (inp[3]) ? node126 : 1'b1;
									assign node126 = (inp[7]) ? 1'b0 : node127;
										assign node127 = (inp[0]) ? node129 : 1'b1;
											assign node129 = (inp[1]) ? 1'b0 : 1'b1;
							assign node133 = (inp[11]) ? node143 : node134;
								assign node134 = (inp[7]) ? node136 : 1'b1;
									assign node136 = (inp[1]) ? node138 : 1'b1;
										assign node138 = (inp[8]) ? 1'b0 : node139;
											assign node139 = (inp[0]) ? 1'b0 : 1'b1;
								assign node143 = (inp[3]) ? 1'b0 : node144;
									assign node144 = (inp[1]) ? 1'b0 : 1'b1;
					assign node148 = (inp[1]) ? node168 : node149;
						assign node149 = (inp[9]) ? node155 : node150;
							assign node150 = (inp[7]) ? node152 : 1'b1;
								assign node152 = (inp[11]) ? 1'b0 : 1'b1;
							assign node155 = (inp[3]) ? node163 : node156;
								assign node156 = (inp[7]) ? node158 : 1'b1;
									assign node158 = (inp[0]) ? 1'b0 : node159;
										assign node159 = (inp[11]) ? 1'b0 : 1'b1;
								assign node163 = (inp[11]) ? 1'b0 : node164;
									assign node164 = (inp[2]) ? 1'b0 : 1'b1;
						assign node168 = (inp[3]) ? node182 : node169;
							assign node169 = (inp[9]) ? node177 : node170;
								assign node170 = (inp[8]) ? node172 : 1'b1;
									assign node172 = (inp[12]) ? 1'b0 : node173;
										assign node173 = (inp[2]) ? 1'b0 : 1'b1;
								assign node177 = (inp[12]) ? 1'b0 : node178;
									assign node178 = (inp[7]) ? 1'b0 : 1'b1;
							assign node182 = (inp[2]) ? 1'b0 : node183;
								assign node183 = (inp[9]) ? node187 : node184;
									assign node184 = (inp[12]) ? 1'b0 : 1'b1;
									assign node187 = (inp[0]) ? 1'b0 : node188;
										assign node188 = (inp[8]) ? 1'b0 : 1'b1;
				assign node193 = (inp[7]) ? node235 : node194;
					assign node194 = (inp[2]) ? node216 : node195;
						assign node195 = (inp[3]) ? node207 : node196;
							assign node196 = (inp[8]) ? node198 : 1'b1;
								assign node198 = (inp[1]) ? node200 : 1'b1;
									assign node200 = (inp[12]) ? node202 : 1'b1;
										assign node202 = (inp[11]) ? 1'b0 : node203;
											assign node203 = (inp[9]) ? 1'b0 : 1'b1;
							assign node207 = (inp[8]) ? 1'b0 : node208;
								assign node208 = (inp[6]) ? node210 : 1'b1;
									assign node210 = (inp[11]) ? 1'b0 : node211;
										assign node211 = (inp[9]) ? 1'b0 : 1'b1;
						assign node216 = (inp[12]) ? node228 : node217;
							assign node217 = (inp[11]) ? node221 : node218;
								assign node218 = (inp[0]) ? 1'b0 : 1'b1;
								assign node221 = (inp[9]) ? 1'b0 : node222;
									assign node222 = (inp[1]) ? node224 : 1'b1;
										assign node224 = (inp[8]) ? 1'b0 : 1'b1;
							assign node228 = (inp[8]) ? 1'b0 : node229;
								assign node229 = (inp[3]) ? 1'b0 : node230;
									assign node230 = (inp[6]) ? 1'b0 : 1'b1;
					assign node235 = (inp[3]) ? node255 : node236;
						assign node236 = (inp[0]) ? node248 : node237;
							assign node237 = (inp[6]) ? node243 : node238;
								assign node238 = (inp[8]) ? node240 : 1'b1;
									assign node240 = (inp[9]) ? 1'b0 : 1'b1;
								assign node243 = (inp[2]) ? 1'b0 : node244;
									assign node244 = (inp[11]) ? 1'b0 : 1'b1;
							assign node248 = (inp[8]) ? 1'b0 : node249;
								assign node249 = (inp[6]) ? 1'b0 : node250;
									assign node250 = (inp[12]) ? 1'b0 : 1'b1;
						assign node255 = (inp[8]) ? 1'b0 : node256;
							assign node256 = (inp[2]) ? 1'b0 : node257;
								assign node257 = (inp[11]) ? 1'b1 : 1'b0;
		assign node262 = (inp[6]) ? node378 : node263;
			assign node263 = (inp[8]) ? node323 : node264;
				assign node264 = (inp[12]) ? node290 : node265;
					assign node265 = (inp[1]) ? node273 : node266;
						assign node266 = (inp[7]) ? node268 : 1'b1;
							assign node268 = (inp[3]) ? node270 : 1'b1;
								assign node270 = (inp[2]) ? 1'b0 : 1'b1;
						assign node273 = (inp[11]) ? node279 : node274;
							assign node274 = (inp[5]) ? node276 : 1'b1;
								assign node276 = (inp[3]) ? 1'b0 : 1'b1;
							assign node279 = (inp[5]) ? node285 : node280;
								assign node280 = (inp[0]) ? node282 : 1'b1;
									assign node282 = (inp[3]) ? 1'b0 : 1'b1;
								assign node285 = (inp[2]) ? 1'b0 : node286;
									assign node286 = (inp[3]) ? 1'b0 : 1'b1;
					assign node290 = (inp[0]) ? node304 : node291;
						assign node291 = (inp[1]) ? node293 : 1'b1;
							assign node293 = (inp[7]) ? node299 : node294;
								assign node294 = (inp[4]) ? node296 : 1'b1;
									assign node296 = (inp[2]) ? 1'b0 : 1'b1;
								assign node299 = (inp[2]) ? 1'b0 : node300;
									assign node300 = (inp[11]) ? 1'b0 : 1'b1;
						assign node304 = (inp[11]) ? node316 : node305;
							assign node305 = (inp[4]) ? node311 : node306;
								assign node306 = (inp[1]) ? 1'b1 : node307;
									assign node307 = (inp[2]) ? 1'b0 : 1'b1;
								assign node311 = (inp[1]) ? 1'b0 : node312;
									assign node312 = (inp[7]) ? 1'b0 : 1'b1;
							assign node316 = (inp[9]) ? 1'b0 : node317;
								assign node317 = (inp[3]) ? 1'b0 : node318;
									assign node318 = (inp[2]) ? 1'b0 : 1'b1;
				assign node323 = (inp[4]) ? node363 : node324;
					assign node324 = (inp[9]) ? node344 : node325;
						assign node325 = (inp[5]) ? node331 : node326;
							assign node326 = (inp[12]) ? node328 : 1'b1;
								assign node328 = (inp[3]) ? 1'b0 : 1'b1;
							assign node331 = (inp[1]) ? node339 : node332;
								assign node332 = (inp[11]) ? node334 : 1'b1;
									assign node334 = (inp[7]) ? 1'b0 : node335;
										assign node335 = (inp[0]) ? 1'b0 : 1'b1;
								assign node339 = (inp[0]) ? 1'b0 : node340;
									assign node340 = (inp[7]) ? 1'b0 : 1'b1;
						assign node344 = (inp[0]) ? node356 : node345;
							assign node345 = (inp[2]) ? node351 : node346;
								assign node346 = (inp[11]) ? node348 : 1'b1;
									assign node348 = (inp[1]) ? 1'b0 : 1'b1;
								assign node351 = (inp[5]) ? 1'b0 : node352;
									assign node352 = (inp[1]) ? 1'b0 : 1'b1;
							assign node356 = (inp[11]) ? 1'b0 : node357;
								assign node357 = (inp[12]) ? 1'b0 : node358;
									assign node358 = (inp[2]) ? 1'b0 : 1'b1;
					assign node363 = (inp[5]) ? 1'b0 : node364;
						assign node364 = (inp[7]) ? node372 : node365;
							assign node365 = (inp[12]) ? node367 : 1'b1;
								assign node367 = (inp[1]) ? 1'b0 : node368;
									assign node368 = (inp[2]) ? 1'b0 : 1'b1;
							assign node372 = (inp[12]) ? 1'b0 : node373;
								assign node373 = (inp[2]) ? 1'b0 : 1'b1;
			assign node378 = (inp[2]) ? node446 : node379;
				assign node379 = (inp[7]) ? node417 : node380;
					assign node380 = (inp[5]) ? node402 : node381;
						assign node381 = (inp[9]) ? node391 : node382;
							assign node382 = (inp[3]) ? node384 : 1'b1;
								assign node384 = (inp[12]) ? node386 : 1'b1;
									assign node386 = (inp[1]) ? 1'b0 : node387;
										assign node387 = (inp[8]) ? 1'b0 : 1'b1;
							assign node391 = (inp[8]) ? node397 : node392;
								assign node392 = (inp[1]) ? node394 : 1'b1;
									assign node394 = (inp[0]) ? 1'b0 : 1'b1;
								assign node397 = (inp[0]) ? 1'b0 : node398;
									assign node398 = (inp[1]) ? 1'b0 : 1'b1;
						assign node402 = (inp[12]) ? node408 : node403;
							assign node403 = (inp[1]) ? node405 : 1'b1;
								assign node405 = (inp[8]) ? 1'b1 : 1'b0;
							assign node408 = (inp[3]) ? 1'b0 : node409;
								assign node409 = (inp[1]) ? 1'b0 : node410;
									assign node410 = (inp[11]) ? 1'b0 : node411;
										assign node411 = (inp[9]) ? 1'b0 : 1'b1;
					assign node417 = (inp[1]) ? node437 : node418;
						assign node418 = (inp[3]) ? node430 : node419;
							assign node419 = (inp[9]) ? node421 : 1'b1;
								assign node421 = (inp[8]) ? node423 : 1'b1;
									assign node423 = (inp[0]) ? 1'b0 : node424;
										assign node424 = (inp[11]) ? 1'b0 : node425;
											assign node425 = (inp[12]) ? 1'b0 : 1'b1;
							assign node430 = (inp[11]) ? 1'b0 : node431;
								assign node431 = (inp[4]) ? 1'b0 : node432;
									assign node432 = (inp[8]) ? 1'b0 : 1'b1;
						assign node437 = (inp[4]) ? 1'b0 : node438;
							assign node438 = (inp[12]) ? 1'b0 : node439;
								assign node439 = (inp[8]) ? 1'b0 : node440;
									assign node440 = (inp[0]) ? 1'b0 : 1'b1;
				assign node446 = (inp[5]) ? node476 : node447;
					assign node447 = (inp[3]) ? node467 : node448;
						assign node448 = (inp[12]) ? node458 : node449;
							assign node449 = (inp[9]) ? node451 : 1'b1;
								assign node451 = (inp[4]) ? 1'b0 : node452;
									assign node452 = (inp[8]) ? node454 : 1'b1;
										assign node454 = (inp[7]) ? 1'b0 : 1'b1;
							assign node458 = (inp[4]) ? 1'b0 : node459;
								assign node459 = (inp[1]) ? 1'b0 : node460;
									assign node460 = (inp[7]) ? node462 : 1'b1;
										assign node462 = (inp[8]) ? 1'b0 : 1'b1;
						assign node467 = (inp[9]) ? 1'b0 : node468;
							assign node468 = (inp[0]) ? 1'b0 : node469;
								assign node469 = (inp[7]) ? 1'b0 : node470;
									assign node470 = (inp[8]) ? 1'b0 : 1'b1;
					assign node476 = (inp[8]) ? 1'b0 : node477;
						assign node477 = (inp[11]) ? 1'b0 : node478;
							assign node478 = (inp[0]) ? node486 : node479;
								assign node479 = (inp[3]) ? 1'b0 : node480;
									assign node480 = (inp[9]) ? node482 : 1'b1;
										assign node482 = (inp[7]) ? 1'b1 : 1'b0;
								assign node486 = (inp[7]) ? 1'b0 : node487;
									assign node487 = (inp[9]) ? 1'b0 : node488;
										assign node488 = (inp[4]) ? 1'b0 : 1'b1;

endmodule