module dtc_split33_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;

	assign outp = (inp[2]) ? node90 : node1;
		assign node1 = (inp[3]) ? node49 : node2;
			assign node2 = (inp[10]) ? node26 : node3;
				assign node3 = (inp[4]) ? node17 : node4;
					assign node4 = (inp[5]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[9]) ? node10 : 3'b111;
								assign node10 = (inp[1]) ? 3'b110 : node11;
									assign node11 = (inp[6]) ? node13 : 3'b111;
										assign node13 = (inp[11]) ? 3'b110 : 3'b111;
					assign node17 = (inp[5]) ? 3'b111 : node18;
						assign node18 = (inp[7]) ? node20 : 3'b110;
							assign node20 = (inp[8]) ? node22 : 3'b110;
								assign node22 = (inp[9]) ? 3'b111 : 3'b110;
				assign node26 = (inp[9]) ? node40 : node27;
					assign node27 = (inp[5]) ? 3'b110 : node28;
						assign node28 = (inp[4]) ? node30 : 3'b110;
							assign node30 = (inp[7]) ? 3'b110 : node31;
								assign node31 = (inp[8]) ? node33 : 3'b111;
									assign node33 = (inp[6]) ? node35 : 3'b111;
										assign node35 = (inp[11]) ? 3'b110 : 3'b111;
					assign node40 = (inp[5]) ? node42 : 3'b110;
						assign node42 = (inp[4]) ? 3'b011 : node43;
							assign node43 = (inp[8]) ? node45 : 3'b110;
								assign node45 = (inp[7]) ? 3'b111 : 3'b110;
			assign node49 = (inp[4]) ? node63 : node50;
				assign node50 = (inp[10]) ? node58 : node51;
					assign node51 = (inp[7]) ? node53 : 3'b111;
						assign node53 = (inp[5]) ? node55 : 3'b111;
							assign node55 = (inp[9]) ? 3'b110 : 3'b111;
					assign node58 = (inp[9]) ? node60 : 3'b110;
						assign node60 = (inp[5]) ? 3'b011 : 3'b110;
				assign node63 = (inp[5]) ? node81 : node64;
					assign node64 = (inp[9]) ? node66 : 3'b011;
						assign node66 = (inp[10]) ? node74 : node67;
							assign node67 = (inp[7]) ? 3'b010 : node68;
								assign node68 = (inp[11]) ? node70 : 3'b011;
									assign node70 = (inp[6]) ? 3'b010 : 3'b011;
							assign node74 = (inp[6]) ? node76 : 3'b011;
								assign node76 = (inp[11]) ? node78 : 3'b011;
									assign node78 = (inp[8]) ? 3'b010 : 3'b011;
					assign node81 = (inp[9]) ? node83 : 3'b010;
						assign node83 = (inp[10]) ? 3'b010 : node84;
							assign node84 = (inp[8]) ? node86 : 3'b010;
								assign node86 = (inp[7]) ? 3'b011 : 3'b010;
		assign node90 = (inp[4]) ? node136 : node91;
			assign node91 = (inp[10]) ? node115 : node92;
				assign node92 = (inp[5]) ? node104 : node93;
					assign node93 = (inp[3]) ? node95 : 3'b011;
						assign node95 = (inp[9]) ? 3'b010 : node96;
							assign node96 = (inp[8]) ? node98 : 3'b011;
								assign node98 = (inp[0]) ? 3'b011 : node99;
									assign node99 = (inp[11]) ? 3'b010 : 3'b011;
					assign node104 = (inp[7]) ? 3'b010 : node105;
						assign node105 = (inp[9]) ? 3'b010 : node106;
							assign node106 = (inp[3]) ? 3'b010 : node107;
								assign node107 = (inp[6]) ? node109 : 3'b011;
									assign node109 = (inp[1]) ? 3'b010 : 3'b011;
				assign node115 = (inp[3]) ? node125 : node116;
					assign node116 = (inp[5]) ? 3'b011 : node117;
						assign node117 = (inp[9]) ? node119 : 3'b010;
							assign node119 = (inp[7]) ? node121 : 3'b010;
								assign node121 = (inp[8]) ? 3'b011 : 3'b010;
					assign node125 = (inp[5]) ? node127 : 3'b111;
						assign node127 = (inp[9]) ? 3'b110 : node128;
							assign node128 = (inp[6]) ? node130 : 3'b111;
								assign node130 = (inp[11]) ? node132 : 3'b111;
									assign node132 = (inp[7]) ? 3'b110 : 3'b111;
			assign node136 = (inp[3]) ? node160 : node137;
				assign node137 = (inp[5]) ? node151 : node138;
					assign node138 = (inp[10]) ? node140 : 3'b101;
						assign node140 = (inp[9]) ? node142 : 3'b101;
							assign node142 = (inp[7]) ? 3'b100 : node143;
								assign node143 = (inp[1]) ? 3'b101 : node144;
									assign node144 = (inp[11]) ? node146 : 3'b101;
										assign node146 = (inp[6]) ? 3'b100 : 3'b101;
					assign node151 = (inp[9]) ? node153 : 3'b100;
						assign node153 = (inp[10]) ? 3'b001 : node154;
							assign node154 = (inp[8]) ? node156 : 3'b100;
								assign node156 = (inp[7]) ? 3'b101 : 3'b100;
				assign node160 = (inp[10]) ? node184 : node161;
					assign node161 = (inp[9]) ? node177 : node162;
						assign node162 = (inp[7]) ? node170 : node163;
							assign node163 = (inp[5]) ? 3'b001 : node164;
								assign node164 = (inp[6]) ? node166 : 3'b001;
									assign node166 = (inp[11]) ? 3'b000 : 3'b001;
							assign node170 = (inp[5]) ? node172 : 3'b000;
								assign node172 = (inp[6]) ? node174 : 3'b001;
									assign node174 = (inp[8]) ? 3'b000 : 3'b001;
						assign node177 = (inp[5]) ? 3'b000 : node178;
							assign node178 = (inp[7]) ? node180 : 3'b000;
								assign node180 = (inp[8]) ? 3'b001 : 3'b000;
					assign node184 = (inp[5]) ? node200 : node185;
						assign node185 = (inp[9]) ? node195 : node186;
							assign node186 = (inp[11]) ? node188 : 3'b101;
								assign node188 = (inp[0]) ? 3'b101 : node189;
									assign node189 = (inp[8]) ? node191 : 3'b101;
										assign node191 = (inp[7]) ? 3'b100 : 3'b101;
							assign node195 = (inp[8]) ? node197 : 3'b100;
								assign node197 = (inp[7]) ? 3'b101 : 3'b100;
						assign node200 = (inp[9]) ? node210 : node201;
							assign node201 = (inp[7]) ? 3'b100 : node202;
								assign node202 = (inp[6]) ? node204 : 3'b101;
									assign node204 = (inp[8]) ? node206 : 3'b101;
										assign node206 = (inp[11]) ? 3'b100 : 3'b101;
							assign node210 = (inp[7]) ? node218 : node211;
								assign node211 = (inp[11]) ? node213 : 3'b001;
									assign node213 = (inp[6]) ? node215 : 3'b001;
										assign node215 = (inp[8]) ? 3'b000 : 3'b001;
								assign node218 = (inp[11]) ? 3'b000 : node219;
									assign node219 = (inp[8]) ? 3'b001 : 3'b000;

endmodule