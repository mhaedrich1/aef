module dtc_split25_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node11;
	wire [14-1:0] node13;
	wire [14-1:0] node14;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node26;
	wire [14-1:0] node27;
	wire [14-1:0] node31;
	wire [14-1:0] node34;
	wire [14-1:0] node35;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node43;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node46;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node53;
	wire [14-1:0] node57;
	wire [14-1:0] node58;
	wire [14-1:0] node59;
	wire [14-1:0] node62;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node77;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node87;
	wire [14-1:0] node89;
	wire [14-1:0] node92;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node95;
	wire [14-1:0] node98;
	wire [14-1:0] node100;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node111;
	wire [14-1:0] node113;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node119;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node127;
	wire [14-1:0] node129;
	wire [14-1:0] node130;
	wire [14-1:0] node134;
	wire [14-1:0] node135;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node142;
	wire [14-1:0] node145;
	wire [14-1:0] node146;
	wire [14-1:0] node150;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node157;
	wire [14-1:0] node159;
	wire [14-1:0] node162;
	wire [14-1:0] node163;
	wire [14-1:0] node166;
	wire [14-1:0] node167;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node175;
	wire [14-1:0] node176;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node181;
	wire [14-1:0] node182;
	wire [14-1:0] node186;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node191;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node198;
	wire [14-1:0] node201;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node216;
	wire [14-1:0] node218;
	wire [14-1:0] node221;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node229;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node233;
	wire [14-1:0] node236;
	wire [14-1:0] node237;
	wire [14-1:0] node242;
	wire [14-1:0] node243;
	wire [14-1:0] node246;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node257;
	wire [14-1:0] node258;
	wire [14-1:0] node259;
	wire [14-1:0] node261;
	wire [14-1:0] node266;
	wire [14-1:0] node267;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node273;
	wire [14-1:0] node276;
	wire [14-1:0] node278;
	wire [14-1:0] node279;
	wire [14-1:0] node282;
	wire [14-1:0] node284;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node293;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node298;
	wire [14-1:0] node302;
	wire [14-1:0] node304;
	wire [14-1:0] node305;
	wire [14-1:0] node307;
	wire [14-1:0] node310;
	wire [14-1:0] node313;
	wire [14-1:0] node314;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node320;
	wire [14-1:0] node323;
	wire [14-1:0] node327;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node333;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node342;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node349;
	wire [14-1:0] node352;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node359;
	wire [14-1:0] node361;
	wire [14-1:0] node364;
	wire [14-1:0] node365;
	wire [14-1:0] node366;
	wire [14-1:0] node367;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node374;
	wire [14-1:0] node376;
	wire [14-1:0] node379;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node384;
	wire [14-1:0] node386;
	wire [14-1:0] node389;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node395;
	wire [14-1:0] node398;
	wire [14-1:0] node400;
	wire [14-1:0] node401;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node407;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node416;
	wire [14-1:0] node417;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node425;
	wire [14-1:0] node427;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node434;
	wire [14-1:0] node438;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node443;
	wire [14-1:0] node445;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node453;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node459;
	wire [14-1:0] node460;
	wire [14-1:0] node462;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node470;
	wire [14-1:0] node471;
	wire [14-1:0] node472;
	wire [14-1:0] node475;
	wire [14-1:0] node476;
	wire [14-1:0] node478;
	wire [14-1:0] node482;
	wire [14-1:0] node483;
	wire [14-1:0] node486;
	wire [14-1:0] node488;
	wire [14-1:0] node491;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node495;
	wire [14-1:0] node497;
	wire [14-1:0] node500;
	wire [14-1:0] node502;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node509;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node520;
	wire [14-1:0] node522;
	wire [14-1:0] node523;
	wire [14-1:0] node527;
	wire [14-1:0] node529;
	wire [14-1:0] node532;
	wire [14-1:0] node534;
	wire [14-1:0] node535;
	wire [14-1:0] node538;
	wire [14-1:0] node541;
	wire [14-1:0] node543;
	wire [14-1:0] node544;
	wire [14-1:0] node547;
	wire [14-1:0] node548;
	wire [14-1:0] node552;
	wire [14-1:0] node553;
	wire [14-1:0] node554;
	wire [14-1:0] node556;
	wire [14-1:0] node557;
	wire [14-1:0] node560;
	wire [14-1:0] node562;
	wire [14-1:0] node565;
	wire [14-1:0] node566;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node576;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node584;
	wire [14-1:0] node587;
	wire [14-1:0] node589;
	wire [14-1:0] node590;
	wire [14-1:0] node594;
	wire [14-1:0] node595;
	wire [14-1:0] node598;
	wire [14-1:0] node600;
	wire [14-1:0] node603;
	wire [14-1:0] node604;
	wire [14-1:0] node605;
	wire [14-1:0] node606;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node613;
	wire [14-1:0] node616;
	wire [14-1:0] node619;
	wire [14-1:0] node620;
	wire [14-1:0] node621;
	wire [14-1:0] node624;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node630;
	wire [14-1:0] node631;
	wire [14-1:0] node633;
	wire [14-1:0] node634;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node644;
	wire [14-1:0] node648;
	wire [14-1:0] node652;
	wire [14-1:0] node653;
	wire [14-1:0] node654;
	wire [14-1:0] node655;
	wire [14-1:0] node659;
	wire [14-1:0] node662;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node668;
	wire [14-1:0] node669;
	wire [14-1:0] node671;
	wire [14-1:0] node675;
	wire [14-1:0] node676;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node680;
	wire [14-1:0] node683;
	wire [14-1:0] node684;
	wire [14-1:0] node685;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node692;
	wire [14-1:0] node693;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node701;
	wire [14-1:0] node703;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node711;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node719;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node728;
	wire [14-1:0] node729;
	wire [14-1:0] node732;
	wire [14-1:0] node734;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node740;
	wire [14-1:0] node742;
	wire [14-1:0] node745;
	wire [14-1:0] node746;
	wire [14-1:0] node749;
	wire [14-1:0] node751;
	wire [14-1:0] node753;
	wire [14-1:0] node755;
	wire [14-1:0] node758;
	wire [14-1:0] node759;
	wire [14-1:0] node760;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node763;
	wire [14-1:0] node764;
	wire [14-1:0] node766;
	wire [14-1:0] node767;
	wire [14-1:0] node769;
	wire [14-1:0] node770;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node777;
	wire [14-1:0] node778;
	wire [14-1:0] node780;
	wire [14-1:0] node784;
	wire [14-1:0] node787;
	wire [14-1:0] node789;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node798;
	wire [14-1:0] node801;
	wire [14-1:0] node802;
	wire [14-1:0] node803;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node816;
	wire [14-1:0] node819;
	wire [14-1:0] node820;
	wire [14-1:0] node821;
	wire [14-1:0] node822;
	wire [14-1:0] node823;
	wire [14-1:0] node826;
	wire [14-1:0] node829;
	wire [14-1:0] node832;
	wire [14-1:0] node833;
	wire [14-1:0] node836;
	wire [14-1:0] node837;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node847;
	wire [14-1:0] node849;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node858;
	wire [14-1:0] node859;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node864;
	wire [14-1:0] node868;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node878;
	wire [14-1:0] node881;
	wire [14-1:0] node884;
	wire [14-1:0] node885;
	wire [14-1:0] node888;
	wire [14-1:0] node891;
	wire [14-1:0] node892;
	wire [14-1:0] node894;
	wire [14-1:0] node897;
	wire [14-1:0] node898;
	wire [14-1:0] node902;
	wire [14-1:0] node903;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node907;
	wire [14-1:0] node910;
	wire [14-1:0] node911;
	wire [14-1:0] node915;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node921;
	wire [14-1:0] node923;
	wire [14-1:0] node925;
	wire [14-1:0] node927;
	wire [14-1:0] node930;
	wire [14-1:0] node931;
	wire [14-1:0] node932;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node939;
	wire [14-1:0] node941;
	wire [14-1:0] node944;
	wire [14-1:0] node947;
	wire [14-1:0] node948;
	wire [14-1:0] node949;
	wire [14-1:0] node950;
	wire [14-1:0] node951;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node955;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node963;
	wire [14-1:0] node964;
	wire [14-1:0] node967;
	wire [14-1:0] node970;
	wire [14-1:0] node971;
	wire [14-1:0] node972;
	wire [14-1:0] node976;
	wire [14-1:0] node979;
	wire [14-1:0] node980;
	wire [14-1:0] node981;
	wire [14-1:0] node983;
	wire [14-1:0] node986;
	wire [14-1:0] node987;
	wire [14-1:0] node991;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node998;
	wire [14-1:0] node999;
	wire [14-1:0] node1000;
	wire [14-1:0] node1002;
	wire [14-1:0] node1003;
	wire [14-1:0] node1004;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1012;
	wire [14-1:0] node1015;
	wire [14-1:0] node1018;
	wire [14-1:0] node1019;
	wire [14-1:0] node1021;
	wire [14-1:0] node1024;
	wire [14-1:0] node1026;
	wire [14-1:0] node1028;
	wire [14-1:0] node1031;
	wire [14-1:0] node1032;
	wire [14-1:0] node1033;
	wire [14-1:0] node1034;
	wire [14-1:0] node1036;
	wire [14-1:0] node1037;
	wire [14-1:0] node1042;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1047;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1056;
	wire [14-1:0] node1057;
	wire [14-1:0] node1058;
	wire [14-1:0] node1062;
	wire [14-1:0] node1064;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1069;
	wire [14-1:0] node1070;
	wire [14-1:0] node1073;
	wire [14-1:0] node1075;
	wire [14-1:0] node1078;
	wire [14-1:0] node1079;
	wire [14-1:0] node1081;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1087;
	wire [14-1:0] node1090;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1096;
	wire [14-1:0] node1098;
	wire [14-1:0] node1101;
	wire [14-1:0] node1102;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1108;
	wire [14-1:0] node1109;
	wire [14-1:0] node1110;
	wire [14-1:0] node1111;
	wire [14-1:0] node1112;
	wire [14-1:0] node1115;
	wire [14-1:0] node1116;
	wire [14-1:0] node1118;
	wire [14-1:0] node1122;
	wire [14-1:0] node1123;
	wire [14-1:0] node1124;
	wire [14-1:0] node1127;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1133;
	wire [14-1:0] node1134;
	wire [14-1:0] node1137;
	wire [14-1:0] node1140;
	wire [14-1:0] node1141;
	wire [14-1:0] node1142;
	wire [14-1:0] node1147;
	wire [14-1:0] node1150;
	wire [14-1:0] node1151;
	wire [14-1:0] node1152;
	wire [14-1:0] node1153;
	wire [14-1:0] node1156;
	wire [14-1:0] node1158;
	wire [14-1:0] node1161;
	wire [14-1:0] node1163;
	wire [14-1:0] node1164;
	wire [14-1:0] node1167;
	wire [14-1:0] node1170;
	wire [14-1:0] node1171;
	wire [14-1:0] node1172;
	wire [14-1:0] node1174;
	wire [14-1:0] node1177;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1183;
	wire [14-1:0] node1185;
	wire [14-1:0] node1188;
	wire [14-1:0] node1191;
	wire [14-1:0] node1192;
	wire [14-1:0] node1193;
	wire [14-1:0] node1194;
	wire [14-1:0] node1197;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1201;
	wire [14-1:0] node1203;
	wire [14-1:0] node1208;
	wire [14-1:0] node1209;
	wire [14-1:0] node1211;
	wire [14-1:0] node1212;
	wire [14-1:0] node1216;
	wire [14-1:0] node1218;
	wire [14-1:0] node1219;
	wire [14-1:0] node1220;
	wire [14-1:0] node1223;
	wire [14-1:0] node1226;
	wire [14-1:0] node1227;
	wire [14-1:0] node1231;
	wire [14-1:0] node1232;
	wire [14-1:0] node1233;
	wire [14-1:0] node1235;
	wire [14-1:0] node1236;
	wire [14-1:0] node1240;
	wire [14-1:0] node1241;
	wire [14-1:0] node1242;
	wire [14-1:0] node1243;
	wire [14-1:0] node1247;
	wire [14-1:0] node1249;
	wire [14-1:0] node1252;
	wire [14-1:0] node1253;
	wire [14-1:0] node1257;
	wire [14-1:0] node1258;
	wire [14-1:0] node1259;
	wire [14-1:0] node1261;
	wire [14-1:0] node1264;
	wire [14-1:0] node1267;
	wire [14-1:0] node1269;
	wire [14-1:0] node1272;
	wire [14-1:0] node1273;
	wire [14-1:0] node1274;
	wire [14-1:0] node1275;
	wire [14-1:0] node1276;
	wire [14-1:0] node1277;
	wire [14-1:0] node1279;
	wire [14-1:0] node1283;
	wire [14-1:0] node1284;
	wire [14-1:0] node1286;
	wire [14-1:0] node1290;
	wire [14-1:0] node1291;
	wire [14-1:0] node1292;
	wire [14-1:0] node1296;
	wire [14-1:0] node1297;
	wire [14-1:0] node1301;
	wire [14-1:0] node1302;
	wire [14-1:0] node1303;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1308;
	wire [14-1:0] node1312;
	wire [14-1:0] node1314;
	wire [14-1:0] node1317;
	wire [14-1:0] node1318;
	wire [14-1:0] node1319;
	wire [14-1:0] node1321;
	wire [14-1:0] node1324;
	wire [14-1:0] node1326;
	wire [14-1:0] node1327;
	wire [14-1:0] node1331;
	wire [14-1:0] node1333;
	wire [14-1:0] node1336;
	wire [14-1:0] node1337;
	wire [14-1:0] node1338;
	wire [14-1:0] node1339;
	wire [14-1:0] node1340;
	wire [14-1:0] node1341;
	wire [14-1:0] node1344;
	wire [14-1:0] node1347;
	wire [14-1:0] node1348;
	wire [14-1:0] node1352;
	wire [14-1:0] node1353;
	wire [14-1:0] node1357;
	wire [14-1:0] node1358;
	wire [14-1:0] node1359;
	wire [14-1:0] node1361;
	wire [14-1:0] node1362;
	wire [14-1:0] node1366;
	wire [14-1:0] node1367;
	wire [14-1:0] node1371;
	wire [14-1:0] node1372;
	wire [14-1:0] node1374;
	wire [14-1:0] node1375;
	wire [14-1:0] node1379;
	wire [14-1:0] node1381;
	wire [14-1:0] node1384;
	wire [14-1:0] node1385;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1392;
	wire [14-1:0] node1395;
	wire [14-1:0] node1397;
	wire [14-1:0] node1399;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1404;
	wire [14-1:0] node1408;
	wire [14-1:0] node1409;
	wire [14-1:0] node1410;
	wire [14-1:0] node1413;
	wire [14-1:0] node1416;
	wire [14-1:0] node1418;
	wire [14-1:0] node1421;
	wire [14-1:0] node1422;
	wire [14-1:0] node1423;
	wire [14-1:0] node1424;
	wire [14-1:0] node1425;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1428;
	wire [14-1:0] node1429;
	wire [14-1:0] node1431;
	wire [14-1:0] node1434;
	wire [14-1:0] node1435;
	wire [14-1:0] node1437;
	wire [14-1:0] node1441;
	wire [14-1:0] node1442;
	wire [14-1:0] node1443;
	wire [14-1:0] node1446;
	wire [14-1:0] node1448;
	wire [14-1:0] node1451;
	wire [14-1:0] node1452;
	wire [14-1:0] node1456;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1460;
	wire [14-1:0] node1463;
	wire [14-1:0] node1464;
	wire [14-1:0] node1466;
	wire [14-1:0] node1467;
	wire [14-1:0] node1471;
	wire [14-1:0] node1473;
	wire [14-1:0] node1476;
	wire [14-1:0] node1477;
	wire [14-1:0] node1479;
	wire [14-1:0] node1481;
	wire [14-1:0] node1482;
	wire [14-1:0] node1486;
	wire [14-1:0] node1487;
	wire [14-1:0] node1488;
	wire [14-1:0] node1492;
	wire [14-1:0] node1495;
	wire [14-1:0] node1496;
	wire [14-1:0] node1497;
	wire [14-1:0] node1498;
	wire [14-1:0] node1499;
	wire [14-1:0] node1500;
	wire [14-1:0] node1505;
	wire [14-1:0] node1507;
	wire [14-1:0] node1508;
	wire [14-1:0] node1512;
	wire [14-1:0] node1514;
	wire [14-1:0] node1515;
	wire [14-1:0] node1519;
	wire [14-1:0] node1520;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1527;
	wire [14-1:0] node1528;
	wire [14-1:0] node1529;
	wire [14-1:0] node1532;
	wire [14-1:0] node1535;
	wire [14-1:0] node1537;
	wire [14-1:0] node1540;
	wire [14-1:0] node1541;
	wire [14-1:0] node1542;
	wire [14-1:0] node1543;
	wire [14-1:0] node1544;
	wire [14-1:0] node1546;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1554;
	wire [14-1:0] node1555;
	wire [14-1:0] node1556;
	wire [14-1:0] node1557;
	wire [14-1:0] node1559;
	wire [14-1:0] node1563;
	wire [14-1:0] node1565;
	wire [14-1:0] node1569;
	wire [14-1:0] node1570;
	wire [14-1:0] node1571;
	wire [14-1:0] node1573;
	wire [14-1:0] node1576;
	wire [14-1:0] node1577;
	wire [14-1:0] node1578;
	wire [14-1:0] node1580;
	wire [14-1:0] node1584;
	wire [14-1:0] node1587;
	wire [14-1:0] node1589;
	wire [14-1:0] node1592;
	wire [14-1:0] node1593;
	wire [14-1:0] node1594;
	wire [14-1:0] node1595;
	wire [14-1:0] node1596;
	wire [14-1:0] node1600;
	wire [14-1:0] node1601;
	wire [14-1:0] node1605;
	wire [14-1:0] node1606;
	wire [14-1:0] node1607;
	wire [14-1:0] node1610;
	wire [14-1:0] node1611;
	wire [14-1:0] node1615;
	wire [14-1:0] node1618;
	wire [14-1:0] node1619;
	wire [14-1:0] node1620;
	wire [14-1:0] node1622;
	wire [14-1:0] node1625;
	wire [14-1:0] node1627;
	wire [14-1:0] node1630;
	wire [14-1:0] node1632;
	wire [14-1:0] node1635;
	wire [14-1:0] node1636;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1639;
	wire [14-1:0] node1640;
	wire [14-1:0] node1643;
	wire [14-1:0] node1644;
	wire [14-1:0] node1645;
	wire [14-1:0] node1649;
	wire [14-1:0] node1652;
	wire [14-1:0] node1653;
	wire [14-1:0] node1655;
	wire [14-1:0] node1659;
	wire [14-1:0] node1660;
	wire [14-1:0] node1663;
	wire [14-1:0] node1666;
	wire [14-1:0] node1667;
	wire [14-1:0] node1668;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1672;
	wire [14-1:0] node1675;
	wire [14-1:0] node1678;
	wire [14-1:0] node1679;
	wire [14-1:0] node1680;
	wire [14-1:0] node1685;
	wire [14-1:0] node1686;
	wire [14-1:0] node1687;
	wire [14-1:0] node1691;
	wire [14-1:0] node1692;
	wire [14-1:0] node1695;
	wire [14-1:0] node1698;
	wire [14-1:0] node1699;
	wire [14-1:0] node1700;
	wire [14-1:0] node1701;
	wire [14-1:0] node1702;
	wire [14-1:0] node1704;
	wire [14-1:0] node1709;
	wire [14-1:0] node1712;
	wire [14-1:0] node1714;
	wire [14-1:0] node1717;
	wire [14-1:0] node1718;
	wire [14-1:0] node1719;
	wire [14-1:0] node1720;
	wire [14-1:0] node1721;
	wire [14-1:0] node1722;
	wire [14-1:0] node1723;
	wire [14-1:0] node1727;
	wire [14-1:0] node1730;
	wire [14-1:0] node1731;
	wire [14-1:0] node1735;
	wire [14-1:0] node1736;
	wire [14-1:0] node1737;
	wire [14-1:0] node1741;
	wire [14-1:0] node1744;
	wire [14-1:0] node1745;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1750;
	wire [14-1:0] node1751;
	wire [14-1:0] node1755;
	wire [14-1:0] node1757;
	wire [14-1:0] node1760;
	wire [14-1:0] node1761;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1767;
	wire [14-1:0] node1768;
	wire [14-1:0] node1769;
	wire [14-1:0] node1773;
	wire [14-1:0] node1774;
	wire [14-1:0] node1778;
	wire [14-1:0] node1780;
	wire [14-1:0] node1782;
	wire [14-1:0] node1784;
	wire [14-1:0] node1787;
	wire [14-1:0] node1788;
	wire [14-1:0] node1789;
	wire [14-1:0] node1790;
	wire [14-1:0] node1794;
	wire [14-1:0] node1796;
	wire [14-1:0] node1799;
	wire [14-1:0] node1800;
	wire [14-1:0] node1802;
	wire [14-1:0] node1805;
	wire [14-1:0] node1806;
	wire [14-1:0] node1807;
	wire [14-1:0] node1812;
	wire [14-1:0] node1813;
	wire [14-1:0] node1814;
	wire [14-1:0] node1815;
	wire [14-1:0] node1816;
	wire [14-1:0] node1817;
	wire [14-1:0] node1818;
	wire [14-1:0] node1820;
	wire [14-1:0] node1823;
	wire [14-1:0] node1824;
	wire [14-1:0] node1828;
	wire [14-1:0] node1829;
	wire [14-1:0] node1830;
	wire [14-1:0] node1832;
	wire [14-1:0] node1835;
	wire [14-1:0] node1836;
	wire [14-1:0] node1837;
	wire [14-1:0] node1842;
	wire [14-1:0] node1843;
	wire [14-1:0] node1847;
	wire [14-1:0] node1848;
	wire [14-1:0] node1849;
	wire [14-1:0] node1852;
	wire [14-1:0] node1855;
	wire [14-1:0] node1856;
	wire [14-1:0] node1857;
	wire [14-1:0] node1861;
	wire [14-1:0] node1862;
	wire [14-1:0] node1865;
	wire [14-1:0] node1866;
	wire [14-1:0] node1870;
	wire [14-1:0] node1871;
	wire [14-1:0] node1872;
	wire [14-1:0] node1873;
	wire [14-1:0] node1874;
	wire [14-1:0] node1878;
	wire [14-1:0] node1879;
	wire [14-1:0] node1882;
	wire [14-1:0] node1885;
	wire [14-1:0] node1887;
	wire [14-1:0] node1888;
	wire [14-1:0] node1892;
	wire [14-1:0] node1893;
	wire [14-1:0] node1894;
	wire [14-1:0] node1897;
	wire [14-1:0] node1898;
	wire [14-1:0] node1899;
	wire [14-1:0] node1903;
	wire [14-1:0] node1906;
	wire [14-1:0] node1907;
	wire [14-1:0] node1908;
	wire [14-1:0] node1912;
	wire [14-1:0] node1913;
	wire [14-1:0] node1917;
	wire [14-1:0] node1918;
	wire [14-1:0] node1919;
	wire [14-1:0] node1920;
	wire [14-1:0] node1921;
	wire [14-1:0] node1925;
	wire [14-1:0] node1926;
	wire [14-1:0] node1928;
	wire [14-1:0] node1931;
	wire [14-1:0] node1932;
	wire [14-1:0] node1936;
	wire [14-1:0] node1937;
	wire [14-1:0] node1938;
	wire [14-1:0] node1939;
	wire [14-1:0] node1942;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1950;
	wire [14-1:0] node1951;
	wire [14-1:0] node1953;
	wire [14-1:0] node1954;
	wire [14-1:0] node1957;
	wire [14-1:0] node1958;
	wire [14-1:0] node1963;
	wire [14-1:0] node1964;
	wire [14-1:0] node1965;
	wire [14-1:0] node1966;
	wire [14-1:0] node1967;
	wire [14-1:0] node1969;
	wire [14-1:0] node1973;
	wire [14-1:0] node1976;
	wire [14-1:0] node1977;
	wire [14-1:0] node1978;
	wire [14-1:0] node1979;
	wire [14-1:0] node1983;
	wire [14-1:0] node1986;
	wire [14-1:0] node1987;
	wire [14-1:0] node1991;
	wire [14-1:0] node1992;
	wire [14-1:0] node1993;
	wire [14-1:0] node1994;
	wire [14-1:0] node1998;
	wire [14-1:0] node1999;
	wire [14-1:0] node2002;
	wire [14-1:0] node2003;
	wire [14-1:0] node2007;
	wire [14-1:0] node2008;
	wire [14-1:0] node2009;
	wire [14-1:0] node2010;
	wire [14-1:0] node2015;
	wire [14-1:0] node2017;
	wire [14-1:0] node2020;
	wire [14-1:0] node2021;
	wire [14-1:0] node2022;
	wire [14-1:0] node2023;
	wire [14-1:0] node2024;
	wire [14-1:0] node2025;
	wire [14-1:0] node2029;
	wire [14-1:0] node2030;
	wire [14-1:0] node2032;
	wire [14-1:0] node2035;
	wire [14-1:0] node2036;
	wire [14-1:0] node2040;
	wire [14-1:0] node2041;
	wire [14-1:0] node2042;
	wire [14-1:0] node2044;
	wire [14-1:0] node2048;
	wire [14-1:0] node2050;
	wire [14-1:0] node2053;
	wire [14-1:0] node2054;
	wire [14-1:0] node2055;
	wire [14-1:0] node2056;
	wire [14-1:0] node2058;
	wire [14-1:0] node2059;
	wire [14-1:0] node2061;
	wire [14-1:0] node2065;
	wire [14-1:0] node2067;
	wire [14-1:0] node2070;
	wire [14-1:0] node2071;
	wire [14-1:0] node2073;
	wire [14-1:0] node2076;
	wire [14-1:0] node2078;
	wire [14-1:0] node2081;
	wire [14-1:0] node2082;
	wire [14-1:0] node2083;
	wire [14-1:0] node2084;
	wire [14-1:0] node2087;
	wire [14-1:0] node2089;
	wire [14-1:0] node2093;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2100;
	wire [14-1:0] node2101;
	wire [14-1:0] node2102;
	wire [14-1:0] node2103;
	wire [14-1:0] node2105;
	wire [14-1:0] node2106;
	wire [14-1:0] node2107;
	wire [14-1:0] node2109;
	wire [14-1:0] node2114;
	wire [14-1:0] node2115;
	wire [14-1:0] node2117;
	wire [14-1:0] node2119;
	wire [14-1:0] node2120;
	wire [14-1:0] node2124;
	wire [14-1:0] node2127;
	wire [14-1:0] node2128;
	wire [14-1:0] node2130;
	wire [14-1:0] node2131;
	wire [14-1:0] node2132;
	wire [14-1:0] node2137;
	wire [14-1:0] node2139;
	wire [14-1:0] node2141;
	wire [14-1:0] node2144;
	wire [14-1:0] node2145;
	wire [14-1:0] node2146;
	wire [14-1:0] node2147;
	wire [14-1:0] node2148;
	wire [14-1:0] node2149;
	wire [14-1:0] node2153;
	wire [14-1:0] node2155;
	wire [14-1:0] node2157;
	wire [14-1:0] node2161;
	wire [14-1:0] node2162;
	wire [14-1:0] node2163;
	wire [14-1:0] node2167;
	wire [14-1:0] node2169;
	wire [14-1:0] node2170;
	wire [14-1:0] node2172;
	wire [14-1:0] node2175;
	wire [14-1:0] node2178;
	wire [14-1:0] node2179;
	wire [14-1:0] node2180;
	wire [14-1:0] node2183;
	wire [14-1:0] node2185;
	wire [14-1:0] node2188;
	wire [14-1:0] node2189;
	wire [14-1:0] node2190;
	wire [14-1:0] node2192;
	wire [14-1:0] node2195;
	wire [14-1:0] node2199;
	wire [14-1:0] node2200;
	wire [14-1:0] node2201;
	wire [14-1:0] node2202;
	wire [14-1:0] node2203;
	wire [14-1:0] node2204;
	wire [14-1:0] node2205;
	wire [14-1:0] node2206;
	wire [14-1:0] node2207;
	wire [14-1:0] node2211;
	wire [14-1:0] node2212;
	wire [14-1:0] node2214;
	wire [14-1:0] node2215;
	wire [14-1:0] node2220;
	wire [14-1:0] node2221;
	wire [14-1:0] node2222;
	wire [14-1:0] node2225;
	wire [14-1:0] node2228;
	wire [14-1:0] node2229;
	wire [14-1:0] node2233;
	wire [14-1:0] node2234;
	wire [14-1:0] node2235;
	wire [14-1:0] node2238;
	wire [14-1:0] node2239;
	wire [14-1:0] node2243;
	wire [14-1:0] node2245;
	wire [14-1:0] node2247;
	wire [14-1:0] node2250;
	wire [14-1:0] node2251;
	wire [14-1:0] node2252;
	wire [14-1:0] node2253;
	wire [14-1:0] node2255;
	wire [14-1:0] node2258;
	wire [14-1:0] node2259;
	wire [14-1:0] node2260;
	wire [14-1:0] node2265;
	wire [14-1:0] node2266;
	wire [14-1:0] node2267;
	wire [14-1:0] node2268;
	wire [14-1:0] node2272;
	wire [14-1:0] node2275;
	wire [14-1:0] node2276;
	wire [14-1:0] node2278;
	wire [14-1:0] node2281;
	wire [14-1:0] node2284;
	wire [14-1:0] node2285;
	wire [14-1:0] node2286;
	wire [14-1:0] node2287;
	wire [14-1:0] node2289;
	wire [14-1:0] node2293;
	wire [14-1:0] node2296;
	wire [14-1:0] node2298;
	wire [14-1:0] node2299;
	wire [14-1:0] node2301;
	wire [14-1:0] node2302;
	wire [14-1:0] node2306;
	wire [14-1:0] node2309;
	wire [14-1:0] node2310;
	wire [14-1:0] node2311;
	wire [14-1:0] node2312;
	wire [14-1:0] node2313;
	wire [14-1:0] node2315;
	wire [14-1:0] node2318;
	wire [14-1:0] node2321;
	wire [14-1:0] node2322;
	wire [14-1:0] node2323;
	wire [14-1:0] node2326;
	wire [14-1:0] node2329;
	wire [14-1:0] node2332;
	wire [14-1:0] node2333;
	wire [14-1:0] node2334;
	wire [14-1:0] node2337;
	wire [14-1:0] node2338;
	wire [14-1:0] node2342;
	wire [14-1:0] node2343;
	wire [14-1:0] node2346;
	wire [14-1:0] node2347;
	wire [14-1:0] node2348;
	wire [14-1:0] node2353;
	wire [14-1:0] node2354;
	wire [14-1:0] node2355;
	wire [14-1:0] node2356;
	wire [14-1:0] node2358;
	wire [14-1:0] node2361;
	wire [14-1:0] node2362;
	wire [14-1:0] node2366;
	wire [14-1:0] node2367;
	wire [14-1:0] node2369;
	wire [14-1:0] node2372;
	wire [14-1:0] node2374;
	wire [14-1:0] node2377;
	wire [14-1:0] node2378;
	wire [14-1:0] node2379;
	wire [14-1:0] node2381;
	wire [14-1:0] node2384;
	wire [14-1:0] node2387;
	wire [14-1:0] node2389;
	wire [14-1:0] node2390;
	wire [14-1:0] node2393;
	wire [14-1:0] node2394;
	wire [14-1:0] node2396;
	wire [14-1:0] node2399;
	wire [14-1:0] node2400;
	wire [14-1:0] node2404;
	wire [14-1:0] node2405;
	wire [14-1:0] node2406;
	wire [14-1:0] node2407;
	wire [14-1:0] node2408;
	wire [14-1:0] node2410;
	wire [14-1:0] node2411;
	wire [14-1:0] node2414;
	wire [14-1:0] node2417;
	wire [14-1:0] node2419;
	wire [14-1:0] node2420;
	wire [14-1:0] node2421;
	wire [14-1:0] node2425;
	wire [14-1:0] node2428;
	wire [14-1:0] node2429;
	wire [14-1:0] node2430;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2436;
	wire [14-1:0] node2438;
	wire [14-1:0] node2441;
	wire [14-1:0] node2442;
	wire [14-1:0] node2446;
	wire [14-1:0] node2447;
	wire [14-1:0] node2448;
	wire [14-1:0] node2451;
	wire [14-1:0] node2455;
	wire [14-1:0] node2456;
	wire [14-1:0] node2457;
	wire [14-1:0] node2458;
	wire [14-1:0] node2459;
	wire [14-1:0] node2462;
	wire [14-1:0] node2466;
	wire [14-1:0] node2467;
	wire [14-1:0] node2470;
	wire [14-1:0] node2471;
	wire [14-1:0] node2474;
	wire [14-1:0] node2477;
	wire [14-1:0] node2478;
	wire [14-1:0] node2479;
	wire [14-1:0] node2480;
	wire [14-1:0] node2483;
	wire [14-1:0] node2486;
	wire [14-1:0] node2489;
	wire [14-1:0] node2490;
	wire [14-1:0] node2492;
	wire [14-1:0] node2495;
	wire [14-1:0] node2498;
	wire [14-1:0] node2499;
	wire [14-1:0] node2500;
	wire [14-1:0] node2501;
	wire [14-1:0] node2502;
	wire [14-1:0] node2503;
	wire [14-1:0] node2508;
	wire [14-1:0] node2509;
	wire [14-1:0] node2513;
	wire [14-1:0] node2514;
	wire [14-1:0] node2515;
	wire [14-1:0] node2516;
	wire [14-1:0] node2519;
	wire [14-1:0] node2522;
	wire [14-1:0] node2523;
	wire [14-1:0] node2524;
	wire [14-1:0] node2529;
	wire [14-1:0] node2530;
	wire [14-1:0] node2532;
	wire [14-1:0] node2535;
	wire [14-1:0] node2537;
	wire [14-1:0] node2540;
	wire [14-1:0] node2541;
	wire [14-1:0] node2542;
	wire [14-1:0] node2543;
	wire [14-1:0] node2544;
	wire [14-1:0] node2547;
	wire [14-1:0] node2550;
	wire [14-1:0] node2552;
	wire [14-1:0] node2554;
	wire [14-1:0] node2557;
	wire [14-1:0] node2558;
	wire [14-1:0] node2560;
	wire [14-1:0] node2562;
	wire [14-1:0] node2566;
	wire [14-1:0] node2567;
	wire [14-1:0] node2568;
	wire [14-1:0] node2569;
	wire [14-1:0] node2574;
	wire [14-1:0] node2575;
	wire [14-1:0] node2576;
	wire [14-1:0] node2579;
	wire [14-1:0] node2583;
	wire [14-1:0] node2584;
	wire [14-1:0] node2585;
	wire [14-1:0] node2586;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2590;
	wire [14-1:0] node2591;
	wire [14-1:0] node2592;
	wire [14-1:0] node2593;
	wire [14-1:0] node2597;
	wire [14-1:0] node2601;
	wire [14-1:0] node2602;
	wire [14-1:0] node2604;
	wire [14-1:0] node2607;
	wire [14-1:0] node2609;
	wire [14-1:0] node2612;
	wire [14-1:0] node2613;
	wire [14-1:0] node2614;
	wire [14-1:0] node2616;
	wire [14-1:0] node2617;
	wire [14-1:0] node2622;
	wire [14-1:0] node2624;
	wire [14-1:0] node2627;
	wire [14-1:0] node2628;
	wire [14-1:0] node2629;
	wire [14-1:0] node2630;
	wire [14-1:0] node2633;
	wire [14-1:0] node2634;
	wire [14-1:0] node2637;
	wire [14-1:0] node2639;
	wire [14-1:0] node2642;
	wire [14-1:0] node2643;
	wire [14-1:0] node2645;
	wire [14-1:0] node2647;
	wire [14-1:0] node2650;
	wire [14-1:0] node2651;
	wire [14-1:0] node2655;
	wire [14-1:0] node2656;
	wire [14-1:0] node2657;
	wire [14-1:0] node2661;
	wire [14-1:0] node2663;
	wire [14-1:0] node2665;
	wire [14-1:0] node2668;
	wire [14-1:0] node2669;
	wire [14-1:0] node2670;
	wire [14-1:0] node2671;
	wire [14-1:0] node2672;
	wire [14-1:0] node2673;
	wire [14-1:0] node2676;
	wire [14-1:0] node2679;
	wire [14-1:0] node2680;
	wire [14-1:0] node2683;
	wire [14-1:0] node2686;
	wire [14-1:0] node2687;
	wire [14-1:0] node2689;
	wire [14-1:0] node2691;
	wire [14-1:0] node2694;
	wire [14-1:0] node2695;
	wire [14-1:0] node2696;
	wire [14-1:0] node2701;
	wire [14-1:0] node2702;
	wire [14-1:0] node2703;
	wire [14-1:0] node2706;
	wire [14-1:0] node2707;
	wire [14-1:0] node2709;
	wire [14-1:0] node2712;
	wire [14-1:0] node2713;
	wire [14-1:0] node2714;
	wire [14-1:0] node2719;
	wire [14-1:0] node2720;
	wire [14-1:0] node2722;
	wire [14-1:0] node2725;
	wire [14-1:0] node2728;
	wire [14-1:0] node2729;
	wire [14-1:0] node2730;
	wire [14-1:0] node2732;
	wire [14-1:0] node2733;
	wire [14-1:0] node2734;
	wire [14-1:0] node2739;
	wire [14-1:0] node2740;
	wire [14-1:0] node2744;
	wire [14-1:0] node2745;
	wire [14-1:0] node2746;
	wire [14-1:0] node2747;
	wire [14-1:0] node2748;
	wire [14-1:0] node2752;
	wire [14-1:0] node2755;
	wire [14-1:0] node2756;
	wire [14-1:0] node2759;
	wire [14-1:0] node2762;
	wire [14-1:0] node2763;
	wire [14-1:0] node2766;
	wire [14-1:0] node2767;
	wire [14-1:0] node2771;
	wire [14-1:0] node2772;
	wire [14-1:0] node2773;
	wire [14-1:0] node2774;
	wire [14-1:0] node2775;
	wire [14-1:0] node2776;
	wire [14-1:0] node2778;
	wire [14-1:0] node2781;
	wire [14-1:0] node2782;
	wire [14-1:0] node2785;
	wire [14-1:0] node2788;
	wire [14-1:0] node2789;
	wire [14-1:0] node2791;
	wire [14-1:0] node2795;
	wire [14-1:0] node2796;
	wire [14-1:0] node2798;
	wire [14-1:0] node2800;
	wire [14-1:0] node2802;
	wire [14-1:0] node2805;
	wire [14-1:0] node2806;
	wire [14-1:0] node2809;
	wire [14-1:0] node2812;
	wire [14-1:0] node2813;
	wire [14-1:0] node2814;
	wire [14-1:0] node2815;
	wire [14-1:0] node2818;
	wire [14-1:0] node2821;
	wire [14-1:0] node2822;
	wire [14-1:0] node2823;
	wire [14-1:0] node2826;
	wire [14-1:0] node2828;
	wire [14-1:0] node2829;
	wire [14-1:0] node2833;
	wire [14-1:0] node2834;
	wire [14-1:0] node2836;
	wire [14-1:0] node2838;
	wire [14-1:0] node2842;
	wire [14-1:0] node2843;
	wire [14-1:0] node2844;
	wire [14-1:0] node2847;
	wire [14-1:0] node2848;
	wire [14-1:0] node2852;
	wire [14-1:0] node2853;
	wire [14-1:0] node2857;
	wire [14-1:0] node2858;
	wire [14-1:0] node2859;
	wire [14-1:0] node2860;
	wire [14-1:0] node2861;
	wire [14-1:0] node2863;
	wire [14-1:0] node2866;
	wire [14-1:0] node2867;
	wire [14-1:0] node2868;
	wire [14-1:0] node2870;
	wire [14-1:0] node2875;
	wire [14-1:0] node2876;
	wire [14-1:0] node2877;
	wire [14-1:0] node2879;
	wire [14-1:0] node2880;
	wire [14-1:0] node2885;
	wire [14-1:0] node2887;
	wire [14-1:0] node2889;
	wire [14-1:0] node2892;
	wire [14-1:0] node2893;
	wire [14-1:0] node2894;
	wire [14-1:0] node2896;
	wire [14-1:0] node2899;
	wire [14-1:0] node2900;
	wire [14-1:0] node2903;
	wire [14-1:0] node2906;
	wire [14-1:0] node2907;
	wire [14-1:0] node2909;
	wire [14-1:0] node2910;
	wire [14-1:0] node2914;
	wire [14-1:0] node2915;
	wire [14-1:0] node2916;
	wire [14-1:0] node2920;
	wire [14-1:0] node2923;
	wire [14-1:0] node2924;
	wire [14-1:0] node2925;
	wire [14-1:0] node2926;
	wire [14-1:0] node2927;
	wire [14-1:0] node2930;
	wire [14-1:0] node2931;
	wire [14-1:0] node2935;
	wire [14-1:0] node2936;
	wire [14-1:0] node2940;
	wire [14-1:0] node2941;
	wire [14-1:0] node2942;
	wire [14-1:0] node2945;
	wire [14-1:0] node2946;
	wire [14-1:0] node2950;
	wire [14-1:0] node2952;
	wire [14-1:0] node2955;
	wire [14-1:0] node2956;
	wire [14-1:0] node2957;
	wire [14-1:0] node2959;
	wire [14-1:0] node2962;
	wire [14-1:0] node2963;
	wire [14-1:0] node2967;
	wire [14-1:0] node2968;
	wire [14-1:0] node2969;
	wire [14-1:0] node2972;
	wire [14-1:0] node2974;
	wire [14-1:0] node2977;
	wire [14-1:0] node2978;
	wire [14-1:0] node2980;
	wire [14-1:0] node2984;
	wire [14-1:0] node2985;
	wire [14-1:0] node2986;
	wire [14-1:0] node2987;
	wire [14-1:0] node2988;
	wire [14-1:0] node2989;
	wire [14-1:0] node2990;
	wire [14-1:0] node2991;
	wire [14-1:0] node2992;
	wire [14-1:0] node2993;
	wire [14-1:0] node2994;
	wire [14-1:0] node2998;
	wire [14-1:0] node3000;
	wire [14-1:0] node3001;
	wire [14-1:0] node3005;
	wire [14-1:0] node3006;
	wire [14-1:0] node3008;
	wire [14-1:0] node3011;
	wire [14-1:0] node3012;
	wire [14-1:0] node3016;
	wire [14-1:0] node3017;
	wire [14-1:0] node3018;
	wire [14-1:0] node3019;
	wire [14-1:0] node3022;
	wire [14-1:0] node3023;
	wire [14-1:0] node3027;
	wire [14-1:0] node3028;
	wire [14-1:0] node3032;
	wire [14-1:0] node3033;
	wire [14-1:0] node3034;
	wire [14-1:0] node3037;
	wire [14-1:0] node3040;
	wire [14-1:0] node3042;
	wire [14-1:0] node3043;
	wire [14-1:0] node3045;
	wire [14-1:0] node3049;
	wire [14-1:0] node3050;
	wire [14-1:0] node3051;
	wire [14-1:0] node3052;
	wire [14-1:0] node3055;
	wire [14-1:0] node3056;
	wire [14-1:0] node3059;
	wire [14-1:0] node3060;
	wire [14-1:0] node3064;
	wire [14-1:0] node3067;
	wire [14-1:0] node3068;
	wire [14-1:0] node3069;
	wire [14-1:0] node3070;
	wire [14-1:0] node3074;
	wire [14-1:0] node3075;
	wire [14-1:0] node3076;
	wire [14-1:0] node3081;
	wire [14-1:0] node3082;
	wire [14-1:0] node3083;
	wire [14-1:0] node3084;
	wire [14-1:0] node3088;
	wire [14-1:0] node3091;
	wire [14-1:0] node3092;
	wire [14-1:0] node3095;
	wire [14-1:0] node3098;
	wire [14-1:0] node3099;
	wire [14-1:0] node3100;
	wire [14-1:0] node3101;
	wire [14-1:0] node3102;
	wire [14-1:0] node3104;
	wire [14-1:0] node3107;
	wire [14-1:0] node3110;
	wire [14-1:0] node3111;
	wire [14-1:0] node3112;
	wire [14-1:0] node3116;
	wire [14-1:0] node3118;
	wire [14-1:0] node3121;
	wire [14-1:0] node3122;
	wire [14-1:0] node3123;
	wire [14-1:0] node3124;
	wire [14-1:0] node3128;
	wire [14-1:0] node3129;
	wire [14-1:0] node3133;
	wire [14-1:0] node3134;
	wire [14-1:0] node3135;
	wire [14-1:0] node3136;
	wire [14-1:0] node3140;
	wire [14-1:0] node3143;
	wire [14-1:0] node3146;
	wire [14-1:0] node3147;
	wire [14-1:0] node3148;
	wire [14-1:0] node3149;
	wire [14-1:0] node3150;
	wire [14-1:0] node3151;
	wire [14-1:0] node3156;
	wire [14-1:0] node3158;
	wire [14-1:0] node3160;
	wire [14-1:0] node3161;
	wire [14-1:0] node3165;
	wire [14-1:0] node3166;
	wire [14-1:0] node3168;
	wire [14-1:0] node3170;
	wire [14-1:0] node3173;
	wire [14-1:0] node3174;
	wire [14-1:0] node3178;
	wire [14-1:0] node3179;
	wire [14-1:0] node3182;
	wire [14-1:0] node3184;
	wire [14-1:0] node3185;
	wire [14-1:0] node3189;
	wire [14-1:0] node3190;
	wire [14-1:0] node3191;
	wire [14-1:0] node3192;
	wire [14-1:0] node3193;
	wire [14-1:0] node3195;
	wire [14-1:0] node3196;
	wire [14-1:0] node3198;
	wire [14-1:0] node3199;
	wire [14-1:0] node3203;
	wire [14-1:0] node3206;
	wire [14-1:0] node3207;
	wire [14-1:0] node3208;
	wire [14-1:0] node3209;
	wire [14-1:0] node3214;
	wire [14-1:0] node3215;
	wire [14-1:0] node3219;
	wire [14-1:0] node3220;
	wire [14-1:0] node3221;
	wire [14-1:0] node3222;
	wire [14-1:0] node3223;
	wire [14-1:0] node3225;
	wire [14-1:0] node3229;
	wire [14-1:0] node3232;
	wire [14-1:0] node3233;
	wire [14-1:0] node3234;
	wire [14-1:0] node3238;
	wire [14-1:0] node3241;
	wire [14-1:0] node3242;
	wire [14-1:0] node3244;
	wire [14-1:0] node3245;
	wire [14-1:0] node3247;
	wire [14-1:0] node3250;
	wire [14-1:0] node3252;
	wire [14-1:0] node3256;
	wire [14-1:0] node3257;
	wire [14-1:0] node3258;
	wire [14-1:0] node3259;
	wire [14-1:0] node3260;
	wire [14-1:0] node3263;
	wire [14-1:0] node3266;
	wire [14-1:0] node3267;
	wire [14-1:0] node3270;
	wire [14-1:0] node3273;
	wire [14-1:0] node3274;
	wire [14-1:0] node3275;
	wire [14-1:0] node3278;
	wire [14-1:0] node3281;
	wire [14-1:0] node3282;
	wire [14-1:0] node3285;
	wire [14-1:0] node3288;
	wire [14-1:0] node3289;
	wire [14-1:0] node3290;
	wire [14-1:0] node3291;
	wire [14-1:0] node3295;
	wire [14-1:0] node3296;
	wire [14-1:0] node3297;
	wire [14-1:0] node3299;
	wire [14-1:0] node3302;
	wire [14-1:0] node3306;
	wire [14-1:0] node3307;
	wire [14-1:0] node3309;
	wire [14-1:0] node3312;
	wire [14-1:0] node3315;
	wire [14-1:0] node3316;
	wire [14-1:0] node3317;
	wire [14-1:0] node3319;
	wire [14-1:0] node3320;
	wire [14-1:0] node3323;
	wire [14-1:0] node3324;
	wire [14-1:0] node3326;
	wire [14-1:0] node3330;
	wire [14-1:0] node3331;
	wire [14-1:0] node3332;
	wire [14-1:0] node3334;
	wire [14-1:0] node3335;
	wire [14-1:0] node3337;
	wire [14-1:0] node3341;
	wire [14-1:0] node3342;
	wire [14-1:0] node3346;
	wire [14-1:0] node3349;
	wire [14-1:0] node3350;
	wire [14-1:0] node3351;
	wire [14-1:0] node3352;
	wire [14-1:0] node3353;
	wire [14-1:0] node3354;
	wire [14-1:0] node3356;
	wire [14-1:0] node3361;
	wire [14-1:0] node3362;
	wire [14-1:0] node3366;
	wire [14-1:0] node3367;
	wire [14-1:0] node3368;
	wire [14-1:0] node3369;
	wire [14-1:0] node3371;
	wire [14-1:0] node3375;
	wire [14-1:0] node3378;
	wire [14-1:0] node3381;
	wire [14-1:0] node3382;
	wire [14-1:0] node3383;
	wire [14-1:0] node3386;
	wire [14-1:0] node3388;
	wire [14-1:0] node3390;
	wire [14-1:0] node3393;
	wire [14-1:0] node3394;
	wire [14-1:0] node3397;
	wire [14-1:0] node3398;
	wire [14-1:0] node3401;
	wire [14-1:0] node3402;
	wire [14-1:0] node3406;
	wire [14-1:0] node3407;
	wire [14-1:0] node3408;
	wire [14-1:0] node3409;
	wire [14-1:0] node3410;
	wire [14-1:0] node3411;
	wire [14-1:0] node3412;
	wire [14-1:0] node3413;
	wire [14-1:0] node3417;
	wire [14-1:0] node3418;
	wire [14-1:0] node3419;
	wire [14-1:0] node3423;
	wire [14-1:0] node3424;
	wire [14-1:0] node3428;
	wire [14-1:0] node3429;
	wire [14-1:0] node3432;
	wire [14-1:0] node3434;
	wire [14-1:0] node3437;
	wire [14-1:0] node3438;
	wire [14-1:0] node3439;
	wire [14-1:0] node3441;
	wire [14-1:0] node3444;
	wire [14-1:0] node3446;
	wire [14-1:0] node3449;
	wire [14-1:0] node3451;
	wire [14-1:0] node3452;
	wire [14-1:0] node3456;
	wire [14-1:0] node3457;
	wire [14-1:0] node3458;
	wire [14-1:0] node3459;
	wire [14-1:0] node3460;
	wire [14-1:0] node3462;
	wire [14-1:0] node3466;
	wire [14-1:0] node3469;
	wire [14-1:0] node3470;
	wire [14-1:0] node3472;
	wire [14-1:0] node3475;
	wire [14-1:0] node3478;
	wire [14-1:0] node3479;
	wire [14-1:0] node3480;
	wire [14-1:0] node3483;
	wire [14-1:0] node3485;
	wire [14-1:0] node3487;
	wire [14-1:0] node3488;
	wire [14-1:0] node3492;
	wire [14-1:0] node3494;
	wire [14-1:0] node3495;
	wire [14-1:0] node3496;
	wire [14-1:0] node3498;
	wire [14-1:0] node3503;
	wire [14-1:0] node3504;
	wire [14-1:0] node3505;
	wire [14-1:0] node3506;
	wire [14-1:0] node3508;
	wire [14-1:0] node3509;
	wire [14-1:0] node3511;
	wire [14-1:0] node3514;
	wire [14-1:0] node3517;
	wire [14-1:0] node3518;
	wire [14-1:0] node3519;
	wire [14-1:0] node3522;
	wire [14-1:0] node3526;
	wire [14-1:0] node3527;
	wire [14-1:0] node3529;
	wire [14-1:0] node3530;
	wire [14-1:0] node3534;
	wire [14-1:0] node3535;
	wire [14-1:0] node3537;
	wire [14-1:0] node3540;
	wire [14-1:0] node3542;
	wire [14-1:0] node3545;
	wire [14-1:0] node3546;
	wire [14-1:0] node3547;
	wire [14-1:0] node3548;
	wire [14-1:0] node3552;
	wire [14-1:0] node3553;
	wire [14-1:0] node3554;
	wire [14-1:0] node3558;
	wire [14-1:0] node3559;
	wire [14-1:0] node3562;
	wire [14-1:0] node3564;
	wire [14-1:0] node3567;
	wire [14-1:0] node3568;
	wire [14-1:0] node3569;
	wire [14-1:0] node3571;
	wire [14-1:0] node3574;
	wire [14-1:0] node3577;
	wire [14-1:0] node3579;
	wire [14-1:0] node3582;
	wire [14-1:0] node3583;
	wire [14-1:0] node3584;
	wire [14-1:0] node3585;
	wire [14-1:0] node3586;
	wire [14-1:0] node3587;
	wire [14-1:0] node3589;
	wire [14-1:0] node3590;
	wire [14-1:0] node3591;
	wire [14-1:0] node3596;
	wire [14-1:0] node3598;
	wire [14-1:0] node3600;
	wire [14-1:0] node3601;
	wire [14-1:0] node3605;
	wire [14-1:0] node3606;
	wire [14-1:0] node3607;
	wire [14-1:0] node3611;
	wire [14-1:0] node3613;
	wire [14-1:0] node3616;
	wire [14-1:0] node3617;
	wire [14-1:0] node3618;
	wire [14-1:0] node3619;
	wire [14-1:0] node3622;
	wire [14-1:0] node3624;
	wire [14-1:0] node3625;
	wire [14-1:0] node3629;
	wire [14-1:0] node3631;
	wire [14-1:0] node3634;
	wire [14-1:0] node3635;
	wire [14-1:0] node3636;
	wire [14-1:0] node3639;
	wire [14-1:0] node3641;
	wire [14-1:0] node3644;
	wire [14-1:0] node3645;
	wire [14-1:0] node3648;
	wire [14-1:0] node3651;
	wire [14-1:0] node3652;
	wire [14-1:0] node3653;
	wire [14-1:0] node3654;
	wire [14-1:0] node3655;
	wire [14-1:0] node3657;
	wire [14-1:0] node3661;
	wire [14-1:0] node3663;
	wire [14-1:0] node3665;
	wire [14-1:0] node3668;
	wire [14-1:0] node3669;
	wire [14-1:0] node3672;
	wire [14-1:0] node3674;
	wire [14-1:0] node3677;
	wire [14-1:0] node3678;
	wire [14-1:0] node3680;
	wire [14-1:0] node3681;
	wire [14-1:0] node3685;
	wire [14-1:0] node3686;
	wire [14-1:0] node3687;
	wire [14-1:0] node3688;
	wire [14-1:0] node3692;
	wire [14-1:0] node3695;
	wire [14-1:0] node3697;
	wire [14-1:0] node3700;
	wire [14-1:0] node3701;
	wire [14-1:0] node3702;
	wire [14-1:0] node3703;
	wire [14-1:0] node3704;
	wire [14-1:0] node3706;
	wire [14-1:0] node3708;
	wire [14-1:0] node3711;
	wire [14-1:0] node3714;
	wire [14-1:0] node3715;
	wire [14-1:0] node3718;
	wire [14-1:0] node3720;
	wire [14-1:0] node3723;
	wire [14-1:0] node3724;
	wire [14-1:0] node3725;
	wire [14-1:0] node3726;
	wire [14-1:0] node3731;
	wire [14-1:0] node3732;
	wire [14-1:0] node3733;
	wire [14-1:0] node3737;
	wire [14-1:0] node3738;
	wire [14-1:0] node3739;
	wire [14-1:0] node3743;
	wire [14-1:0] node3744;
	wire [14-1:0] node3748;
	wire [14-1:0] node3749;
	wire [14-1:0] node3750;
	wire [14-1:0] node3751;
	wire [14-1:0] node3752;
	wire [14-1:0] node3755;
	wire [14-1:0] node3757;
	wire [14-1:0] node3758;
	wire [14-1:0] node3762;
	wire [14-1:0] node3763;
	wire [14-1:0] node3766;
	wire [14-1:0] node3767;
	wire [14-1:0] node3771;
	wire [14-1:0] node3772;
	wire [14-1:0] node3774;
	wire [14-1:0] node3775;
	wire [14-1:0] node3777;
	wire [14-1:0] node3781;
	wire [14-1:0] node3782;
	wire [14-1:0] node3786;
	wire [14-1:0] node3787;
	wire [14-1:0] node3789;
	wire [14-1:0] node3791;
	wire [14-1:0] node3793;
	wire [14-1:0] node3796;
	wire [14-1:0] node3797;
	wire [14-1:0] node3798;
	wire [14-1:0] node3802;
	wire [14-1:0] node3804;
	wire [14-1:0] node3807;
	wire [14-1:0] node3808;
	wire [14-1:0] node3809;
	wire [14-1:0] node3810;
	wire [14-1:0] node3811;
	wire [14-1:0] node3812;
	wire [14-1:0] node3813;
	wire [14-1:0] node3815;
	wire [14-1:0] node3816;
	wire [14-1:0] node3820;
	wire [14-1:0] node3821;
	wire [14-1:0] node3824;
	wire [14-1:0] node3825;
	wire [14-1:0] node3827;
	wire [14-1:0] node3830;
	wire [14-1:0] node3833;
	wire [14-1:0] node3834;
	wire [14-1:0] node3835;
	wire [14-1:0] node3839;
	wire [14-1:0] node3840;
	wire [14-1:0] node3841;
	wire [14-1:0] node3845;
	wire [14-1:0] node3846;
	wire [14-1:0] node3850;
	wire [14-1:0] node3851;
	wire [14-1:0] node3852;
	wire [14-1:0] node3854;
	wire [14-1:0] node3855;
	wire [14-1:0] node3856;
	wire [14-1:0] node3861;
	wire [14-1:0] node3863;
	wire [14-1:0] node3864;
	wire [14-1:0] node3865;
	wire [14-1:0] node3869;
	wire [14-1:0] node3871;
	wire [14-1:0] node3874;
	wire [14-1:0] node3875;
	wire [14-1:0] node3876;
	wire [14-1:0] node3878;
	wire [14-1:0] node3881;
	wire [14-1:0] node3883;
	wire [14-1:0] node3886;
	wire [14-1:0] node3887;
	wire [14-1:0] node3888;
	wire [14-1:0] node3889;
	wire [14-1:0] node3893;
	wire [14-1:0] node3895;
	wire [14-1:0] node3898;
	wire [14-1:0] node3899;
	wire [14-1:0] node3903;
	wire [14-1:0] node3904;
	wire [14-1:0] node3905;
	wire [14-1:0] node3906;
	wire [14-1:0] node3907;
	wire [14-1:0] node3908;
	wire [14-1:0] node3911;
	wire [14-1:0] node3913;
	wire [14-1:0] node3916;
	wire [14-1:0] node3917;
	wire [14-1:0] node3920;
	wire [14-1:0] node3922;
	wire [14-1:0] node3923;
	wire [14-1:0] node3927;
	wire [14-1:0] node3928;
	wire [14-1:0] node3930;
	wire [14-1:0] node3933;
	wire [14-1:0] node3934;
	wire [14-1:0] node3938;
	wire [14-1:0] node3939;
	wire [14-1:0] node3942;
	wire [14-1:0] node3944;
	wire [14-1:0] node3945;
	wire [14-1:0] node3949;
	wire [14-1:0] node3950;
	wire [14-1:0] node3951;
	wire [14-1:0] node3952;
	wire [14-1:0] node3954;
	wire [14-1:0] node3957;
	wire [14-1:0] node3958;
	wire [14-1:0] node3961;
	wire [14-1:0] node3964;
	wire [14-1:0] node3966;
	wire [14-1:0] node3968;
	wire [14-1:0] node3971;
	wire [14-1:0] node3972;
	wire [14-1:0] node3973;
	wire [14-1:0] node3975;
	wire [14-1:0] node3976;
	wire [14-1:0] node3977;
	wire [14-1:0] node3982;
	wire [14-1:0] node3983;
	wire [14-1:0] node3984;
	wire [14-1:0] node3988;
	wire [14-1:0] node3990;
	wire [14-1:0] node3992;
	wire [14-1:0] node3995;
	wire [14-1:0] node3996;
	wire [14-1:0] node3998;
	wire [14-1:0] node3999;
	wire [14-1:0] node4001;
	wire [14-1:0] node4005;
	wire [14-1:0] node4006;
	wire [14-1:0] node4007;
	wire [14-1:0] node4011;
	wire [14-1:0] node4014;
	wire [14-1:0] node4015;
	wire [14-1:0] node4016;
	wire [14-1:0] node4017;
	wire [14-1:0] node4018;
	wire [14-1:0] node4019;
	wire [14-1:0] node4020;
	wire [14-1:0] node4024;
	wire [14-1:0] node4025;
	wire [14-1:0] node4029;
	wire [14-1:0] node4030;
	wire [14-1:0] node4031;
	wire [14-1:0] node4032;
	wire [14-1:0] node4034;
	wire [14-1:0] node4037;
	wire [14-1:0] node4042;
	wire [14-1:0] node4043;
	wire [14-1:0] node4045;
	wire [14-1:0] node4046;
	wire [14-1:0] node4050;
	wire [14-1:0] node4051;
	wire [14-1:0] node4054;
	wire [14-1:0] node4057;
	wire [14-1:0] node4058;
	wire [14-1:0] node4059;
	wire [14-1:0] node4060;
	wire [14-1:0] node4061;
	wire [14-1:0] node4066;
	wire [14-1:0] node4067;
	wire [14-1:0] node4070;
	wire [14-1:0] node4072;
	wire [14-1:0] node4075;
	wire [14-1:0] node4076;
	wire [14-1:0] node4077;
	wire [14-1:0] node4079;
	wire [14-1:0] node4081;
	wire [14-1:0] node4082;
	wire [14-1:0] node4086;
	wire [14-1:0] node4088;
	wire [14-1:0] node4091;
	wire [14-1:0] node4092;
	wire [14-1:0] node4093;
	wire [14-1:0] node4096;
	wire [14-1:0] node4097;
	wire [14-1:0] node4101;
	wire [14-1:0] node4104;
	wire [14-1:0] node4105;
	wire [14-1:0] node4106;
	wire [14-1:0] node4107;
	wire [14-1:0] node4109;
	wire [14-1:0] node4110;
	wire [14-1:0] node4112;
	wire [14-1:0] node4113;
	wire [14-1:0] node4118;
	wire [14-1:0] node4119;
	wire [14-1:0] node4121;
	wire [14-1:0] node4125;
	wire [14-1:0] node4126;
	wire [14-1:0] node4127;
	wire [14-1:0] node4129;
	wire [14-1:0] node4132;
	wire [14-1:0] node4135;
	wire [14-1:0] node4136;
	wire [14-1:0] node4138;
	wire [14-1:0] node4141;
	wire [14-1:0] node4144;
	wire [14-1:0] node4145;
	wire [14-1:0] node4146;
	wire [14-1:0] node4147;
	wire [14-1:0] node4149;
	wire [14-1:0] node4151;
	wire [14-1:0] node4152;
	wire [14-1:0] node4156;
	wire [14-1:0] node4157;
	wire [14-1:0] node4158;
	wire [14-1:0] node4162;
	wire [14-1:0] node4165;
	wire [14-1:0] node4166;
	wire [14-1:0] node4169;
	wire [14-1:0] node4170;
	wire [14-1:0] node4173;
	wire [14-1:0] node4175;
	wire [14-1:0] node4178;
	wire [14-1:0] node4179;
	wire [14-1:0] node4180;
	wire [14-1:0] node4181;
	wire [14-1:0] node4185;
	wire [14-1:0] node4187;
	wire [14-1:0] node4190;
	wire [14-1:0] node4192;
	wire [14-1:0] node4194;
	wire [14-1:0] node4197;
	wire [14-1:0] node4198;
	wire [14-1:0] node4199;
	wire [14-1:0] node4200;
	wire [14-1:0] node4201;
	wire [14-1:0] node4202;
	wire [14-1:0] node4203;
	wire [14-1:0] node4204;
	wire [14-1:0] node4206;
	wire [14-1:0] node4211;
	wire [14-1:0] node4212;
	wire [14-1:0] node4213;
	wire [14-1:0] node4215;
	wire [14-1:0] node4219;
	wire [14-1:0] node4220;
	wire [14-1:0] node4222;
	wire [14-1:0] node4223;
	wire [14-1:0] node4228;
	wire [14-1:0] node4229;
	wire [14-1:0] node4231;
	wire [14-1:0] node4234;
	wire [14-1:0] node4236;
	wire [14-1:0] node4238;
	wire [14-1:0] node4241;
	wire [14-1:0] node4242;
	wire [14-1:0] node4243;
	wire [14-1:0] node4244;
	wire [14-1:0] node4246;
	wire [14-1:0] node4250;
	wire [14-1:0] node4252;
	wire [14-1:0] node4253;
	wire [14-1:0] node4257;
	wire [14-1:0] node4258;
	wire [14-1:0] node4259;
	wire [14-1:0] node4260;
	wire [14-1:0] node4264;
	wire [14-1:0] node4265;
	wire [14-1:0] node4267;
	wire [14-1:0] node4268;
	wire [14-1:0] node4272;
	wire [14-1:0] node4275;
	wire [14-1:0] node4276;
	wire [14-1:0] node4277;
	wire [14-1:0] node4278;
	wire [14-1:0] node4283;
	wire [14-1:0] node4284;
	wire [14-1:0] node4287;
	wire [14-1:0] node4290;
	wire [14-1:0] node4291;
	wire [14-1:0] node4292;
	wire [14-1:0] node4293;
	wire [14-1:0] node4296;
	wire [14-1:0] node4297;
	wire [14-1:0] node4298;
	wire [14-1:0] node4302;
	wire [14-1:0] node4303;
	wire [14-1:0] node4307;
	wire [14-1:0] node4308;
	wire [14-1:0] node4309;
	wire [14-1:0] node4311;
	wire [14-1:0] node4315;
	wire [14-1:0] node4316;
	wire [14-1:0] node4317;
	wire [14-1:0] node4321;
	wire [14-1:0] node4322;
	wire [14-1:0] node4325;
	wire [14-1:0] node4326;
	wire [14-1:0] node4330;
	wire [14-1:0] node4331;
	wire [14-1:0] node4332;
	wire [14-1:0] node4333;
	wire [14-1:0] node4336;
	wire [14-1:0] node4338;
	wire [14-1:0] node4340;
	wire [14-1:0] node4343;
	wire [14-1:0] node4344;
	wire [14-1:0] node4345;
	wire [14-1:0] node4349;
	wire [14-1:0] node4350;
	wire [14-1:0] node4353;
	wire [14-1:0] node4354;
	wire [14-1:0] node4358;
	wire [14-1:0] node4359;
	wire [14-1:0] node4360;
	wire [14-1:0] node4362;
	wire [14-1:0] node4363;
	wire [14-1:0] node4366;
	wire [14-1:0] node4370;
	wire [14-1:0] node4371;
	wire [14-1:0] node4374;
	wire [14-1:0] node4376;
	wire [14-1:0] node4377;
	wire [14-1:0] node4381;
	wire [14-1:0] node4382;
	wire [14-1:0] node4383;
	wire [14-1:0] node4384;
	wire [14-1:0] node4385;
	wire [14-1:0] node4386;
	wire [14-1:0] node4387;
	wire [14-1:0] node4391;
	wire [14-1:0] node4393;
	wire [14-1:0] node4396;
	wire [14-1:0] node4397;
	wire [14-1:0] node4399;
	wire [14-1:0] node4403;
	wire [14-1:0] node4404;
	wire [14-1:0] node4405;
	wire [14-1:0] node4406;
	wire [14-1:0] node4409;
	wire [14-1:0] node4412;
	wire [14-1:0] node4413;
	wire [14-1:0] node4414;
	wire [14-1:0] node4418;
	wire [14-1:0] node4421;
	wire [14-1:0] node4422;
	wire [14-1:0] node4423;
	wire [14-1:0] node4427;
	wire [14-1:0] node4428;
	wire [14-1:0] node4431;
	wire [14-1:0] node4432;
	wire [14-1:0] node4436;
	wire [14-1:0] node4437;
	wire [14-1:0] node4438;
	wire [14-1:0] node4439;
	wire [14-1:0] node4440;
	wire [14-1:0] node4443;
	wire [14-1:0] node4446;
	wire [14-1:0] node4447;
	wire [14-1:0] node4451;
	wire [14-1:0] node4453;
	wire [14-1:0] node4455;
	wire [14-1:0] node4458;
	wire [14-1:0] node4459;
	wire [14-1:0] node4460;
	wire [14-1:0] node4464;
	wire [14-1:0] node4465;
	wire [14-1:0] node4466;
	wire [14-1:0] node4467;
	wire [14-1:0] node4471;
	wire [14-1:0] node4472;
	wire [14-1:0] node4476;
	wire [14-1:0] node4479;
	wire [14-1:0] node4480;
	wire [14-1:0] node4481;
	wire [14-1:0] node4482;
	wire [14-1:0] node4485;
	wire [14-1:0] node4486;
	wire [14-1:0] node4488;
	wire [14-1:0] node4490;
	wire [14-1:0] node4493;
	wire [14-1:0] node4494;
	wire [14-1:0] node4498;
	wire [14-1:0] node4499;
	wire [14-1:0] node4501;
	wire [14-1:0] node4502;
	wire [14-1:0] node4505;
	wire [14-1:0] node4507;
	wire [14-1:0] node4510;
	wire [14-1:0] node4511;
	wire [14-1:0] node4514;
	wire [14-1:0] node4515;
	wire [14-1:0] node4516;
	wire [14-1:0] node4518;
	wire [14-1:0] node4522;
	wire [14-1:0] node4525;
	wire [14-1:0] node4526;
	wire [14-1:0] node4527;
	wire [14-1:0] node4528;
	wire [14-1:0] node4531;
	wire [14-1:0] node4534;
	wire [14-1:0] node4535;
	wire [14-1:0] node4536;
	wire [14-1:0] node4539;
	wire [14-1:0] node4542;
	wire [14-1:0] node4543;
	wire [14-1:0] node4546;
	wire [14-1:0] node4548;
	wire [14-1:0] node4551;
	wire [14-1:0] node4552;
	wire [14-1:0] node4553;
	wire [14-1:0] node4556;
	wire [14-1:0] node4558;
	wire [14-1:0] node4561;
	wire [14-1:0] node4562;
	wire [14-1:0] node4564;
	wire [14-1:0] node4565;
	wire [14-1:0] node4569;
	wire [14-1:0] node4571;
	wire [14-1:0] node4573;
	wire [14-1:0] node4576;
	wire [14-1:0] node4577;
	wire [14-1:0] node4578;
	wire [14-1:0] node4579;
	wire [14-1:0] node4580;
	wire [14-1:0] node4581;
	wire [14-1:0] node4582;
	wire [14-1:0] node4583;
	wire [14-1:0] node4584;
	wire [14-1:0] node4586;
	wire [14-1:0] node4590;
	wire [14-1:0] node4591;
	wire [14-1:0] node4592;
	wire [14-1:0] node4593;
	wire [14-1:0] node4597;
	wire [14-1:0] node4600;
	wire [14-1:0] node4603;
	wire [14-1:0] node4604;
	wire [14-1:0] node4605;
	wire [14-1:0] node4607;
	wire [14-1:0] node4609;
	wire [14-1:0] node4612;
	wire [14-1:0] node4613;
	wire [14-1:0] node4616;
	wire [14-1:0] node4619;
	wire [14-1:0] node4620;
	wire [14-1:0] node4622;
	wire [14-1:0] node4625;
	wire [14-1:0] node4626;
	wire [14-1:0] node4630;
	wire [14-1:0] node4631;
	wire [14-1:0] node4632;
	wire [14-1:0] node4633;
	wire [14-1:0] node4636;
	wire [14-1:0] node4637;
	wire [14-1:0] node4641;
	wire [14-1:0] node4642;
	wire [14-1:0] node4643;
	wire [14-1:0] node4647;
	wire [14-1:0] node4648;
	wire [14-1:0] node4649;
	wire [14-1:0] node4650;
	wire [14-1:0] node4655;
	wire [14-1:0] node4657;
	wire [14-1:0] node4660;
	wire [14-1:0] node4661;
	wire [14-1:0] node4663;
	wire [14-1:0] node4664;
	wire [14-1:0] node4667;
	wire [14-1:0] node4670;
	wire [14-1:0] node4671;
	wire [14-1:0] node4672;
	wire [14-1:0] node4675;
	wire [14-1:0] node4679;
	wire [14-1:0] node4680;
	wire [14-1:0] node4681;
	wire [14-1:0] node4682;
	wire [14-1:0] node4683;
	wire [14-1:0] node4686;
	wire [14-1:0] node4689;
	wire [14-1:0] node4690;
	wire [14-1:0] node4692;
	wire [14-1:0] node4695;
	wire [14-1:0] node4696;
	wire [14-1:0] node4700;
	wire [14-1:0] node4701;
	wire [14-1:0] node4702;
	wire [14-1:0] node4704;
	wire [14-1:0] node4708;
	wire [14-1:0] node4710;
	wire [14-1:0] node4711;
	wire [14-1:0] node4714;
	wire [14-1:0] node4717;
	wire [14-1:0] node4718;
	wire [14-1:0] node4719;
	wire [14-1:0] node4720;
	wire [14-1:0] node4724;
	wire [14-1:0] node4726;
	wire [14-1:0] node4729;
	wire [14-1:0] node4730;
	wire [14-1:0] node4732;
	wire [14-1:0] node4735;
	wire [14-1:0] node4736;
	wire [14-1:0] node4738;
	wire [14-1:0] node4741;
	wire [14-1:0] node4744;
	wire [14-1:0] node4745;
	wire [14-1:0] node4746;
	wire [14-1:0] node4747;
	wire [14-1:0] node4748;
	wire [14-1:0] node4749;
	wire [14-1:0] node4750;
	wire [14-1:0] node4754;
	wire [14-1:0] node4757;
	wire [14-1:0] node4758;
	wire [14-1:0] node4759;
	wire [14-1:0] node4763;
	wire [14-1:0] node4766;
	wire [14-1:0] node4767;
	wire [14-1:0] node4768;
	wire [14-1:0] node4772;
	wire [14-1:0] node4773;
	wire [14-1:0] node4774;
	wire [14-1:0] node4777;
	wire [14-1:0] node4778;
	wire [14-1:0] node4783;
	wire [14-1:0] node4784;
	wire [14-1:0] node4785;
	wire [14-1:0] node4786;
	wire [14-1:0] node4788;
	wire [14-1:0] node4792;
	wire [14-1:0] node4793;
	wire [14-1:0] node4794;
	wire [14-1:0] node4798;
	wire [14-1:0] node4799;
	wire [14-1:0] node4800;
	wire [14-1:0] node4805;
	wire [14-1:0] node4806;
	wire [14-1:0] node4808;
	wire [14-1:0] node4809;
	wire [14-1:0] node4810;
	wire [14-1:0] node4812;
	wire [14-1:0] node4816;
	wire [14-1:0] node4817;
	wire [14-1:0] node4821;
	wire [14-1:0] node4822;
	wire [14-1:0] node4823;
	wire [14-1:0] node4826;
	wire [14-1:0] node4830;
	wire [14-1:0] node4831;
	wire [14-1:0] node4832;
	wire [14-1:0] node4833;
	wire [14-1:0] node4834;
	wire [14-1:0] node4837;
	wire [14-1:0] node4838;
	wire [14-1:0] node4842;
	wire [14-1:0] node4843;
	wire [14-1:0] node4845;
	wire [14-1:0] node4848;
	wire [14-1:0] node4851;
	wire [14-1:0] node4852;
	wire [14-1:0] node4853;
	wire [14-1:0] node4856;
	wire [14-1:0] node4858;
	wire [14-1:0] node4861;
	wire [14-1:0] node4862;
	wire [14-1:0] node4865;
	wire [14-1:0] node4868;
	wire [14-1:0] node4869;
	wire [14-1:0] node4870;
	wire [14-1:0] node4871;
	wire [14-1:0] node4873;
	wire [14-1:0] node4877;
	wire [14-1:0] node4878;
	wire [14-1:0] node4879;
	wire [14-1:0] node4882;
	wire [14-1:0] node4885;
	wire [14-1:0] node4886;
	wire [14-1:0] node4887;
	wire [14-1:0] node4892;
	wire [14-1:0] node4894;
	wire [14-1:0] node4895;
	wire [14-1:0] node4896;
	wire [14-1:0] node4899;
	wire [14-1:0] node4900;
	wire [14-1:0] node4904;
	wire [14-1:0] node4905;
	wire [14-1:0] node4909;
	wire [14-1:0] node4910;
	wire [14-1:0] node4911;
	wire [14-1:0] node4912;
	wire [14-1:0] node4913;
	wire [14-1:0] node4914;
	wire [14-1:0] node4915;
	wire [14-1:0] node4918;
	wire [14-1:0] node4920;
	wire [14-1:0] node4921;
	wire [14-1:0] node4925;
	wire [14-1:0] node4926;
	wire [14-1:0] node4927;
	wire [14-1:0] node4929;
	wire [14-1:0] node4933;
	wire [14-1:0] node4934;
	wire [14-1:0] node4938;
	wire [14-1:0] node4939;
	wire [14-1:0] node4940;
	wire [14-1:0] node4941;
	wire [14-1:0] node4944;
	wire [14-1:0] node4946;
	wire [14-1:0] node4950;
	wire [14-1:0] node4951;
	wire [14-1:0] node4952;
	wire [14-1:0] node4956;
	wire [14-1:0] node4959;
	wire [14-1:0] node4960;
	wire [14-1:0] node4961;
	wire [14-1:0] node4962;
	wire [14-1:0] node4965;
	wire [14-1:0] node4966;
	wire [14-1:0] node4970;
	wire [14-1:0] node4971;
	wire [14-1:0] node4975;
	wire [14-1:0] node4976;
	wire [14-1:0] node4977;
	wire [14-1:0] node4978;
	wire [14-1:0] node4980;
	wire [14-1:0] node4983;
	wire [14-1:0] node4987;
	wire [14-1:0] node4989;
	wire [14-1:0] node4992;
	wire [14-1:0] node4993;
	wire [14-1:0] node4994;
	wire [14-1:0] node4995;
	wire [14-1:0] node4996;
	wire [14-1:0] node4998;
	wire [14-1:0] node5000;
	wire [14-1:0] node5003;
	wire [14-1:0] node5004;
	wire [14-1:0] node5007;
	wire [14-1:0] node5010;
	wire [14-1:0] node5011;
	wire [14-1:0] node5015;
	wire [14-1:0] node5016;
	wire [14-1:0] node5017;
	wire [14-1:0] node5019;
	wire [14-1:0] node5022;
	wire [14-1:0] node5023;
	wire [14-1:0] node5026;
	wire [14-1:0] node5029;
	wire [14-1:0] node5030;
	wire [14-1:0] node5031;
	wire [14-1:0] node5032;
	wire [14-1:0] node5036;
	wire [14-1:0] node5039;
	wire [14-1:0] node5042;
	wire [14-1:0] node5043;
	wire [14-1:0] node5044;
	wire [14-1:0] node5045;
	wire [14-1:0] node5049;
	wire [14-1:0] node5050;
	wire [14-1:0] node5051;
	wire [14-1:0] node5052;
	wire [14-1:0] node5056;
	wire [14-1:0] node5059;
	wire [14-1:0] node5060;
	wire [14-1:0] node5061;
	wire [14-1:0] node5066;
	wire [14-1:0] node5067;
	wire [14-1:0] node5069;
	wire [14-1:0] node5070;
	wire [14-1:0] node5073;
	wire [14-1:0] node5074;
	wire [14-1:0] node5078;
	wire [14-1:0] node5080;
	wire [14-1:0] node5082;
	wire [14-1:0] node5084;
	wire [14-1:0] node5086;
	wire [14-1:0] node5089;
	wire [14-1:0] node5090;
	wire [14-1:0] node5091;
	wire [14-1:0] node5092;
	wire [14-1:0] node5093;
	wire [14-1:0] node5094;
	wire [14-1:0] node5096;
	wire [14-1:0] node5100;
	wire [14-1:0] node5102;
	wire [14-1:0] node5105;
	wire [14-1:0] node5106;
	wire [14-1:0] node5107;
	wire [14-1:0] node5109;
	wire [14-1:0] node5111;
	wire [14-1:0] node5112;
	wire [14-1:0] node5116;
	wire [14-1:0] node5117;
	wire [14-1:0] node5118;
	wire [14-1:0] node5123;
	wire [14-1:0] node5125;
	wire [14-1:0] node5128;
	wire [14-1:0] node5129;
	wire [14-1:0] node5130;
	wire [14-1:0] node5131;
	wire [14-1:0] node5134;
	wire [14-1:0] node5135;
	wire [14-1:0] node5138;
	wire [14-1:0] node5140;
	wire [14-1:0] node5143;
	wire [14-1:0] node5144;
	wire [14-1:0] node5146;
	wire [14-1:0] node5150;
	wire [14-1:0] node5151;
	wire [14-1:0] node5152;
	wire [14-1:0] node5153;
	wire [14-1:0] node5157;
	wire [14-1:0] node5158;
	wire [14-1:0] node5162;
	wire [14-1:0] node5164;
	wire [14-1:0] node5165;
	wire [14-1:0] node5168;
	wire [14-1:0] node5171;
	wire [14-1:0] node5172;
	wire [14-1:0] node5173;
	wire [14-1:0] node5174;
	wire [14-1:0] node5175;
	wire [14-1:0] node5176;
	wire [14-1:0] node5177;
	wire [14-1:0] node5179;
	wire [14-1:0] node5184;
	wire [14-1:0] node5186;
	wire [14-1:0] node5188;
	wire [14-1:0] node5191;
	wire [14-1:0] node5194;
	wire [14-1:0] node5195;
	wire [14-1:0] node5196;
	wire [14-1:0] node5198;
	wire [14-1:0] node5201;
	wire [14-1:0] node5202;
	wire [14-1:0] node5205;
	wire [14-1:0] node5208;
	wire [14-1:0] node5210;
	wire [14-1:0] node5212;
	wire [14-1:0] node5215;
	wire [14-1:0] node5216;
	wire [14-1:0] node5217;
	wire [14-1:0] node5219;
	wire [14-1:0] node5220;
	wire [14-1:0] node5222;
	wire [14-1:0] node5223;
	wire [14-1:0] node5228;
	wire [14-1:0] node5229;
	wire [14-1:0] node5230;
	wire [14-1:0] node5232;
	wire [14-1:0] node5237;
	wire [14-1:0] node5238;
	wire [14-1:0] node5239;
	wire [14-1:0] node5241;
	wire [14-1:0] node5242;
	wire [14-1:0] node5246;
	wire [14-1:0] node5247;
	wire [14-1:0] node5251;
	wire [14-1:0] node5253;
	wire [14-1:0] node5254;
	wire [14-1:0] node5258;
	wire [14-1:0] node5259;
	wire [14-1:0] node5260;
	wire [14-1:0] node5261;
	wire [14-1:0] node5262;
	wire [14-1:0] node5263;
	wire [14-1:0] node5264;
	wire [14-1:0] node5265;
	wire [14-1:0] node5266;
	wire [14-1:0] node5268;
	wire [14-1:0] node5269;
	wire [14-1:0] node5275;
	wire [14-1:0] node5276;
	wire [14-1:0] node5278;
	wire [14-1:0] node5279;
	wire [14-1:0] node5283;
	wire [14-1:0] node5286;
	wire [14-1:0] node5287;
	wire [14-1:0] node5289;
	wire [14-1:0] node5292;
	wire [14-1:0] node5294;
	wire [14-1:0] node5296;
	wire [14-1:0] node5299;
	wire [14-1:0] node5300;
	wire [14-1:0] node5301;
	wire [14-1:0] node5302;
	wire [14-1:0] node5305;
	wire [14-1:0] node5306;
	wire [14-1:0] node5307;
	wire [14-1:0] node5312;
	wire [14-1:0] node5313;
	wire [14-1:0] node5314;
	wire [14-1:0] node5318;
	wire [14-1:0] node5319;
	wire [14-1:0] node5323;
	wire [14-1:0] node5324;
	wire [14-1:0] node5325;
	wire [14-1:0] node5326;
	wire [14-1:0] node5329;
	wire [14-1:0] node5331;
	wire [14-1:0] node5334;
	wire [14-1:0] node5335;
	wire [14-1:0] node5339;
	wire [14-1:0] node5340;
	wire [14-1:0] node5343;
	wire [14-1:0] node5345;
	wire [14-1:0] node5348;
	wire [14-1:0] node5349;
	wire [14-1:0] node5350;
	wire [14-1:0] node5351;
	wire [14-1:0] node5352;
	wire [14-1:0] node5354;
	wire [14-1:0] node5357;
	wire [14-1:0] node5358;
	wire [14-1:0] node5362;
	wire [14-1:0] node5363;
	wire [14-1:0] node5366;
	wire [14-1:0] node5369;
	wire [14-1:0] node5370;
	wire [14-1:0] node5371;
	wire [14-1:0] node5372;
	wire [14-1:0] node5375;
	wire [14-1:0] node5377;
	wire [14-1:0] node5380;
	wire [14-1:0] node5382;
	wire [14-1:0] node5385;
	wire [14-1:0] node5387;
	wire [14-1:0] node5389;
	wire [14-1:0] node5391;
	wire [14-1:0] node5394;
	wire [14-1:0] node5395;
	wire [14-1:0] node5396;
	wire [14-1:0] node5397;
	wire [14-1:0] node5398;
	wire [14-1:0] node5401;
	wire [14-1:0] node5404;
	wire [14-1:0] node5405;
	wire [14-1:0] node5409;
	wire [14-1:0] node5411;
	wire [14-1:0] node5412;
	wire [14-1:0] node5416;
	wire [14-1:0] node5417;
	wire [14-1:0] node5420;
	wire [14-1:0] node5421;
	wire [14-1:0] node5423;
	wire [14-1:0] node5426;
	wire [14-1:0] node5427;
	wire [14-1:0] node5430;
	wire [14-1:0] node5432;
	wire [14-1:0] node5435;
	wire [14-1:0] node5436;
	wire [14-1:0] node5437;
	wire [14-1:0] node5438;
	wire [14-1:0] node5439;
	wire [14-1:0] node5441;
	wire [14-1:0] node5442;
	wire [14-1:0] node5444;
	wire [14-1:0] node5448;
	wire [14-1:0] node5449;
	wire [14-1:0] node5450;
	wire [14-1:0] node5454;
	wire [14-1:0] node5457;
	wire [14-1:0] node5458;
	wire [14-1:0] node5460;
	wire [14-1:0] node5461;
	wire [14-1:0] node5464;
	wire [14-1:0] node5467;
	wire [14-1:0] node5468;
	wire [14-1:0] node5470;
	wire [14-1:0] node5473;
	wire [14-1:0] node5474;
	wire [14-1:0] node5478;
	wire [14-1:0] node5479;
	wire [14-1:0] node5480;
	wire [14-1:0] node5481;
	wire [14-1:0] node5484;
	wire [14-1:0] node5486;
	wire [14-1:0] node5487;
	wire [14-1:0] node5489;
	wire [14-1:0] node5493;
	wire [14-1:0] node5494;
	wire [14-1:0] node5496;
	wire [14-1:0] node5500;
	wire [14-1:0] node5501;
	wire [14-1:0] node5502;
	wire [14-1:0] node5504;
	wire [14-1:0] node5506;
	wire [14-1:0] node5509;
	wire [14-1:0] node5511;
	wire [14-1:0] node5514;
	wire [14-1:0] node5516;
	wire [14-1:0] node5517;
	wire [14-1:0] node5519;
	wire [14-1:0] node5520;
	wire [14-1:0] node5525;
	wire [14-1:0] node5526;
	wire [14-1:0] node5527;
	wire [14-1:0] node5528;
	wire [14-1:0] node5529;
	wire [14-1:0] node5530;
	wire [14-1:0] node5533;
	wire [14-1:0] node5535;
	wire [14-1:0] node5538;
	wire [14-1:0] node5540;
	wire [14-1:0] node5543;
	wire [14-1:0] node5544;
	wire [14-1:0] node5545;
	wire [14-1:0] node5549;
	wire [14-1:0] node5552;
	wire [14-1:0] node5553;
	wire [14-1:0] node5554;
	wire [14-1:0] node5558;
	wire [14-1:0] node5559;
	wire [14-1:0] node5562;
	wire [14-1:0] node5563;
	wire [14-1:0] node5566;
	wire [14-1:0] node5569;
	wire [14-1:0] node5570;
	wire [14-1:0] node5571;
	wire [14-1:0] node5572;
	wire [14-1:0] node5575;
	wire [14-1:0] node5576;
	wire [14-1:0] node5579;
	wire [14-1:0] node5582;
	wire [14-1:0] node5583;
	wire [14-1:0] node5584;
	wire [14-1:0] node5586;
	wire [14-1:0] node5591;
	wire [14-1:0] node5592;
	wire [14-1:0] node5593;
	wire [14-1:0] node5595;
	wire [14-1:0] node5598;
	wire [14-1:0] node5599;
	wire [14-1:0] node5600;
	wire [14-1:0] node5604;
	wire [14-1:0] node5607;
	wire [14-1:0] node5608;
	wire [14-1:0] node5609;
	wire [14-1:0] node5613;
	wire [14-1:0] node5615;
	wire [14-1:0] node5616;
	wire [14-1:0] node5620;
	wire [14-1:0] node5621;
	wire [14-1:0] node5622;
	wire [14-1:0] node5623;
	wire [14-1:0] node5624;
	wire [14-1:0] node5625;
	wire [14-1:0] node5626;
	wire [14-1:0] node5628;
	wire [14-1:0] node5632;
	wire [14-1:0] node5633;
	wire [14-1:0] node5634;
	wire [14-1:0] node5637;
	wire [14-1:0] node5640;
	wire [14-1:0] node5641;
	wire [14-1:0] node5643;
	wire [14-1:0] node5646;
	wire [14-1:0] node5648;
	wire [14-1:0] node5651;
	wire [14-1:0] node5652;
	wire [14-1:0] node5654;
	wire [14-1:0] node5655;
	wire [14-1:0] node5658;
	wire [14-1:0] node5660;
	wire [14-1:0] node5663;
	wire [14-1:0] node5665;
	wire [14-1:0] node5668;
	wire [14-1:0] node5669;
	wire [14-1:0] node5670;
	wire [14-1:0] node5671;
	wire [14-1:0] node5672;
	wire [14-1:0] node5676;
	wire [14-1:0] node5677;
	wire [14-1:0] node5680;
	wire [14-1:0] node5683;
	wire [14-1:0] node5684;
	wire [14-1:0] node5686;
	wire [14-1:0] node5689;
	wire [14-1:0] node5691;
	wire [14-1:0] node5693;
	wire [14-1:0] node5696;
	wire [14-1:0] node5697;
	wire [14-1:0] node5698;
	wire [14-1:0] node5700;
	wire [14-1:0] node5701;
	wire [14-1:0] node5705;
	wire [14-1:0] node5706;
	wire [14-1:0] node5707;
	wire [14-1:0] node5711;
	wire [14-1:0] node5714;
	wire [14-1:0] node5715;
	wire [14-1:0] node5718;
	wire [14-1:0] node5721;
	wire [14-1:0] node5722;
	wire [14-1:0] node5723;
	wire [14-1:0] node5724;
	wire [14-1:0] node5725;
	wire [14-1:0] node5728;
	wire [14-1:0] node5729;
	wire [14-1:0] node5730;
	wire [14-1:0] node5735;
	wire [14-1:0] node5737;
	wire [14-1:0] node5738;
	wire [14-1:0] node5742;
	wire [14-1:0] node5743;
	wire [14-1:0] node5744;
	wire [14-1:0] node5745;
	wire [14-1:0] node5746;
	wire [14-1:0] node5748;
	wire [14-1:0] node5753;
	wire [14-1:0] node5756;
	wire [14-1:0] node5757;
	wire [14-1:0] node5760;
	wire [14-1:0] node5762;
	wire [14-1:0] node5763;
	wire [14-1:0] node5765;
	wire [14-1:0] node5769;
	wire [14-1:0] node5770;
	wire [14-1:0] node5771;
	wire [14-1:0] node5772;
	wire [14-1:0] node5774;
	wire [14-1:0] node5776;
	wire [14-1:0] node5778;
	wire [14-1:0] node5782;
	wire [14-1:0] node5783;
	wire [14-1:0] node5785;
	wire [14-1:0] node5787;
	wire [14-1:0] node5791;
	wire [14-1:0] node5792;
	wire [14-1:0] node5793;
	wire [14-1:0] node5794;
	wire [14-1:0] node5797;
	wire [14-1:0] node5801;
	wire [14-1:0] node5802;
	wire [14-1:0] node5804;
	wire [14-1:0] node5807;
	wire [14-1:0] node5808;
	wire [14-1:0] node5811;
	wire [14-1:0] node5813;
	wire [14-1:0] node5816;
	wire [14-1:0] node5817;
	wire [14-1:0] node5818;
	wire [14-1:0] node5819;
	wire [14-1:0] node5820;
	wire [14-1:0] node5821;
	wire [14-1:0] node5822;
	wire [14-1:0] node5827;
	wire [14-1:0] node5828;
	wire [14-1:0] node5831;
	wire [14-1:0] node5833;
	wire [14-1:0] node5834;
	wire [14-1:0] node5838;
	wire [14-1:0] node5839;
	wire [14-1:0] node5840;
	wire [14-1:0] node5841;
	wire [14-1:0] node5845;
	wire [14-1:0] node5846;
	wire [14-1:0] node5847;
	wire [14-1:0] node5851;
	wire [14-1:0] node5854;
	wire [14-1:0] node5855;
	wire [14-1:0] node5857;
	wire [14-1:0] node5860;
	wire [14-1:0] node5861;
	wire [14-1:0] node5865;
	wire [14-1:0] node5866;
	wire [14-1:0] node5867;
	wire [14-1:0] node5868;
	wire [14-1:0] node5869;
	wire [14-1:0] node5871;
	wire [14-1:0] node5875;
	wire [14-1:0] node5876;
	wire [14-1:0] node5877;
	wire [14-1:0] node5881;
	wire [14-1:0] node5884;
	wire [14-1:0] node5885;
	wire [14-1:0] node5886;
	wire [14-1:0] node5887;
	wire [14-1:0] node5892;
	wire [14-1:0] node5893;
	wire [14-1:0] node5896;
	wire [14-1:0] node5898;
	wire [14-1:0] node5899;
	wire [14-1:0] node5903;
	wire [14-1:0] node5904;
	wire [14-1:0] node5905;
	wire [14-1:0] node5906;
	wire [14-1:0] node5908;
	wire [14-1:0] node5912;
	wire [14-1:0] node5914;
	wire [14-1:0] node5917;
	wire [14-1:0] node5918;
	wire [14-1:0] node5920;
	wire [14-1:0] node5922;
	wire [14-1:0] node5925;
	wire [14-1:0] node5927;
	wire [14-1:0] node5929;
	wire [14-1:0] node5932;
	wire [14-1:0] node5933;
	wire [14-1:0] node5934;
	wire [14-1:0] node5935;
	wire [14-1:0] node5936;
	wire [14-1:0] node5938;
	wire [14-1:0] node5942;
	wire [14-1:0] node5944;
	wire [14-1:0] node5945;
	wire [14-1:0] node5949;
	wire [14-1:0] node5950;
	wire [14-1:0] node5951;
	wire [14-1:0] node5952;
	wire [14-1:0] node5956;
	wire [14-1:0] node5958;
	wire [14-1:0] node5961;
	wire [14-1:0] node5962;
	wire [14-1:0] node5963;
	wire [14-1:0] node5967;
	wire [14-1:0] node5968;
	wire [14-1:0] node5970;
	wire [14-1:0] node5974;
	wire [14-1:0] node5975;
	wire [14-1:0] node5976;
	wire [14-1:0] node5977;
	wire [14-1:0] node5979;
	wire [14-1:0] node5982;
	wire [14-1:0] node5983;
	wire [14-1:0] node5987;
	wire [14-1:0] node5988;
	wire [14-1:0] node5989;
	wire [14-1:0] node5992;
	wire [14-1:0] node5994;
	wire [14-1:0] node5995;
	wire [14-1:0] node5999;
	wire [14-1:0] node6000;
	wire [14-1:0] node6003;
	wire [14-1:0] node6005;
	wire [14-1:0] node6008;
	wire [14-1:0] node6009;
	wire [14-1:0] node6010;
	wire [14-1:0] node6012;
	wire [14-1:0] node6014;
	wire [14-1:0] node6017;
	wire [14-1:0] node6018;
	wire [14-1:0] node6021;
	wire [14-1:0] node6023;
	wire [14-1:0] node6026;
	wire [14-1:0] node6027;
	wire [14-1:0] node6028;
	wire [14-1:0] node6031;
	wire [14-1:0] node6032;
	wire [14-1:0] node6034;
	wire [14-1:0] node6037;
	wire [14-1:0] node6038;
	wire [14-1:0] node6042;
	wire [14-1:0] node6043;
	wire [14-1:0] node6046;
	wire [14-1:0] node6047;
	wire [14-1:0] node6049;

	assign outp = (inp[4]) ? node2984 : node1;
		assign node1 = (inp[10]) ? node1421 : node2;
			assign node2 = (inp[8]) ? node758 : node3;
				assign node3 = (inp[5]) ? node405 : node4;
					assign node4 = (inp[13]) ? node224 : node5;
						assign node5 = (inp[1]) ? node123 : node6;
							assign node6 = (inp[0]) ? node66 : node7;
								assign node7 = (inp[12]) ? node43 : node8;
									assign node8 = (inp[6]) ? node18 : node9;
										assign node9 = (inp[11]) ? node11 : 14'b00111111111111;
											assign node11 = (inp[7]) ? node13 : 14'b00111111111111;
												assign node13 = (inp[2]) ? 14'b00011111111111 : node14;
													assign node14 = (inp[9]) ? 14'b00011111111111 : 14'b00111111111111;
										assign node18 = (inp[2]) ? node34 : node19;
											assign node19 = (inp[9]) ? node31 : node20;
												assign node20 = (inp[11]) ? node26 : node21;
													assign node21 = (inp[3]) ? 14'b00111111111111 : node22;
														assign node22 = (inp[7]) ? 14'b00111111111111 : 14'b01111111111111;
													assign node26 = (inp[7]) ? 14'b00011111111111 : node27;
														assign node27 = (inp[3]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node31 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node34 = (inp[3]) ? 14'b00000111111111 : node35;
												assign node35 = (inp[11]) ? node37 : 14'b00011111111111;
													assign node37 = (inp[7]) ? 14'b00001111111111 : node38;
														assign node38 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node43 = (inp[11]) ? node57 : node44;
										assign node44 = (inp[6]) ? node50 : node45;
											assign node45 = (inp[9]) ? 14'b00011111111111 : node46;
												assign node46 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node50 = (inp[7]) ? 14'b00001111111111 : node51;
												assign node51 = (inp[2]) ? node53 : 14'b00011111111111;
													assign node53 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node57 = (inp[7]) ? 14'b00000111111111 : node58;
											assign node58 = (inp[2]) ? node62 : node59;
												assign node59 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node62 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node66 = (inp[11]) ? node92 : node67;
									assign node67 = (inp[12]) ? node81 : node68;
										assign node68 = (inp[6]) ? node74 : node69;
											assign node69 = (inp[3]) ? 14'b00011111111111 : node70;
												assign node70 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node74 = (inp[3]) ? 14'b00001111111111 : node75;
												assign node75 = (inp[2]) ? node77 : 14'b00011111111111;
													assign node77 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node81 = (inp[2]) ? node87 : node82;
											assign node82 = (inp[9]) ? 14'b00001111111111 : node83;
												assign node83 = (inp[6]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node87 = (inp[7]) ? node89 : 14'b00001111111111;
												assign node89 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node92 = (inp[2]) ? node110 : node93;
										assign node93 = (inp[6]) ? node103 : node94;
											assign node94 = (inp[12]) ? node98 : node95;
												assign node95 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node98 = (inp[7]) ? node100 : 14'b00001111111111;
													assign node100 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node103 = (inp[9]) ? node107 : node104;
												assign node104 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node107 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node110 = (inp[3]) ? node116 : node111;
											assign node111 = (inp[9]) ? node113 : 14'b00000111111111;
												assign node113 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node116 = (inp[6]) ? 14'b00000011111111 : node117;
												assign node117 = (inp[7]) ? node119 : 14'b00000111111111;
													assign node119 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node123 = (inp[7]) ? node175 : node124;
								assign node124 = (inp[3]) ? node150 : node125;
									assign node125 = (inp[12]) ? node139 : node126;
										assign node126 = (inp[9]) ? node134 : node127;
											assign node127 = (inp[11]) ? node129 : 14'b00111111111111;
												assign node129 = (inp[6]) ? 14'b00001111111111 : node130;
													assign node130 = (inp[0]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node134 = (inp[2]) ? 14'b00001111111111 : node135;
												assign node135 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node139 = (inp[11]) ? node145 : node140;
											assign node140 = (inp[9]) ? node142 : 14'b00011111111111;
												assign node142 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node145 = (inp[2]) ? 14'b00000111111111 : node146;
												assign node146 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node150 = (inp[11]) ? node162 : node151;
										assign node151 = (inp[2]) ? node157 : node152;
											assign node152 = (inp[6]) ? 14'b00001111111111 : node153;
												assign node153 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node157 = (inp[6]) ? node159 : 14'b00001111111111;
												assign node159 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node162 = (inp[6]) ? node166 : node163;
											assign node163 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node166 = (inp[9]) ? node170 : node167;
												assign node167 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node170 = (inp[12]) ? 14'b00000001111111 : node171;
													assign node171 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node175 = (inp[12]) ? node195 : node176;
									assign node176 = (inp[6]) ? node186 : node177;
										assign node177 = (inp[11]) ? node181 : node178;
											assign node178 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node181 = (inp[3]) ? 14'b00000111111111 : node182;
												assign node182 = (inp[9]) ? 14'b00000111111111 : 14'b00011111111111;
										assign node186 = (inp[0]) ? node188 : 14'b00000111111111;
											assign node188 = (inp[9]) ? 14'b00000011111111 : node189;
												assign node189 = (inp[11]) ? node191 : 14'b00001111111111;
													assign node191 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node195 = (inp[11]) ? node215 : node196;
										assign node196 = (inp[6]) ? node204 : node197;
											assign node197 = (inp[2]) ? node201 : node198;
												assign node198 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node201 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node204 = (inp[3]) ? node212 : node205;
												assign node205 = (inp[9]) ? node207 : 14'b00000111111111;
													assign node207 = (inp[2]) ? 14'b00000011111111 : node208;
														assign node208 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node212 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node215 = (inp[9]) ? node221 : node216;
											assign node216 = (inp[2]) ? node218 : 14'b00000011111111;
												assign node218 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node221 = (inp[6]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node224 = (inp[3]) ? node336 : node225;
							assign node225 = (inp[11]) ? node287 : node226;
								assign node226 = (inp[0]) ? node266 : node227;
									assign node227 = (inp[1]) ? node249 : node228;
										assign node228 = (inp[6]) ? node242 : node229;
											assign node229 = (inp[12]) ? 14'b00011111111111 : node230;
												assign node230 = (inp[7]) ? node236 : node231;
													assign node231 = (inp[9]) ? node233 : 14'b00111111111111;
														assign node233 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
													assign node236 = (inp[2]) ? 14'b00011111111111 : node237;
														assign node237 = (inp[9]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node242 = (inp[2]) ? node246 : node243;
												assign node243 = (inp[12]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node246 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node249 = (inp[9]) ? node257 : node250;
											assign node250 = (inp[2]) ? node252 : 14'b00001111111111;
												assign node252 = (inp[7]) ? 14'b00001111111111 : node253;
													assign node253 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node257 = (inp[12]) ? 14'b00000011111111 : node258;
												assign node258 = (inp[6]) ? 14'b00000111111111 : node259;
													assign node259 = (inp[2]) ? node261 : 14'b00011111111111;
														assign node261 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node266 = (inp[2]) ? node276 : node267;
										assign node267 = (inp[1]) ? node273 : node268;
											assign node268 = (inp[6]) ? 14'b00001111111111 : node269;
												assign node269 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node273 = (inp[9]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node276 = (inp[7]) ? node278 : 14'b00000111111111;
											assign node278 = (inp[6]) ? node282 : node279;
												assign node279 = (inp[9]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node282 = (inp[9]) ? node284 : 14'b00000011111111;
													assign node284 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node287 = (inp[1]) ? node313 : node288;
									assign node288 = (inp[0]) ? node296 : node289;
										assign node289 = (inp[6]) ? node293 : node290;
											assign node290 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node293 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node296 = (inp[7]) ? node302 : node297;
											assign node297 = (inp[2]) ? 14'b00000111111111 : node298;
												assign node298 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node302 = (inp[6]) ? node304 : 14'b00000111111111;
												assign node304 = (inp[9]) ? node310 : node305;
													assign node305 = (inp[12]) ? node307 : 14'b00000011111111;
														assign node307 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
													assign node310 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node313 = (inp[6]) ? node327 : node314;
										assign node314 = (inp[7]) ? node316 : 14'b00000111111111;
											assign node316 = (inp[2]) ? 14'b00000001111111 : node317;
												assign node317 = (inp[12]) ? node323 : node318;
													assign node318 = (inp[9]) ? node320 : 14'b00000111111111;
														assign node320 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
													assign node323 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node327 = (inp[2]) ? node333 : node328;
											assign node328 = (inp[0]) ? 14'b00000011111111 : node329;
												assign node329 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node333 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node336 = (inp[9]) ? node364 : node337;
								assign node337 = (inp[11]) ? node345 : node338;
									assign node338 = (inp[6]) ? node342 : node339;
										assign node339 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node342 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node345 = (inp[0]) ? node355 : node346;
										assign node346 = (inp[2]) ? node352 : node347;
											assign node347 = (inp[1]) ? node349 : 14'b00000111111111;
												assign node349 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node352 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node355 = (inp[2]) ? node359 : node356;
											assign node356 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node359 = (inp[6]) ? node361 : 14'b00000001111111;
												assign node361 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node364 = (inp[6]) ? node382 : node365;
									assign node365 = (inp[0]) ? node371 : node366;
										assign node366 = (inp[12]) ? 14'b00000011111111 : node367;
											assign node367 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node371 = (inp[1]) ? node379 : node372;
											assign node372 = (inp[12]) ? node374 : 14'b00000111111111;
												assign node374 = (inp[11]) ? node376 : 14'b00000011111111;
													assign node376 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node379 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node382 = (inp[12]) ? node392 : node383;
										assign node383 = (inp[2]) ? node389 : node384;
											assign node384 = (inp[1]) ? node386 : 14'b00000011111111;
												assign node386 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node389 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node392 = (inp[7]) ? node398 : node393;
											assign node393 = (inp[0]) ? node395 : 14'b00000011111111;
												assign node395 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node398 = (inp[0]) ? node400 : 14'b00000000111111;
												assign node400 = (inp[1]) ? 14'b00000000011111 : node401;
													assign node401 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node405 = (inp[1]) ? node603 : node406;
						assign node406 = (inp[6]) ? node516 : node407;
							assign node407 = (inp[7]) ? node457 : node408;
								assign node408 = (inp[3]) ? node430 : node409;
									assign node409 = (inp[9]) ? node425 : node410;
										assign node410 = (inp[11]) ? node416 : node411;
											assign node411 = (inp[2]) ? 14'b00011111111111 : node412;
												assign node412 = (inp[12]) ? 14'b00111111111111 : 14'b01111111111111;
											assign node416 = (inp[2]) ? 14'b00000111111111 : node417;
												assign node417 = (inp[0]) ? node419 : 14'b00011111111111;
													assign node419 = (inp[13]) ? 14'b00001111111111 : node420;
														assign node420 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node425 = (inp[11]) ? node427 : 14'b00001111111111;
											assign node427 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node430 = (inp[0]) ? node450 : node431;
										assign node431 = (inp[2]) ? node441 : node432;
											assign node432 = (inp[12]) ? node438 : node433;
												assign node433 = (inp[9]) ? 14'b00001111111111 : node434;
													assign node434 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node438 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node441 = (inp[12]) ? 14'b00000111111111 : node442;
												assign node442 = (inp[13]) ? 14'b00000111111111 : node443;
													assign node443 = (inp[11]) ? node445 : 14'b00001111111111;
														assign node445 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node450 = (inp[13]) ? 14'b00000111111111 : node451;
											assign node451 = (inp[12]) ? node453 : 14'b00000011111111;
												assign node453 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node457 = (inp[2]) ? node491 : node458;
									assign node458 = (inp[11]) ? node470 : node459;
										assign node459 = (inp[3]) ? node465 : node460;
											assign node460 = (inp[0]) ? node462 : 14'b00001111111111;
												assign node462 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node465 = (inp[13]) ? 14'b00000111111111 : node466;
												assign node466 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node470 = (inp[0]) ? node482 : node471;
											assign node471 = (inp[12]) ? node475 : node472;
												assign node472 = (inp[9]) ? 14'b00001111111111 : 14'b00000111111111;
												assign node475 = (inp[9]) ? 14'b00000011111111 : node476;
													assign node476 = (inp[13]) ? node478 : 14'b00000111111111;
														assign node478 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node482 = (inp[9]) ? node486 : node483;
												assign node483 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node486 = (inp[13]) ? node488 : 14'b00000011111111;
													assign node488 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node491 = (inp[3]) ? node505 : node492;
										assign node492 = (inp[12]) ? node500 : node493;
											assign node493 = (inp[11]) ? node495 : 14'b00001111111111;
												assign node495 = (inp[13]) ? node497 : 14'b00000111111111;
													assign node497 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node500 = (inp[0]) ? node502 : 14'b00000111111111;
												assign node502 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node505 = (inp[13]) ? node509 : node506;
											assign node506 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node509 = (inp[9]) ? node513 : node510;
												assign node510 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node513 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node516 = (inp[12]) ? node552 : node517;
								assign node517 = (inp[9]) ? node541 : node518;
									assign node518 = (inp[13]) ? node532 : node519;
										assign node519 = (inp[3]) ? node527 : node520;
											assign node520 = (inp[0]) ? node522 : 14'b00111111111111;
												assign node522 = (inp[11]) ? 14'b00001111111111 : node523;
													assign node523 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node527 = (inp[0]) ? node529 : 14'b00001111111111;
												assign node529 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node532 = (inp[7]) ? node534 : 14'b00000111111111;
											assign node534 = (inp[2]) ? node538 : node535;
												assign node535 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node538 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node541 = (inp[13]) ? node543 : 14'b00000011111111;
										assign node543 = (inp[3]) ? node547 : node544;
											assign node544 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node547 = (inp[11]) ? 14'b00000001111111 : node548;
												assign node548 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node552 = (inp[2]) ? node580 : node553;
									assign node553 = (inp[13]) ? node565 : node554;
										assign node554 = (inp[3]) ? node556 : 14'b00000111111111;
											assign node556 = (inp[0]) ? node560 : node557;
												assign node557 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node560 = (inp[11]) ? node562 : 14'b00000011111111;
													assign node562 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node565 = (inp[7]) ? node569 : node566;
											assign node566 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node569 = (inp[0]) ? node573 : node570;
												assign node570 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node573 = (inp[11]) ? 14'b00000000111111 : node574;
													assign node574 = (inp[9]) ? node576 : 14'b00000001111111;
														assign node576 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node580 = (inp[7]) ? node594 : node581;
										assign node581 = (inp[13]) ? node587 : node582;
											assign node582 = (inp[9]) ? node584 : 14'b00000011111111;
												assign node584 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node587 = (inp[11]) ? node589 : 14'b00000011111111;
												assign node589 = (inp[3]) ? 14'b00000000111111 : node590;
													assign node590 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node594 = (inp[0]) ? node598 : node595;
											assign node595 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node598 = (inp[3]) ? node600 : 14'b00000001111111;
												assign node600 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node603 = (inp[11]) ? node675 : node604;
							assign node604 = (inp[12]) ? node628 : node605;
								assign node605 = (inp[3]) ? node619 : node606;
									assign node606 = (inp[9]) ? node616 : node607;
										assign node607 = (inp[2]) ? node613 : node608;
											assign node608 = (inp[6]) ? 14'b00001111111111 : node609;
												assign node609 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node613 = (inp[6]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node616 = (inp[7]) ? 14'b00000011111111 : 14'b00001111111111;
									assign node619 = (inp[2]) ? 14'b00000011111111 : node620;
										assign node620 = (inp[13]) ? node624 : node621;
											assign node621 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node624 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node628 = (inp[2]) ? node652 : node629;
									assign node629 = (inp[0]) ? node639 : node630;
										assign node630 = (inp[13]) ? 14'b00000011111111 : node631;
											assign node631 = (inp[7]) ? node633 : 14'b00000111111111;
												assign node633 = (inp[3]) ? 14'b00000011111111 : node634;
													assign node634 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node639 = (inp[9]) ? 14'b00000001111111 : node640;
											assign node640 = (inp[3]) ? node648 : node641;
												assign node641 = (inp[13]) ? 14'b00000011111111 : node642;
													assign node642 = (inp[7]) ? node644 : 14'b00000111111111;
														assign node644 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node648 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node652 = (inp[0]) ? node662 : node653;
										assign node653 = (inp[7]) ? node659 : node654;
											assign node654 = (inp[9]) ? 14'b00000011111111 : node655;
												assign node655 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node659 = (inp[6]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node662 = (inp[6]) ? node664 : 14'b00000001111111;
											assign node664 = (inp[9]) ? node668 : node665;
												assign node665 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node668 = (inp[7]) ? 14'b00000000011111 : node669;
													assign node669 = (inp[3]) ? node671 : 14'b00000000111111;
														assign node671 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node675 = (inp[7]) ? node711 : node676;
								assign node676 = (inp[13]) ? node690 : node677;
									assign node677 = (inp[6]) ? node683 : node678;
										assign node678 = (inp[0]) ? node680 : 14'b00000111111111;
											assign node680 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node683 = (inp[3]) ? 14'b00000011111111 : node684;
											assign node684 = (inp[2]) ? 14'b00000011111111 : node685;
												assign node685 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node690 = (inp[0]) ? node700 : node691;
										assign node691 = (inp[2]) ? node697 : node692;
											assign node692 = (inp[6]) ? 14'b00000011111111 : node693;
												assign node693 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node697 = (inp[6]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node700 = (inp[2]) ? node706 : node701;
											assign node701 = (inp[3]) ? node703 : 14'b00000011111111;
												assign node703 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node706 = (inp[3]) ? 14'b00000000111111 : node707;
												assign node707 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node711 = (inp[0]) ? node737 : node712;
									assign node712 = (inp[3]) ? node728 : node713;
										assign node713 = (inp[13]) ? node723 : node714;
											assign node714 = (inp[6]) ? node716 : 14'b00000011111111;
												assign node716 = (inp[12]) ? 14'b00000001111111 : node717;
													assign node717 = (inp[9]) ? node719 : 14'b00000011111111;
														assign node719 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node723 = (inp[2]) ? 14'b00000000111111 : node724;
												assign node724 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node728 = (inp[13]) ? node732 : node729;
											assign node729 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node732 = (inp[12]) ? node734 : 14'b00000000111111;
												assign node734 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node737 = (inp[12]) ? node745 : node738;
										assign node738 = (inp[2]) ? node740 : 14'b00000001111111;
											assign node740 = (inp[3]) ? node742 : 14'b00000000111111;
												assign node742 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node745 = (inp[6]) ? node749 : node746;
											assign node746 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node749 = (inp[3]) ? node751 : 14'b00000000011111;
												assign node751 = (inp[9]) ? node753 : 14'b00000000011111;
													assign node753 = (inp[2]) ? node755 : 14'b00000000001111;
														assign node755 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node758 = (inp[12]) ? node1106 : node759;
					assign node759 = (inp[2]) ? node947 : node760;
						assign node760 = (inp[13]) ? node858 : node761;
							assign node761 = (inp[5]) ? node819 : node762;
								assign node762 = (inp[0]) ? node792 : node763;
									assign node763 = (inp[9]) ? node775 : node764;
										assign node764 = (inp[6]) ? node766 : 14'b00011111111111;
											assign node766 = (inp[3]) ? 14'b00001111111111 : node767;
												assign node767 = (inp[11]) ? node769 : 14'b00011111111111;
													assign node769 = (inp[7]) ? 14'b00001111111111 : node770;
														assign node770 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node775 = (inp[3]) ? node787 : node776;
											assign node776 = (inp[11]) ? node784 : node777;
												assign node777 = (inp[1]) ? 14'b00001111111111 : node778;
													assign node778 = (inp[6]) ? node780 : 14'b00011111111111;
														assign node780 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node784 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node787 = (inp[6]) ? node789 : 14'b00001111111111;
												assign node789 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node792 = (inp[7]) ? node808 : node793;
										assign node793 = (inp[9]) ? node801 : node794;
											assign node794 = (inp[3]) ? node798 : node795;
												assign node795 = (inp[6]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node798 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node801 = (inp[6]) ? 14'b00000111111111 : node802;
												assign node802 = (inp[3]) ? 14'b00000111111111 : node803;
													assign node803 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node808 = (inp[9]) ? node816 : node809;
											assign node809 = (inp[1]) ? 14'b00000111111111 : node810;
												assign node810 = (inp[6]) ? 14'b00000111111111 : node811;
													assign node811 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node816 = (inp[11]) ? 14'b00000001111111 : 14'b00000111111111;
								assign node819 = (inp[0]) ? node841 : node820;
									assign node820 = (inp[9]) ? node832 : node821;
										assign node821 = (inp[7]) ? node829 : node822;
											assign node822 = (inp[6]) ? node826 : node823;
												assign node823 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node826 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node829 = (inp[11]) ? 14'b00001111111111 : 14'b00000111111111;
										assign node832 = (inp[1]) ? node836 : node833;
											assign node833 = (inp[7]) ? 14'b00000111111111 : 14'b00011111111111;
											assign node836 = (inp[7]) ? 14'b00000011111111 : node837;
												assign node837 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node841 = (inp[1]) ? node847 : node842;
										assign node842 = (inp[6]) ? 14'b00000011111111 : node843;
											assign node843 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node847 = (inp[7]) ? node849 : 14'b00000011111111;
											assign node849 = (inp[3]) ? node853 : node850;
												assign node850 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node853 = (inp[6]) ? 14'b00000000011111 : node854;
													assign node854 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node858 = (inp[6]) ? node902 : node859;
								assign node859 = (inp[3]) ? node875 : node860;
									assign node860 = (inp[11]) ? node868 : node861;
										assign node861 = (inp[5]) ? 14'b00000011111111 : node862;
											assign node862 = (inp[7]) ? node864 : 14'b00001111111111;
												assign node864 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node868 = (inp[1]) ? 14'b00000111111111 : node869;
											assign node869 = (inp[7]) ? 14'b00000111111111 : node870;
												assign node870 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node875 = (inp[5]) ? node891 : node876;
										assign node876 = (inp[1]) ? node884 : node877;
											assign node877 = (inp[9]) ? node881 : node878;
												assign node878 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node881 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node884 = (inp[0]) ? node888 : node885;
												assign node885 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node888 = (inp[7]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node891 = (inp[7]) ? node897 : node892;
											assign node892 = (inp[1]) ? node894 : 14'b00000011111111;
												assign node894 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node897 = (inp[1]) ? 14'b00000000111111 : node898;
												assign node898 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node902 = (inp[5]) ? node930 : node903;
									assign node903 = (inp[11]) ? node915 : node904;
										assign node904 = (inp[1]) ? node910 : node905;
											assign node905 = (inp[9]) ? node907 : 14'b00000111111111;
												assign node907 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node910 = (inp[7]) ? 14'b00000011111111 : node911;
												assign node911 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node915 = (inp[3]) ? node921 : node916;
											assign node916 = (inp[1]) ? 14'b00000001111111 : node917;
												assign node917 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node921 = (inp[7]) ? node923 : 14'b00000011111111;
												assign node923 = (inp[9]) ? node925 : 14'b00000001111111;
													assign node925 = (inp[0]) ? node927 : 14'b00000001111111;
														assign node927 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node930 = (inp[9]) ? node944 : node931;
										assign node931 = (inp[3]) ? node939 : node932;
											assign node932 = (inp[1]) ? node934 : 14'b00000011111111;
												assign node934 = (inp[0]) ? 14'b00000001111111 : node935;
													assign node935 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node939 = (inp[1]) ? node941 : 14'b00000001111111;
												assign node941 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node944 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node947 = (inp[9]) ? node1031 : node948;
							assign node948 = (inp[0]) ? node998 : node949;
								assign node949 = (inp[7]) ? node979 : node950;
									assign node950 = (inp[11]) ? node970 : node951;
										assign node951 = (inp[13]) ? node963 : node952;
											assign node952 = (inp[1]) ? node958 : node953;
												assign node953 = (inp[5]) ? node955 : 14'b00011111111111;
													assign node955 = (inp[6]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node958 = (inp[6]) ? 14'b00000111111111 : node959;
													assign node959 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node963 = (inp[5]) ? node967 : node964;
												assign node964 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node967 = (inp[1]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node970 = (inp[6]) ? node976 : node971;
											assign node971 = (inp[13]) ? 14'b00000111111111 : node972;
												assign node972 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node976 = (inp[5]) ? 14'b00000011111111 : 14'b00000001111111;
									assign node979 = (inp[1]) ? node991 : node980;
										assign node980 = (inp[6]) ? node986 : node981;
											assign node981 = (inp[13]) ? node983 : 14'b00000111111111;
												assign node983 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node986 = (inp[3]) ? 14'b00000011111111 : node987;
												assign node987 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node991 = (inp[5]) ? 14'b00000001111111 : node992;
											assign node992 = (inp[13]) ? 14'b00000011111111 : node993;
												assign node993 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node998 = (inp[3]) ? node1018 : node999;
									assign node999 = (inp[11]) ? node1009 : node1000;
										assign node1000 = (inp[1]) ? node1002 : 14'b00000111111111;
											assign node1002 = (inp[5]) ? 14'b00000001111111 : node1003;
												assign node1003 = (inp[13]) ? 14'b00000011111111 : node1004;
													assign node1004 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1009 = (inp[1]) ? node1015 : node1010;
											assign node1010 = (inp[6]) ? node1012 : 14'b00000011111111;
												assign node1012 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1015 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1018 = (inp[11]) ? node1024 : node1019;
										assign node1019 = (inp[13]) ? node1021 : 14'b00000011111111;
											assign node1021 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1024 = (inp[1]) ? node1026 : 14'b00000001111111;
											assign node1026 = (inp[13]) ? node1028 : 14'b00000000111111;
												assign node1028 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1031 = (inp[6]) ? node1067 : node1032;
								assign node1032 = (inp[7]) ? node1042 : node1033;
									assign node1033 = (inp[11]) ? 14'b00000011111111 : node1034;
										assign node1034 = (inp[3]) ? node1036 : 14'b00000111111111;
											assign node1036 = (inp[1]) ? 14'b00000001111111 : node1037;
												assign node1037 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1042 = (inp[13]) ? node1056 : node1043;
										assign node1043 = (inp[5]) ? node1051 : node1044;
											assign node1044 = (inp[1]) ? 14'b00000111111111 : node1045;
												assign node1045 = (inp[0]) ? node1047 : 14'b00000011111111;
													assign node1047 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1051 = (inp[11]) ? 14'b00000001111111 : node1052;
												assign node1052 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1056 = (inp[0]) ? node1062 : node1057;
											assign node1057 = (inp[11]) ? 14'b00000001111111 : node1058;
												assign node1058 = (inp[5]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1062 = (inp[3]) ? node1064 : 14'b00000001111111;
												assign node1064 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1067 = (inp[5]) ? node1085 : node1068;
									assign node1068 = (inp[3]) ? node1078 : node1069;
										assign node1069 = (inp[11]) ? node1073 : node1070;
											assign node1070 = (inp[7]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node1073 = (inp[1]) ? node1075 : 14'b00000011111111;
												assign node1075 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1078 = (inp[13]) ? 14'b00000000111111 : node1079;
											assign node1079 = (inp[11]) ? node1081 : 14'b00000011111111;
												assign node1081 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1085 = (inp[7]) ? node1093 : node1086;
										assign node1086 = (inp[0]) ? node1090 : node1087;
											assign node1087 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1090 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1093 = (inp[13]) ? node1101 : node1094;
											assign node1094 = (inp[1]) ? node1096 : 14'b00000000111111;
												assign node1096 = (inp[3]) ? node1098 : 14'b00000000111111;
													assign node1098 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1101 = (inp[3]) ? 14'b00000000011111 : node1102;
												assign node1102 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node1106 = (inp[5]) ? node1272 : node1107;
						assign node1107 = (inp[9]) ? node1191 : node1108;
							assign node1108 = (inp[7]) ? node1150 : node1109;
								assign node1109 = (inp[13]) ? node1131 : node1110;
									assign node1110 = (inp[6]) ? node1122 : node1111;
										assign node1111 = (inp[1]) ? node1115 : node1112;
											assign node1112 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1115 = (inp[11]) ? 14'b00000011111111 : node1116;
												assign node1116 = (inp[0]) ? node1118 : 14'b00001111111111;
													assign node1118 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1122 = (inp[11]) ? 14'b00000011111111 : node1123;
											assign node1123 = (inp[3]) ? node1127 : node1124;
												assign node1124 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1127 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1131 = (inp[6]) ? node1147 : node1132;
										assign node1132 = (inp[1]) ? node1140 : node1133;
											assign node1133 = (inp[3]) ? node1137 : node1134;
												assign node1134 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1137 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node1140 = (inp[3]) ? 14'b00000001111111 : node1141;
												assign node1141 = (inp[11]) ? 14'b00000011111111 : node1142;
													assign node1142 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1147 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1150 = (inp[1]) ? node1170 : node1151;
									assign node1151 = (inp[13]) ? node1161 : node1152;
										assign node1152 = (inp[2]) ? node1156 : node1153;
											assign node1153 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1156 = (inp[0]) ? node1158 : 14'b00000011111111;
												assign node1158 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1161 = (inp[6]) ? node1163 : 14'b00000011111111;
											assign node1163 = (inp[11]) ? node1167 : node1164;
												assign node1164 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1167 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1170 = (inp[0]) ? node1180 : node1171;
										assign node1171 = (inp[13]) ? node1177 : node1172;
											assign node1172 = (inp[2]) ? node1174 : 14'b00000011111111;
												assign node1174 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1177 = (inp[11]) ? 14'b00000000111111 : 14'b00000111111111;
										assign node1180 = (inp[13]) ? node1188 : node1181;
											assign node1181 = (inp[3]) ? node1183 : 14'b00000001111111;
												assign node1183 = (inp[6]) ? node1185 : 14'b00000001111111;
													assign node1185 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1188 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1191 = (inp[1]) ? node1231 : node1192;
								assign node1192 = (inp[0]) ? node1208 : node1193;
									assign node1193 = (inp[2]) ? node1197 : node1194;
										assign node1194 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1197 = (inp[6]) ? node1199 : 14'b00000011111111;
											assign node1199 = (inp[3]) ? 14'b00000000111111 : node1200;
												assign node1200 = (inp[7]) ? 14'b00000001111111 : node1201;
													assign node1201 = (inp[13]) ? node1203 : 14'b00000011111111;
														assign node1203 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1208 = (inp[3]) ? node1216 : node1209;
										assign node1209 = (inp[6]) ? node1211 : 14'b00000111111111;
											assign node1211 = (inp[13]) ? 14'b00000001111111 : node1212;
												assign node1212 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1216 = (inp[11]) ? node1218 : 14'b00000001111111;
											assign node1218 = (inp[13]) ? node1226 : node1219;
												assign node1219 = (inp[2]) ? node1223 : node1220;
													assign node1220 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
													assign node1223 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1226 = (inp[6]) ? 14'b00000000111111 : node1227;
													assign node1227 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1231 = (inp[13]) ? node1257 : node1232;
									assign node1232 = (inp[6]) ? node1240 : node1233;
										assign node1233 = (inp[2]) ? node1235 : 14'b00000011111111;
											assign node1235 = (inp[11]) ? 14'b00000001111111 : node1236;
												assign node1236 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1240 = (inp[7]) ? node1252 : node1241;
											assign node1241 = (inp[11]) ? node1247 : node1242;
												assign node1242 = (inp[2]) ? 14'b00000001111111 : node1243;
													assign node1243 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1247 = (inp[3]) ? node1249 : 14'b00000001111111;
													assign node1249 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1252 = (inp[3]) ? 14'b00000000111111 : node1253;
												assign node1253 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1257 = (inp[7]) ? node1267 : node1258;
										assign node1258 = (inp[6]) ? node1264 : node1259;
											assign node1259 = (inp[11]) ? node1261 : 14'b00000001111111;
												assign node1261 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1264 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1267 = (inp[0]) ? node1269 : 14'b00000000111111;
											assign node1269 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node1272 = (inp[6]) ? node1336 : node1273;
							assign node1273 = (inp[1]) ? node1301 : node1274;
								assign node1274 = (inp[13]) ? node1290 : node1275;
									assign node1275 = (inp[2]) ? node1283 : node1276;
										assign node1276 = (inp[11]) ? 14'b00000011111111 : node1277;
											assign node1277 = (inp[7]) ? node1279 : 14'b00000111111111;
												assign node1279 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1283 = (inp[0]) ? 14'b00000001111111 : node1284;
											assign node1284 = (inp[11]) ? node1286 : 14'b00000011111111;
												assign node1286 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1290 = (inp[11]) ? node1296 : node1291;
										assign node1291 = (inp[3]) ? 14'b00000001111111 : node1292;
											assign node1292 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1296 = (inp[7]) ? 14'b00000000111111 : node1297;
											assign node1297 = (inp[0]) ? 14'b00000000111111 : 14'b00000111111111;
								assign node1301 = (inp[9]) ? node1317 : node1302;
									assign node1302 = (inp[7]) ? node1312 : node1303;
										assign node1303 = (inp[13]) ? node1305 : 14'b00000111111111;
											assign node1305 = (inp[11]) ? 14'b00000001111111 : node1306;
												assign node1306 = (inp[3]) ? node1308 : 14'b00000011111111;
													assign node1308 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1312 = (inp[11]) ? node1314 : 14'b00000001111111;
											assign node1314 = (inp[0]) ? 14'b00000000001111 : 14'b00000001111111;
									assign node1317 = (inp[11]) ? node1331 : node1318;
										assign node1318 = (inp[2]) ? node1324 : node1319;
											assign node1319 = (inp[0]) ? node1321 : 14'b00000001111111;
												assign node1321 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1324 = (inp[3]) ? node1326 : 14'b00000001111111;
												assign node1326 = (inp[0]) ? 14'b00000000011111 : node1327;
													assign node1327 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1331 = (inp[13]) ? node1333 : 14'b00000000111111;
											assign node1333 = (inp[3]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node1336 = (inp[13]) ? node1384 : node1337;
								assign node1337 = (inp[2]) ? node1357 : node1338;
									assign node1338 = (inp[0]) ? node1352 : node1339;
										assign node1339 = (inp[3]) ? node1347 : node1340;
											assign node1340 = (inp[11]) ? node1344 : node1341;
												assign node1341 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1344 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1347 = (inp[11]) ? 14'b00000000111111 : node1348;
												assign node1348 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1352 = (inp[3]) ? 14'b00000001111111 : node1353;
											assign node1353 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1357 = (inp[9]) ? node1371 : node1358;
										assign node1358 = (inp[0]) ? node1366 : node1359;
											assign node1359 = (inp[1]) ? node1361 : 14'b00000011111111;
												assign node1361 = (inp[7]) ? 14'b00000001111111 : node1362;
													assign node1362 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1366 = (inp[1]) ? 14'b00000000111111 : node1367;
												assign node1367 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1371 = (inp[7]) ? node1379 : node1372;
											assign node1372 = (inp[3]) ? node1374 : 14'b00000000111111;
												assign node1374 = (inp[11]) ? 14'b00000000011111 : node1375;
													assign node1375 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1379 = (inp[11]) ? node1381 : 14'b00000000011111;
												assign node1381 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node1384 = (inp[1]) ? node1402 : node1385;
									assign node1385 = (inp[3]) ? node1395 : node1386;
										assign node1386 = (inp[11]) ? node1392 : node1387;
											assign node1387 = (inp[2]) ? 14'b00000001111111 : node1388;
												assign node1388 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1392 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1395 = (inp[7]) ? node1397 : 14'b00000000111111;
											assign node1397 = (inp[11]) ? node1399 : 14'b00000000011111;
												assign node1399 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node1402 = (inp[2]) ? node1408 : node1403;
										assign node1403 = (inp[9]) ? 14'b00000000011111 : node1404;
											assign node1404 = (inp[11]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node1408 = (inp[3]) ? node1416 : node1409;
											assign node1409 = (inp[0]) ? node1413 : node1410;
												assign node1410 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1413 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node1416 = (inp[0]) ? node1418 : 14'b00000000001111;
												assign node1418 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
			assign node1421 = (inp[13]) ? node2199 : node1422;
				assign node1422 = (inp[0]) ? node1812 : node1423;
					assign node1423 = (inp[9]) ? node1635 : node1424;
						assign node1424 = (inp[2]) ? node1540 : node1425;
							assign node1425 = (inp[1]) ? node1495 : node1426;
								assign node1426 = (inp[3]) ? node1456 : node1427;
									assign node1427 = (inp[7]) ? node1441 : node1428;
										assign node1428 = (inp[8]) ? node1434 : node1429;
											assign node1429 = (inp[6]) ? node1431 : 14'b00011111111111;
												assign node1431 = (inp[11]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node1434 = (inp[6]) ? 14'b00001111111111 : node1435;
												assign node1435 = (inp[5]) ? node1437 : 14'b00011111111111;
													assign node1437 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node1441 = (inp[6]) ? node1451 : node1442;
											assign node1442 = (inp[8]) ? node1446 : node1443;
												assign node1443 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1446 = (inp[5]) ? node1448 : 14'b00001111111111;
													assign node1448 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1451 = (inp[8]) ? 14'b00000011111111 : node1452;
												assign node1452 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node1456 = (inp[6]) ? node1476 : node1457;
										assign node1457 = (inp[8]) ? node1463 : node1458;
											assign node1458 = (inp[5]) ? node1460 : 14'b00001111111111;
												assign node1460 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1463 = (inp[5]) ? node1471 : node1464;
												assign node1464 = (inp[11]) ? node1466 : 14'b00011111111111;
													assign node1466 = (inp[12]) ? 14'b00000111111111 : node1467;
														assign node1467 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1471 = (inp[11]) ? node1473 : 14'b00000111111111;
													assign node1473 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1476 = (inp[11]) ? node1486 : node1477;
											assign node1477 = (inp[12]) ? node1479 : 14'b00001111111111;
												assign node1479 = (inp[8]) ? node1481 : 14'b00000111111111;
													assign node1481 = (inp[5]) ? 14'b00000011111111 : node1482;
														assign node1482 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1486 = (inp[8]) ? node1492 : node1487;
												assign node1487 = (inp[12]) ? 14'b00000011111111 : node1488;
													assign node1488 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1492 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1495 = (inp[5]) ? node1519 : node1496;
									assign node1496 = (inp[6]) ? node1512 : node1497;
										assign node1497 = (inp[8]) ? node1505 : node1498;
											assign node1498 = (inp[11]) ? 14'b00001111111111 : node1499;
												assign node1499 = (inp[3]) ? 14'b00011111111111 : node1500;
													assign node1500 = (inp[12]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node1505 = (inp[3]) ? node1507 : 14'b00000011111111;
												assign node1507 = (inp[7]) ? 14'b00000111111111 : node1508;
													assign node1508 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1512 = (inp[3]) ? node1514 : 14'b00000111111111;
											assign node1514 = (inp[8]) ? 14'b00000001111111 : node1515;
												assign node1515 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1519 = (inp[12]) ? node1527 : node1520;
										assign node1520 = (inp[3]) ? node1522 : 14'b00000111111111;
											assign node1522 = (inp[7]) ? 14'b00000011111111 : node1523;
												assign node1523 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1527 = (inp[11]) ? node1535 : node1528;
											assign node1528 = (inp[3]) ? node1532 : node1529;
												assign node1529 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1532 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1535 = (inp[8]) ? node1537 : 14'b00000011111111;
												assign node1537 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1540 = (inp[7]) ? node1592 : node1541;
								assign node1541 = (inp[6]) ? node1569 : node1542;
									assign node1542 = (inp[1]) ? node1554 : node1543;
										assign node1543 = (inp[12]) ? node1549 : node1544;
											assign node1544 = (inp[11]) ? node1546 : 14'b00011111111111;
												assign node1546 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1549 = (inp[3]) ? 14'b00000111111111 : node1550;
												assign node1550 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1554 = (inp[3]) ? 14'b00000011111111 : node1555;
											assign node1555 = (inp[5]) ? node1563 : node1556;
												assign node1556 = (inp[12]) ? 14'b00000111111111 : node1557;
													assign node1557 = (inp[11]) ? node1559 : 14'b00001111111111;
														assign node1559 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1563 = (inp[11]) ? node1565 : 14'b00000111111111;
													assign node1565 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1569 = (inp[11]) ? node1587 : node1570;
										assign node1570 = (inp[3]) ? node1576 : node1571;
											assign node1571 = (inp[5]) ? node1573 : 14'b00001111111111;
												assign node1573 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1576 = (inp[12]) ? node1584 : node1577;
												assign node1577 = (inp[5]) ? 14'b00000011111111 : node1578;
													assign node1578 = (inp[8]) ? node1580 : 14'b00000111111111;
														assign node1580 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1584 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1587 = (inp[12]) ? node1589 : 14'b00000011111111;
											assign node1589 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1592 = (inp[1]) ? node1618 : node1593;
									assign node1593 = (inp[5]) ? node1605 : node1594;
										assign node1594 = (inp[8]) ? node1600 : node1595;
											assign node1595 = (inp[12]) ? 14'b00000001111111 : node1596;
												assign node1596 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1600 = (inp[6]) ? 14'b00000011111111 : node1601;
												assign node1601 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1605 = (inp[12]) ? node1615 : node1606;
											assign node1606 = (inp[11]) ? node1610 : node1607;
												assign node1607 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1610 = (inp[3]) ? 14'b00000001111111 : node1611;
													assign node1611 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1615 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1618 = (inp[6]) ? node1630 : node1619;
										assign node1619 = (inp[5]) ? node1625 : node1620;
											assign node1620 = (inp[11]) ? node1622 : 14'b00000011111111;
												assign node1622 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1625 = (inp[8]) ? node1627 : 14'b00000001111111;
												assign node1627 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1630 = (inp[8]) ? node1632 : 14'b00000001111111;
											assign node1632 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node1635 = (inp[1]) ? node1717 : node1636;
							assign node1636 = (inp[8]) ? node1666 : node1637;
								assign node1637 = (inp[11]) ? node1659 : node1638;
									assign node1638 = (inp[5]) ? node1652 : node1639;
										assign node1639 = (inp[2]) ? node1643 : node1640;
											assign node1640 = (inp[3]) ? 14'b00011111111111 : 14'b00001111111111;
											assign node1643 = (inp[6]) ? node1649 : node1644;
												assign node1644 = (inp[12]) ? 14'b00000111111111 : node1645;
													assign node1645 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1649 = (inp[12]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node1652 = (inp[6]) ? 14'b00000011111111 : node1653;
											assign node1653 = (inp[3]) ? node1655 : 14'b00001111111111;
												assign node1655 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1659 = (inp[7]) ? node1663 : node1660;
										assign node1660 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1663 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
								assign node1666 = (inp[5]) ? node1698 : node1667;
									assign node1667 = (inp[3]) ? node1685 : node1668;
										assign node1668 = (inp[7]) ? node1678 : node1669;
											assign node1669 = (inp[6]) ? node1675 : node1670;
												assign node1670 = (inp[12]) ? node1672 : 14'b00001111111111;
													assign node1672 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1675 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1678 = (inp[2]) ? 14'b00000011111111 : node1679;
												assign node1679 = (inp[12]) ? 14'b00000011111111 : node1680;
													assign node1680 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1685 = (inp[6]) ? node1691 : node1686;
											assign node1686 = (inp[11]) ? 14'b00000011111111 : node1687;
												assign node1687 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1691 = (inp[12]) ? node1695 : node1692;
												assign node1692 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1695 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1698 = (inp[6]) ? node1712 : node1699;
										assign node1699 = (inp[7]) ? node1709 : node1700;
											assign node1700 = (inp[12]) ? 14'b00000001111111 : node1701;
												assign node1701 = (inp[3]) ? 14'b00000011111111 : node1702;
													assign node1702 = (inp[2]) ? node1704 : 14'b00000111111111;
														assign node1704 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1709 = (inp[12]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node1712 = (inp[11]) ? node1714 : 14'b00000001111111;
											assign node1714 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1717 = (inp[6]) ? node1765 : node1718;
								assign node1718 = (inp[11]) ? node1744 : node1719;
									assign node1719 = (inp[8]) ? node1735 : node1720;
										assign node1720 = (inp[12]) ? node1730 : node1721;
											assign node1721 = (inp[5]) ? node1727 : node1722;
												assign node1722 = (inp[3]) ? 14'b00000111111111 : node1723;
													assign node1723 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1727 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1730 = (inp[7]) ? 14'b00000011111111 : node1731;
												assign node1731 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1735 = (inp[5]) ? node1741 : node1736;
											assign node1736 = (inp[7]) ? 14'b00000011111111 : node1737;
												assign node1737 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1741 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node1744 = (inp[5]) ? node1760 : node1745;
										assign node1745 = (inp[12]) ? node1755 : node1746;
											assign node1746 = (inp[3]) ? node1750 : node1747;
												assign node1747 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1750 = (inp[8]) ? 14'b00000001111111 : node1751;
													assign node1751 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1755 = (inp[2]) ? node1757 : 14'b00000001111111;
												assign node1757 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1760 = (inp[3]) ? 14'b00000000011111 : node1761;
											assign node1761 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1765 = (inp[7]) ? node1787 : node1766;
									assign node1766 = (inp[12]) ? node1778 : node1767;
										assign node1767 = (inp[8]) ? node1773 : node1768;
											assign node1768 = (inp[5]) ? 14'b00000011111111 : node1769;
												assign node1769 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node1773 = (inp[11]) ? 14'b00000000111111 : node1774;
												assign node1774 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1778 = (inp[5]) ? node1780 : 14'b00000001111111;
											assign node1780 = (inp[3]) ? node1782 : 14'b00000001111111;
												assign node1782 = (inp[11]) ? node1784 : 14'b00000000111111;
													assign node1784 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1787 = (inp[3]) ? node1799 : node1788;
										assign node1788 = (inp[5]) ? node1794 : node1789;
											assign node1789 = (inp[12]) ? 14'b00000000111111 : node1790;
												assign node1790 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1794 = (inp[8]) ? node1796 : 14'b00000000111111;
												assign node1796 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1799 = (inp[2]) ? node1805 : node1800;
											assign node1800 = (inp[11]) ? node1802 : 14'b00000000111111;
												assign node1802 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1805 = (inp[8]) ? 14'b00000000001111 : node1806;
												assign node1806 = (inp[11]) ? 14'b00000000011111 : node1807;
													assign node1807 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node1812 = (inp[8]) ? node2020 : node1813;
						assign node1813 = (inp[7]) ? node1917 : node1814;
							assign node1814 = (inp[9]) ? node1870 : node1815;
								assign node1815 = (inp[3]) ? node1847 : node1816;
									assign node1816 = (inp[11]) ? node1828 : node1817;
										assign node1817 = (inp[12]) ? node1823 : node1818;
											assign node1818 = (inp[6]) ? node1820 : 14'b00011111111111;
												assign node1820 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1823 = (inp[1]) ? 14'b00000111111111 : node1824;
												assign node1824 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1828 = (inp[12]) ? node1842 : node1829;
											assign node1829 = (inp[6]) ? node1835 : node1830;
												assign node1830 = (inp[1]) ? node1832 : 14'b00001111111111;
													assign node1832 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1835 = (inp[1]) ? 14'b00000011111111 : node1836;
													assign node1836 = (inp[5]) ? 14'b00000111111111 : node1837;
														assign node1837 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1842 = (inp[6]) ? 14'b00000011111111 : node1843;
												assign node1843 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1847 = (inp[2]) ? node1855 : node1848;
										assign node1848 = (inp[5]) ? node1852 : node1849;
											assign node1849 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1852 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1855 = (inp[6]) ? node1861 : node1856;
											assign node1856 = (inp[1]) ? 14'b00000011111111 : node1857;
												assign node1857 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node1861 = (inp[11]) ? node1865 : node1862;
												assign node1862 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1865 = (inp[1]) ? 14'b00000001111111 : node1866;
													assign node1866 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1870 = (inp[5]) ? node1892 : node1871;
									assign node1871 = (inp[3]) ? node1885 : node1872;
										assign node1872 = (inp[1]) ? node1878 : node1873;
											assign node1873 = (inp[12]) ? 14'b00000111111111 : node1874;
												assign node1874 = (inp[11]) ? 14'b00000111111111 : 14'b00011111111111;
											assign node1878 = (inp[11]) ? node1882 : node1879;
												assign node1879 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1882 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1885 = (inp[6]) ? node1887 : 14'b00000011111111;
											assign node1887 = (inp[1]) ? 14'b00000000111111 : node1888;
												assign node1888 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1892 = (inp[6]) ? node1906 : node1893;
										assign node1893 = (inp[11]) ? node1897 : node1894;
											assign node1894 = (inp[12]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node1897 = (inp[2]) ? node1903 : node1898;
												assign node1898 = (inp[1]) ? 14'b00000001111111 : node1899;
													assign node1899 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1903 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1906 = (inp[1]) ? node1912 : node1907;
											assign node1907 = (inp[2]) ? 14'b00000000111111 : node1908;
												assign node1908 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1912 = (inp[12]) ? 14'b00000000011111 : node1913;
												assign node1913 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1917 = (inp[1]) ? node1963 : node1918;
								assign node1918 = (inp[11]) ? node1936 : node1919;
									assign node1919 = (inp[6]) ? node1925 : node1920;
										assign node1920 = (inp[5]) ? 14'b00000011111111 : node1921;
											assign node1921 = (inp[9]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node1925 = (inp[9]) ? node1931 : node1926;
											assign node1926 = (inp[2]) ? node1928 : 14'b00000011111111;
												assign node1928 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1931 = (inp[5]) ? 14'b00000000111111 : node1932;
												assign node1932 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1936 = (inp[6]) ? node1950 : node1937;
										assign node1937 = (inp[9]) ? node1945 : node1938;
											assign node1938 = (inp[5]) ? node1942 : node1939;
												assign node1939 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1942 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1945 = (inp[2]) ? 14'b00000001111111 : node1946;
												assign node1946 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1950 = (inp[9]) ? 14'b00000000111111 : node1951;
											assign node1951 = (inp[2]) ? node1953 : 14'b00000111111111;
												assign node1953 = (inp[5]) ? node1957 : node1954;
													assign node1954 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
													assign node1957 = (inp[12]) ? 14'b00000000111111 : node1958;
														assign node1958 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1963 = (inp[3]) ? node1991 : node1964;
									assign node1964 = (inp[2]) ? node1976 : node1965;
										assign node1965 = (inp[5]) ? node1973 : node1966;
											assign node1966 = (inp[12]) ? 14'b00000011111111 : node1967;
												assign node1967 = (inp[9]) ? node1969 : 14'b00001111111111;
													assign node1969 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1973 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1976 = (inp[9]) ? node1986 : node1977;
											assign node1977 = (inp[6]) ? node1983 : node1978;
												assign node1978 = (inp[12]) ? 14'b00000001111111 : node1979;
													assign node1979 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1983 = (inp[5]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node1986 = (inp[5]) ? 14'b00000000011111 : node1987;
												assign node1987 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1991 = (inp[6]) ? node2007 : node1992;
										assign node1992 = (inp[2]) ? node1998 : node1993;
											assign node1993 = (inp[11]) ? 14'b00000000111111 : node1994;
												assign node1994 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1998 = (inp[5]) ? node2002 : node1999;
												assign node1999 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2002 = (inp[12]) ? 14'b00000000011111 : node2003;
													assign node2003 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2007 = (inp[12]) ? node2015 : node2008;
											assign node2008 = (inp[2]) ? 14'b00000000011111 : node2009;
												assign node2009 = (inp[9]) ? 14'b00000000111111 : node2010;
													assign node2010 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2015 = (inp[2]) ? node2017 : 14'b00000000011111;
												assign node2017 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2020 = (inp[9]) ? node2100 : node2021;
							assign node2021 = (inp[2]) ? node2053 : node2022;
								assign node2022 = (inp[3]) ? node2040 : node2023;
									assign node2023 = (inp[12]) ? node2029 : node2024;
										assign node2024 = (inp[5]) ? 14'b00000011111111 : node2025;
											assign node2025 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2029 = (inp[1]) ? node2035 : node2030;
											assign node2030 = (inp[7]) ? node2032 : 14'b00000111111111;
												assign node2032 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2035 = (inp[6]) ? 14'b00000001111111 : node2036;
												assign node2036 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2040 = (inp[6]) ? node2048 : node2041;
										assign node2041 = (inp[11]) ? 14'b00000001111111 : node2042;
											assign node2042 = (inp[12]) ? node2044 : 14'b00000011111111;
												assign node2044 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2048 = (inp[7]) ? node2050 : 14'b00000001111111;
											assign node2050 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2053 = (inp[12]) ? node2081 : node2054;
									assign node2054 = (inp[6]) ? node2070 : node2055;
										assign node2055 = (inp[7]) ? node2065 : node2056;
											assign node2056 = (inp[3]) ? node2058 : 14'b00000011111111;
												assign node2058 = (inp[11]) ? 14'b00000001111111 : node2059;
													assign node2059 = (inp[5]) ? node2061 : 14'b00000011111111;
														assign node2061 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2065 = (inp[1]) ? node2067 : 14'b00000011111111;
												assign node2067 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2070 = (inp[3]) ? node2076 : node2071;
											assign node2071 = (inp[11]) ? node2073 : 14'b00000011111111;
												assign node2073 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2076 = (inp[5]) ? node2078 : 14'b00000000111111;
												assign node2078 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2081 = (inp[3]) ? node2093 : node2082;
										assign node2082 = (inp[1]) ? 14'b00000000111111 : node2083;
											assign node2083 = (inp[5]) ? node2087 : node2084;
												assign node2084 = (inp[11]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node2087 = (inp[7]) ? node2089 : 14'b00000001111111;
													assign node2089 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2093 = (inp[6]) ? 14'b00000000001111 : node2094;
											assign node2094 = (inp[1]) ? 14'b00000000011111 : node2095;
												assign node2095 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2100 = (inp[1]) ? node2144 : node2101;
								assign node2101 = (inp[11]) ? node2127 : node2102;
									assign node2102 = (inp[7]) ? node2114 : node2103;
										assign node2103 = (inp[5]) ? node2105 : 14'b00000011111111;
											assign node2105 = (inp[3]) ? 14'b00000001111111 : node2106;
												assign node2106 = (inp[12]) ? 14'b00000001111111 : node2107;
													assign node2107 = (inp[2]) ? node2109 : 14'b00000011111111;
														assign node2109 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2114 = (inp[2]) ? node2124 : node2115;
											assign node2115 = (inp[5]) ? node2117 : 14'b00000011111111;
												assign node2117 = (inp[6]) ? node2119 : 14'b00000001111111;
													assign node2119 = (inp[3]) ? 14'b00000000111111 : node2120;
														assign node2120 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2124 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2127 = (inp[5]) ? node2137 : node2128;
										assign node2128 = (inp[6]) ? node2130 : 14'b00000001111111;
											assign node2130 = (inp[3]) ? 14'b00000000111111 : node2131;
												assign node2131 = (inp[12]) ? 14'b00000000111111 : node2132;
													assign node2132 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2137 = (inp[7]) ? node2139 : 14'b00000000111111;
											assign node2139 = (inp[3]) ? node2141 : 14'b00000000111111;
												assign node2141 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2144 = (inp[7]) ? node2178 : node2145;
									assign node2145 = (inp[12]) ? node2161 : node2146;
										assign node2146 = (inp[2]) ? 14'b00000000111111 : node2147;
											assign node2147 = (inp[3]) ? node2153 : node2148;
												assign node2148 = (inp[11]) ? 14'b00000001111111 : node2149;
													assign node2149 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2153 = (inp[5]) ? node2155 : 14'b00000001111111;
													assign node2155 = (inp[6]) ? node2157 : 14'b00000000111111;
														assign node2157 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2161 = (inp[5]) ? node2167 : node2162;
											assign node2162 = (inp[3]) ? 14'b00000000111111 : node2163;
												assign node2163 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2167 = (inp[6]) ? node2169 : 14'b00000000111111;
												assign node2169 = (inp[2]) ? node2175 : node2170;
													assign node2170 = (inp[11]) ? node2172 : 14'b00000000011111;
														assign node2172 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
													assign node2175 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node2178 = (inp[5]) ? node2188 : node2179;
										assign node2179 = (inp[2]) ? node2183 : node2180;
											assign node2180 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2183 = (inp[11]) ? node2185 : 14'b00000000011111;
												assign node2185 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2188 = (inp[2]) ? 14'b00000000000111 : node2189;
											assign node2189 = (inp[3]) ? node2195 : node2190;
												assign node2190 = (inp[6]) ? node2192 : 14'b00000000011111;
													assign node2192 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2195 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node2199 = (inp[8]) ? node2583 : node2200;
					assign node2200 = (inp[9]) ? node2404 : node2201;
						assign node2201 = (inp[12]) ? node2309 : node2202;
							assign node2202 = (inp[1]) ? node2250 : node2203;
								assign node2203 = (inp[3]) ? node2233 : node2204;
									assign node2204 = (inp[7]) ? node2220 : node2205;
										assign node2205 = (inp[0]) ? node2211 : node2206;
											assign node2206 = (inp[5]) ? 14'b00001111111111 : node2207;
												assign node2207 = (inp[6]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node2211 = (inp[11]) ? 14'b00000111111111 : node2212;
												assign node2212 = (inp[5]) ? node2214 : 14'b00001111111111;
													assign node2214 = (inp[2]) ? 14'b00000111111111 : node2215;
														assign node2215 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node2220 = (inp[11]) ? node2228 : node2221;
											assign node2221 = (inp[5]) ? node2225 : node2222;
												assign node2222 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2225 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2228 = (inp[5]) ? 14'b00000000111111 : node2229;
												assign node2229 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node2233 = (inp[6]) ? node2243 : node2234;
										assign node2234 = (inp[7]) ? node2238 : node2235;
											assign node2235 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2238 = (inp[0]) ? 14'b00000011111111 : node2239;
												assign node2239 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2243 = (inp[2]) ? node2245 : 14'b00000011111111;
											assign node2245 = (inp[5]) ? node2247 : 14'b00000011111111;
												assign node2247 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2250 = (inp[7]) ? node2284 : node2251;
									assign node2251 = (inp[11]) ? node2265 : node2252;
										assign node2252 = (inp[5]) ? node2258 : node2253;
											assign node2253 = (inp[0]) ? node2255 : 14'b00001111111111;
												assign node2255 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2258 = (inp[0]) ? 14'b00000001111111 : node2259;
												assign node2259 = (inp[2]) ? 14'b00000011111111 : node2260;
													assign node2260 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2265 = (inp[2]) ? node2275 : node2266;
											assign node2266 = (inp[0]) ? node2272 : node2267;
												assign node2267 = (inp[6]) ? 14'b00000011111111 : node2268;
													assign node2268 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2272 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2275 = (inp[6]) ? node2281 : node2276;
												assign node2276 = (inp[3]) ? node2278 : 14'b00000011111111;
													assign node2278 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2281 = (inp[5]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node2284 = (inp[2]) ? node2296 : node2285;
										assign node2285 = (inp[3]) ? node2293 : node2286;
											assign node2286 = (inp[0]) ? 14'b00000011111111 : node2287;
												assign node2287 = (inp[11]) ? node2289 : 14'b00000111111111;
													assign node2289 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2293 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2296 = (inp[11]) ? node2298 : 14'b00000001111111;
											assign node2298 = (inp[3]) ? node2306 : node2299;
												assign node2299 = (inp[5]) ? node2301 : 14'b00000001111111;
													assign node2301 = (inp[0]) ? 14'b00000000111111 : node2302;
														assign node2302 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2306 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2309 = (inp[5]) ? node2353 : node2310;
								assign node2310 = (inp[6]) ? node2332 : node2311;
									assign node2311 = (inp[0]) ? node2321 : node2312;
										assign node2312 = (inp[7]) ? node2318 : node2313;
											assign node2313 = (inp[2]) ? node2315 : 14'b00001111111111;
												assign node2315 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2318 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2321 = (inp[3]) ? node2329 : node2322;
											assign node2322 = (inp[1]) ? node2326 : node2323;
												assign node2323 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2326 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2329 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2332 = (inp[1]) ? node2342 : node2333;
										assign node2333 = (inp[7]) ? node2337 : node2334;
											assign node2334 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2337 = (inp[3]) ? 14'b00000001111111 : node2338;
												assign node2338 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2342 = (inp[0]) ? node2346 : node2343;
											assign node2343 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2346 = (inp[11]) ? 14'b00000000011111 : node2347;
												assign node2347 = (inp[3]) ? 14'b00000000111111 : node2348;
													assign node2348 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2353 = (inp[1]) ? node2377 : node2354;
									assign node2354 = (inp[2]) ? node2366 : node2355;
										assign node2355 = (inp[11]) ? node2361 : node2356;
											assign node2356 = (inp[0]) ? node2358 : 14'b00000111111111;
												assign node2358 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2361 = (inp[3]) ? 14'b00000001111111 : node2362;
												assign node2362 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2366 = (inp[0]) ? node2372 : node2367;
											assign node2367 = (inp[7]) ? node2369 : 14'b00000011111111;
												assign node2369 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2372 = (inp[11]) ? node2374 : 14'b00000000111111;
												assign node2374 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2377 = (inp[3]) ? node2387 : node2378;
										assign node2378 = (inp[2]) ? node2384 : node2379;
											assign node2379 = (inp[7]) ? node2381 : 14'b00000011111111;
												assign node2381 = (inp[11]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node2384 = (inp[0]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node2387 = (inp[0]) ? node2389 : 14'b00000000111111;
											assign node2389 = (inp[11]) ? node2393 : node2390;
												assign node2390 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2393 = (inp[7]) ? node2399 : node2394;
													assign node2394 = (inp[6]) ? node2396 : 14'b00000000011111;
														assign node2396 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
													assign node2399 = (inp[2]) ? 14'b00000000001111 : node2400;
														assign node2400 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2404 = (inp[11]) ? node2498 : node2405;
							assign node2405 = (inp[2]) ? node2455 : node2406;
								assign node2406 = (inp[5]) ? node2428 : node2407;
									assign node2407 = (inp[1]) ? node2417 : node2408;
										assign node2408 = (inp[3]) ? node2410 : 14'b00000111111111;
											assign node2410 = (inp[6]) ? node2414 : node2411;
												assign node2411 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2414 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2417 = (inp[6]) ? node2419 : 14'b00000011111111;
											assign node2419 = (inp[0]) ? node2425 : node2420;
												assign node2420 = (inp[3]) ? 14'b00000001111111 : node2421;
													assign node2421 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2425 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2428 = (inp[7]) ? node2446 : node2429;
										assign node2429 = (inp[12]) ? node2433 : node2430;
											assign node2430 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node2433 = (inp[1]) ? node2441 : node2434;
												assign node2434 = (inp[3]) ? node2436 : 14'b00000001111111;
													assign node2436 = (inp[6]) ? node2438 : 14'b00000001111111;
														assign node2438 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2441 = (inp[0]) ? 14'b00000001111111 : node2442;
													assign node2442 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2446 = (inp[6]) ? 14'b00000000111111 : node2447;
											assign node2447 = (inp[1]) ? node2451 : node2448;
												assign node2448 = (inp[12]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node2451 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2455 = (inp[3]) ? node2477 : node2456;
									assign node2456 = (inp[12]) ? node2466 : node2457;
										assign node2457 = (inp[1]) ? 14'b00000001111111 : node2458;
											assign node2458 = (inp[0]) ? node2462 : node2459;
												assign node2459 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2462 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2466 = (inp[6]) ? node2470 : node2467;
											assign node2467 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2470 = (inp[0]) ? node2474 : node2471;
												assign node2471 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2474 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2477 = (inp[6]) ? node2489 : node2478;
										assign node2478 = (inp[12]) ? node2486 : node2479;
											assign node2479 = (inp[0]) ? node2483 : node2480;
												assign node2480 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2483 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2486 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2489 = (inp[5]) ? node2495 : node2490;
											assign node2490 = (inp[7]) ? node2492 : 14'b00000000111111;
												assign node2492 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2495 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2498 = (inp[6]) ? node2540 : node2499;
								assign node2499 = (inp[3]) ? node2513 : node2500;
									assign node2500 = (inp[2]) ? node2508 : node2501;
										assign node2501 = (inp[5]) ? 14'b00000001111111 : node2502;
											assign node2502 = (inp[0]) ? 14'b00000011111111 : node2503;
												assign node2503 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2508 = (inp[0]) ? 14'b00000000111111 : node2509;
											assign node2509 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2513 = (inp[12]) ? node2529 : node2514;
										assign node2514 = (inp[1]) ? node2522 : node2515;
											assign node2515 = (inp[0]) ? node2519 : node2516;
												assign node2516 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2519 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2522 = (inp[5]) ? 14'b00000000111111 : node2523;
												assign node2523 = (inp[0]) ? 14'b00000000111111 : node2524;
													assign node2524 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2529 = (inp[0]) ? node2535 : node2530;
											assign node2530 = (inp[5]) ? node2532 : 14'b00000001111111;
												assign node2532 = (inp[7]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node2535 = (inp[5]) ? node2537 : 14'b00000000011111;
												assign node2537 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2540 = (inp[1]) ? node2566 : node2541;
									assign node2541 = (inp[0]) ? node2557 : node2542;
										assign node2542 = (inp[5]) ? node2550 : node2543;
											assign node2543 = (inp[2]) ? node2547 : node2544;
												assign node2544 = (inp[7]) ? 14'b00000011111111 : 14'b00000001111111;
												assign node2547 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2550 = (inp[3]) ? node2552 : 14'b00000000111111;
												assign node2552 = (inp[12]) ? node2554 : 14'b00000000111111;
													assign node2554 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2557 = (inp[5]) ? 14'b00000000011111 : node2558;
											assign node2558 = (inp[7]) ? node2560 : 14'b00000000111111;
												assign node2560 = (inp[2]) ? node2562 : 14'b00000000111111;
													assign node2562 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2566 = (inp[12]) ? node2574 : node2567;
										assign node2567 = (inp[2]) ? 14'b00000000011111 : node2568;
											assign node2568 = (inp[3]) ? 14'b00000000111111 : node2569;
												assign node2569 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2574 = (inp[3]) ? 14'b00000000001111 : node2575;
											assign node2575 = (inp[7]) ? node2579 : node2576;
												assign node2576 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2579 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node2583 = (inp[7]) ? node2771 : node2584;
						assign node2584 = (inp[2]) ? node2668 : node2585;
							assign node2585 = (inp[11]) ? node2627 : node2586;
								assign node2586 = (inp[5]) ? node2612 : node2587;
									assign node2587 = (inp[1]) ? node2601 : node2588;
										assign node2588 = (inp[9]) ? node2590 : 14'b00000111111111;
											assign node2590 = (inp[6]) ? 14'b00000011111111 : node2591;
												assign node2591 = (inp[0]) ? node2597 : node2592;
													assign node2592 = (inp[12]) ? 14'b00000111111111 : node2593;
														assign node2593 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
													assign node2597 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2601 = (inp[0]) ? node2607 : node2602;
											assign node2602 = (inp[9]) ? node2604 : 14'b00000011111111;
												assign node2604 = (inp[3]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node2607 = (inp[12]) ? node2609 : 14'b00000011111111;
												assign node2609 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2612 = (inp[6]) ? node2622 : node2613;
										assign node2613 = (inp[0]) ? 14'b00000001111111 : node2614;
											assign node2614 = (inp[3]) ? node2616 : 14'b00000011111111;
												assign node2616 = (inp[1]) ? 14'b00000001111111 : node2617;
													assign node2617 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2622 = (inp[3]) ? node2624 : 14'b00000001111111;
											assign node2624 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2627 = (inp[3]) ? node2655 : node2628;
									assign node2628 = (inp[12]) ? node2642 : node2629;
										assign node2629 = (inp[1]) ? node2633 : node2630;
											assign node2630 = (inp[6]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node2633 = (inp[6]) ? node2637 : node2634;
												assign node2634 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2637 = (inp[9]) ? node2639 : 14'b00000001111111;
													assign node2639 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2642 = (inp[0]) ? node2650 : node2643;
											assign node2643 = (inp[9]) ? node2645 : 14'b00000001111111;
												assign node2645 = (inp[1]) ? node2647 : 14'b00000001111111;
													assign node2647 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2650 = (inp[9]) ? 14'b00000000011111 : node2651;
												assign node2651 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2655 = (inp[5]) ? node2661 : node2656;
										assign node2656 = (inp[6]) ? 14'b00000000111111 : node2657;
											assign node2657 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2661 = (inp[0]) ? node2663 : 14'b00000000111111;
											assign node2663 = (inp[6]) ? node2665 : 14'b00000000011111;
												assign node2665 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2668 = (inp[6]) ? node2728 : node2669;
								assign node2669 = (inp[1]) ? node2701 : node2670;
									assign node2670 = (inp[5]) ? node2686 : node2671;
										assign node2671 = (inp[0]) ? node2679 : node2672;
											assign node2672 = (inp[3]) ? node2676 : node2673;
												assign node2673 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2676 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2679 = (inp[12]) ? node2683 : node2680;
												assign node2680 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2683 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2686 = (inp[9]) ? node2694 : node2687;
											assign node2687 = (inp[3]) ? node2689 : 14'b00000001111111;
												assign node2689 = (inp[12]) ? node2691 : 14'b00000001111111;
													assign node2691 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2694 = (inp[3]) ? 14'b00000000111111 : node2695;
												assign node2695 = (inp[0]) ? 14'b00000000111111 : node2696;
													assign node2696 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2701 = (inp[3]) ? node2719 : node2702;
										assign node2702 = (inp[12]) ? node2706 : node2703;
											assign node2703 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2706 = (inp[0]) ? node2712 : node2707;
												assign node2707 = (inp[9]) ? node2709 : 14'b00000001111111;
													assign node2709 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2712 = (inp[9]) ? 14'b00000000011111 : node2713;
													assign node2713 = (inp[11]) ? 14'b00000000111111 : node2714;
														assign node2714 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2719 = (inp[0]) ? node2725 : node2720;
											assign node2720 = (inp[5]) ? node2722 : 14'b00000000111111;
												assign node2722 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2725 = (inp[5]) ? 14'b00000000001111 : 14'b00000001111111;
								assign node2728 = (inp[3]) ? node2744 : node2729;
									assign node2729 = (inp[5]) ? node2739 : node2730;
										assign node2730 = (inp[12]) ? node2732 : 14'b00000001111111;
											assign node2732 = (inp[1]) ? 14'b00000000111111 : node2733;
												assign node2733 = (inp[9]) ? 14'b00000000111111 : node2734;
													assign node2734 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2739 = (inp[11]) ? 14'b00000000011111 : node2740;
											assign node2740 = (inp[1]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node2744 = (inp[0]) ? node2762 : node2745;
										assign node2745 = (inp[9]) ? node2755 : node2746;
											assign node2746 = (inp[11]) ? node2752 : node2747;
												assign node2747 = (inp[5]) ? 14'b00000000111111 : node2748;
													assign node2748 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2752 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2755 = (inp[12]) ? node2759 : node2756;
												assign node2756 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2759 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2762 = (inp[11]) ? node2766 : node2763;
											assign node2763 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2766 = (inp[9]) ? 14'b00000000000111 : node2767;
												assign node2767 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2771 = (inp[3]) ? node2857 : node2772;
							assign node2772 = (inp[1]) ? node2812 : node2773;
								assign node2773 = (inp[2]) ? node2795 : node2774;
									assign node2774 = (inp[5]) ? node2788 : node2775;
										assign node2775 = (inp[12]) ? node2781 : node2776;
											assign node2776 = (inp[9]) ? node2778 : 14'b00000111111111;
												assign node2778 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2781 = (inp[0]) ? node2785 : node2782;
												assign node2782 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2785 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2788 = (inp[12]) ? 14'b00000000111111 : node2789;
											assign node2789 = (inp[11]) ? node2791 : 14'b00000001111111;
												assign node2791 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2795 = (inp[6]) ? node2805 : node2796;
										assign node2796 = (inp[9]) ? node2798 : 14'b00000001111111;
											assign node2798 = (inp[11]) ? node2800 : 14'b00000001111111;
												assign node2800 = (inp[5]) ? node2802 : 14'b00000000111111;
													assign node2802 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2805 = (inp[5]) ? node2809 : node2806;
											assign node2806 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2809 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2812 = (inp[11]) ? node2842 : node2813;
									assign node2813 = (inp[6]) ? node2821 : node2814;
										assign node2814 = (inp[9]) ? node2818 : node2815;
											assign node2815 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2818 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2821 = (inp[2]) ? node2833 : node2822;
											assign node2822 = (inp[12]) ? node2826 : node2823;
												assign node2823 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2826 = (inp[9]) ? node2828 : 14'b00000000111111;
													assign node2828 = (inp[0]) ? 14'b00000000011111 : node2829;
														assign node2829 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2833 = (inp[9]) ? 14'b00000000001111 : node2834;
												assign node2834 = (inp[0]) ? node2836 : 14'b00000000111111;
													assign node2836 = (inp[12]) ? node2838 : 14'b00000000011111;
														assign node2838 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2842 = (inp[9]) ? node2852 : node2843;
										assign node2843 = (inp[5]) ? node2847 : node2844;
											assign node2844 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2847 = (inp[6]) ? 14'b00000000011111 : node2848;
												assign node2848 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2852 = (inp[5]) ? 14'b00000000000111 : node2853;
											assign node2853 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2857 = (inp[9]) ? node2923 : node2858;
								assign node2858 = (inp[11]) ? node2892 : node2859;
									assign node2859 = (inp[2]) ? node2875 : node2860;
										assign node2860 = (inp[0]) ? node2866 : node2861;
											assign node2861 = (inp[5]) ? node2863 : 14'b00000001111111;
												assign node2863 = (inp[6]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node2866 = (inp[1]) ? 14'b00000000111111 : node2867;
												assign node2867 = (inp[5]) ? 14'b00000000111111 : node2868;
													assign node2868 = (inp[6]) ? node2870 : 14'b00000001111111;
														assign node2870 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2875 = (inp[12]) ? node2885 : node2876;
											assign node2876 = (inp[0]) ? 14'b00000000011111 : node2877;
												assign node2877 = (inp[6]) ? node2879 : 14'b00000001111111;
													assign node2879 = (inp[5]) ? 14'b00000000111111 : node2880;
														assign node2880 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2885 = (inp[0]) ? node2887 : 14'b00000000011111;
												assign node2887 = (inp[1]) ? node2889 : 14'b00000000001111;
													assign node2889 = (inp[5]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node2892 = (inp[1]) ? node2906 : node2893;
										assign node2893 = (inp[0]) ? node2899 : node2894;
											assign node2894 = (inp[12]) ? node2896 : 14'b00000001111111;
												assign node2896 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2899 = (inp[6]) ? node2903 : node2900;
												assign node2900 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2903 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2906 = (inp[12]) ? node2914 : node2907;
											assign node2907 = (inp[6]) ? node2909 : 14'b00000000011111;
												assign node2909 = (inp[0]) ? 14'b00000000001111 : node2910;
													assign node2910 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2914 = (inp[2]) ? node2920 : node2915;
												assign node2915 = (inp[5]) ? 14'b00000000001111 : node2916;
													assign node2916 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2920 = (inp[5]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node2923 = (inp[2]) ? node2955 : node2924;
									assign node2924 = (inp[11]) ? node2940 : node2925;
										assign node2925 = (inp[5]) ? node2935 : node2926;
											assign node2926 = (inp[0]) ? node2930 : node2927;
												assign node2927 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2930 = (inp[6]) ? 14'b00000000011111 : node2931;
													assign node2931 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2935 = (inp[12]) ? 14'b00000000001111 : node2936;
												assign node2936 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2940 = (inp[0]) ? node2950 : node2941;
											assign node2941 = (inp[12]) ? node2945 : node2942;
												assign node2942 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2945 = (inp[1]) ? 14'b00000000001111 : node2946;
													assign node2946 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2950 = (inp[1]) ? node2952 : 14'b00000000001111;
												assign node2952 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node2955 = (inp[6]) ? node2967 : node2956;
										assign node2956 = (inp[11]) ? node2962 : node2957;
											assign node2957 = (inp[1]) ? node2959 : 14'b00000000011111;
												assign node2959 = (inp[12]) ? 14'b00000000011111 : 14'b00000000001111;
											assign node2962 = (inp[5]) ? 14'b00000000001111 : node2963;
												assign node2963 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2967 = (inp[0]) ? node2977 : node2968;
											assign node2968 = (inp[12]) ? node2972 : node2969;
												assign node2969 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2972 = (inp[1]) ? node2974 : 14'b00000000001111;
													assign node2974 = (inp[5]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node2977 = (inp[5]) ? 14'b00000000000111 : node2978;
												assign node2978 = (inp[1]) ? node2980 : 14'b00000000001111;
													assign node2980 = (inp[12]) ? 14'b00000000000011 : 14'b00000000001111;
		assign node2984 = (inp[10]) ? node4576 : node2985;
			assign node2985 = (inp[12]) ? node3807 : node2986;
				assign node2986 = (inp[9]) ? node3406 : node2987;
					assign node2987 = (inp[6]) ? node3189 : node2988;
						assign node2988 = (inp[0]) ? node3098 : node2989;
							assign node2989 = (inp[3]) ? node3049 : node2990;
								assign node2990 = (inp[13]) ? node3016 : node2991;
									assign node2991 = (inp[8]) ? node3005 : node2992;
										assign node2992 = (inp[2]) ? node2998 : node2993;
											assign node2993 = (inp[1]) ? 14'b00001111111111 : node2994;
												assign node2994 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node2998 = (inp[11]) ? node3000 : 14'b00011111111111;
												assign node3000 = (inp[5]) ? 14'b00001111111111 : node3001;
													assign node3001 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node3005 = (inp[1]) ? node3011 : node3006;
											assign node3006 = (inp[2]) ? node3008 : 14'b00011111111111;
												assign node3008 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3011 = (inp[2]) ? 14'b00000111111111 : node3012;
												assign node3012 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node3016 = (inp[2]) ? node3032 : node3017;
										assign node3017 = (inp[5]) ? node3027 : node3018;
											assign node3018 = (inp[11]) ? node3022 : node3019;
												assign node3019 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3022 = (inp[7]) ? 14'b00000111111111 : node3023;
													assign node3023 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3027 = (inp[1]) ? 14'b00000111111111 : node3028;
												assign node3028 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3032 = (inp[1]) ? node3040 : node3033;
											assign node3033 = (inp[5]) ? node3037 : node3034;
												assign node3034 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3037 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3040 = (inp[8]) ? node3042 : 14'b00000011111111;
												assign node3042 = (inp[5]) ? 14'b00000001111111 : node3043;
													assign node3043 = (inp[11]) ? node3045 : 14'b00000011111111;
														assign node3045 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node3049 = (inp[2]) ? node3067 : node3050;
									assign node3050 = (inp[1]) ? node3064 : node3051;
										assign node3051 = (inp[8]) ? node3055 : node3052;
											assign node3052 = (inp[11]) ? 14'b00001111111111 : 14'b00000111111111;
											assign node3055 = (inp[5]) ? node3059 : node3056;
												assign node3056 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3059 = (inp[13]) ? 14'b00000011111111 : node3060;
													assign node3060 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3064 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node3067 = (inp[7]) ? node3081 : node3068;
										assign node3068 = (inp[8]) ? node3074 : node3069;
											assign node3069 = (inp[11]) ? 14'b00000111111111 : node3070;
												assign node3070 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node3074 = (inp[13]) ? 14'b00000001111111 : node3075;
												assign node3075 = (inp[1]) ? 14'b00000011111111 : node3076;
													assign node3076 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3081 = (inp[5]) ? node3091 : node3082;
											assign node3082 = (inp[13]) ? node3088 : node3083;
												assign node3083 = (inp[1]) ? 14'b00000011111111 : node3084;
													assign node3084 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3088 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3091 = (inp[13]) ? node3095 : node3092;
												assign node3092 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3095 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
							assign node3098 = (inp[8]) ? node3146 : node3099;
								assign node3099 = (inp[13]) ? node3121 : node3100;
									assign node3100 = (inp[1]) ? node3110 : node3101;
										assign node3101 = (inp[3]) ? node3107 : node3102;
											assign node3102 = (inp[7]) ? node3104 : 14'b00001111111111;
												assign node3104 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3107 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3110 = (inp[5]) ? node3116 : node3111;
											assign node3111 = (inp[3]) ? 14'b00000111111111 : node3112;
												assign node3112 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3116 = (inp[7]) ? node3118 : 14'b00000111111111;
												assign node3118 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node3121 = (inp[11]) ? node3133 : node3122;
										assign node3122 = (inp[5]) ? node3128 : node3123;
											assign node3123 = (inp[7]) ? 14'b00000111111111 : node3124;
												assign node3124 = (inp[1]) ? 14'b00000111111111 : 14'b00011111111111;
											assign node3128 = (inp[2]) ? 14'b00000011111111 : node3129;
												assign node3129 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3133 = (inp[3]) ? node3143 : node3134;
											assign node3134 = (inp[1]) ? node3140 : node3135;
												assign node3135 = (inp[5]) ? 14'b00000011111111 : node3136;
													assign node3136 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3140 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3143 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node3146 = (inp[5]) ? node3178 : node3147;
									assign node3147 = (inp[7]) ? node3165 : node3148;
										assign node3148 = (inp[1]) ? node3156 : node3149;
											assign node3149 = (inp[3]) ? 14'b00000011111111 : node3150;
												assign node3150 = (inp[11]) ? 14'b00000011111111 : node3151;
													assign node3151 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3156 = (inp[2]) ? node3158 : 14'b00000011111111;
												assign node3158 = (inp[13]) ? node3160 : 14'b00000011111111;
													assign node3160 = (inp[11]) ? 14'b00000001111111 : node3161;
														assign node3161 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3165 = (inp[11]) ? node3173 : node3166;
											assign node3166 = (inp[2]) ? node3168 : 14'b00000011111111;
												assign node3168 = (inp[13]) ? node3170 : 14'b00000011111111;
													assign node3170 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3173 = (inp[2]) ? 14'b00000001111111 : node3174;
												assign node3174 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3178 = (inp[2]) ? node3182 : node3179;
										assign node3179 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3182 = (inp[11]) ? node3184 : 14'b00000001111111;
											assign node3184 = (inp[13]) ? 14'b00000000111111 : node3185;
												assign node3185 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node3189 = (inp[7]) ? node3315 : node3190;
							assign node3190 = (inp[0]) ? node3256 : node3191;
								assign node3191 = (inp[11]) ? node3219 : node3192;
									assign node3192 = (inp[8]) ? node3206 : node3193;
										assign node3193 = (inp[1]) ? node3195 : 14'b00001111111111;
											assign node3195 = (inp[2]) ? node3203 : node3196;
												assign node3196 = (inp[13]) ? node3198 : 14'b00001111111111;
													assign node3198 = (inp[3]) ? 14'b00000111111111 : node3199;
														assign node3199 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3203 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3206 = (inp[13]) ? node3214 : node3207;
											assign node3207 = (inp[1]) ? 14'b00000011111111 : node3208;
												assign node3208 = (inp[3]) ? 14'b00000111111111 : node3209;
													assign node3209 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3214 = (inp[5]) ? 14'b00000011111111 : node3215;
												assign node3215 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node3219 = (inp[2]) ? node3241 : node3220;
										assign node3220 = (inp[5]) ? node3232 : node3221;
											assign node3221 = (inp[3]) ? node3229 : node3222;
												assign node3222 = (inp[1]) ? 14'b00000111111111 : node3223;
													assign node3223 = (inp[13]) ? node3225 : 14'b00001111111111;
														assign node3225 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3229 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3232 = (inp[1]) ? node3238 : node3233;
												assign node3233 = (inp[13]) ? 14'b00000011111111 : node3234;
													assign node3234 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3238 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3241 = (inp[3]) ? 14'b00000001111111 : node3242;
											assign node3242 = (inp[8]) ? node3244 : 14'b00000011111111;
												assign node3244 = (inp[5]) ? node3250 : node3245;
													assign node3245 = (inp[13]) ? node3247 : 14'b00000011111111;
														assign node3247 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
													assign node3250 = (inp[1]) ? node3252 : 14'b00000001111111;
														assign node3252 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node3256 = (inp[5]) ? node3288 : node3257;
									assign node3257 = (inp[8]) ? node3273 : node3258;
										assign node3258 = (inp[13]) ? node3266 : node3259;
											assign node3259 = (inp[11]) ? node3263 : node3260;
												assign node3260 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3263 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3266 = (inp[11]) ? node3270 : node3267;
												assign node3267 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3270 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3273 = (inp[13]) ? node3281 : node3274;
											assign node3274 = (inp[1]) ? node3278 : node3275;
												assign node3275 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3278 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3281 = (inp[11]) ? node3285 : node3282;
												assign node3282 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3285 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3288 = (inp[11]) ? node3306 : node3289;
										assign node3289 = (inp[3]) ? node3295 : node3290;
											assign node3290 = (inp[13]) ? 14'b00000011111111 : node3291;
												assign node3291 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3295 = (inp[2]) ? 14'b00000000111111 : node3296;
												assign node3296 = (inp[1]) ? node3302 : node3297;
													assign node3297 = (inp[13]) ? node3299 : 14'b00000011111111;
														assign node3299 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
													assign node3302 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3306 = (inp[13]) ? node3312 : node3307;
											assign node3307 = (inp[8]) ? node3309 : 14'b00000001111111;
												assign node3309 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3312 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node3315 = (inp[13]) ? node3349 : node3316;
								assign node3316 = (inp[11]) ? node3330 : node3317;
									assign node3317 = (inp[5]) ? node3319 : 14'b00000011111111;
										assign node3319 = (inp[0]) ? node3323 : node3320;
											assign node3320 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3323 = (inp[3]) ? 14'b00000001111111 : node3324;
												assign node3324 = (inp[1]) ? node3326 : 14'b00000111111111;
													assign node3326 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3330 = (inp[2]) ? node3346 : node3331;
										assign node3331 = (inp[0]) ? node3341 : node3332;
											assign node3332 = (inp[5]) ? node3334 : 14'b00000111111111;
												assign node3334 = (inp[1]) ? 14'b00000001111111 : node3335;
													assign node3335 = (inp[3]) ? node3337 : 14'b00000011111111;
														assign node3337 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3341 = (inp[1]) ? 14'b00000001111111 : node3342;
												assign node3342 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3346 = (inp[1]) ? 14'b00000000111111 : 14'b00000000011111;
								assign node3349 = (inp[1]) ? node3381 : node3350;
									assign node3350 = (inp[0]) ? node3366 : node3351;
										assign node3351 = (inp[8]) ? node3361 : node3352;
											assign node3352 = (inp[5]) ? 14'b00000001111111 : node3353;
												assign node3353 = (inp[3]) ? 14'b00000011111111 : node3354;
													assign node3354 = (inp[11]) ? node3356 : 14'b00000111111111;
														assign node3356 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3361 = (inp[5]) ? 14'b00000001111111 : node3362;
												assign node3362 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3366 = (inp[11]) ? node3378 : node3367;
											assign node3367 = (inp[5]) ? node3375 : node3368;
												assign node3368 = (inp[3]) ? 14'b00000001111111 : node3369;
													assign node3369 = (inp[2]) ? node3371 : 14'b00000011111111;
														assign node3371 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3375 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3378 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3381 = (inp[5]) ? node3393 : node3382;
										assign node3382 = (inp[0]) ? node3386 : node3383;
											assign node3383 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3386 = (inp[3]) ? node3388 : 14'b00000000111111;
												assign node3388 = (inp[2]) ? node3390 : 14'b00000000111111;
													assign node3390 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3393 = (inp[8]) ? node3397 : node3394;
											assign node3394 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node3397 = (inp[0]) ? node3401 : node3398;
												assign node3398 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3401 = (inp[11]) ? 14'b00000000001111 : node3402;
													assign node3402 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node3406 = (inp[2]) ? node3582 : node3407;
						assign node3407 = (inp[13]) ? node3503 : node3408;
							assign node3408 = (inp[5]) ? node3456 : node3409;
								assign node3409 = (inp[1]) ? node3437 : node3410;
									assign node3410 = (inp[7]) ? node3428 : node3411;
										assign node3411 = (inp[0]) ? node3417 : node3412;
											assign node3412 = (inp[8]) ? 14'b00001111111111 : node3413;
												assign node3413 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node3417 = (inp[6]) ? node3423 : node3418;
												assign node3418 = (inp[11]) ? 14'b00001111111111 : node3419;
													assign node3419 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3423 = (inp[11]) ? 14'b00000111111111 : node3424;
													assign node3424 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3428 = (inp[0]) ? node3432 : node3429;
											assign node3429 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3432 = (inp[6]) ? node3434 : 14'b00000111111111;
												assign node3434 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3437 = (inp[3]) ? node3449 : node3438;
										assign node3438 = (inp[0]) ? node3444 : node3439;
											assign node3439 = (inp[7]) ? node3441 : 14'b00000111111111;
												assign node3441 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3444 = (inp[7]) ? node3446 : 14'b00000011111111;
												assign node3446 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3449 = (inp[8]) ? node3451 : 14'b00000011111111;
											assign node3451 = (inp[7]) ? 14'b00000000111111 : node3452;
												assign node3452 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node3456 = (inp[0]) ? node3478 : node3457;
									assign node3457 = (inp[7]) ? node3469 : node3458;
										assign node3458 = (inp[6]) ? node3466 : node3459;
											assign node3459 = (inp[8]) ? 14'b00000111111111 : node3460;
												assign node3460 = (inp[1]) ? node3462 : 14'b00001111111111;
													assign node3462 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3466 = (inp[11]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node3469 = (inp[8]) ? node3475 : node3470;
											assign node3470 = (inp[1]) ? node3472 : 14'b00000011111111;
												assign node3472 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3475 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3478 = (inp[7]) ? node3492 : node3479;
										assign node3479 = (inp[3]) ? node3483 : node3480;
											assign node3480 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3483 = (inp[1]) ? node3485 : 14'b00000111111111;
												assign node3485 = (inp[8]) ? node3487 : 14'b00000001111111;
													assign node3487 = (inp[11]) ? 14'b00000000111111 : node3488;
														assign node3488 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3492 = (inp[11]) ? node3494 : 14'b00000001111111;
											assign node3494 = (inp[3]) ? 14'b00000000011111 : node3495;
												assign node3495 = (inp[1]) ? 14'b00000000111111 : node3496;
													assign node3496 = (inp[8]) ? node3498 : 14'b00000001111111;
														assign node3498 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node3503 = (inp[8]) ? node3545 : node3504;
								assign node3504 = (inp[6]) ? node3526 : node3505;
									assign node3505 = (inp[11]) ? node3517 : node3506;
										assign node3506 = (inp[5]) ? node3508 : 14'b00000111111111;
											assign node3508 = (inp[3]) ? node3514 : node3509;
												assign node3509 = (inp[7]) ? node3511 : 14'b00000111111111;
													assign node3511 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3514 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3517 = (inp[3]) ? 14'b00000001111111 : node3518;
											assign node3518 = (inp[7]) ? node3522 : node3519;
												assign node3519 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3522 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3526 = (inp[0]) ? node3534 : node3527;
										assign node3527 = (inp[11]) ? node3529 : 14'b00000011111111;
											assign node3529 = (inp[5]) ? 14'b00000001111111 : node3530;
												assign node3530 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3534 = (inp[7]) ? node3540 : node3535;
											assign node3535 = (inp[3]) ? node3537 : 14'b00000001111111;
												assign node3537 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3540 = (inp[1]) ? node3542 : 14'b00000011111111;
												assign node3542 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3545 = (inp[7]) ? node3567 : node3546;
									assign node3546 = (inp[11]) ? node3552 : node3547;
										assign node3547 = (inp[0]) ? 14'b00000001111111 : node3548;
											assign node3548 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3552 = (inp[0]) ? node3558 : node3553;
											assign node3553 = (inp[6]) ? 14'b00000000111111 : node3554;
												assign node3554 = (inp[1]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node3558 = (inp[5]) ? node3562 : node3559;
												assign node3559 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3562 = (inp[1]) ? node3564 : 14'b00000000111111;
													assign node3564 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3567 = (inp[6]) ? node3577 : node3568;
										assign node3568 = (inp[0]) ? node3574 : node3569;
											assign node3569 = (inp[5]) ? node3571 : 14'b00000001111111;
												assign node3571 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3574 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3577 = (inp[5]) ? node3579 : 14'b00000000011111;
											assign node3579 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node3582 = (inp[6]) ? node3700 : node3583;
							assign node3583 = (inp[13]) ? node3651 : node3584;
								assign node3584 = (inp[7]) ? node3616 : node3585;
									assign node3585 = (inp[0]) ? node3605 : node3586;
										assign node3586 = (inp[1]) ? node3596 : node3587;
											assign node3587 = (inp[11]) ? node3589 : 14'b00011111111111;
												assign node3589 = (inp[3]) ? 14'b00000111111111 : node3590;
													assign node3590 = (inp[8]) ? 14'b00000111111111 : node3591;
														assign node3591 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3596 = (inp[5]) ? node3598 : 14'b00000111111111;
												assign node3598 = (inp[11]) ? node3600 : 14'b00000011111111;
													assign node3600 = (inp[8]) ? 14'b00000001111111 : node3601;
														assign node3601 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3605 = (inp[3]) ? node3611 : node3606;
											assign node3606 = (inp[5]) ? 14'b00000011111111 : node3607;
												assign node3607 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3611 = (inp[5]) ? node3613 : 14'b00000001111111;
												assign node3613 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3616 = (inp[5]) ? node3634 : node3617;
										assign node3617 = (inp[11]) ? node3629 : node3618;
											assign node3618 = (inp[0]) ? node3622 : node3619;
												assign node3619 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3622 = (inp[1]) ? node3624 : 14'b00000011111111;
													assign node3624 = (inp[3]) ? 14'b00000001111111 : node3625;
														assign node3625 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3629 = (inp[0]) ? node3631 : 14'b00000001111111;
												assign node3631 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3634 = (inp[8]) ? node3644 : node3635;
											assign node3635 = (inp[1]) ? node3639 : node3636;
												assign node3636 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3639 = (inp[0]) ? node3641 : 14'b00000001111111;
													assign node3641 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3644 = (inp[1]) ? node3648 : node3645;
												assign node3645 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3648 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3651 = (inp[1]) ? node3677 : node3652;
									assign node3652 = (inp[8]) ? node3668 : node3653;
										assign node3653 = (inp[3]) ? node3661 : node3654;
											assign node3654 = (inp[11]) ? 14'b00000001111111 : node3655;
												assign node3655 = (inp[5]) ? node3657 : 14'b00000011111111;
													assign node3657 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3661 = (inp[11]) ? node3663 : 14'b00000001111111;
												assign node3663 = (inp[7]) ? node3665 : 14'b00000001111111;
													assign node3665 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3668 = (inp[0]) ? node3672 : node3669;
											assign node3669 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3672 = (inp[11]) ? node3674 : 14'b00000000111111;
												assign node3674 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3677 = (inp[5]) ? node3685 : node3678;
										assign node3678 = (inp[0]) ? node3680 : 14'b00000001111111;
											assign node3680 = (inp[8]) ? 14'b00000000111111 : node3681;
												assign node3681 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3685 = (inp[8]) ? node3695 : node3686;
											assign node3686 = (inp[11]) ? node3692 : node3687;
												assign node3687 = (inp[3]) ? 14'b00000000111111 : node3688;
													assign node3688 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3692 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node3695 = (inp[7]) ? node3697 : 14'b00000000011111;
												assign node3697 = (inp[0]) ? 14'b00000000000111 : 14'b00000000011111;
							assign node3700 = (inp[5]) ? node3748 : node3701;
								assign node3701 = (inp[1]) ? node3723 : node3702;
									assign node3702 = (inp[13]) ? node3714 : node3703;
										assign node3703 = (inp[7]) ? node3711 : node3704;
											assign node3704 = (inp[11]) ? node3706 : 14'b00000011111111;
												assign node3706 = (inp[8]) ? node3708 : 14'b00000011111111;
													assign node3708 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3711 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3714 = (inp[7]) ? node3718 : node3715;
											assign node3715 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3718 = (inp[11]) ? node3720 : 14'b00000000111111;
												assign node3720 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3723 = (inp[7]) ? node3731 : node3724;
										assign node3724 = (inp[13]) ? 14'b00000000111111 : node3725;
											assign node3725 = (inp[0]) ? 14'b00000000111111 : node3726;
												assign node3726 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3731 = (inp[3]) ? node3737 : node3732;
											assign node3732 = (inp[0]) ? 14'b00000000111111 : node3733;
												assign node3733 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3737 = (inp[0]) ? node3743 : node3738;
												assign node3738 = (inp[11]) ? 14'b00000000011111 : node3739;
													assign node3739 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3743 = (inp[13]) ? 14'b00000000000111 : node3744;
													assign node3744 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node3748 = (inp[8]) ? node3786 : node3749;
									assign node3749 = (inp[3]) ? node3771 : node3750;
										assign node3750 = (inp[13]) ? node3762 : node3751;
											assign node3751 = (inp[7]) ? node3755 : node3752;
												assign node3752 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3755 = (inp[0]) ? node3757 : 14'b00000001111111;
													assign node3757 = (inp[11]) ? 14'b00000000111111 : node3758;
														assign node3758 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3762 = (inp[1]) ? node3766 : node3763;
												assign node3763 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3766 = (inp[11]) ? 14'b00000000011111 : node3767;
													assign node3767 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3771 = (inp[7]) ? node3781 : node3772;
											assign node3772 = (inp[11]) ? node3774 : 14'b00000000111111;
												assign node3774 = (inp[13]) ? 14'b00000000011111 : node3775;
													assign node3775 = (inp[1]) ? node3777 : 14'b00000000111111;
														assign node3777 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3781 = (inp[0]) ? 14'b00000000011111 : node3782;
												assign node3782 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3786 = (inp[0]) ? node3796 : node3787;
										assign node3787 = (inp[7]) ? node3789 : 14'b00000000111111;
											assign node3789 = (inp[1]) ? node3791 : 14'b00000000111111;
												assign node3791 = (inp[11]) ? node3793 : 14'b00000000011111;
													assign node3793 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3796 = (inp[1]) ? node3802 : node3797;
											assign node3797 = (inp[13]) ? 14'b00000000011111 : node3798;
												assign node3798 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3802 = (inp[11]) ? node3804 : 14'b00000000011111;
												assign node3804 = (inp[3]) ? 14'b00000000001111 : 14'b00000000000111;
				assign node3807 = (inp[7]) ? node4197 : node3808;
					assign node3808 = (inp[3]) ? node4014 : node3809;
						assign node3809 = (inp[11]) ? node3903 : node3810;
							assign node3810 = (inp[2]) ? node3850 : node3811;
								assign node3811 = (inp[0]) ? node3833 : node3812;
									assign node3812 = (inp[13]) ? node3820 : node3813;
										assign node3813 = (inp[1]) ? node3815 : 14'b00001111111111;
											assign node3815 = (inp[9]) ? 14'b00000111111111 : node3816;
												assign node3816 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3820 = (inp[6]) ? node3824 : node3821;
											assign node3821 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3824 = (inp[9]) ? node3830 : node3825;
												assign node3825 = (inp[5]) ? node3827 : 14'b00000111111111;
													assign node3827 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3830 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3833 = (inp[6]) ? node3839 : node3834;
										assign node3834 = (inp[9]) ? 14'b00000011111111 : node3835;
											assign node3835 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3839 = (inp[1]) ? node3845 : node3840;
											assign node3840 = (inp[8]) ? 14'b00000001111111 : node3841;
												assign node3841 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3845 = (inp[5]) ? 14'b00000001111111 : node3846;
												assign node3846 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node3850 = (inp[13]) ? node3874 : node3851;
									assign node3851 = (inp[5]) ? node3861 : node3852;
										assign node3852 = (inp[9]) ? node3854 : 14'b00000111111111;
											assign node3854 = (inp[6]) ? 14'b00000011111111 : node3855;
												assign node3855 = (inp[8]) ? 14'b00000111111111 : node3856;
													assign node3856 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3861 = (inp[1]) ? node3863 : 14'b00000011111111;
											assign node3863 = (inp[6]) ? node3869 : node3864;
												assign node3864 = (inp[8]) ? 14'b00000001111111 : node3865;
													assign node3865 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3869 = (inp[8]) ? node3871 : 14'b00000000111111;
													assign node3871 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3874 = (inp[1]) ? node3886 : node3875;
										assign node3875 = (inp[5]) ? node3881 : node3876;
											assign node3876 = (inp[6]) ? node3878 : 14'b00000011111111;
												assign node3878 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3881 = (inp[6]) ? node3883 : 14'b00000001111111;
												assign node3883 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node3886 = (inp[6]) ? node3898 : node3887;
											assign node3887 = (inp[5]) ? node3893 : node3888;
												assign node3888 = (inp[0]) ? 14'b00000001111111 : node3889;
													assign node3889 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3893 = (inp[0]) ? node3895 : 14'b00000001111111;
													assign node3895 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3898 = (inp[0]) ? 14'b00000000011111 : node3899;
												assign node3899 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node3903 = (inp[8]) ? node3949 : node3904;
								assign node3904 = (inp[13]) ? node3938 : node3905;
									assign node3905 = (inp[6]) ? node3927 : node3906;
										assign node3906 = (inp[5]) ? node3916 : node3907;
											assign node3907 = (inp[2]) ? node3911 : node3908;
												assign node3908 = (inp[1]) ? 14'b00001111111111 : 14'b00000111111111;
												assign node3911 = (inp[1]) ? node3913 : 14'b00000111111111;
													assign node3913 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3916 = (inp[0]) ? node3920 : node3917;
												assign node3917 = (inp[2]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node3920 = (inp[2]) ? node3922 : 14'b00000011111111;
													assign node3922 = (inp[1]) ? 14'b00000001111111 : node3923;
														assign node3923 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3927 = (inp[2]) ? node3933 : node3928;
											assign node3928 = (inp[9]) ? node3930 : 14'b00000011111111;
												assign node3930 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3933 = (inp[1]) ? 14'b00000000111111 : node3934;
												assign node3934 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3938 = (inp[5]) ? node3942 : node3939;
										assign node3939 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3942 = (inp[0]) ? node3944 : 14'b00000001111111;
											assign node3944 = (inp[6]) ? 14'b00000000011111 : node3945;
												assign node3945 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node3949 = (inp[1]) ? node3971 : node3950;
									assign node3950 = (inp[9]) ? node3964 : node3951;
										assign node3951 = (inp[6]) ? node3957 : node3952;
											assign node3952 = (inp[13]) ? node3954 : 14'b00000011111111;
												assign node3954 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3957 = (inp[5]) ? node3961 : node3958;
												assign node3958 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3961 = (inp[0]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node3964 = (inp[5]) ? node3966 : 14'b00000001111111;
											assign node3966 = (inp[2]) ? node3968 : 14'b00000000111111;
												assign node3968 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3971 = (inp[9]) ? node3995 : node3972;
										assign node3972 = (inp[2]) ? node3982 : node3973;
											assign node3973 = (inp[6]) ? node3975 : 14'b00000111111111;
												assign node3975 = (inp[13]) ? 14'b00000001111111 : node3976;
													assign node3976 = (inp[0]) ? 14'b00000001111111 : node3977;
														assign node3977 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3982 = (inp[13]) ? node3988 : node3983;
												assign node3983 = (inp[0]) ? 14'b00000000111111 : node3984;
													assign node3984 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3988 = (inp[6]) ? node3990 : 14'b00000000111111;
													assign node3990 = (inp[0]) ? node3992 : 14'b00000000011111;
														assign node3992 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3995 = (inp[6]) ? node4005 : node3996;
											assign node3996 = (inp[5]) ? node3998 : 14'b00000000111111;
												assign node3998 = (inp[2]) ? 14'b00000000011111 : node3999;
													assign node3999 = (inp[13]) ? node4001 : 14'b00000000111111;
														assign node4001 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4005 = (inp[2]) ? node4011 : node4006;
												assign node4006 = (inp[13]) ? 14'b00000000011111 : node4007;
													assign node4007 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4011 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
						assign node4014 = (inp[8]) ? node4104 : node4015;
							assign node4015 = (inp[0]) ? node4057 : node4016;
								assign node4016 = (inp[5]) ? node4042 : node4017;
									assign node4017 = (inp[11]) ? node4029 : node4018;
										assign node4018 = (inp[1]) ? node4024 : node4019;
											assign node4019 = (inp[6]) ? 14'b00000111111111 : node4020;
												assign node4020 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4024 = (inp[9]) ? 14'b00000011111111 : node4025;
												assign node4025 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4029 = (inp[9]) ? 14'b00000001111111 : node4030;
											assign node4030 = (inp[2]) ? 14'b00000001111111 : node4031;
												assign node4031 = (inp[1]) ? node4037 : node4032;
													assign node4032 = (inp[6]) ? node4034 : 14'b00000111111111;
														assign node4034 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
													assign node4037 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4042 = (inp[1]) ? node4050 : node4043;
										assign node4043 = (inp[9]) ? node4045 : 14'b00000011111111;
											assign node4045 = (inp[13]) ? 14'b00000001111111 : node4046;
												assign node4046 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4050 = (inp[2]) ? node4054 : node4051;
											assign node4051 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4054 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4057 = (inp[13]) ? node4075 : node4058;
									assign node4058 = (inp[6]) ? node4066 : node4059;
										assign node4059 = (inp[11]) ? 14'b00000011111111 : node4060;
											assign node4060 = (inp[9]) ? 14'b00000001111111 : node4061;
												assign node4061 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4066 = (inp[9]) ? node4070 : node4067;
											assign node4067 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4070 = (inp[5]) ? node4072 : 14'b00000000111111;
												assign node4072 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4075 = (inp[6]) ? node4091 : node4076;
										assign node4076 = (inp[11]) ? node4086 : node4077;
											assign node4077 = (inp[1]) ? node4079 : 14'b00000001111111;
												assign node4079 = (inp[2]) ? node4081 : 14'b00000001111111;
													assign node4081 = (inp[5]) ? 14'b00000000111111 : node4082;
														assign node4082 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4086 = (inp[5]) ? node4088 : 14'b00000000111111;
												assign node4088 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4091 = (inp[11]) ? node4101 : node4092;
											assign node4092 = (inp[9]) ? node4096 : node4093;
												assign node4093 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4096 = (inp[2]) ? 14'b00000000011111 : node4097;
													assign node4097 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4101 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
							assign node4104 = (inp[13]) ? node4144 : node4105;
								assign node4105 = (inp[1]) ? node4125 : node4106;
									assign node4106 = (inp[5]) ? node4118 : node4107;
										assign node4107 = (inp[11]) ? node4109 : 14'b00000011111111;
											assign node4109 = (inp[6]) ? 14'b00000000111111 : node4110;
												assign node4110 = (inp[0]) ? node4112 : 14'b00000011111111;
													assign node4112 = (inp[2]) ? 14'b00000001111111 : node4113;
														assign node4113 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4118 = (inp[11]) ? 14'b00000000111111 : node4119;
											assign node4119 = (inp[6]) ? node4121 : 14'b00000001111111;
												assign node4121 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4125 = (inp[2]) ? node4135 : node4126;
										assign node4126 = (inp[9]) ? node4132 : node4127;
											assign node4127 = (inp[0]) ? node4129 : 14'b00000001111111;
												assign node4129 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4132 = (inp[11]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node4135 = (inp[11]) ? node4141 : node4136;
											assign node4136 = (inp[5]) ? node4138 : 14'b00000000111111;
												assign node4138 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4141 = (inp[9]) ? 14'b00000000011111 : 14'b00000000001111;
								assign node4144 = (inp[1]) ? node4178 : node4145;
									assign node4145 = (inp[2]) ? node4165 : node4146;
										assign node4146 = (inp[5]) ? node4156 : node4147;
											assign node4147 = (inp[6]) ? node4149 : 14'b00000001111111;
												assign node4149 = (inp[9]) ? node4151 : 14'b00000001111111;
													assign node4151 = (inp[0]) ? 14'b00000000111111 : node4152;
														assign node4152 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4156 = (inp[9]) ? node4162 : node4157;
												assign node4157 = (inp[0]) ? 14'b00000000111111 : node4158;
													assign node4158 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4162 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4165 = (inp[6]) ? node4169 : node4166;
											assign node4166 = (inp[5]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node4169 = (inp[11]) ? node4173 : node4170;
												assign node4170 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4173 = (inp[0]) ? node4175 : 14'b00000000011111;
													assign node4175 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node4178 = (inp[2]) ? node4190 : node4179;
										assign node4179 = (inp[9]) ? node4185 : node4180;
											assign node4180 = (inp[6]) ? 14'b00000000111111 : node4181;
												assign node4181 = (inp[0]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node4185 = (inp[5]) ? node4187 : 14'b00000000011111;
												assign node4187 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4190 = (inp[11]) ? node4192 : 14'b00000000011111;
											assign node4192 = (inp[0]) ? node4194 : 14'b00000000011111;
												assign node4194 = (inp[6]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node4197 = (inp[6]) ? node4381 : node4198;
						assign node4198 = (inp[1]) ? node4290 : node4199;
							assign node4199 = (inp[11]) ? node4241 : node4200;
								assign node4200 = (inp[9]) ? node4228 : node4201;
									assign node4201 = (inp[13]) ? node4211 : node4202;
										assign node4202 = (inp[5]) ? 14'b00000011111111 : node4203;
											assign node4203 = (inp[2]) ? 14'b00000111111111 : node4204;
												assign node4204 = (inp[0]) ? node4206 : 14'b00011111111111;
													assign node4206 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node4211 = (inp[2]) ? node4219 : node4212;
											assign node4212 = (inp[3]) ? 14'b00000011111111 : node4213;
												assign node4213 = (inp[8]) ? node4215 : 14'b00001111111111;
													assign node4215 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4219 = (inp[8]) ? 14'b00000001111111 : node4220;
												assign node4220 = (inp[3]) ? node4222 : 14'b00000011111111;
													assign node4222 = (inp[0]) ? 14'b00000001111111 : node4223;
														assign node4223 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4228 = (inp[2]) ? node4234 : node4229;
										assign node4229 = (inp[13]) ? node4231 : 14'b00000011111111;
											assign node4231 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4234 = (inp[13]) ? node4236 : 14'b00000001111111;
											assign node4236 = (inp[5]) ? node4238 : 14'b00000000111111;
												assign node4238 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4241 = (inp[13]) ? node4257 : node4242;
									assign node4242 = (inp[0]) ? node4250 : node4243;
										assign node4243 = (inp[2]) ? 14'b00000001111111 : node4244;
											assign node4244 = (inp[8]) ? node4246 : 14'b00000011111111;
												assign node4246 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4250 = (inp[5]) ? node4252 : 14'b00000001111111;
											assign node4252 = (inp[8]) ? 14'b00000000011111 : node4253;
												assign node4253 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4257 = (inp[8]) ? node4275 : node4258;
										assign node4258 = (inp[3]) ? node4264 : node4259;
											assign node4259 = (inp[5]) ? 14'b00000001111111 : node4260;
												assign node4260 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4264 = (inp[9]) ? node4272 : node4265;
												assign node4265 = (inp[5]) ? node4267 : 14'b00000011111111;
													assign node4267 = (inp[0]) ? 14'b00000000111111 : node4268;
														assign node4268 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4272 = (inp[0]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node4275 = (inp[0]) ? node4283 : node4276;
											assign node4276 = (inp[5]) ? 14'b00000000111111 : node4277;
												assign node4277 = (inp[2]) ? 14'b00000000111111 : node4278;
													assign node4278 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4283 = (inp[5]) ? node4287 : node4284;
												assign node4284 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4287 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node4290 = (inp[3]) ? node4330 : node4291;
								assign node4291 = (inp[5]) ? node4307 : node4292;
									assign node4292 = (inp[8]) ? node4296 : node4293;
										assign node4293 = (inp[9]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node4296 = (inp[0]) ? node4302 : node4297;
											assign node4297 = (inp[9]) ? 14'b00000001111111 : node4298;
												assign node4298 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4302 = (inp[13]) ? 14'b00000000111111 : node4303;
												assign node4303 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4307 = (inp[11]) ? node4315 : node4308;
										assign node4308 = (inp[2]) ? 14'b00000000111111 : node4309;
											assign node4309 = (inp[13]) ? node4311 : 14'b00000001111111;
												assign node4311 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4315 = (inp[9]) ? node4321 : node4316;
											assign node4316 = (inp[2]) ? 14'b00000000011111 : node4317;
												assign node4317 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4321 = (inp[8]) ? node4325 : node4322;
												assign node4322 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4325 = (inp[0]) ? 14'b00000000001111 : node4326;
													assign node4326 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node4330 = (inp[2]) ? node4358 : node4331;
									assign node4331 = (inp[13]) ? node4343 : node4332;
										assign node4332 = (inp[5]) ? node4336 : node4333;
											assign node4333 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4336 = (inp[0]) ? node4338 : 14'b00000001111111;
												assign node4338 = (inp[8]) ? node4340 : 14'b00000000111111;
													assign node4340 = (inp[11]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node4343 = (inp[11]) ? node4349 : node4344;
											assign node4344 = (inp[0]) ? 14'b00000000111111 : node4345;
												assign node4345 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4349 = (inp[0]) ? node4353 : node4350;
												assign node4350 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4353 = (inp[5]) ? 14'b00000000001111 : node4354;
													assign node4354 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4358 = (inp[0]) ? node4370 : node4359;
										assign node4359 = (inp[11]) ? 14'b00000000011111 : node4360;
											assign node4360 = (inp[13]) ? node4362 : 14'b00000001111111;
												assign node4362 = (inp[9]) ? node4366 : node4363;
													assign node4363 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
													assign node4366 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4370 = (inp[11]) ? node4374 : node4371;
											assign node4371 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4374 = (inp[9]) ? node4376 : 14'b00000000011111;
												assign node4376 = (inp[5]) ? 14'b00000000000111 : node4377;
													assign node4377 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node4381 = (inp[11]) ? node4479 : node4382;
							assign node4382 = (inp[2]) ? node4436 : node4383;
								assign node4383 = (inp[8]) ? node4403 : node4384;
									assign node4384 = (inp[9]) ? node4396 : node4385;
										assign node4385 = (inp[13]) ? node4391 : node4386;
											assign node4386 = (inp[0]) ? 14'b00000001111111 : node4387;
												assign node4387 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4391 = (inp[0]) ? node4393 : 14'b00000001111111;
												assign node4393 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4396 = (inp[1]) ? 14'b00000000111111 : node4397;
											assign node4397 = (inp[13]) ? node4399 : 14'b00000001111111;
												assign node4399 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node4403 = (inp[1]) ? node4421 : node4404;
										assign node4404 = (inp[9]) ? node4412 : node4405;
											assign node4405 = (inp[3]) ? node4409 : node4406;
												assign node4406 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4409 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4412 = (inp[13]) ? node4418 : node4413;
												assign node4413 = (inp[5]) ? 14'b00000000111111 : node4414;
													assign node4414 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4418 = (inp[3]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node4421 = (inp[5]) ? node4427 : node4422;
											assign node4422 = (inp[9]) ? 14'b00000000011111 : node4423;
												assign node4423 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4427 = (inp[3]) ? node4431 : node4428;
												assign node4428 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4431 = (inp[13]) ? 14'b00000000001111 : node4432;
													assign node4432 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node4436 = (inp[8]) ? node4458 : node4437;
									assign node4437 = (inp[1]) ? node4451 : node4438;
										assign node4438 = (inp[0]) ? node4446 : node4439;
											assign node4439 = (inp[5]) ? node4443 : node4440;
												assign node4440 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4443 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4446 = (inp[13]) ? 14'b00000000111111 : node4447;
												assign node4447 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4451 = (inp[13]) ? node4453 : 14'b00000000111111;
											assign node4453 = (inp[0]) ? node4455 : 14'b00000000011111;
												assign node4455 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node4458 = (inp[5]) ? node4464 : node4459;
										assign node4459 = (inp[1]) ? 14'b00000000011111 : node4460;
											assign node4460 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4464 = (inp[13]) ? node4476 : node4465;
											assign node4465 = (inp[3]) ? node4471 : node4466;
												assign node4466 = (inp[9]) ? 14'b00000000011111 : node4467;
													assign node4467 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4471 = (inp[1]) ? 14'b00000000001111 : node4472;
													assign node4472 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4476 = (inp[1]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node4479 = (inp[3]) ? node4525 : node4480;
								assign node4480 = (inp[0]) ? node4498 : node4481;
									assign node4481 = (inp[5]) ? node4485 : node4482;
										assign node4482 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4485 = (inp[2]) ? node4493 : node4486;
											assign node4486 = (inp[13]) ? node4488 : 14'b00000000111111;
												assign node4488 = (inp[9]) ? node4490 : 14'b00000000111111;
													assign node4490 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4493 = (inp[8]) ? 14'b00000000001111 : node4494;
												assign node4494 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4498 = (inp[13]) ? node4510 : node4499;
										assign node4499 = (inp[2]) ? node4501 : 14'b00000000111111;
											assign node4501 = (inp[5]) ? node4505 : node4502;
												assign node4502 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4505 = (inp[1]) ? node4507 : 14'b00000000011111;
													assign node4507 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4510 = (inp[8]) ? node4514 : node4511;
											assign node4511 = (inp[9]) ? 14'b00000000111111 : 14'b00000000011111;
											assign node4514 = (inp[1]) ? node4522 : node4515;
												assign node4515 = (inp[9]) ? 14'b00000000000111 : node4516;
													assign node4516 = (inp[2]) ? node4518 : 14'b00000000011111;
														assign node4518 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node4522 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node4525 = (inp[1]) ? node4551 : node4526;
									assign node4526 = (inp[13]) ? node4534 : node4527;
										assign node4527 = (inp[5]) ? node4531 : node4528;
											assign node4528 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node4531 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4534 = (inp[5]) ? node4542 : node4535;
											assign node4535 = (inp[9]) ? node4539 : node4536;
												assign node4536 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4539 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4542 = (inp[2]) ? node4546 : node4543;
												assign node4543 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node4546 = (inp[8]) ? node4548 : 14'b00000000000111;
													assign node4548 = (inp[9]) ? 14'b00000000000011 : 14'b00000000000111;
									assign node4551 = (inp[8]) ? node4561 : node4552;
										assign node4552 = (inp[9]) ? node4556 : node4553;
											assign node4553 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4556 = (inp[0]) ? node4558 : 14'b00000000001111;
												assign node4558 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node4561 = (inp[13]) ? node4569 : node4562;
											assign node4562 = (inp[0]) ? node4564 : 14'b00000000001111;
												assign node4564 = (inp[9]) ? 14'b00000000000111 : node4565;
													assign node4565 = (inp[5]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node4569 = (inp[0]) ? node4571 : 14'b00000000000111;
												assign node4571 = (inp[9]) ? node4573 : 14'b00000000000011;
													assign node4573 = (inp[5]) ? 14'b00000000000001 : 14'b00000000000011;
			assign node4576 = (inp[5]) ? node5258 : node4577;
				assign node4577 = (inp[8]) ? node4909 : node4578;
					assign node4578 = (inp[0]) ? node4744 : node4579;
						assign node4579 = (inp[9]) ? node4679 : node4580;
							assign node4580 = (inp[13]) ? node4630 : node4581;
								assign node4581 = (inp[11]) ? node4603 : node4582;
									assign node4582 = (inp[3]) ? node4590 : node4583;
										assign node4583 = (inp[1]) ? 14'b00000111111111 : node4584;
											assign node4584 = (inp[7]) ? node4586 : 14'b00011111111111;
												assign node4586 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node4590 = (inp[2]) ? node4600 : node4591;
											assign node4591 = (inp[12]) ? node4597 : node4592;
												assign node4592 = (inp[6]) ? 14'b00000111111111 : node4593;
													assign node4593 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4597 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4600 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4603 = (inp[3]) ? node4619 : node4604;
										assign node4604 = (inp[2]) ? node4612 : node4605;
											assign node4605 = (inp[12]) ? node4607 : 14'b00011111111111;
												assign node4607 = (inp[6]) ? node4609 : 14'b00000111111111;
													assign node4609 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4612 = (inp[7]) ? node4616 : node4613;
												assign node4613 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4616 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4619 = (inp[1]) ? node4625 : node4620;
											assign node4620 = (inp[6]) ? node4622 : 14'b00000011111111;
												assign node4622 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4625 = (inp[7]) ? 14'b00000001111111 : node4626;
												assign node4626 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node4630 = (inp[1]) ? node4660 : node4631;
									assign node4631 = (inp[12]) ? node4641 : node4632;
										assign node4632 = (inp[3]) ? node4636 : node4633;
											assign node4633 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4636 = (inp[7]) ? 14'b00000011111111 : node4637;
												assign node4637 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4641 = (inp[3]) ? node4647 : node4642;
											assign node4642 = (inp[11]) ? 14'b00000011111111 : node4643;
												assign node4643 = (inp[6]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node4647 = (inp[6]) ? node4655 : node4648;
												assign node4648 = (inp[2]) ? 14'b00000001111111 : node4649;
													assign node4649 = (inp[11]) ? 14'b00000011111111 : node4650;
														assign node4650 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4655 = (inp[2]) ? node4657 : 14'b00000001111111;
													assign node4657 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4660 = (inp[11]) ? node4670 : node4661;
										assign node4661 = (inp[6]) ? node4663 : 14'b00000011111111;
											assign node4663 = (inp[12]) ? node4667 : node4664;
												assign node4664 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4667 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4670 = (inp[2]) ? 14'b00000000111111 : node4671;
											assign node4671 = (inp[12]) ? node4675 : node4672;
												assign node4672 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4675 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node4679 = (inp[7]) ? node4717 : node4680;
								assign node4680 = (inp[13]) ? node4700 : node4681;
									assign node4681 = (inp[12]) ? node4689 : node4682;
										assign node4682 = (inp[11]) ? node4686 : node4683;
											assign node4683 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node4686 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4689 = (inp[11]) ? node4695 : node4690;
											assign node4690 = (inp[1]) ? node4692 : 14'b00000011111111;
												assign node4692 = (inp[6]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node4695 = (inp[6]) ? 14'b00000001111111 : node4696;
												assign node4696 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4700 = (inp[3]) ? node4708 : node4701;
										assign node4701 = (inp[12]) ? 14'b00000001111111 : node4702;
											assign node4702 = (inp[6]) ? node4704 : 14'b00000111111111;
												assign node4704 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4708 = (inp[11]) ? node4710 : 14'b00000001111111;
											assign node4710 = (inp[6]) ? node4714 : node4711;
												assign node4711 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4714 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4717 = (inp[3]) ? node4729 : node4718;
									assign node4718 = (inp[1]) ? node4724 : node4719;
										assign node4719 = (inp[6]) ? 14'b00000001111111 : node4720;
											assign node4720 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4724 = (inp[11]) ? node4726 : 14'b00000001111111;
											assign node4726 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4729 = (inp[12]) ? node4735 : node4730;
										assign node4730 = (inp[2]) ? node4732 : 14'b00000001111111;
											assign node4732 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4735 = (inp[13]) ? node4741 : node4736;
											assign node4736 = (inp[6]) ? node4738 : 14'b00000000111111;
												assign node4738 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4741 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node4744 = (inp[1]) ? node4830 : node4745;
							assign node4745 = (inp[7]) ? node4783 : node4746;
								assign node4746 = (inp[13]) ? node4766 : node4747;
									assign node4747 = (inp[11]) ? node4757 : node4748;
										assign node4748 = (inp[3]) ? node4754 : node4749;
											assign node4749 = (inp[2]) ? 14'b00000111111111 : node4750;
												assign node4750 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4754 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4757 = (inp[9]) ? node4763 : node4758;
											assign node4758 = (inp[3]) ? 14'b00000011111111 : node4759;
												assign node4759 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4763 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4766 = (inp[6]) ? node4772 : node4767;
										assign node4767 = (inp[3]) ? 14'b00000001111111 : node4768;
											assign node4768 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node4772 = (inp[3]) ? 14'b00000000111111 : node4773;
											assign node4773 = (inp[2]) ? node4777 : node4774;
												assign node4774 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4777 = (inp[9]) ? 14'b00000000111111 : node4778;
													assign node4778 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4783 = (inp[3]) ? node4805 : node4784;
									assign node4784 = (inp[13]) ? node4792 : node4785;
										assign node4785 = (inp[6]) ? 14'b00000001111111 : node4786;
											assign node4786 = (inp[11]) ? node4788 : 14'b00000011111111;
												assign node4788 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4792 = (inp[9]) ? node4798 : node4793;
											assign node4793 = (inp[2]) ? 14'b00000001111111 : node4794;
												assign node4794 = (inp[11]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node4798 = (inp[11]) ? 14'b00000001111111 : node4799;
												assign node4799 = (inp[12]) ? 14'b00000000111111 : node4800;
													assign node4800 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4805 = (inp[9]) ? node4821 : node4806;
										assign node4806 = (inp[2]) ? node4808 : 14'b00000001111111;
											assign node4808 = (inp[11]) ? node4816 : node4809;
												assign node4809 = (inp[12]) ? 14'b00000000111111 : node4810;
													assign node4810 = (inp[6]) ? node4812 : 14'b00000001111111;
														assign node4812 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4816 = (inp[12]) ? 14'b00000000001111 : node4817;
													assign node4817 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4821 = (inp[13]) ? 14'b00000000011111 : node4822;
											assign node4822 = (inp[2]) ? node4826 : node4823;
												assign node4823 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4826 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node4830 = (inp[3]) ? node4868 : node4831;
								assign node4831 = (inp[2]) ? node4851 : node4832;
									assign node4832 = (inp[6]) ? node4842 : node4833;
										assign node4833 = (inp[13]) ? node4837 : node4834;
											assign node4834 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4837 = (inp[7]) ? 14'b00000001111111 : node4838;
												assign node4838 = (inp[9]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node4842 = (inp[9]) ? node4848 : node4843;
											assign node4843 = (inp[7]) ? node4845 : 14'b00000011111111;
												assign node4845 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4848 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4851 = (inp[12]) ? node4861 : node4852;
										assign node4852 = (inp[11]) ? node4856 : node4853;
											assign node4853 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4856 = (inp[13]) ? node4858 : 14'b00000000111111;
												assign node4858 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node4861 = (inp[9]) ? node4865 : node4862;
											assign node4862 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4865 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node4868 = (inp[12]) ? node4892 : node4869;
									assign node4869 = (inp[6]) ? node4877 : node4870;
										assign node4870 = (inp[7]) ? 14'b00000000111111 : node4871;
											assign node4871 = (inp[9]) ? node4873 : 14'b00000001111111;
												assign node4873 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4877 = (inp[2]) ? node4885 : node4878;
											assign node4878 = (inp[7]) ? node4882 : node4879;
												assign node4879 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4882 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4885 = (inp[11]) ? 14'b00000000001111 : node4886;
												assign node4886 = (inp[9]) ? 14'b00000000011111 : node4887;
													assign node4887 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4892 = (inp[7]) ? node4894 : 14'b00000000011111;
										assign node4894 = (inp[2]) ? node4904 : node4895;
											assign node4895 = (inp[11]) ? node4899 : node4896;
												assign node4896 = (inp[13]) ? 14'b00000000111111 : 14'b00000000011111;
												assign node4899 = (inp[6]) ? 14'b00000000001111 : node4900;
													assign node4900 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4904 = (inp[13]) ? 14'b00000000001111 : node4905;
												assign node4905 = (inp[6]) ? 14'b00000000011111 : 14'b00000000001111;
					assign node4909 = (inp[2]) ? node5089 : node4910;
						assign node4910 = (inp[13]) ? node4992 : node4911;
							assign node4911 = (inp[12]) ? node4959 : node4912;
								assign node4912 = (inp[1]) ? node4938 : node4913;
									assign node4913 = (inp[3]) ? node4925 : node4914;
										assign node4914 = (inp[11]) ? node4918 : node4915;
											assign node4915 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4918 = (inp[9]) ? node4920 : 14'b00000111111111;
												assign node4920 = (inp[0]) ? 14'b00000011111111 : node4921;
													assign node4921 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4925 = (inp[9]) ? node4933 : node4926;
											assign node4926 = (inp[7]) ? 14'b00000011111111 : node4927;
												assign node4927 = (inp[11]) ? node4929 : 14'b00000111111111;
													assign node4929 = (inp[6]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4933 = (inp[6]) ? 14'b00000001111111 : node4934;
												assign node4934 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4938 = (inp[3]) ? node4950 : node4939;
										assign node4939 = (inp[11]) ? 14'b00000001111111 : node4940;
											assign node4940 = (inp[9]) ? node4944 : node4941;
												assign node4941 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4944 = (inp[7]) ? node4946 : 14'b00000011111111;
													assign node4946 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4950 = (inp[11]) ? node4956 : node4951;
											assign node4951 = (inp[0]) ? 14'b00000001111111 : node4952;
												assign node4952 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4956 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4959 = (inp[1]) ? node4975 : node4960;
									assign node4960 = (inp[9]) ? node4970 : node4961;
										assign node4961 = (inp[11]) ? node4965 : node4962;
											assign node4962 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4965 = (inp[3]) ? 14'b00000000111111 : node4966;
												assign node4966 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4970 = (inp[7]) ? 14'b00000001111111 : node4971;
											assign node4971 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4975 = (inp[7]) ? node4987 : node4976;
										assign node4976 = (inp[6]) ? 14'b00000000111111 : node4977;
											assign node4977 = (inp[11]) ? node4983 : node4978;
												assign node4978 = (inp[9]) ? node4980 : 14'b00000111111111;
													assign node4980 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4983 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4987 = (inp[9]) ? node4989 : 14'b00000000111111;
											assign node4989 = (inp[0]) ? 14'b00000000111111 : 14'b00000000011111;
							assign node4992 = (inp[1]) ? node5042 : node4993;
								assign node4993 = (inp[7]) ? node5015 : node4994;
									assign node4994 = (inp[11]) ? node5010 : node4995;
										assign node4995 = (inp[12]) ? node5003 : node4996;
											assign node4996 = (inp[6]) ? node4998 : 14'b00000011111111;
												assign node4998 = (inp[9]) ? node5000 : 14'b00000011111111;
													assign node5000 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5003 = (inp[0]) ? node5007 : node5004;
												assign node5004 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5007 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5010 = (inp[3]) ? 14'b00000000111111 : node5011;
											assign node5011 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5015 = (inp[3]) ? node5029 : node5016;
										assign node5016 = (inp[0]) ? node5022 : node5017;
											assign node5017 = (inp[9]) ? node5019 : 14'b00000001111111;
												assign node5019 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5022 = (inp[9]) ? node5026 : node5023;
												assign node5023 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5026 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5029 = (inp[0]) ? node5039 : node5030;
											assign node5030 = (inp[6]) ? node5036 : node5031;
												assign node5031 = (inp[9]) ? 14'b00000000111111 : node5032;
													assign node5032 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5036 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5039 = (inp[6]) ? 14'b00000000111111 : 14'b00000000011111;
								assign node5042 = (inp[12]) ? node5066 : node5043;
									assign node5043 = (inp[6]) ? node5049 : node5044;
										assign node5044 = (inp[11]) ? 14'b00000000111111 : node5045;
											assign node5045 = (inp[7]) ? 14'b00000001111111 : 14'b00000000111111;
										assign node5049 = (inp[9]) ? node5059 : node5050;
											assign node5050 = (inp[7]) ? node5056 : node5051;
												assign node5051 = (inp[0]) ? 14'b00000000111111 : node5052;
													assign node5052 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5056 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5059 = (inp[7]) ? 14'b00000000011111 : node5060;
												assign node5060 = (inp[0]) ? 14'b00000000011111 : node5061;
													assign node5061 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5066 = (inp[9]) ? node5078 : node5067;
										assign node5067 = (inp[7]) ? node5069 : 14'b00000000111111;
											assign node5069 = (inp[6]) ? node5073 : node5070;
												assign node5070 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5073 = (inp[0]) ? 14'b00000000001111 : node5074;
													assign node5074 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5078 = (inp[3]) ? node5080 : 14'b00000000011111;
											assign node5080 = (inp[11]) ? node5082 : 14'b00000000001111;
												assign node5082 = (inp[0]) ? node5084 : 14'b00000000000111;
													assign node5084 = (inp[6]) ? node5086 : 14'b00000000000111;
														assign node5086 = (inp[7]) ? 14'b00000000000011 : 14'b00000000000111;
						assign node5089 = (inp[0]) ? node5171 : node5090;
							assign node5090 = (inp[12]) ? node5128 : node5091;
								assign node5091 = (inp[3]) ? node5105 : node5092;
									assign node5092 = (inp[1]) ? node5100 : node5093;
										assign node5093 = (inp[7]) ? 14'b00000000111111 : node5094;
											assign node5094 = (inp[11]) ? node5096 : 14'b00000011111111;
												assign node5096 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5100 = (inp[6]) ? node5102 : 14'b00000001111111;
											assign node5102 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5105 = (inp[13]) ? node5123 : node5106;
										assign node5106 = (inp[7]) ? node5116 : node5107;
											assign node5107 = (inp[1]) ? node5109 : 14'b00000011111111;
												assign node5109 = (inp[11]) ? node5111 : 14'b00000001111111;
													assign node5111 = (inp[6]) ? 14'b00000000111111 : node5112;
														assign node5112 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5116 = (inp[1]) ? 14'b00000000111111 : node5117;
												assign node5117 = (inp[11]) ? 14'b00000000111111 : node5118;
													assign node5118 = (inp[6]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5123 = (inp[7]) ? node5125 : 14'b00000000111111;
											assign node5125 = (inp[11]) ? 14'b00000000011111 : 14'b00000000001111;
								assign node5128 = (inp[7]) ? node5150 : node5129;
									assign node5129 = (inp[6]) ? node5143 : node5130;
										assign node5130 = (inp[9]) ? node5134 : node5131;
											assign node5131 = (inp[3]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node5134 = (inp[1]) ? node5138 : node5135;
												assign node5135 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5138 = (inp[13]) ? node5140 : 14'b00000000111111;
													assign node5140 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5143 = (inp[9]) ? 14'b00000000011111 : node5144;
											assign node5144 = (inp[1]) ? node5146 : 14'b00000000111111;
												assign node5146 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5150 = (inp[1]) ? node5162 : node5151;
										assign node5151 = (inp[3]) ? node5157 : node5152;
											assign node5152 = (inp[11]) ? 14'b00000000111111 : node5153;
												assign node5153 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5157 = (inp[13]) ? 14'b00000000011111 : node5158;
												assign node5158 = (inp[9]) ? 14'b00000000111111 : 14'b00000000011111;
										assign node5162 = (inp[9]) ? node5164 : 14'b00000000011111;
											assign node5164 = (inp[11]) ? node5168 : node5165;
												assign node5165 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5168 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node5171 = (inp[9]) ? node5215 : node5172;
								assign node5172 = (inp[7]) ? node5194 : node5173;
									assign node5173 = (inp[13]) ? node5191 : node5174;
										assign node5174 = (inp[6]) ? node5184 : node5175;
											assign node5175 = (inp[1]) ? 14'b00000000111111 : node5176;
												assign node5176 = (inp[3]) ? 14'b00000001111111 : node5177;
													assign node5177 = (inp[12]) ? node5179 : 14'b00000111111111;
														assign node5179 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5184 = (inp[12]) ? node5186 : 14'b00000001111111;
												assign node5186 = (inp[3]) ? node5188 : 14'b00000000111111;
													assign node5188 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5191 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5194 = (inp[12]) ? node5208 : node5195;
										assign node5195 = (inp[11]) ? node5201 : node5196;
											assign node5196 = (inp[13]) ? node5198 : 14'b00000000111111;
												assign node5198 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5201 = (inp[3]) ? node5205 : node5202;
												assign node5202 = (inp[6]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5205 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5208 = (inp[6]) ? node5210 : 14'b00000000111111;
											assign node5210 = (inp[13]) ? node5212 : 14'b00000000001111;
												assign node5212 = (inp[11]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node5215 = (inp[6]) ? node5237 : node5216;
									assign node5216 = (inp[12]) ? node5228 : node5217;
										assign node5217 = (inp[13]) ? node5219 : 14'b00000000001111;
											assign node5219 = (inp[11]) ? 14'b00000000011111 : node5220;
												assign node5220 = (inp[7]) ? node5222 : 14'b00000000111111;
													assign node5222 = (inp[3]) ? 14'b00000000011111 : node5223;
														assign node5223 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5228 = (inp[13]) ? 14'b00000000001111 : node5229;
											assign node5229 = (inp[7]) ? 14'b00000000011111 : node5230;
												assign node5230 = (inp[11]) ? node5232 : 14'b00000000011111;
													assign node5232 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5237 = (inp[1]) ? node5251 : node5238;
										assign node5238 = (inp[12]) ? node5246 : node5239;
											assign node5239 = (inp[11]) ? node5241 : 14'b00000000111111;
												assign node5241 = (inp[3]) ? 14'b00000000001111 : node5242;
													assign node5242 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5246 = (inp[11]) ? 14'b00000000000111 : node5247;
												assign node5247 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5251 = (inp[7]) ? node5253 : 14'b00000000001111;
											assign node5253 = (inp[12]) ? 14'b00000000000111 : node5254;
												assign node5254 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node5258 = (inp[6]) ? node5620 : node5259;
					assign node5259 = (inp[1]) ? node5435 : node5260;
						assign node5260 = (inp[7]) ? node5348 : node5261;
							assign node5261 = (inp[0]) ? node5299 : node5262;
								assign node5262 = (inp[9]) ? node5286 : node5263;
									assign node5263 = (inp[8]) ? node5275 : node5264;
										assign node5264 = (inp[2]) ? 14'b00000011111111 : node5265;
											assign node5265 = (inp[3]) ? 14'b00000111111111 : node5266;
												assign node5266 = (inp[11]) ? node5268 : 14'b00001111111111;
													assign node5268 = (inp[12]) ? 14'b00000111111111 : node5269;
														assign node5269 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node5275 = (inp[11]) ? node5283 : node5276;
											assign node5276 = (inp[13]) ? node5278 : 14'b00000111111111;
												assign node5278 = (inp[3]) ? 14'b00000011111111 : node5279;
													assign node5279 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5283 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node5286 = (inp[13]) ? node5292 : node5287;
										assign node5287 = (inp[3]) ? node5289 : 14'b00000011111111;
											assign node5289 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5292 = (inp[8]) ? node5294 : 14'b00000111111111;
											assign node5294 = (inp[12]) ? node5296 : 14'b00000001111111;
												assign node5296 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5299 = (inp[13]) ? node5323 : node5300;
									assign node5300 = (inp[3]) ? node5312 : node5301;
										assign node5301 = (inp[8]) ? node5305 : node5302;
											assign node5302 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5305 = (inp[12]) ? 14'b00000001111111 : node5306;
												assign node5306 = (inp[2]) ? 14'b00000011111111 : node5307;
													assign node5307 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5312 = (inp[2]) ? node5318 : node5313;
											assign node5313 = (inp[8]) ? 14'b00000001111111 : node5314;
												assign node5314 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5318 = (inp[11]) ? 14'b00000000011111 : node5319;
												assign node5319 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5323 = (inp[9]) ? node5339 : node5324;
										assign node5324 = (inp[12]) ? node5334 : node5325;
											assign node5325 = (inp[3]) ? node5329 : node5326;
												assign node5326 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5329 = (inp[8]) ? node5331 : 14'b00000001111111;
													assign node5331 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5334 = (inp[11]) ? 14'b00000000111111 : node5335;
												assign node5335 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node5339 = (inp[11]) ? node5343 : node5340;
											assign node5340 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5343 = (inp[2]) ? node5345 : 14'b00000000011111;
												assign node5345 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node5348 = (inp[11]) ? node5394 : node5349;
								assign node5349 = (inp[3]) ? node5369 : node5350;
									assign node5350 = (inp[12]) ? node5362 : node5351;
										assign node5351 = (inp[13]) ? node5357 : node5352;
											assign node5352 = (inp[0]) ? node5354 : 14'b00000011111111;
												assign node5354 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5357 = (inp[0]) ? 14'b00000000111111 : node5358;
												assign node5358 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5362 = (inp[0]) ? node5366 : node5363;
											assign node5363 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5366 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node5369 = (inp[9]) ? node5385 : node5370;
										assign node5370 = (inp[2]) ? node5380 : node5371;
											assign node5371 = (inp[8]) ? node5375 : node5372;
												assign node5372 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5375 = (inp[0]) ? node5377 : 14'b00000001111111;
													assign node5377 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5380 = (inp[0]) ? node5382 : 14'b00000000111111;
												assign node5382 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5385 = (inp[12]) ? node5387 : 14'b00000000111111;
											assign node5387 = (inp[13]) ? node5389 : 14'b00000000011111;
												assign node5389 = (inp[0]) ? node5391 : 14'b00000000001111;
													assign node5391 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node5394 = (inp[2]) ? node5416 : node5395;
									assign node5395 = (inp[9]) ? node5409 : node5396;
										assign node5396 = (inp[8]) ? node5404 : node5397;
											assign node5397 = (inp[13]) ? node5401 : node5398;
												assign node5398 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5401 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5404 = (inp[12]) ? 14'b00000000011111 : node5405;
												assign node5405 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5409 = (inp[3]) ? node5411 : 14'b00000000111111;
											assign node5411 = (inp[8]) ? 14'b00000000001111 : node5412;
												assign node5412 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5416 = (inp[12]) ? node5420 : node5417;
										assign node5417 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5420 = (inp[9]) ? node5426 : node5421;
											assign node5421 = (inp[3]) ? node5423 : 14'b00000000011111;
												assign node5423 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5426 = (inp[3]) ? node5430 : node5427;
												assign node5427 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5430 = (inp[8]) ? node5432 : 14'b00000000001111;
													assign node5432 = (inp[13]) ? 14'b00000000000011 : 14'b00000000000111;
						assign node5435 = (inp[0]) ? node5525 : node5436;
							assign node5436 = (inp[13]) ? node5478 : node5437;
								assign node5437 = (inp[11]) ? node5457 : node5438;
									assign node5438 = (inp[2]) ? node5448 : node5439;
										assign node5439 = (inp[3]) ? node5441 : 14'b00000011111111;
											assign node5441 = (inp[8]) ? 14'b00000001111111 : node5442;
												assign node5442 = (inp[9]) ? node5444 : 14'b00000011111111;
													assign node5444 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5448 = (inp[7]) ? node5454 : node5449;
											assign node5449 = (inp[8]) ? 14'b00000001111111 : node5450;
												assign node5450 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5454 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5457 = (inp[7]) ? node5467 : node5458;
										assign node5458 = (inp[8]) ? node5460 : 14'b00000001111111;
											assign node5460 = (inp[2]) ? node5464 : node5461;
												assign node5461 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5464 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5467 = (inp[8]) ? node5473 : node5468;
											assign node5468 = (inp[12]) ? node5470 : 14'b00000000111111;
												assign node5470 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5473 = (inp[3]) ? 14'b00000000001111 : node5474;
												assign node5474 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node5478 = (inp[3]) ? node5500 : node5479;
									assign node5479 = (inp[12]) ? node5493 : node5480;
										assign node5480 = (inp[8]) ? node5484 : node5481;
											assign node5481 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5484 = (inp[7]) ? node5486 : 14'b00000001111111;
												assign node5486 = (inp[11]) ? 14'b00000000011111 : node5487;
													assign node5487 = (inp[9]) ? node5489 : 14'b00000000111111;
														assign node5489 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5493 = (inp[9]) ? 14'b00000000000111 : node5494;
											assign node5494 = (inp[2]) ? node5496 : 14'b00000000111111;
												assign node5496 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5500 = (inp[7]) ? node5514 : node5501;
										assign node5501 = (inp[11]) ? node5509 : node5502;
											assign node5502 = (inp[8]) ? node5504 : 14'b00000001111111;
												assign node5504 = (inp[12]) ? node5506 : 14'b00000000111111;
													assign node5506 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5509 = (inp[12]) ? node5511 : 14'b00000000011111;
												assign node5511 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5514 = (inp[9]) ? node5516 : 14'b00000000011111;
											assign node5516 = (inp[12]) ? 14'b00000000001111 : node5517;
												assign node5517 = (inp[8]) ? node5519 : 14'b00000000011111;
													assign node5519 = (inp[2]) ? 14'b00000000001111 : node5520;
														assign node5520 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node5525 = (inp[3]) ? node5569 : node5526;
								assign node5526 = (inp[11]) ? node5552 : node5527;
									assign node5527 = (inp[8]) ? node5543 : node5528;
										assign node5528 = (inp[2]) ? node5538 : node5529;
											assign node5529 = (inp[9]) ? node5533 : node5530;
												assign node5530 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5533 = (inp[13]) ? node5535 : 14'b00000001111111;
													assign node5535 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5538 = (inp[12]) ? node5540 : 14'b00000000111111;
												assign node5540 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node5543 = (inp[9]) ? node5549 : node5544;
											assign node5544 = (inp[12]) ? 14'b00000000111111 : node5545;
												assign node5545 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5549 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5552 = (inp[12]) ? node5558 : node5553;
										assign node5553 = (inp[2]) ? 14'b00000000011111 : node5554;
											assign node5554 = (inp[13]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node5558 = (inp[2]) ? node5562 : node5559;
											assign node5559 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5562 = (inp[9]) ? node5566 : node5563;
												assign node5563 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5566 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node5569 = (inp[9]) ? node5591 : node5570;
									assign node5570 = (inp[7]) ? node5582 : node5571;
										assign node5571 = (inp[12]) ? node5575 : node5572;
											assign node5572 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node5575 = (inp[8]) ? node5579 : node5576;
												assign node5576 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5579 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5582 = (inp[12]) ? 14'b00000000001111 : node5583;
											assign node5583 = (inp[13]) ? 14'b00000000011111 : node5584;
												assign node5584 = (inp[8]) ? node5586 : 14'b00000000011111;
													assign node5586 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5591 = (inp[13]) ? node5607 : node5592;
										assign node5592 = (inp[11]) ? node5598 : node5593;
											assign node5593 = (inp[7]) ? node5595 : 14'b00000000011111;
												assign node5595 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5598 = (inp[12]) ? node5604 : node5599;
												assign node5599 = (inp[7]) ? 14'b00000000001111 : node5600;
													assign node5600 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5604 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node5607 = (inp[8]) ? node5613 : node5608;
											assign node5608 = (inp[7]) ? 14'b00000000000011 : node5609;
												assign node5609 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5613 = (inp[7]) ? node5615 : 14'b00000000000111;
												assign node5615 = (inp[11]) ? 14'b00000000000111 : node5616;
													assign node5616 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node5620 = (inp[0]) ? node5816 : node5621;
						assign node5621 = (inp[13]) ? node5721 : node5622;
							assign node5622 = (inp[3]) ? node5668 : node5623;
								assign node5623 = (inp[2]) ? node5651 : node5624;
									assign node5624 = (inp[8]) ? node5632 : node5625;
										assign node5625 = (inp[12]) ? 14'b00000001111111 : node5626;
											assign node5626 = (inp[9]) ? node5628 : 14'b00000111111111;
												assign node5628 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5632 = (inp[7]) ? node5640 : node5633;
											assign node5633 = (inp[11]) ? node5637 : node5634;
												assign node5634 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5637 = (inp[12]) ? 14'b00000001111111 : 14'b00000000111111;
											assign node5640 = (inp[12]) ? node5646 : node5641;
												assign node5641 = (inp[11]) ? node5643 : 14'b00000001111111;
													assign node5643 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5646 = (inp[11]) ? node5648 : 14'b00000000111111;
													assign node5648 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5651 = (inp[8]) ? node5663 : node5652;
										assign node5652 = (inp[7]) ? node5654 : 14'b00000001111111;
											assign node5654 = (inp[12]) ? node5658 : node5655;
												assign node5655 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5658 = (inp[11]) ? node5660 : 14'b00000000111111;
													assign node5660 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5663 = (inp[11]) ? node5665 : 14'b00000000111111;
											assign node5665 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5668 = (inp[8]) ? node5696 : node5669;
									assign node5669 = (inp[7]) ? node5683 : node5670;
										assign node5670 = (inp[12]) ? node5676 : node5671;
											assign node5671 = (inp[11]) ? 14'b00000001111111 : node5672;
												assign node5672 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5676 = (inp[9]) ? node5680 : node5677;
												assign node5677 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5680 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5683 = (inp[1]) ? node5689 : node5684;
											assign node5684 = (inp[12]) ? node5686 : 14'b00000000111111;
												assign node5686 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5689 = (inp[11]) ? node5691 : 14'b00000000011111;
												assign node5691 = (inp[9]) ? node5693 : 14'b00000000001111;
													assign node5693 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node5696 = (inp[12]) ? node5714 : node5697;
										assign node5697 = (inp[7]) ? node5705 : node5698;
											assign node5698 = (inp[11]) ? node5700 : 14'b00000000111111;
												assign node5700 = (inp[2]) ? 14'b00000000001111 : node5701;
													assign node5701 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5705 = (inp[2]) ? node5711 : node5706;
												assign node5706 = (inp[9]) ? 14'b00000000011111 : node5707;
													assign node5707 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5711 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5714 = (inp[9]) ? node5718 : node5715;
											assign node5715 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5718 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node5721 = (inp[12]) ? node5769 : node5722;
								assign node5722 = (inp[7]) ? node5742 : node5723;
									assign node5723 = (inp[8]) ? node5735 : node5724;
										assign node5724 = (inp[1]) ? node5728 : node5725;
											assign node5725 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5728 = (inp[9]) ? 14'b00000000111111 : node5729;
												assign node5729 = (inp[2]) ? 14'b00000000111111 : node5730;
													assign node5730 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5735 = (inp[2]) ? node5737 : 14'b00000000111111;
											assign node5737 = (inp[11]) ? 14'b00000000001111 : node5738;
												assign node5738 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5742 = (inp[9]) ? node5756 : node5743;
										assign node5743 = (inp[3]) ? node5753 : node5744;
											assign node5744 = (inp[8]) ? 14'b00000000111111 : node5745;
												assign node5745 = (inp[1]) ? 14'b00000000111111 : node5746;
													assign node5746 = (inp[11]) ? node5748 : 14'b00000001111111;
														assign node5748 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5753 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5756 = (inp[2]) ? node5760 : node5757;
											assign node5757 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5760 = (inp[8]) ? node5762 : 14'b00000000011111;
												assign node5762 = (inp[11]) ? 14'b00000000000111 : node5763;
													assign node5763 = (inp[3]) ? node5765 : 14'b00000000001111;
														assign node5765 = (inp[1]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node5769 = (inp[11]) ? node5791 : node5770;
									assign node5770 = (inp[2]) ? node5782 : node5771;
										assign node5771 = (inp[8]) ? 14'b00000000011111 : node5772;
											assign node5772 = (inp[1]) ? node5774 : 14'b00000000111111;
												assign node5774 = (inp[9]) ? node5776 : 14'b00000000111111;
													assign node5776 = (inp[3]) ? node5778 : 14'b00000000011111;
														assign node5778 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5782 = (inp[3]) ? 14'b00000000000011 : node5783;
											assign node5783 = (inp[1]) ? node5785 : 14'b00000000011111;
												assign node5785 = (inp[7]) ? node5787 : 14'b00000000011111;
													assign node5787 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node5791 = (inp[8]) ? node5801 : node5792;
										assign node5792 = (inp[7]) ? 14'b00000000001111 : node5793;
											assign node5793 = (inp[2]) ? node5797 : node5794;
												assign node5794 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5797 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5801 = (inp[3]) ? node5807 : node5802;
											assign node5802 = (inp[2]) ? node5804 : 14'b00000000001111;
												assign node5804 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node5807 = (inp[9]) ? node5811 : node5808;
												assign node5808 = (inp[2]) ? 14'b00000000000011 : 14'b00000000001111;
												assign node5811 = (inp[2]) ? node5813 : 14'b00000000000011;
													assign node5813 = (inp[7]) ? 14'b00000000000001 : 14'b00000000000011;
						assign node5816 = (inp[9]) ? node5932 : node5817;
							assign node5817 = (inp[7]) ? node5865 : node5818;
								assign node5818 = (inp[2]) ? node5838 : node5819;
									assign node5819 = (inp[8]) ? node5827 : node5820;
										assign node5820 = (inp[3]) ? 14'b00000000111111 : node5821;
											assign node5821 = (inp[1]) ? 14'b00000001111111 : node5822;
												assign node5822 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5827 = (inp[1]) ? node5831 : node5828;
											assign node5828 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5831 = (inp[13]) ? node5833 : 14'b00000000111111;
												assign node5833 = (inp[11]) ? 14'b00000000011111 : node5834;
													assign node5834 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5838 = (inp[8]) ? node5854 : node5839;
										assign node5839 = (inp[13]) ? node5845 : node5840;
											assign node5840 = (inp[1]) ? 14'b00000000111111 : node5841;
												assign node5841 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node5845 = (inp[3]) ? node5851 : node5846;
												assign node5846 = (inp[12]) ? 14'b00000000011111 : node5847;
													assign node5847 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5851 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5854 = (inp[1]) ? node5860 : node5855;
											assign node5855 = (inp[13]) ? node5857 : 14'b00000000011111;
												assign node5857 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5860 = (inp[11]) ? 14'b00000000001111 : node5861;
												assign node5861 = (inp[13]) ? 14'b00000000011111 : 14'b00000000001111;
								assign node5865 = (inp[11]) ? node5903 : node5866;
									assign node5866 = (inp[1]) ? node5884 : node5867;
										assign node5867 = (inp[12]) ? node5875 : node5868;
											assign node5868 = (inp[8]) ? 14'b00000000111111 : node5869;
												assign node5869 = (inp[3]) ? node5871 : 14'b00000001111111;
													assign node5871 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5875 = (inp[8]) ? node5881 : node5876;
												assign node5876 = (inp[13]) ? 14'b00000000011111 : node5877;
													assign node5877 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5881 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5884 = (inp[2]) ? node5892 : node5885;
											assign node5885 = (inp[13]) ? 14'b00000000001111 : node5886;
												assign node5886 = (inp[3]) ? 14'b00000000011111 : node5887;
													assign node5887 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5892 = (inp[3]) ? node5896 : node5893;
												assign node5893 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5896 = (inp[8]) ? node5898 : 14'b00000000001111;
													assign node5898 = (inp[13]) ? 14'b00000000000111 : node5899;
														assign node5899 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node5903 = (inp[2]) ? node5917 : node5904;
										assign node5904 = (inp[8]) ? node5912 : node5905;
											assign node5905 = (inp[12]) ? 14'b00000000001111 : node5906;
												assign node5906 = (inp[3]) ? node5908 : 14'b00000000011111;
													assign node5908 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5912 = (inp[13]) ? node5914 : 14'b00000000001111;
												assign node5914 = (inp[1]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node5917 = (inp[12]) ? node5925 : node5918;
											assign node5918 = (inp[13]) ? node5920 : 14'b00000000011111;
												assign node5920 = (inp[1]) ? node5922 : 14'b00000000001111;
													assign node5922 = (inp[8]) ? 14'b00000000000011 : 14'b00000000000111;
											assign node5925 = (inp[13]) ? node5927 : 14'b00000000000111;
												assign node5927 = (inp[1]) ? node5929 : 14'b00000000000111;
													assign node5929 = (inp[3]) ? 14'b00000000000001 : 14'b00000000000011;
							assign node5932 = (inp[12]) ? node5974 : node5933;
								assign node5933 = (inp[2]) ? node5949 : node5934;
									assign node5934 = (inp[11]) ? node5942 : node5935;
										assign node5935 = (inp[7]) ? 14'b00000000011111 : node5936;
											assign node5936 = (inp[1]) ? node5938 : 14'b00000001111111;
												assign node5938 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5942 = (inp[13]) ? node5944 : 14'b00000000011111;
											assign node5944 = (inp[3]) ? 14'b00000000001111 : node5945;
												assign node5945 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node5949 = (inp[8]) ? node5961 : node5950;
										assign node5950 = (inp[7]) ? node5956 : node5951;
											assign node5951 = (inp[1]) ? 14'b00000000011111 : node5952;
												assign node5952 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5956 = (inp[11]) ? node5958 : 14'b00000000001111;
												assign node5958 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node5961 = (inp[1]) ? node5967 : node5962;
											assign node5962 = (inp[3]) ? 14'b00000000000111 : node5963;
												assign node5963 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5967 = (inp[7]) ? 14'b00000000000011 : node5968;
												assign node5968 = (inp[3]) ? node5970 : 14'b00000000000111;
													assign node5970 = (inp[13]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node5974 = (inp[13]) ? node6008 : node5975;
									assign node5975 = (inp[1]) ? node5987 : node5976;
										assign node5976 = (inp[7]) ? node5982 : node5977;
											assign node5977 = (inp[11]) ? node5979 : 14'b00000000011111;
												assign node5979 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5982 = (inp[2]) ? 14'b00000000001111 : node5983;
												assign node5983 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5987 = (inp[2]) ? node5999 : node5988;
											assign node5988 = (inp[3]) ? node5992 : node5989;
												assign node5989 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5992 = (inp[7]) ? node5994 : 14'b00000000001111;
													assign node5994 = (inp[8]) ? 14'b00000000000111 : node5995;
														assign node5995 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node5999 = (inp[11]) ? node6003 : node6000;
												assign node6000 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node6003 = (inp[8]) ? node6005 : 14'b00000000000111;
													assign node6005 = (inp[3]) ? 14'b00000000000011 : 14'b00000000000111;
									assign node6008 = (inp[8]) ? node6026 : node6009;
										assign node6009 = (inp[7]) ? node6017 : node6010;
											assign node6010 = (inp[11]) ? node6012 : 14'b00000000011111;
												assign node6012 = (inp[2]) ? node6014 : 14'b00000000001111;
													assign node6014 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node6017 = (inp[11]) ? node6021 : node6018;
												assign node6018 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node6021 = (inp[3]) ? node6023 : 14'b00000000000111;
													assign node6023 = (inp[1]) ? 14'b00000000000011 : 14'b00000000000111;
										assign node6026 = (inp[2]) ? node6042 : node6027;
											assign node6027 = (inp[3]) ? node6031 : node6028;
												assign node6028 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node6031 = (inp[1]) ? node6037 : node6032;
													assign node6032 = (inp[7]) ? node6034 : 14'b00000000000111;
														assign node6034 = (inp[11]) ? 14'b00000000000011 : 14'b00000000000111;
													assign node6037 = (inp[7]) ? 14'b00000000000011 : node6038;
														assign node6038 = (inp[11]) ? 14'b00000000000011 : 14'b00000000000111;
											assign node6042 = (inp[7]) ? node6046 : node6043;
												assign node6043 = (inp[11]) ? 14'b00000000000011 : 14'b00000000000111;
												assign node6046 = (inp[11]) ? 14'b00000000000001 : node6047;
													assign node6047 = (inp[1]) ? node6049 : 14'b00000000000011;
														assign node6049 = (inp[3]) ? 14'b00000000000001 : 14'b00000000000011;

endmodule