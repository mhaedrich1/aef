module dtc_split875_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node336;

	assign outp = (inp[3]) ? node250 : node1;
		assign node1 = (inp[9]) ? node117 : node2;
			assign node2 = (inp[4]) ? node40 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[6]) ? 3'b000 : node5;
						assign node5 = (inp[1]) ? 3'b001 : node6;
							assign node6 = (inp[5]) ? 3'b000 : 3'b001;
					assign node11 = (inp[6]) ? 3'b001 : node12;
						assign node12 = (inp[5]) ? node26 : node13;
							assign node13 = (inp[1]) ? 3'b000 : node14;
								assign node14 = (inp[11]) ? node20 : node15;
									assign node15 = (inp[2]) ? node17 : 3'b000;
										assign node17 = (inp[8]) ? 3'b001 : 3'b000;
									assign node20 = (inp[8]) ? 3'b000 : node21;
										assign node21 = (inp[2]) ? 3'b000 : 3'b001;
							assign node26 = (inp[1]) ? 3'b001 : node27;
								assign node27 = (inp[11]) ? node33 : node28;
									assign node28 = (inp[8]) ? node30 : 3'b000;
										assign node30 = (inp[2]) ? 3'b001 : 3'b000;
									assign node33 = (inp[8]) ? 3'b000 : node34;
										assign node34 = (inp[2]) ? 3'b000 : 3'b001;
				assign node40 = (inp[0]) ? node42 : 3'b000;
					assign node42 = (inp[10]) ? node98 : node43;
						assign node43 = (inp[7]) ? node67 : node44;
							assign node44 = (inp[8]) ? node56 : node45;
								assign node45 = (inp[6]) ? node51 : node46;
									assign node46 = (inp[5]) ? 3'b000 : node47;
										assign node47 = (inp[1]) ? 3'b001 : 3'b000;
									assign node51 = (inp[5]) ? node53 : 3'b000;
										assign node53 = (inp[1]) ? 3'b000 : 3'b001;
								assign node56 = (inp[5]) ? node62 : node57;
									assign node57 = (inp[6]) ? 3'b000 : node58;
										assign node58 = (inp[1]) ? 3'b001 : 3'b000;
									assign node62 = (inp[6]) ? node64 : 3'b000;
										assign node64 = (inp[1]) ? 3'b000 : 3'b001;
							assign node67 = (inp[11]) ? node87 : node68;
								assign node68 = (inp[2]) ? node76 : node69;
									assign node69 = (inp[5]) ? node71 : 3'b000;
										assign node71 = (inp[1]) ? 3'b000 : node72;
											assign node72 = (inp[6]) ? 3'b001 : 3'b000;
									assign node76 = (inp[1]) ? node82 : node77;
										assign node77 = (inp[6]) ? node79 : 3'b000;
											assign node79 = (inp[5]) ? 3'b001 : 3'b000;
										assign node82 = (inp[5]) ? 3'b000 : node83;
											assign node83 = (inp[6]) ? 3'b000 : 3'b001;
								assign node87 = (inp[5]) ? node93 : node88;
									assign node88 = (inp[6]) ? 3'b000 : node89;
										assign node89 = (inp[1]) ? 3'b001 : 3'b000;
									assign node93 = (inp[6]) ? node95 : 3'b000;
										assign node95 = (inp[1]) ? 3'b000 : 3'b001;
						assign node98 = (inp[6]) ? node112 : node99;
							assign node99 = (inp[5]) ? node107 : node100;
								assign node100 = (inp[1]) ? 3'b001 : node101;
									assign node101 = (inp[2]) ? node103 : 3'b000;
										assign node103 = (inp[7]) ? 3'b001 : 3'b000;
								assign node107 = (inp[7]) ? node109 : 3'b000;
									assign node109 = (inp[1]) ? 3'b000 : 3'b001;
							assign node112 = (inp[5]) ? node114 : 3'b000;
								assign node114 = (inp[1]) ? 3'b000 : 3'b001;
			assign node117 = (inp[6]) ? node199 : node118;
				assign node118 = (inp[4]) ? node170 : node119;
					assign node119 = (inp[0]) ? node129 : node120;
						assign node120 = (inp[5]) ? node126 : node121;
							assign node121 = (inp[7]) ? 3'b110 : node122;
								assign node122 = (inp[1]) ? 3'b110 : 3'b010;
							assign node126 = (inp[1]) ? 3'b010 : 3'b100;
						assign node129 = (inp[5]) ? node157 : node130;
							assign node130 = (inp[7]) ? node144 : node131;
								assign node131 = (inp[1]) ? 3'b001 : node132;
									assign node132 = (inp[2]) ? node138 : node133;
										assign node133 = (inp[11]) ? node135 : 3'b001;
											assign node135 = (inp[10]) ? 3'b110 : 3'b001;
										assign node138 = (inp[8]) ? node140 : 3'b001;
											assign node140 = (inp[11]) ? 3'b001 : 3'b110;
								assign node144 = (inp[1]) ? 3'b101 : node145;
									assign node145 = (inp[8]) ? node151 : node146;
										assign node146 = (inp[11]) ? node148 : 3'b001;
											assign node148 = (inp[2]) ? 3'b001 : 3'b110;
										assign node151 = (inp[11]) ? 3'b001 : node152;
											assign node152 = (inp[2]) ? 3'b110 : 3'b001;
							assign node157 = (inp[1]) ? 3'b110 : node158;
								assign node158 = (inp[2]) ? node164 : node159;
									assign node159 = (inp[8]) ? 3'b001 : node160;
										assign node160 = (inp[11]) ? 3'b110 : 3'b001;
									assign node164 = (inp[8]) ? node166 : 3'b001;
										assign node166 = (inp[11]) ? 3'b001 : 3'b110;
					assign node170 = (inp[0]) ? node182 : node171;
						assign node171 = (inp[5]) ? 3'b000 : node172;
							assign node172 = (inp[7]) ? 3'b000 : node173;
								assign node173 = (inp[1]) ? node175 : 3'b000;
									assign node175 = (inp[10]) ? node177 : 3'b000;
										assign node177 = (inp[2]) ? 3'b100 : 3'b000;
						assign node182 = (inp[5]) ? node192 : node183;
							assign node183 = (inp[1]) ? 3'b010 : node184;
								assign node184 = (inp[2]) ? node186 : 3'b100;
									assign node186 = (inp[10]) ? node188 : 3'b100;
										assign node188 = (inp[7]) ? 3'b010 : 3'b100;
							assign node192 = (inp[10]) ? node194 : 3'b100;
								assign node194 = (inp[7]) ? node196 : 3'b100;
									assign node196 = (inp[1]) ? 3'b100 : 3'b010;
				assign node199 = (inp[0]) ? node215 : node200;
					assign node200 = (inp[10]) ? node202 : 3'b001;
						assign node202 = (inp[7]) ? node204 : 3'b001;
							assign node204 = (inp[1]) ? node206 : 3'b001;
								assign node206 = (inp[2]) ? node208 : 3'b001;
									assign node208 = (inp[5]) ? 3'b001 : node209;
										assign node209 = (inp[4]) ? 3'b001 : node210;
											assign node210 = (inp[8]) ? 3'b011 : 3'b001;
					assign node215 = (inp[4]) ? node233 : node216;
						assign node216 = (inp[5]) ? node226 : node217;
							assign node217 = (inp[1]) ? 3'b111 : node218;
								assign node218 = (inp[7]) ? node220 : 3'b011;
									assign node220 = (inp[2]) ? node222 : 3'b011;
										assign node222 = (inp[10]) ? 3'b111 : 3'b011;
							assign node226 = (inp[1]) ? 3'b011 : node227;
								assign node227 = (inp[10]) ? node229 : 3'b011;
									assign node229 = (inp[7]) ? 3'b111 : 3'b011;
						assign node233 = (inp[5]) ? node243 : node234;
							assign node234 = (inp[1]) ? 3'b101 : node235;
								assign node235 = (inp[7]) ? node237 : 3'b001;
									assign node237 = (inp[2]) ? node239 : 3'b001;
										assign node239 = (inp[10]) ? 3'b101 : 3'b001;
							assign node243 = (inp[1]) ? 3'b001 : node244;
								assign node244 = (inp[7]) ? node246 : 3'b010;
									assign node246 = (inp[10]) ? 3'b110 : 3'b010;
		assign node250 = (inp[6]) ? node252 : 3'b000;
			assign node252 = (inp[0]) ? node268 : node253;
				assign node253 = (inp[4]) ? node257 : node254;
					assign node254 = (inp[9]) ? 3'b100 : 3'b000;
					assign node257 = (inp[9]) ? 3'b000 : node258;
						assign node258 = (inp[1]) ? node260 : 3'b010;
							assign node260 = (inp[10]) ? node262 : 3'b010;
								assign node262 = (inp[5]) ? 3'b100 : node263;
									assign node263 = (inp[2]) ? 3'b100 : 3'b010;
				assign node268 = (inp[4]) ? node286 : node269;
					assign node269 = (inp[9]) ? node271 : 3'b001;
						assign node271 = (inp[5]) ? 3'b010 : node272;
							assign node272 = (inp[11]) ? node274 : 3'b010;
								assign node274 = (inp[10]) ? node276 : 3'b010;
									assign node276 = (inp[8]) ? node278 : 3'b010;
										assign node278 = (inp[7]) ? node280 : 3'b010;
											assign node280 = (inp[2]) ? node282 : 3'b010;
												assign node282 = (inp[1]) ? 3'b110 : 3'b010;
					assign node286 = (inp[9]) ? node322 : node287;
						assign node287 = (inp[1]) ? node297 : node288;
							assign node288 = (inp[10]) ? 3'b010 : node289;
								assign node289 = (inp[7]) ? node291 : 3'b010;
									assign node291 = (inp[11]) ? node293 : 3'b110;
										assign node293 = (inp[2]) ? 3'b110 : 3'b010;
							assign node297 = (inp[7]) ? node299 : 3'b110;
								assign node299 = (inp[10]) ? node311 : node300;
									assign node300 = (inp[2]) ? node306 : node301;
										assign node301 = (inp[8]) ? 3'b110 : node302;
											assign node302 = (inp[11]) ? 3'b010 : 3'b110;
										assign node306 = (inp[11]) ? 3'b110 : node307;
											assign node307 = (inp[8]) ? 3'b001 : 3'b110;
									assign node311 = (inp[2]) ? node317 : node312;
										assign node312 = (inp[8]) ? 3'b010 : node313;
											assign node313 = (inp[11]) ? 3'b110 : 3'b010;
										assign node317 = (inp[11]) ? 3'b010 : node318;
											assign node318 = (inp[8]) ? 3'b110 : 3'b010;
						assign node322 = (inp[10]) ? 3'b000 : node323;
							assign node323 = (inp[7]) ? node325 : 3'b000;
								assign node325 = (inp[11]) ? node333 : node326;
									assign node326 = (inp[2]) ? node328 : 3'b100;
										assign node328 = (inp[8]) ? node330 : 3'b100;
											assign node330 = (inp[1]) ? 3'b010 : 3'b100;
									assign node333 = (inp[1]) ? node335 : 3'b000;
										assign node335 = (inp[2]) ? 3'b100 : node336;
											assign node336 = (inp[8]) ? 3'b100 : 3'b000;

endmodule