module dtc_split25_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node150 : node3;
			assign node3 = (inp[4]) ? node65 : node4;
				assign node4 = (inp[11]) ? node32 : node5;
					assign node5 = (inp[1]) ? node27 : node6;
						assign node6 = (inp[9]) ? node14 : node7;
							assign node7 = (inp[8]) ? 3'b100 : node8;
								assign node8 = (inp[3]) ? node10 : 3'b100;
									assign node10 = (inp[5]) ? 3'b100 : 3'b000;
							assign node14 = (inp[8]) ? node22 : node15;
								assign node15 = (inp[2]) ? 3'b000 : node16;
									assign node16 = (inp[5]) ? node18 : 3'b000;
										assign node18 = (inp[3]) ? 3'b100 : 3'b000;
								assign node22 = (inp[10]) ? 3'b100 : node23;
									assign node23 = (inp[3]) ? 3'b000 : 3'b100;
						assign node27 = (inp[9]) ? node29 : 3'b000;
							assign node29 = (inp[8]) ? 3'b000 : 3'b100;
					assign node32 = (inp[9]) ? node42 : node33;
						assign node33 = (inp[8]) ? node35 : 3'b000;
							assign node35 = (inp[1]) ? 3'b000 : node36;
								assign node36 = (inp[7]) ? node38 : 3'b100;
									assign node38 = (inp[10]) ? 3'b100 : 3'b000;
						assign node42 = (inp[1]) ? node58 : node43;
							assign node43 = (inp[7]) ? node49 : node44;
								assign node44 = (inp[8]) ? 3'b000 : node45;
									assign node45 = (inp[5]) ? 3'b100 : 3'b000;
								assign node49 = (inp[3]) ? 3'b100 : node50;
									assign node50 = (inp[5]) ? node52 : 3'b000;
										assign node52 = (inp[10]) ? 3'b100 : node53;
											assign node53 = (inp[2]) ? 3'b000 : 3'b100;
							assign node58 = (inp[10]) ? node60 : 3'b100;
								assign node60 = (inp[8]) ? node62 : 3'b100;
									assign node62 = (inp[2]) ? 3'b000 : 3'b100;
				assign node65 = (inp[9]) ? node85 : node66;
					assign node66 = (inp[1]) ? node68 : 3'b100;
						assign node68 = (inp[11]) ? node76 : node69;
							assign node69 = (inp[3]) ? node71 : 3'b100;
								assign node71 = (inp[8]) ? 3'b100 : node72;
									assign node72 = (inp[10]) ? 3'b100 : 3'b000;
							assign node76 = (inp[8]) ? node78 : 3'b000;
								assign node78 = (inp[7]) ? 3'b000 : node79;
									assign node79 = (inp[3]) ? node81 : 3'b100;
										assign node81 = (inp[10]) ? 3'b100 : 3'b000;
					assign node85 = (inp[1]) ? node121 : node86;
						assign node86 = (inp[8]) ? node108 : node87;
							assign node87 = (inp[10]) ? node95 : node88;
								assign node88 = (inp[7]) ? 3'b001 : node89;
									assign node89 = (inp[11]) ? node91 : 3'b001;
										assign node91 = (inp[5]) ? 3'b001 : 3'b100;
								assign node95 = (inp[3]) ? node101 : node96;
									assign node96 = (inp[7]) ? 3'b101 : node97;
										assign node97 = (inp[5]) ? 3'b101 : 3'b001;
									assign node101 = (inp[11]) ? node103 : 3'b101;
										assign node103 = (inp[2]) ? 3'b001 : node104;
											assign node104 = (inp[7]) ? 3'b001 : 3'b101;
							assign node108 = (inp[2]) ? node118 : node109;
								assign node109 = (inp[10]) ? node113 : node110;
									assign node110 = (inp[11]) ? 3'b100 : 3'b000;
									assign node113 = (inp[7]) ? node115 : 3'b111;
										assign node115 = (inp[11]) ? 3'b010 : 3'b011;
								assign node118 = (inp[10]) ? 3'b000 : 3'b001;
						assign node121 = (inp[8]) ? node135 : node122;
							assign node122 = (inp[10]) ? node128 : node123;
								assign node123 = (inp[3]) ? node125 : 3'b100;
									assign node125 = (inp[11]) ? 3'b000 : 3'b100;
								assign node128 = (inp[11]) ? node132 : node129;
									assign node129 = (inp[2]) ? 3'b101 : 3'b001;
									assign node132 = (inp[2]) ? 3'b001 : 3'b100;
							assign node135 = (inp[2]) ? node145 : node136;
								assign node136 = (inp[10]) ? node142 : node137;
									assign node137 = (inp[3]) ? 3'b101 : node138;
										assign node138 = (inp[11]) ? 3'b001 : 3'b101;
									assign node142 = (inp[5]) ? 3'b110 : 3'b011;
								assign node145 = (inp[11]) ? node147 : 3'b000;
									assign node147 = (inp[3]) ? 3'b000 : 3'b100;
			assign node150 = (inp[9]) ? node152 : 3'b000;
				assign node152 = (inp[1]) ? node220 : node153;
					assign node153 = (inp[4]) ? node169 : node154;
						assign node154 = (inp[8]) ? node162 : node155;
							assign node155 = (inp[11]) ? 3'b000 : node156;
								assign node156 = (inp[3]) ? node158 : 3'b100;
									assign node158 = (inp[7]) ? 3'b000 : 3'b100;
							assign node162 = (inp[3]) ? node164 : 3'b100;
								assign node164 = (inp[11]) ? node166 : 3'b100;
									assign node166 = (inp[2]) ? 3'b000 : 3'b100;
						assign node169 = (inp[8]) ? node197 : node170;
							assign node170 = (inp[5]) ? node184 : node171;
								assign node171 = (inp[2]) ? node173 : 3'b000;
									assign node173 = (inp[3]) ? 3'b000 : node174;
										assign node174 = (inp[7]) ? node176 : 3'b000;
											assign node176 = (inp[11]) ? node180 : node177;
												assign node177 = (inp[10]) ? 3'b100 : 3'b000;
												assign node180 = (inp[10]) ? 3'b000 : 3'b100;
								assign node184 = (inp[3]) ? 3'b100 : node185;
									assign node185 = (inp[7]) ? node191 : node186;
										assign node186 = (inp[11]) ? 3'b000 : node187;
											assign node187 = (inp[10]) ? 3'b100 : 3'b000;
										assign node191 = (inp[10]) ? 3'b100 : node192;
											assign node192 = (inp[11]) ? 3'b100 : 3'b000;
							assign node197 = (inp[11]) ? node209 : node198;
								assign node198 = (inp[10]) ? node204 : node199;
									assign node199 = (inp[3]) ? 3'b001 : node200;
										assign node200 = (inp[2]) ? 3'b101 : 3'b001;
									assign node204 = (inp[2]) ? 3'b000 : node205;
										assign node205 = (inp[3]) ? 3'b001 : 3'b101;
								assign node209 = (inp[2]) ? node217 : node210;
									assign node210 = (inp[7]) ? node212 : 3'b100;
										assign node212 = (inp[5]) ? node214 : 3'b000;
											assign node214 = (inp[10]) ? 3'b000 : 3'b100;
									assign node217 = (inp[3]) ? 3'b001 : 3'b101;
					assign node220 = (inp[4]) ? node222 : 3'b000;
						assign node222 = (inp[11]) ? node244 : node223;
							assign node223 = (inp[8]) ? node229 : node224;
								assign node224 = (inp[3]) ? node226 : 3'b100;
									assign node226 = (inp[10]) ? 3'b100 : 3'b000;
								assign node229 = (inp[10]) ? node239 : node230;
									assign node230 = (inp[7]) ? 3'b100 : node231;
										assign node231 = (inp[2]) ? node235 : node232;
											assign node232 = (inp[5]) ? 3'b000 : 3'b100;
											assign node235 = (inp[3]) ? 3'b000 : 3'b100;
									assign node239 = (inp[2]) ? 3'b000 : node240;
										assign node240 = (inp[3]) ? 3'b001 : 3'b101;
							assign node244 = (inp[8]) ? node246 : 3'b000;
								assign node246 = (inp[2]) ? 3'b000 : node247;
									assign node247 = (inp[7]) ? 3'b000 : 3'b100;

endmodule