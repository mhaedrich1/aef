module dtc_split33_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node229;

	assign outp = (inp[3]) ? node168 : node1;
		assign node1 = (inp[9]) ? node49 : node2;
			assign node2 = (inp[4]) ? node32 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[6]) ? 3'b000 : node5;
						assign node5 = (inp[1]) ? 3'b001 : node6;
							assign node6 = (inp[5]) ? 3'b000 : 3'b001;
					assign node11 = (inp[6]) ? 3'b001 : node12;
						assign node12 = (inp[5]) ? node24 : node13;
							assign node13 = (inp[1]) ? 3'b000 : node14;
								assign node14 = (inp[2]) ? node18 : node15;
									assign node15 = (inp[8]) ? 3'b000 : 3'b001;
									assign node18 = (inp[7]) ? 3'b000 : node19;
										assign node19 = (inp[8]) ? 3'b001 : 3'b000;
							assign node24 = (inp[1]) ? 3'b001 : node25;
								assign node25 = (inp[7]) ? 3'b000 : node26;
									assign node26 = (inp[8]) ? 3'b000 : 3'b001;
				assign node32 = (inp[0]) ? node34 : 3'b000;
					assign node34 = (inp[6]) ? node44 : node35;
						assign node35 = (inp[1]) ? node41 : node36;
							assign node36 = (inp[7]) ? node38 : 3'b000;
								assign node38 = (inp[10]) ? 3'b001 : 3'b000;
							assign node41 = (inp[5]) ? 3'b000 : 3'b001;
						assign node44 = (inp[1]) ? 3'b000 : node45;
							assign node45 = (inp[5]) ? 3'b001 : 3'b000;
			assign node49 = (inp[6]) ? node125 : node50;
				assign node50 = (inp[4]) ? node96 : node51;
					assign node51 = (inp[0]) ? node61 : node52;
						assign node52 = (inp[5]) ? node58 : node53;
							assign node53 = (inp[7]) ? 3'b110 : node54;
								assign node54 = (inp[1]) ? 3'b110 : 3'b010;
							assign node58 = (inp[1]) ? 3'b010 : 3'b100;
						assign node61 = (inp[5]) ? node77 : node62;
							assign node62 = (inp[1]) ? node74 : node63;
								assign node63 = (inp[7]) ? 3'b001 : node64;
									assign node64 = (inp[10]) ? node66 : 3'b001;
										assign node66 = (inp[2]) ? node70 : node67;
											assign node67 = (inp[11]) ? 3'b000 : 3'b001;
											assign node70 = (inp[8]) ? 3'b000 : 3'b001;
								assign node74 = (inp[7]) ? 3'b101 : 3'b001;
							assign node77 = (inp[1]) ? 3'b110 : node78;
								assign node78 = (inp[10]) ? node88 : node79;
									assign node79 = (inp[8]) ? node83 : node80;
										assign node80 = (inp[11]) ? 3'b110 : 3'b001;
										assign node83 = (inp[11]) ? 3'b001 : node84;
											assign node84 = (inp[2]) ? 3'b110 : 3'b001;
									assign node88 = (inp[7]) ? node90 : 3'b001;
										assign node90 = (inp[8]) ? node92 : 3'b110;
											assign node92 = (inp[2]) ? 3'b110 : 3'b001;
					assign node96 = (inp[0]) ? node106 : node97;
						assign node97 = (inp[7]) ? 3'b000 : node98;
							assign node98 = (inp[10]) ? node100 : 3'b000;
								assign node100 = (inp[5]) ? 3'b000 : node101;
									assign node101 = (inp[8]) ? 3'b000 : 3'b100;
						assign node106 = (inp[5]) ? node116 : node107;
							assign node107 = (inp[1]) ? 3'b010 : node108;
								assign node108 = (inp[2]) ? node110 : 3'b100;
									assign node110 = (inp[10]) ? node112 : 3'b100;
										assign node112 = (inp[7]) ? 3'b010 : 3'b100;
							assign node116 = (inp[7]) ? node118 : 3'b100;
								assign node118 = (inp[2]) ? node120 : 3'b100;
									assign node120 = (inp[10]) ? node122 : 3'b100;
										assign node122 = (inp[1]) ? 3'b100 : 3'b010;
				assign node125 = (inp[0]) ? node139 : node126;
					assign node126 = (inp[1]) ? node128 : 3'b001;
						assign node128 = (inp[11]) ? node130 : 3'b001;
							assign node130 = (inp[2]) ? node132 : 3'b001;
								assign node132 = (inp[4]) ? 3'b001 : node133;
									assign node133 = (inp[5]) ? 3'b001 : node134;
										assign node134 = (inp[7]) ? 3'b011 : 3'b001;
					assign node139 = (inp[4]) ? node153 : node140;
						assign node140 = (inp[1]) ? node150 : node141;
							assign node141 = (inp[10]) ? node143 : 3'b011;
								assign node143 = (inp[7]) ? node145 : 3'b011;
									assign node145 = (inp[2]) ? 3'b111 : node146;
										assign node146 = (inp[5]) ? 3'b111 : 3'b011;
							assign node150 = (inp[5]) ? 3'b011 : 3'b111;
						assign node153 = (inp[1]) ? node165 : node154;
							assign node154 = (inp[5]) ? node160 : node155;
								assign node155 = (inp[7]) ? node157 : 3'b001;
									assign node157 = (inp[2]) ? 3'b101 : 3'b001;
								assign node160 = (inp[7]) ? node162 : 3'b010;
									assign node162 = (inp[10]) ? 3'b110 : 3'b010;
							assign node165 = (inp[5]) ? 3'b001 : 3'b101;
		assign node168 = (inp[6]) ? node170 : 3'b000;
			assign node170 = (inp[0]) ? node184 : node171;
				assign node171 = (inp[4]) ? node175 : node172;
					assign node172 = (inp[9]) ? 3'b100 : 3'b000;
					assign node175 = (inp[9]) ? 3'b000 : node176;
						assign node176 = (inp[1]) ? node178 : 3'b010;
							assign node178 = (inp[10]) ? node180 : 3'b010;
								assign node180 = (inp[5]) ? 3'b100 : 3'b010;
				assign node184 = (inp[4]) ? node196 : node185;
					assign node185 = (inp[9]) ? node187 : 3'b001;
						assign node187 = (inp[2]) ? node189 : 3'b010;
							assign node189 = (inp[1]) ? node191 : 3'b010;
								assign node191 = (inp[8]) ? node193 : 3'b010;
									assign node193 = (inp[11]) ? 3'b110 : 3'b010;
					assign node196 = (inp[9]) ? node218 : node197;
						assign node197 = (inp[1]) ? node207 : node198;
							assign node198 = (inp[10]) ? 3'b010 : node199;
								assign node199 = (inp[7]) ? node201 : 3'b010;
									assign node201 = (inp[11]) ? node203 : 3'b110;
										assign node203 = (inp[2]) ? 3'b110 : 3'b010;
							assign node207 = (inp[7]) ? node209 : 3'b110;
								assign node209 = (inp[10]) ? node213 : node210;
									assign node210 = (inp[2]) ? 3'b001 : 3'b110;
									assign node213 = (inp[11]) ? 3'b010 : node214;
										assign node214 = (inp[8]) ? 3'b110 : 3'b010;
						assign node218 = (inp[10]) ? 3'b000 : node219;
							assign node219 = (inp[7]) ? node221 : 3'b000;
								assign node221 = (inp[11]) ? node227 : node222;
									assign node222 = (inp[1]) ? node224 : 3'b100;
										assign node224 = (inp[8]) ? 3'b010 : 3'b100;
									assign node227 = (inp[8]) ? node229 : 3'b000;
										assign node229 = (inp[1]) ? 3'b100 : 3'b000;

endmodule