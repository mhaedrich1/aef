module dtc_split66_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node27;
	wire [4-1:0] node29;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node45;
	wire [4-1:0] node47;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node55;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node65;
	wire [4-1:0] node67;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node78;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node95;
	wire [4-1:0] node98;
	wire [4-1:0] node100;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node113;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node118;
	wire [4-1:0] node120;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node134;
	wire [4-1:0] node136;
	wire [4-1:0] node138;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node156;
	wire [4-1:0] node158;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node181;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node192;
	wire [4-1:0] node194;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node216;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node271;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node277;
	wire [4-1:0] node280;
	wire [4-1:0] node281;
	wire [4-1:0] node285;
	wire [4-1:0] node286;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node290;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node304;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node317;
	wire [4-1:0] node320;
	wire [4-1:0] node322;
	wire [4-1:0] node325;
	wire [4-1:0] node327;
	wire [4-1:0] node329;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node339;
	wire [4-1:0] node343;
	wire [4-1:0] node345;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node355;
	wire [4-1:0] node356;
	wire [4-1:0] node359;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node365;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node381;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node405;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node430;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node436;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node443;
	wire [4-1:0] node447;
	wire [4-1:0] node449;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node481;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node499;
	wire [4-1:0] node501;
	wire [4-1:0] node502;
	wire [4-1:0] node505;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node520;
	wire [4-1:0] node522;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node532;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node546;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node569;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node587;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node605;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node613;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node626;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node632;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node664;
	wire [4-1:0] node667;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node688;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node694;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node704;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node723;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node728;
	wire [4-1:0] node732;
	wire [4-1:0] node734;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node745;
	wire [4-1:0] node746;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node757;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node768;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node798;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node806;
	wire [4-1:0] node810;
	wire [4-1:0] node812;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node822;
	wire [4-1:0] node826;
	wire [4-1:0] node828;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node836;
	wire [4-1:0] node839;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node877;
	wire [4-1:0] node879;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node886;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node894;
	wire [4-1:0] node896;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node914;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node939;
	wire [4-1:0] node941;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node956;
	wire [4-1:0] node958;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node967;
	wire [4-1:0] node969;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node986;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1007;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1018;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1030;
	wire [4-1:0] node1032;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1058;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1107;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1129;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1139;
	wire [4-1:0] node1141;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1159;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1181;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1195;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1210;
	wire [4-1:0] node1213;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1220;
	wire [4-1:0] node1224;
	wire [4-1:0] node1226;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1234;
	wire [4-1:0] node1237;
	wire [4-1:0] node1239;
	wire [4-1:0] node1242;
	wire [4-1:0] node1244;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1251;
	wire [4-1:0] node1252;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1275;
	wire [4-1:0] node1277;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1298;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1313;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1341;
	wire [4-1:0] node1343;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1353;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1368;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1387;
	wire [4-1:0] node1388;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1418;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1448;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1456;
	wire [4-1:0] node1458;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1465;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1471;
	wire [4-1:0] node1473;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1484;
	wire [4-1:0] node1486;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1503;
	wire [4-1:0] node1504;
	wire [4-1:0] node1507;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1517;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1524;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1538;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1552;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1564;
	wire [4-1:0] node1566;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1573;
	wire [4-1:0] node1576;
	wire [4-1:0] node1577;
	wire [4-1:0] node1579;
	wire [4-1:0] node1582;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1590;
	wire [4-1:0] node1592;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1604;
	wire [4-1:0] node1607;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1618;
	wire [4-1:0] node1621;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1630;
	wire [4-1:0] node1632;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1652;
	wire [4-1:0] node1653;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1667;
	wire [4-1:0] node1670;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1676;
	wire [4-1:0] node1679;
	wire [4-1:0] node1681;
	wire [4-1:0] node1684;
	wire [4-1:0] node1685;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1691;
	wire [4-1:0] node1692;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1702;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1712;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1718;
	wire [4-1:0] node1721;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1734;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1751;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1772;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1783;
	wire [4-1:0] node1784;
	wire [4-1:0] node1787;
	wire [4-1:0] node1788;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1804;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1817;
	wire [4-1:0] node1818;
	wire [4-1:0] node1821;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1827;
	wire [4-1:0] node1830;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1836;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1898;
	wire [4-1:0] node1901;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1909;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1931;
	wire [4-1:0] node1934;
	wire [4-1:0] node1937;
	wire [4-1:0] node1939;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1945;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1955;
	wire [4-1:0] node1957;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1979;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1996;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2017;
	wire [4-1:0] node2018;
	wire [4-1:0] node2019;
	wire [4-1:0] node2020;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2038;
	wire [4-1:0] node2041;
	wire [4-1:0] node2042;
	wire [4-1:0] node2045;
	wire [4-1:0] node2047;
	wire [4-1:0] node2050;
	wire [4-1:0] node2051;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2054;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2063;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2070;
	wire [4-1:0] node2073;
	wire [4-1:0] node2075;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2085;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2108;
	wire [4-1:0] node2109;
	wire [4-1:0] node2112;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2118;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2150;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2160;
	wire [4-1:0] node2161;
	wire [4-1:0] node2164;
	wire [4-1:0] node2167;
	wire [4-1:0] node2168;
	wire [4-1:0] node2170;
	wire [4-1:0] node2173;
	wire [4-1:0] node2175;
	wire [4-1:0] node2178;
	wire [4-1:0] node2179;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2184;
	wire [4-1:0] node2187;
	wire [4-1:0] node2190;
	wire [4-1:0] node2191;
	wire [4-1:0] node2192;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2204;
	wire [4-1:0] node2206;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2218;
	wire [4-1:0] node2221;
	wire [4-1:0] node2222;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2245;
	wire [4-1:0] node2247;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2261;
	wire [4-1:0] node2263;
	wire [4-1:0] node2266;
	wire [4-1:0] node2267;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2273;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2279;
	wire [4-1:0] node2280;
	wire [4-1:0] node2281;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2295;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2311;
	wire [4-1:0] node2312;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2324;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2328;
	wire [4-1:0] node2331;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2343;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2359;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2365;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2374;
	wire [4-1:0] node2375;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2385;
	wire [4-1:0] node2387;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2393;
	wire [4-1:0] node2397;
	wire [4-1:0] node2398;
	wire [4-1:0] node2399;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2414;
	wire [4-1:0] node2416;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2422;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2429;
	wire [4-1:0] node2430;
	wire [4-1:0] node2431;
	wire [4-1:0] node2433;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2439;
	wire [4-1:0] node2441;
	wire [4-1:0] node2444;
	wire [4-1:0] node2446;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2452;
	wire [4-1:0] node2455;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2461;
	wire [4-1:0] node2462;
	wire [4-1:0] node2465;
	wire [4-1:0] node2467;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2473;
	wire [4-1:0] node2476;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2483;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2487;
	wire [4-1:0] node2488;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2495;
	wire [4-1:0] node2497;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2514;
	wire [4-1:0] node2516;
	wire [4-1:0] node2518;
	wire [4-1:0] node2521;
	wire [4-1:0] node2522;
	wire [4-1:0] node2525;
	wire [4-1:0] node2528;
	wire [4-1:0] node2529;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2546;
	wire [4-1:0] node2550;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2560;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2565;
	wire [4-1:0] node2566;
	wire [4-1:0] node2567;
	wire [4-1:0] node2569;
	wire [4-1:0] node2571;
	wire [4-1:0] node2574;
	wire [4-1:0] node2576;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2582;
	wire [4-1:0] node2585;
	wire [4-1:0] node2586;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2594;
	wire [4-1:0] node2597;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2603;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2616;
	wire [4-1:0] node2617;
	wire [4-1:0] node2618;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2635;
	wire [4-1:0] node2638;
	wire [4-1:0] node2640;
	wire [4-1:0] node2643;
	wire [4-1:0] node2644;
	wire [4-1:0] node2645;
	wire [4-1:0] node2648;
	wire [4-1:0] node2651;
	wire [4-1:0] node2652;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2659;
	wire [4-1:0] node2660;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2670;
	wire [4-1:0] node2672;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2681;
	wire [4-1:0] node2684;
	wire [4-1:0] node2685;
	wire [4-1:0] node2689;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2702;
	wire [4-1:0] node2706;
	wire [4-1:0] node2708;
	wire [4-1:0] node2711;
	wire [4-1:0] node2713;
	wire [4-1:0] node2715;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2724;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2729;
	wire [4-1:0] node2733;
	wire [4-1:0] node2735;
	wire [4-1:0] node2738;
	wire [4-1:0] node2739;
	wire [4-1:0] node2741;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2751;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2762;
	wire [4-1:0] node2765;
	wire [4-1:0] node2767;
	wire [4-1:0] node2770;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2783;
	wire [4-1:0] node2784;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2791;
	wire [4-1:0] node2794;
	wire [4-1:0] node2795;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2808;
	wire [4-1:0] node2811;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2816;
	wire [4-1:0] node2820;
	wire [4-1:0] node2821;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2825;
	wire [4-1:0] node2828;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2835;
	wire [4-1:0] node2838;
	wire [4-1:0] node2839;
	wire [4-1:0] node2841;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2849;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2863;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2868;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2875;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2881;
	wire [4-1:0] node2883;
	wire [4-1:0] node2887;
	wire [4-1:0] node2888;
	wire [4-1:0] node2890;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2900;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2906;
	wire [4-1:0] node2909;
	wire [4-1:0] node2910;
	wire [4-1:0] node2913;
	wire [4-1:0] node2916;
	wire [4-1:0] node2917;
	wire [4-1:0] node2918;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2938;
	wire [4-1:0] node2939;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2947;
	wire [4-1:0] node2948;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2959;
	wire [4-1:0] node2961;
	wire [4-1:0] node2964;
	wire [4-1:0] node2966;
	wire [4-1:0] node2968;
	wire [4-1:0] node2971;
	wire [4-1:0] node2972;
	wire [4-1:0] node2973;
	wire [4-1:0] node2974;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2983;
	wire [4-1:0] node2985;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2995;
	wire [4-1:0] node2996;
	wire [4-1:0] node2998;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3008;
	wire [4-1:0] node3010;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3015;
	wire [4-1:0] node3018;
	wire [4-1:0] node3020;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3026;
	wire [4-1:0] node3029;
	wire [4-1:0] node3031;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3038;
	wire [4-1:0] node3041;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3047;
	wire [4-1:0] node3050;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3055;
	wire [4-1:0] node3058;
	wire [4-1:0] node3060;
	wire [4-1:0] node3063;
	wire [4-1:0] node3064;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3072;
	wire [4-1:0] node3073;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3080;
	wire [4-1:0] node3084;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3092;
	wire [4-1:0] node3095;
	wire [4-1:0] node3096;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3107;
	wire [4-1:0] node3109;
	wire [4-1:0] node3110;
	wire [4-1:0] node3114;
	wire [4-1:0] node3115;
	wire [4-1:0] node3118;
	wire [4-1:0] node3120;
	wire [4-1:0] node3123;
	wire [4-1:0] node3124;
	wire [4-1:0] node3125;
	wire [4-1:0] node3126;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3131;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3139;
	wire [4-1:0] node3140;
	wire [4-1:0] node3143;
	wire [4-1:0] node3146;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3153;
	wire [4-1:0] node3154;
	wire [4-1:0] node3155;
	wire [4-1:0] node3160;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3164;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3173;
	wire [4-1:0] node3174;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3180;
	wire [4-1:0] node3182;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3190;
	wire [4-1:0] node3191;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3197;
	wire [4-1:0] node3198;
	wire [4-1:0] node3201;
	wire [4-1:0] node3202;
	wire [4-1:0] node3207;
	wire [4-1:0] node3208;
	wire [4-1:0] node3210;
	wire [4-1:0] node3213;
	wire [4-1:0] node3217;
	wire [4-1:0] node3218;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3222;
	wire [4-1:0] node3223;
	wire [4-1:0] node3224;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3231;
	wire [4-1:0] node3234;
	wire [4-1:0] node3237;
	wire [4-1:0] node3239;
	wire [4-1:0] node3240;
	wire [4-1:0] node3242;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3249;
	wire [4-1:0] node3251;
	wire [4-1:0] node3252;
	wire [4-1:0] node3255;
	wire [4-1:0] node3258;
	wire [4-1:0] node3259;
	wire [4-1:0] node3261;
	wire [4-1:0] node3263;
	wire [4-1:0] node3266;
	wire [4-1:0] node3267;
	wire [4-1:0] node3270;
	wire [4-1:0] node3272;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3278;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3291;
	wire [4-1:0] node3293;
	wire [4-1:0] node3296;
	wire [4-1:0] node3298;
	wire [4-1:0] node3301;
	wire [4-1:0] node3302;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3313;
	wire [4-1:0] node3317;
	wire [4-1:0] node3319;
	wire [4-1:0] node3322;
	wire [4-1:0] node3323;
	wire [4-1:0] node3324;
	wire [4-1:0] node3326;
	wire [4-1:0] node3327;
	wire [4-1:0] node3331;
	wire [4-1:0] node3333;
	wire [4-1:0] node3336;
	wire [4-1:0] node3337;
	wire [4-1:0] node3339;
	wire [4-1:0] node3344;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3351;
	wire [4-1:0] node3352;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3362;
	wire [4-1:0] node3365;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3370;
	wire [4-1:0] node3373;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3379;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3384;
	wire [4-1:0] node3385;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3393;
	wire [4-1:0] node3394;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3402;
	wire [4-1:0] node3403;
	wire [4-1:0] node3405;
	wire [4-1:0] node3408;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3413;
	wire [4-1:0] node3414;
	wire [4-1:0] node3417;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3439;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3459;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3466;
	wire [4-1:0] node3467;
	wire [4-1:0] node3471;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3474;
	wire [4-1:0] node3477;
	wire [4-1:0] node3480;
	wire [4-1:0] node3481;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3489;
	wire [4-1:0] node3491;
	wire [4-1:0] node3494;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3505;
	wire [4-1:0] node3506;
	wire [4-1:0] node3508;
	wire [4-1:0] node3509;
	wire [4-1:0] node3513;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3526;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3532;
	wire [4-1:0] node3534;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3541;
	wire [4-1:0] node3542;
	wire [4-1:0] node3543;
	wire [4-1:0] node3546;
	wire [4-1:0] node3549;
	wire [4-1:0] node3550;
	wire [4-1:0] node3553;
	wire [4-1:0] node3556;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3561;
	wire [4-1:0] node3562;
	wire [4-1:0] node3565;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3579;
	wire [4-1:0] node3582;
	wire [4-1:0] node3584;
	wire [4-1:0] node3587;
	wire [4-1:0] node3588;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3595;
	wire [4-1:0] node3597;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3606;
	wire [4-1:0] node3607;
	wire [4-1:0] node3609;
	wire [4-1:0] node3612;
	wire [4-1:0] node3614;
	wire [4-1:0] node3617;
	wire [4-1:0] node3618;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3631;
	wire [4-1:0] node3632;
	wire [4-1:0] node3636;
	wire [4-1:0] node3637;
	wire [4-1:0] node3640;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3649;
	wire [4-1:0] node3651;
	wire [4-1:0] node3654;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3659;
	wire [4-1:0] node3662;
	wire [4-1:0] node3665;
	wire [4-1:0] node3666;
	wire [4-1:0] node3669;
	wire [4-1:0] node3672;
	wire [4-1:0] node3673;
	wire [4-1:0] node3674;
	wire [4-1:0] node3675;
	wire [4-1:0] node3678;
	wire [4-1:0] node3681;
	wire [4-1:0] node3683;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3691;
	wire [4-1:0] node3694;
	wire [4-1:0] node3695;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3702;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3708;
	wire [4-1:0] node3709;
	wire [4-1:0] node3711;
	wire [4-1:0] node3714;
	wire [4-1:0] node3715;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3723;
	wire [4-1:0] node3726;
	wire [4-1:0] node3727;
	wire [4-1:0] node3728;
	wire [4-1:0] node3732;
	wire [4-1:0] node3733;
	wire [4-1:0] node3735;
	wire [4-1:0] node3738;
	wire [4-1:0] node3741;
	wire [4-1:0] node3742;
	wire [4-1:0] node3743;
	wire [4-1:0] node3744;
	wire [4-1:0] node3746;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3753;
	wire [4-1:0] node3756;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3761;
	wire [4-1:0] node3764;
	wire [4-1:0] node3766;
	wire [4-1:0] node3769;
	wire [4-1:0] node3771;
	wire [4-1:0] node3774;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3786;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3794;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3798;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3806;
	wire [4-1:0] node3807;
	wire [4-1:0] node3809;
	wire [4-1:0] node3812;
	wire [4-1:0] node3815;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3818;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3825;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3838;
	wire [4-1:0] node3841;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3847;
	wire [4-1:0] node3848;
	wire [4-1:0] node3851;
	wire [4-1:0] node3853;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3861;
	wire [4-1:0] node3864;
	wire [4-1:0] node3865;
	wire [4-1:0] node3868;
	wire [4-1:0] node3871;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3881;
	wire [4-1:0] node3882;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3888;
	wire [4-1:0] node3891;
	wire [4-1:0] node3894;
	wire [4-1:0] node3895;
	wire [4-1:0] node3897;
	wire [4-1:0] node3900;
	wire [4-1:0] node3901;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3911;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3920;
	wire [4-1:0] node3922;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3929;
	wire [4-1:0] node3932;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3940;
	wire [4-1:0] node3941;
	wire [4-1:0] node3942;
	wire [4-1:0] node3943;
	wire [4-1:0] node3947;
	wire [4-1:0] node3948;
	wire [4-1:0] node3950;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3965;
	wire [4-1:0] node3968;
	wire [4-1:0] node3969;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3976;
	wire [4-1:0] node3977;
	wire [4-1:0] node3980;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3987;
	wire [4-1:0] node3990;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3997;
	wire [4-1:0] node4000;
	wire [4-1:0] node4003;
	wire [4-1:0] node4005;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4014;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4023;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4031;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4036;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4047;
	wire [4-1:0] node4049;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4060;
	wire [4-1:0] node4063;
	wire [4-1:0] node4065;
	wire [4-1:0] node4069;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4075;
	wire [4-1:0] node4076;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4081;
	wire [4-1:0] node4085;
	wire [4-1:0] node4087;
	wire [4-1:0] node4088;
	wire [4-1:0] node4091;
	wire [4-1:0] node4094;
	wire [4-1:0] node4095;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4107;
	wire [4-1:0] node4108;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4118;
	wire [4-1:0] node4121;
	wire [4-1:0] node4122;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4128;
	wire [4-1:0] node4131;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4136;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4143;
	wire [4-1:0] node4146;
	wire [4-1:0] node4148;
	wire [4-1:0] node4151;
	wire [4-1:0] node4152;
	wire [4-1:0] node4153;
	wire [4-1:0] node4154;
	wire [4-1:0] node4159;
	wire [4-1:0] node4160;
	wire [4-1:0] node4162;
	wire [4-1:0] node4165;
	wire [4-1:0] node4168;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4173;
	wire [4-1:0] node4175;
	wire [4-1:0] node4176;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4185;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4191;
	wire [4-1:0] node4195;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4202;
	wire [4-1:0] node4203;
	wire [4-1:0] node4207;
	wire [4-1:0] node4208;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4216;
	wire [4-1:0] node4217;
	wire [4-1:0] node4218;
	wire [4-1:0] node4220;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4229;
	wire [4-1:0] node4230;
	wire [4-1:0] node4234;
	wire [4-1:0] node4235;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4241;
	wire [4-1:0] node4242;
	wire [4-1:0] node4244;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4251;
	wire [4-1:0] node4252;
	wire [4-1:0] node4256;
	wire [4-1:0] node4257;
	wire [4-1:0] node4258;
	wire [4-1:0] node4260;
	wire [4-1:0] node4263;
	wire [4-1:0] node4266;
	wire [4-1:0] node4268;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4274;
	wire [4-1:0] node4277;
	wire [4-1:0] node4278;
	wire [4-1:0] node4283;
	wire [4-1:0] node4285;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4294;
	wire [4-1:0] node4298;
	wire [4-1:0] node4301;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4311;
	wire [4-1:0] node4312;
	wire [4-1:0] node4315;
	wire [4-1:0] node4317;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4324;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4330;
	wire [4-1:0] node4331;
	wire [4-1:0] node4334;
	wire [4-1:0] node4335;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4341;
	wire [4-1:0] node4344;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4368;
	wire [4-1:0] node4370;
	wire [4-1:0] node4373;
	wire [4-1:0] node4374;
	wire [4-1:0] node4376;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4384;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4391;
	wire [4-1:0] node4392;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4401;
	wire [4-1:0] node4402;
	wire [4-1:0] node4403;
	wire [4-1:0] node4405;
	wire [4-1:0] node4408;
	wire [4-1:0] node4409;
	wire [4-1:0] node4413;
	wire [4-1:0] node4414;
	wire [4-1:0] node4417;
	wire [4-1:0] node4418;
	wire [4-1:0] node4423;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4428;
	wire [4-1:0] node4430;
	wire [4-1:0] node4431;
	wire [4-1:0] node4435;
	wire [4-1:0] node4436;
	wire [4-1:0] node4437;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4446;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4449;
	wire [4-1:0] node4452;
	wire [4-1:0] node4455;
	wire [4-1:0] node4457;
	wire [4-1:0] node4460;
	wire [4-1:0] node4463;
	wire [4-1:0] node4464;
	wire [4-1:0] node4465;
	wire [4-1:0] node4466;
	wire [4-1:0] node4467;
	wire [4-1:0] node4468;
	wire [4-1:0] node4471;
	wire [4-1:0] node4474;
	wire [4-1:0] node4475;
	wire [4-1:0] node4479;
	wire [4-1:0] node4480;
	wire [4-1:0] node4483;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4493;
	wire [4-1:0] node4496;
	wire [4-1:0] node4498;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4507;
	wire [4-1:0] node4510;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4520;
	wire [4-1:0] node4523;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4531;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4541;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4545;
	wire [4-1:0] node4548;
	wire [4-1:0] node4549;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4557;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4562;
	wire [4-1:0] node4563;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4573;
	wire [4-1:0] node4576;
	wire [4-1:0] node4579;
	wire [4-1:0] node4580;
	wire [4-1:0] node4585;
	wire [4-1:0] node4586;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4593;
	wire [4-1:0] node4595;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4602;
	wire [4-1:0] node4603;
	wire [4-1:0] node4607;
	wire [4-1:0] node4608;
	wire [4-1:0] node4610;
	wire [4-1:0] node4612;
	wire [4-1:0] node4615;
	wire [4-1:0] node4616;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4628;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4634;
	wire [4-1:0] node4638;
	wire [4-1:0] node4639;
	wire [4-1:0] node4641;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4652;
	wire [4-1:0] node4654;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4661;
	wire [4-1:0] node4662;
	wire [4-1:0] node4666;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4671;
	wire [4-1:0] node4674;
	wire [4-1:0] node4676;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4682;
	wire [4-1:0] node4683;
	wire [4-1:0] node4684;
	wire [4-1:0] node4685;
	wire [4-1:0] node4686;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4691;
	wire [4-1:0] node4692;
	wire [4-1:0] node4694;
	wire [4-1:0] node4698;
	wire [4-1:0] node4699;
	wire [4-1:0] node4701;
	wire [4-1:0] node4705;
	wire [4-1:0] node4706;
	wire [4-1:0] node4707;
	wire [4-1:0] node4709;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4716;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4723;
	wire [4-1:0] node4726;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4733;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4739;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4744;
	wire [4-1:0] node4748;
	wire [4-1:0] node4749;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4757;
	wire [4-1:0] node4758;
	wire [4-1:0] node4759;
	wire [4-1:0] node4763;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4772;
	wire [4-1:0] node4775;
	wire [4-1:0] node4776;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4782;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4791;
	wire [4-1:0] node4792;
	wire [4-1:0] node4793;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4798;
	wire [4-1:0] node4801;
	wire [4-1:0] node4803;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4811;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4814;
	wire [4-1:0] node4817;
	wire [4-1:0] node4820;
	wire [4-1:0] node4822;
	wire [4-1:0] node4825;
	wire [4-1:0] node4826;
	wire [4-1:0] node4830;
	wire [4-1:0] node4831;
	wire [4-1:0] node4832;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4838;
	wire [4-1:0] node4841;
	wire [4-1:0] node4842;
	wire [4-1:0] node4845;
	wire [4-1:0] node4848;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4855;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4861;
	wire [4-1:0] node4864;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4878;
	wire [4-1:0] node4879;
	wire [4-1:0] node4880;
	wire [4-1:0] node4881;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4892;
	wire [4-1:0] node4894;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4899;
	wire [4-1:0] node4900;
	wire [4-1:0] node4904;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4911;
	wire [4-1:0] node4915;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4922;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4926;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4938;
	wire [4-1:0] node4942;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4957;
	wire [4-1:0] node4959;
	wire [4-1:0] node4962;
	wire [4-1:0] node4963;
	wire [4-1:0] node4964;
	wire [4-1:0] node4968;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4990;
	wire [4-1:0] node4992;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node4997;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5004;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5015;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5024;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5035;
	wire [4-1:0] node5038;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5042;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5054;
	wire [4-1:0] node5055;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5063;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5066;
	wire [4-1:0] node5069;
	wire [4-1:0] node5073;
	wire [4-1:0] node5075;
	wire [4-1:0] node5076;
	wire [4-1:0] node5079;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5089;
	wire [4-1:0] node5092;
	wire [4-1:0] node5093;
	wire [4-1:0] node5097;
	wire [4-1:0] node5098;
	wire [4-1:0] node5103;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5110;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5117;
	wire [4-1:0] node5118;
	wire [4-1:0] node5119;
	wire [4-1:0] node5122;
	wire [4-1:0] node5123;
	wire [4-1:0] node5127;
	wire [4-1:0] node5129;
	wire [4-1:0] node5130;
	wire [4-1:0] node5133;
	wire [4-1:0] node5136;
	wire [4-1:0] node5137;
	wire [4-1:0] node5138;
	wire [4-1:0] node5139;
	wire [4-1:0] node5141;
	wire [4-1:0] node5144;
	wire [4-1:0] node5146;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5153;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5163;
	wire [4-1:0] node5164;
	wire [4-1:0] node5167;
	wire [4-1:0] node5170;
	wire [4-1:0] node5171;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5178;
	wire [4-1:0] node5179;
	wire [4-1:0] node5183;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5187;
	wire [4-1:0] node5188;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5198;
	wire [4-1:0] node5200;
	wire [4-1:0] node5203;
	wire [4-1:0] node5206;
	wire [4-1:0] node5207;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5213;
	wire [4-1:0] node5214;
	wire [4-1:0] node5215;
	wire [4-1:0] node5220;
	wire [4-1:0] node5221;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5233;
	wire [4-1:0] node5235;
	wire [4-1:0] node5236;
	wire [4-1:0] node5240;
	wire [4-1:0] node5241;
	wire [4-1:0] node5244;
	wire [4-1:0] node5247;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5251;
	wire [4-1:0] node5254;
	wire [4-1:0] node5256;
	wire [4-1:0] node5259;
	wire [4-1:0] node5260;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5271;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5278;
	wire [4-1:0] node5281;
	wire [4-1:0] node5284;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5290;
	wire [4-1:0] node5291;
	wire [4-1:0] node5293;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5300;
	wire [4-1:0] node5304;
	wire [4-1:0] node5305;
	wire [4-1:0] node5306;
	wire [4-1:0] node5307;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5316;
	wire [4-1:0] node5321;
	wire [4-1:0] node5322;
	wire [4-1:0] node5323;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5330;
	wire [4-1:0] node5333;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5339;
	wire [4-1:0] node5340;
	wire [4-1:0] node5343;
	wire [4-1:0] node5347;
	wire [4-1:0] node5348;
	wire [4-1:0] node5349;
	wire [4-1:0] node5351;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5360;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5364;
	wire [4-1:0] node5367;
	wire [4-1:0] node5368;
	wire [4-1:0] node5369;
	wire [4-1:0] node5373;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5379;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5384;
	wire [4-1:0] node5387;
	wire [4-1:0] node5389;
	wire [4-1:0] node5392;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5398;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5406;
	wire [4-1:0] node5407;
	wire [4-1:0] node5410;
	wire [4-1:0] node5413;
	wire [4-1:0] node5415;
	wire [4-1:0] node5418;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5425;
	wire [4-1:0] node5426;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5433;
	wire [4-1:0] node5434;
	wire [4-1:0] node5439;
	wire [4-1:0] node5440;
	wire [4-1:0] node5442;
	wire [4-1:0] node5446;
	wire [4-1:0] node5447;
	wire [4-1:0] node5449;
	wire [4-1:0] node5450;
	wire [4-1:0] node5454;
	wire [4-1:0] node5456;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5470;
	wire [4-1:0] node5473;
	wire [4-1:0] node5477;
	wire [4-1:0] node5478;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5485;
	wire [4-1:0] node5488;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5491;
	wire [4-1:0] node5493;
	wire [4-1:0] node5496;
	wire [4-1:0] node5498;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5508;
	wire [4-1:0] node5511;
	wire [4-1:0] node5514;
	wire [4-1:0] node5516;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5525;
	wire [4-1:0] node5527;
	wire [4-1:0] node5530;
	wire [4-1:0] node5531;
	wire [4-1:0] node5533;
	wire [4-1:0] node5536;
	wire [4-1:0] node5537;
	wire [4-1:0] node5538;
	wire [4-1:0] node5541;
	wire [4-1:0] node5545;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5553;
	wire [4-1:0] node5556;
	wire [4-1:0] node5559;
	wire [4-1:0] node5560;
	wire [4-1:0] node5561;
	wire [4-1:0] node5562;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5570;
	wire [4-1:0] node5572;
	wire [4-1:0] node5576;
	wire [4-1:0] node5577;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5581;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5588;
	wire [4-1:0] node5591;
	wire [4-1:0] node5593;
	wire [4-1:0] node5596;
	wire [4-1:0] node5599;
	wire [4-1:0] node5600;
	wire [4-1:0] node5601;
	wire [4-1:0] node5602;
	wire [4-1:0] node5604;
	wire [4-1:0] node5607;
	wire [4-1:0] node5610;
	wire [4-1:0] node5612;
	wire [4-1:0] node5613;
	wire [4-1:0] node5617;
	wire [4-1:0] node5618;
	wire [4-1:0] node5619;
	wire [4-1:0] node5622;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5629;
	wire [4-1:0] node5631;
	wire [4-1:0] node5634;
	wire [4-1:0] node5635;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5638;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5647;
	wire [4-1:0] node5648;
	wire [4-1:0] node5649;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5660;
	wire [4-1:0] node5663;
	wire [4-1:0] node5665;
	wire [4-1:0] node5668;
	wire [4-1:0] node5669;
	wire [4-1:0] node5673;
	wire [4-1:0] node5674;
	wire [4-1:0] node5675;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5680;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5689;
	wire [4-1:0] node5692;
	wire [4-1:0] node5693;
	wire [4-1:0] node5696;
	wire [4-1:0] node5698;
	wire [4-1:0] node5700;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5705;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5719;
	wire [4-1:0] node5720;
	wire [4-1:0] node5721;
	wire [4-1:0] node5724;
	wire [4-1:0] node5727;
	wire [4-1:0] node5728;
	wire [4-1:0] node5731;
	wire [4-1:0] node5734;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5737;
	wire [4-1:0] node5738;
	wire [4-1:0] node5739;
	wire [4-1:0] node5743;
	wire [4-1:0] node5744;
	wire [4-1:0] node5747;
	wire [4-1:0] node5750;
	wire [4-1:0] node5751;
	wire [4-1:0] node5754;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5759;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5768;
	wire [4-1:0] node5771;
	wire [4-1:0] node5772;
	wire [4-1:0] node5775;
	wire [4-1:0] node5778;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5786;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5795;
	wire [4-1:0] node5797;
	wire [4-1:0] node5800;
	wire [4-1:0] node5801;
	wire [4-1:0] node5802;
	wire [4-1:0] node5806;
	wire [4-1:0] node5807;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5817;
	wire [4-1:0] node5818;
	wire [4-1:0] node5821;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5830;
	wire [4-1:0] node5832;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5841;
	wire [4-1:0] node5846;
	wire [4-1:0] node5847;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5853;
	wire [4-1:0] node5854;
	wire [4-1:0] node5860;
	wire [4-1:0] node5861;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5868;
	wire [4-1:0] node5869;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5875;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5893;
	wire [4-1:0] node5894;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5904;
	wire [4-1:0] node5906;
	wire [4-1:0] node5909;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5913;
	wire [4-1:0] node5917;
	wire [4-1:0] node5920;
	wire [4-1:0] node5921;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5929;
	wire [4-1:0] node5931;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5938;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5945;
	wire [4-1:0] node5947;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5957;
	wire [4-1:0] node5959;
	wire [4-1:0] node5962;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5967;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5975;
	wire [4-1:0] node5976;
	wire [4-1:0] node5977;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5981;
	wire [4-1:0] node5984;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5992;
	wire [4-1:0] node5994;
	wire [4-1:0] node5998;
	wire [4-1:0] node5999;
	wire [4-1:0] node6000;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6007;
	wire [4-1:0] node6008;
	wire [4-1:0] node6011;
	wire [4-1:0] node6016;
	wire [4-1:0] node6017;
	wire [4-1:0] node6018;
	wire [4-1:0] node6019;
	wire [4-1:0] node6020;
	wire [4-1:0] node6021;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6031;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6046;
	wire [4-1:0] node6048;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6060;
	wire [4-1:0] node6061;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6067;
	wire [4-1:0] node6072;
	wire [4-1:0] node6073;
	wire [4-1:0] node6074;
	wire [4-1:0] node6075;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6083;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6092;
	wire [4-1:0] node6093;
	wire [4-1:0] node6094;
	wire [4-1:0] node6095;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6107;
	wire [4-1:0] node6111;
	wire [4-1:0] node6114;
	wire [4-1:0] node6116;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6121;
	wire [4-1:0] node6124;
	wire [4-1:0] node6126;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6132;
	wire [4-1:0] node6135;
	wire [4-1:0] node6138;
	wire [4-1:0] node6139;
	wire [4-1:0] node6141;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6155;
	wire [4-1:0] node6158;
	wire [4-1:0] node6159;
	wire [4-1:0] node6160;
	wire [4-1:0] node6164;
	wire [4-1:0] node6166;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6173;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6180;
	wire [4-1:0] node6184;
	wire [4-1:0] node6185;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6191;
	wire [4-1:0] node6193;
	wire [4-1:0] node6195;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6202;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6213;
	wire [4-1:0] node6215;
	wire [4-1:0] node6218;
	wire [4-1:0] node6219;
	wire [4-1:0] node6220;
	wire [4-1:0] node6224;
	wire [4-1:0] node6225;
	wire [4-1:0] node6229;
	wire [4-1:0] node6230;
	wire [4-1:0] node6232;
	wire [4-1:0] node6235;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6248;
	wire [4-1:0] node6250;
	wire [4-1:0] node6254;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6260;
	wire [4-1:0] node6261;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6272;
	wire [4-1:0] node6276;
	wire [4-1:0] node6278;
	wire [4-1:0] node6281;
	wire [4-1:0] node6282;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6292;
	wire [4-1:0] node6296;
	wire [4-1:0] node6297;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6308;
	wire [4-1:0] node6309;
	wire [4-1:0] node6313;
	wire [4-1:0] node6314;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6321;
	wire [4-1:0] node6322;
	wire [4-1:0] node6326;
	wire [4-1:0] node6327;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6334;
	wire [4-1:0] node6335;
	wire [4-1:0] node6336;
	wire [4-1:0] node6338;
	wire [4-1:0] node6340;
	wire [4-1:0] node6344;
	wire [4-1:0] node6345;
	wire [4-1:0] node6346;
	wire [4-1:0] node6347;
	wire [4-1:0] node6351;
	wire [4-1:0] node6353;
	wire [4-1:0] node6356;
	wire [4-1:0] node6358;
	wire [4-1:0] node6361;
	wire [4-1:0] node6362;
	wire [4-1:0] node6364;
	wire [4-1:0] node6365;
	wire [4-1:0] node6369;
	wire [4-1:0] node6370;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6380;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6389;
	wire [4-1:0] node6390;
	wire [4-1:0] node6391;
	wire [4-1:0] node6394;
	wire [4-1:0] node6396;
	wire [4-1:0] node6399;
	wire [4-1:0] node6401;
	wire [4-1:0] node6404;
	wire [4-1:0] node6405;
	wire [4-1:0] node6406;
	wire [4-1:0] node6408;
	wire [4-1:0] node6412;
	wire [4-1:0] node6414;
	wire [4-1:0] node6417;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6428;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6435;
	wire [4-1:0] node6438;
	wire [4-1:0] node6441;
	wire [4-1:0] node6442;
	wire [4-1:0] node6443;
	wire [4-1:0] node6445;
	wire [4-1:0] node6448;
	wire [4-1:0] node6449;
	wire [4-1:0] node6453;
	wire [4-1:0] node6455;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6463;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6480;
	wire [4-1:0] node6481;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6487;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6494;
	wire [4-1:0] node6495;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6503;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6510;
	wire [4-1:0] node6513;
	wire [4-1:0] node6515;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6527;
	wire [4-1:0] node6529;
	wire [4-1:0] node6533;
	wire [4-1:0] node6535;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6540;
	wire [4-1:0] node6543;
	wire [4-1:0] node6546;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6552;
	wire [4-1:0] node6555;
	wire [4-1:0] node6556;
	wire [4-1:0] node6560;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6564;
	wire [4-1:0] node6565;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6569;
	wire [4-1:0] node6571;
	wire [4-1:0] node6575;
	wire [4-1:0] node6577;
	wire [4-1:0] node6581;
	wire [4-1:0] node6582;
	wire [4-1:0] node6583;
	wire [4-1:0] node6584;
	wire [4-1:0] node6585;
	wire [4-1:0] node6586;
	wire [4-1:0] node6589;
	wire [4-1:0] node6592;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6598;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6604;
	wire [4-1:0] node6607;
	wire [4-1:0] node6609;
	wire [4-1:0] node6612;
	wire [4-1:0] node6613;
	wire [4-1:0] node6614;
	wire [4-1:0] node6617;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6622;
	wire [4-1:0] node6623;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6633;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6638;
	wire [4-1:0] node6640;
	wire [4-1:0] node6643;
	wire [4-1:0] node6647;
	wire [4-1:0] node6648;
	wire [4-1:0] node6649;
	wire [4-1:0] node6653;
	wire [4-1:0] node6654;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6662;
	wire [4-1:0] node6663;
	wire [4-1:0] node6666;
	wire [4-1:0] node6667;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6678;
	wire [4-1:0] node6680;
	wire [4-1:0] node6683;
	wire [4-1:0] node6685;
	wire [4-1:0] node6688;
	wire [4-1:0] node6689;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6701;
	wire [4-1:0] node6703;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6712;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6720;
	wire [4-1:0] node6723;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6727;
	wire [4-1:0] node6730;
	wire [4-1:0] node6733;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6739;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6746;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6752;
	wire [4-1:0] node6756;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6763;
	wire [4-1:0] node6765;
	wire [4-1:0] node6768;
	wire [4-1:0] node6769;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6775;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6784;
	wire [4-1:0] node6785;
	wire [4-1:0] node6786;
	wire [4-1:0] node6788;
	wire [4-1:0] node6791;
	wire [4-1:0] node6793;
	wire [4-1:0] node6794;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6800;
	wire [4-1:0] node6801;
	wire [4-1:0] node6804;
	wire [4-1:0] node6806;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6817;
	wire [4-1:0] node6819;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6835;
	wire [4-1:0] node6836;
	wire [4-1:0] node6837;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6853;
	wire [4-1:0] node6856;
	wire [4-1:0] node6859;
	wire [4-1:0] node6861;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6868;
	wire [4-1:0] node6873;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6878;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6887;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6894;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6901;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6907;
	wire [4-1:0] node6910;
	wire [4-1:0] node6911;
	wire [4-1:0] node6915;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6921;
	wire [4-1:0] node6922;
	wire [4-1:0] node6926;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6932;
	wire [4-1:0] node6935;
	wire [4-1:0] node6936;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6943;
	wire [4-1:0] node6944;
	wire [4-1:0] node6945;
	wire [4-1:0] node6949;
	wire [4-1:0] node6951;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6959;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6969;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6972;
	wire [4-1:0] node6974;
	wire [4-1:0] node6977;
	wire [4-1:0] node6980;
	wire [4-1:0] node6981;
	wire [4-1:0] node6984;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6993;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node6999;
	wire [4-1:0] node7003;
	wire [4-1:0] node7006;
	wire [4-1:0] node7007;
	wire [4-1:0] node7008;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7013;
	wire [4-1:0] node7016;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7024;
	wire [4-1:0] node7027;
	wire [4-1:0] node7028;
	wire [4-1:0] node7030;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7039;
	wire [4-1:0] node7042;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7049;
	wire [4-1:0] node7050;
	wire [4-1:0] node7051;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7054;
	wire [4-1:0] node7057;
	wire [4-1:0] node7058;
	wire [4-1:0] node7060;
	wire [4-1:0] node7064;
	wire [4-1:0] node7065;
	wire [4-1:0] node7068;
	wire [4-1:0] node7070;
	wire [4-1:0] node7072;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7086;
	wire [4-1:0] node7088;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7096;
	wire [4-1:0] node7100;
	wire [4-1:0] node7101;
	wire [4-1:0] node7102;
	wire [4-1:0] node7104;
	wire [4-1:0] node7105;
	wire [4-1:0] node7107;
	wire [4-1:0] node7110;
	wire [4-1:0] node7111;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7125;
	wire [4-1:0] node7126;
	wire [4-1:0] node7129;
	wire [4-1:0] node7132;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7136;
	wire [4-1:0] node7141;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7145;
	wire [4-1:0] node7147;
	wire [4-1:0] node7150;
	wire [4-1:0] node7153;
	wire [4-1:0] node7154;
	wire [4-1:0] node7157;
	wire [4-1:0] node7159;
	wire [4-1:0] node7161;
	wire [4-1:0] node7164;
	wire [4-1:0] node7165;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7171;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7176;
	wire [4-1:0] node7177;
	wire [4-1:0] node7181;
	wire [4-1:0] node7184;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7197;
	wire [4-1:0] node7198;
	wire [4-1:0] node7199;
	wire [4-1:0] node7200;
	wire [4-1:0] node7203;
	wire [4-1:0] node7205;
	wire [4-1:0] node7208;
	wire [4-1:0] node7209;
	wire [4-1:0] node7210;
	wire [4-1:0] node7214;
	wire [4-1:0] node7215;
	wire [4-1:0] node7217;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7228;
	wire [4-1:0] node7231;
	wire [4-1:0] node7235;
	wire [4-1:0] node7236;
	wire [4-1:0] node7238;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7246;
	wire [4-1:0] node7247;
	wire [4-1:0] node7248;
	wire [4-1:0] node7249;
	wire [4-1:0] node7250;
	wire [4-1:0] node7251;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7256;
	wire [4-1:0] node7259;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7270;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7276;
	wire [4-1:0] node7277;
	wire [4-1:0] node7281;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7286;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7297;
	wire [4-1:0] node7299;
	wire [4-1:0] node7302;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7305;
	wire [4-1:0] node7309;
	wire [4-1:0] node7310;
	wire [4-1:0] node7312;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7320;
	wire [4-1:0] node7321;
	wire [4-1:0] node7322;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7328;
	wire [4-1:0] node7331;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7337;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7350;
	wire [4-1:0] node7351;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7358;
	wire [4-1:0] node7361;
	wire [4-1:0] node7364;
	wire [4-1:0] node7365;
	wire [4-1:0] node7366;
	wire [4-1:0] node7369;
	wire [4-1:0] node7370;
	wire [4-1:0] node7374;
	wire [4-1:0] node7375;
	wire [4-1:0] node7376;
	wire [4-1:0] node7380;
	wire [4-1:0] node7382;
	wire [4-1:0] node7385;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7390;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7397;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7403;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7411;
	wire [4-1:0] node7412;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7417;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7425;
	wire [4-1:0] node7426;
	wire [4-1:0] node7427;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7435;
	wire [4-1:0] node7436;
	wire [4-1:0] node7440;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7444;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7453;
	wire [4-1:0] node7455;
	wire [4-1:0] node7458;
	wire [4-1:0] node7459;
	wire [4-1:0] node7460;
	wire [4-1:0] node7464;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7469;
	wire [4-1:0] node7472;
	wire [4-1:0] node7474;
	wire [4-1:0] node7477;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7481;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7489;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7496;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7501;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7508;
	wire [4-1:0] node7511;
	wire [4-1:0] node7513;
	wire [4-1:0] node7516;
	wire [4-1:0] node7517;
	wire [4-1:0] node7518;
	wire [4-1:0] node7519;
	wire [4-1:0] node7520;
	wire [4-1:0] node7523;
	wire [4-1:0] node7526;
	wire [4-1:0] node7527;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7534;
	wire [4-1:0] node7537;
	wire [4-1:0] node7539;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7550;
	wire [4-1:0] node7552;
	wire [4-1:0] node7555;
	wire [4-1:0] node7556;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7560;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7568;
	wire [4-1:0] node7570;
	wire [4-1:0] node7573;
	wire [4-1:0] node7575;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7581;
	wire [4-1:0] node7582;
	wire [4-1:0] node7583;
	wire [4-1:0] node7584;
	wire [4-1:0] node7588;
	wire [4-1:0] node7590;
	wire [4-1:0] node7593;
	wire [4-1:0] node7594;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7599;
	wire [4-1:0] node7603;
	wire [4-1:0] node7604;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7615;
	wire [4-1:0] node7617;
	wire [4-1:0] node7620;
	wire [4-1:0] node7621;
	wire [4-1:0] node7622;
	wire [4-1:0] node7624;
	wire [4-1:0] node7627;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7635;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7645;
	wire [4-1:0] node7646;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7654;
	wire [4-1:0] node7655;
	wire [4-1:0] node7656;
	wire [4-1:0] node7657;
	wire [4-1:0] node7658;
	wire [4-1:0] node7660;
	wire [4-1:0] node7662;
	wire [4-1:0] node7665;
	wire [4-1:0] node7666;
	wire [4-1:0] node7668;
	wire [4-1:0] node7672;
	wire [4-1:0] node7673;
	wire [4-1:0] node7675;
	wire [4-1:0] node7678;
	wire [4-1:0] node7679;
	wire [4-1:0] node7681;
	wire [4-1:0] node7684;
	wire [4-1:0] node7685;
	wire [4-1:0] node7689;
	wire [4-1:0] node7690;
	wire [4-1:0] node7691;
	wire [4-1:0] node7692;
	wire [4-1:0] node7695;
	wire [4-1:0] node7696;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7712;
	wire [4-1:0] node7715;
	wire [4-1:0] node7716;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7723;
	wire [4-1:0] node7725;
	wire [4-1:0] node7728;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7731;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7735;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7744;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7749;
	wire [4-1:0] node7752;
	wire [4-1:0] node7753;
	wire [4-1:0] node7757;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7760;
	wire [4-1:0] node7761;
	wire [4-1:0] node7764;
	wire [4-1:0] node7768;
	wire [4-1:0] node7770;
	wire [4-1:0] node7771;
	wire [4-1:0] node7774;
	wire [4-1:0] node7777;
	wire [4-1:0] node7778;
	wire [4-1:0] node7779;
	wire [4-1:0] node7783;
	wire [4-1:0] node7784;
	wire [4-1:0] node7785;
	wire [4-1:0] node7790;
	wire [4-1:0] node7791;
	wire [4-1:0] node7792;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7807;
	wire [4-1:0] node7811;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7818;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7824;
	wire [4-1:0] node7825;
	wire [4-1:0] node7829;
	wire [4-1:0] node7830;
	wire [4-1:0] node7832;
	wire [4-1:0] node7836;
	wire [4-1:0] node7837;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7844;
	wire [4-1:0] node7845;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7854;
	wire [4-1:0] node7855;
	wire [4-1:0] node7856;
	wire [4-1:0] node7857;
	wire [4-1:0] node7859;
	wire [4-1:0] node7860;
	wire [4-1:0] node7861;
	wire [4-1:0] node7866;
	wire [4-1:0] node7867;
	wire [4-1:0] node7869;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7877;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7881;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7887;
	wire [4-1:0] node7890;
	wire [4-1:0] node7893;
	wire [4-1:0] node7894;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7901;
	wire [4-1:0] node7902;
	wire [4-1:0] node7903;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7912;
	wire [4-1:0] node7915;
	wire [4-1:0] node7917;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7924;
	wire [4-1:0] node7927;
	wire [4-1:0] node7928;
	wire [4-1:0] node7931;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7937;
	wire [4-1:0] node7940;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7946;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7950;
	wire [4-1:0] node7953;
	wire [4-1:0] node7955;
	wire [4-1:0] node7958;
	wire [4-1:0] node7959;
	wire [4-1:0] node7960;
	wire [4-1:0] node7963;
	wire [4-1:0] node7967;
	wire [4-1:0] node7968;
	wire [4-1:0] node7970;
	wire [4-1:0] node7973;
	wire [4-1:0] node7975;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7980;
	wire [4-1:0] node7981;
	wire [4-1:0] node7983;
	wire [4-1:0] node7986;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7992;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8006;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8011;
	wire [4-1:0] node8014;
	wire [4-1:0] node8015;
	wire [4-1:0] node8019;
	wire [4-1:0] node8021;
	wire [4-1:0] node8024;
	wire [4-1:0] node8025;
	wire [4-1:0] node8026;
	wire [4-1:0] node8027;
	wire [4-1:0] node8028;
	wire [4-1:0] node8032;
	wire [4-1:0] node8033;
	wire [4-1:0] node8036;
	wire [4-1:0] node8040;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8058;
	wire [4-1:0] node8060;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8066;
	wire [4-1:0] node8069;
	wire [4-1:0] node8072;
	wire [4-1:0] node8074;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8092;
	wire [4-1:0] node8095;
	wire [4-1:0] node8096;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8103;
	wire [4-1:0] node8106;
	wire [4-1:0] node8109;
	wire [4-1:0] node8110;
	wire [4-1:0] node8111;
	wire [4-1:0] node8113;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8122;
	wire [4-1:0] node8123;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8127;
	wire [4-1:0] node8130;
	wire [4-1:0] node8133;
	wire [4-1:0] node8135;
	wire [4-1:0] node8136;
	wire [4-1:0] node8139;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8151;
	wire [4-1:0] node8154;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8160;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8170;
	wire [4-1:0] node8173;
	wire [4-1:0] node8174;
	wire [4-1:0] node8177;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8183;
	wire [4-1:0] node8187;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8190;
	wire [4-1:0] node8191;
	wire [4-1:0] node8194;
	wire [4-1:0] node8197;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8211;
	wire [4-1:0] node8213;
	wire [4-1:0] node8216;
	wire [4-1:0] node8217;
	wire [4-1:0] node8220;
	wire [4-1:0] node8223;
	wire [4-1:0] node8224;
	wire [4-1:0] node8225;
	wire [4-1:0] node8227;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8237;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8243;
	wire [4-1:0] node8246;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8266;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8276;
	wire [4-1:0] node8277;
	wire [4-1:0] node8280;
	wire [4-1:0] node8283;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8287;
	wire [4-1:0] node8290;
	wire [4-1:0] node8293;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8297;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8305;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8310;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8317;
	wire [4-1:0] node8318;
	wire [4-1:0] node8319;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8332;
	wire [4-1:0] node8335;
	wire [4-1:0] node8336;
	wire [4-1:0] node8340;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8346;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8353;
	wire [4-1:0] node8354;
	wire [4-1:0] node8355;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8361;
	wire [4-1:0] node8364;
	wire [4-1:0] node8365;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8372;
	wire [4-1:0] node8375;
	wire [4-1:0] node8378;
	wire [4-1:0] node8380;
	wire [4-1:0] node8381;
	wire [4-1:0] node8384;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8393;
	wire [4-1:0] node8394;
	wire [4-1:0] node8398;
	wire [4-1:0] node8399;
	wire [4-1:0] node8400;
	wire [4-1:0] node8401;
	wire [4-1:0] node8403;
	wire [4-1:0] node8404;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8413;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8418;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8423;
	wire [4-1:0] node8426;
	wire [4-1:0] node8429;
	wire [4-1:0] node8431;
	wire [4-1:0] node8432;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8438;
	wire [4-1:0] node8441;
	wire [4-1:0] node8444;
	wire [4-1:0] node8446;
	wire [4-1:0] node8448;
	wire [4-1:0] node8451;
	wire [4-1:0] node8452;
	wire [4-1:0] node8453;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8457;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8472;
	wire [4-1:0] node8475;
	wire [4-1:0] node8476;
	wire [4-1:0] node8479;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8485;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8493;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8500;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8513;
	wire [4-1:0] node8515;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8522;
	wire [4-1:0] node8524;
	wire [4-1:0] node8527;
	wire [4-1:0] node8528;
	wire [4-1:0] node8529;
	wire [4-1:0] node8532;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8540;
	wire [4-1:0] node8544;
	wire [4-1:0] node8545;
	wire [4-1:0] node8546;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8552;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8558;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8573;
	wire [4-1:0] node8574;
	wire [4-1:0] node8578;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8587;
	wire [4-1:0] node8590;
	wire [4-1:0] node8593;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8604;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8614;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8619;
	wire [4-1:0] node8623;
	wire [4-1:0] node8624;
	wire [4-1:0] node8628;
	wire [4-1:0] node8629;
	wire [4-1:0] node8630;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8637;
	wire [4-1:0] node8640;
	wire [4-1:0] node8643;
	wire [4-1:0] node8644;
	wire [4-1:0] node8646;
	wire [4-1:0] node8649;
	wire [4-1:0] node8651;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8658;
	wire [4-1:0] node8661;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8670;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8675;
	wire [4-1:0] node8676;
	wire [4-1:0] node8677;
	wire [4-1:0] node8681;
	wire [4-1:0] node8683;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8693;
	wire [4-1:0] node8694;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8700;
	wire [4-1:0] node8702;
	wire [4-1:0] node8705;
	wire [4-1:0] node8708;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8712;
	wire [4-1:0] node8715;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8723;
	wire [4-1:0] node8724;
	wire [4-1:0] node8725;
	wire [4-1:0] node8727;
	wire [4-1:0] node8730;
	wire [4-1:0] node8733;
	wire [4-1:0] node8734;
	wire [4-1:0] node8736;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8746;
	wire [4-1:0] node8747;
	wire [4-1:0] node8749;
	wire [4-1:0] node8752;
	wire [4-1:0] node8755;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8760;
	wire [4-1:0] node8763;
	wire [4-1:0] node8765;
	wire [4-1:0] node8768;
	wire [4-1:0] node8769;
	wire [4-1:0] node8772;
	wire [4-1:0] node8773;
	wire [4-1:0] node8777;
	wire [4-1:0] node8778;
	wire [4-1:0] node8779;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8783;
	wire [4-1:0] node8784;
	wire [4-1:0] node8787;
	wire [4-1:0] node8789;
	wire [4-1:0] node8792;
	wire [4-1:0] node8794;
	wire [4-1:0] node8797;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8804;
	wire [4-1:0] node8806;
	wire [4-1:0] node8809;
	wire [4-1:0] node8810;
	wire [4-1:0] node8812;
	wire [4-1:0] node8814;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8821;
	wire [4-1:0] node8822;
	wire [4-1:0] node8825;
	wire [4-1:0] node8828;
	wire [4-1:0] node8829;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8836;
	wire [4-1:0] node8838;
	wire [4-1:0] node8841;
	wire [4-1:0] node8842;
	wire [4-1:0] node8844;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8851;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8856;
	wire [4-1:0] node8858;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8866;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8872;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8880;
	wire [4-1:0] node8882;
	wire [4-1:0] node8886;
	wire [4-1:0] node8887;
	wire [4-1:0] node8888;
	wire [4-1:0] node8891;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8899;
	wire [4-1:0] node8900;
	wire [4-1:0] node8903;
	wire [4-1:0] node8906;
	wire [4-1:0] node8908;
	wire [4-1:0] node8909;
	wire [4-1:0] node8913;
	wire [4-1:0] node8915;
	wire [4-1:0] node8916;
	wire [4-1:0] node8918;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8930;
	wire [4-1:0] node8932;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8938;
	wire [4-1:0] node8940;
	wire [4-1:0] node8943;
	wire [4-1:0] node8945;
	wire [4-1:0] node8949;
	wire [4-1:0] node8950;
	wire [4-1:0] node8951;
	wire [4-1:0] node8952;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8965;
	wire [4-1:0] node8968;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8973;
	wire [4-1:0] node8975;
	wire [4-1:0] node8978;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8984;
	wire [4-1:0] node8987;
	wire [4-1:0] node8990;
	wire [4-1:0] node8992;
	wire [4-1:0] node8995;
	wire [4-1:0] node8998;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9001;
	wire [4-1:0] node9005;
	wire [4-1:0] node9006;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9015;
	wire [4-1:0] node9018;
	wire [4-1:0] node9020;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9026;
	wire [4-1:0] node9027;
	wire [4-1:0] node9030;
	wire [4-1:0] node9031;
	wire [4-1:0] node9035;
	wire [4-1:0] node9036;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9042;
	wire [4-1:0] node9045;
	wire [4-1:0] node9046;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9061;
	wire [4-1:0] node9063;
	wire [4-1:0] node9064;
	wire [4-1:0] node9068;
	wire [4-1:0] node9069;
	wire [4-1:0] node9070;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9077;
	wire [4-1:0] node9081;
	wire [4-1:0] node9082;
	wire [4-1:0] node9083;
	wire [4-1:0] node9084;
	wire [4-1:0] node9086;
	wire [4-1:0] node9089;
	wire [4-1:0] node9091;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9104;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9108;
	wire [4-1:0] node9109;
	wire [4-1:0] node9111;
	wire [4-1:0] node9114;
	wire [4-1:0] node9116;
	wire [4-1:0] node9119;
	wire [4-1:0] node9120;
	wire [4-1:0] node9121;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9133;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9139;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9146;
	wire [4-1:0] node9149;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9152;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9160;
	wire [4-1:0] node9162;
	wire [4-1:0] node9164;
	wire [4-1:0] node9168;
	wire [4-1:0] node9169;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9177;
	wire [4-1:0] node9179;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9191;
	wire [4-1:0] node9192;
	wire [4-1:0] node9193;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9197;
	wire [4-1:0] node9199;
	wire [4-1:0] node9200;
	wire [4-1:0] node9201;
	wire [4-1:0] node9203;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9211;
	wire [4-1:0] node9213;
	wire [4-1:0] node9214;
	wire [4-1:0] node9217;
	wire [4-1:0] node9219;
	wire [4-1:0] node9222;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9226;
	wire [4-1:0] node9227;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9234;
	wire [4-1:0] node9237;
	wire [4-1:0] node9239;
	wire [4-1:0] node9242;
	wire [4-1:0] node9243;
	wire [4-1:0] node9244;
	wire [4-1:0] node9245;
	wire [4-1:0] node9249;
	wire [4-1:0] node9250;
	wire [4-1:0] node9254;
	wire [4-1:0] node9257;
	wire [4-1:0] node9259;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9263;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9270;
	wire [4-1:0] node9272;
	wire [4-1:0] node9275;
	wire [4-1:0] node9277;
	wire [4-1:0] node9278;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9287;
	wire [4-1:0] node9288;
	wire [4-1:0] node9289;
	wire [4-1:0] node9293;
	wire [4-1:0] node9295;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9300;
	wire [4-1:0] node9304;
	wire [4-1:0] node9306;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9312;
	wire [4-1:0] node9315;
	wire [4-1:0] node9316;
	wire [4-1:0] node9320;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9332;
	wire [4-1:0] node9333;
	wire [4-1:0] node9334;
	wire [4-1:0] node9335;
	wire [4-1:0] node9339;
	wire [4-1:0] node9342;
	wire [4-1:0] node9343;
	wire [4-1:0] node9345;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9358;
	wire [4-1:0] node9359;
	wire [4-1:0] node9363;
	wire [4-1:0] node9364;
	wire [4-1:0] node9365;
	wire [4-1:0] node9367;
	wire [4-1:0] node9371;
	wire [4-1:0] node9372;
	wire [4-1:0] node9374;
	wire [4-1:0] node9378;
	wire [4-1:0] node9379;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9384;
	wire [4-1:0] node9387;
	wire [4-1:0] node9389;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9397;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9404;
	wire [4-1:0] node9405;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9414;
	wire [4-1:0] node9415;
	wire [4-1:0] node9417;
	wire [4-1:0] node9420;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9425;
	wire [4-1:0] node9427;
	wire [4-1:0] node9428;
	wire [4-1:0] node9432;
	wire [4-1:0] node9435;
	wire [4-1:0] node9436;
	wire [4-1:0] node9437;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9446;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9449;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9456;
	wire [4-1:0] node9460;
	wire [4-1:0] node9461;
	wire [4-1:0] node9462;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9470;
	wire [4-1:0] node9473;
	wire [4-1:0] node9474;
	wire [4-1:0] node9475;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9485;
	wire [4-1:0] node9488;
	wire [4-1:0] node9490;
	wire [4-1:0] node9493;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9504;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9518;
	wire [4-1:0] node9519;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9527;
	wire [4-1:0] node9528;
	wire [4-1:0] node9530;
	wire [4-1:0] node9532;
	wire [4-1:0] node9535;
	wire [4-1:0] node9536;
	wire [4-1:0] node9537;
	wire [4-1:0] node9540;
	wire [4-1:0] node9542;
	wire [4-1:0] node9545;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9552;
	wire [4-1:0] node9553;
	wire [4-1:0] node9554;
	wire [4-1:0] node9555;
	wire [4-1:0] node9558;
	wire [4-1:0] node9560;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9567;
	wire [4-1:0] node9568;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9574;
	wire [4-1:0] node9575;
	wire [4-1:0] node9579;
	wire [4-1:0] node9581;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9588;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9595;
	wire [4-1:0] node9597;
	wire [4-1:0] node9599;
	wire [4-1:0] node9600;
	wire [4-1:0] node9601;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9605;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9612;
	wire [4-1:0] node9613;
	wire [4-1:0] node9617;
	wire [4-1:0] node9621;
	wire [4-1:0] node9622;
	wire [4-1:0] node9623;
	wire [4-1:0] node9624;
	wire [4-1:0] node9625;
	wire [4-1:0] node9626;
	wire [4-1:0] node9628;
	wire [4-1:0] node9631;
	wire [4-1:0] node9635;
	wire [4-1:0] node9636;
	wire [4-1:0] node9637;
	wire [4-1:0] node9638;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9648;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9661;
	wire [4-1:0] node9664;
	wire [4-1:0] node9665;
	wire [4-1:0] node9666;
	wire [4-1:0] node9671;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9676;
	wire [4-1:0] node9680;
	wire [4-1:0] node9683;
	wire [4-1:0] node9685;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9696;
	wire [4-1:0] node9697;
	wire [4-1:0] node9698;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9704;
	wire [4-1:0] node9706;
	wire [4-1:0] node9709;
	wire [4-1:0] node9710;
	wire [4-1:0] node9712;
	wire [4-1:0] node9713;
	wire [4-1:0] node9718;
	wire [4-1:0] node9719;
	wire [4-1:0] node9720;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9724;
	wire [4-1:0] node9729;
	wire [4-1:0] node9730;
	wire [4-1:0] node9731;
	wire [4-1:0] node9732;
	wire [4-1:0] node9735;
	wire [4-1:0] node9739;
	wire [4-1:0] node9741;
	wire [4-1:0] node9742;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9752;
	wire [4-1:0] node9755;
	wire [4-1:0] node9757;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9768;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9774;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9777;
	wire [4-1:0] node9779;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9785;
	wire [4-1:0] node9789;
	wire [4-1:0] node9790;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9811;
	wire [4-1:0] node9812;
	wire [4-1:0] node9815;
	wire [4-1:0] node9818;
	wire [4-1:0] node9821;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9824;
	wire [4-1:0] node9825;
	wire [4-1:0] node9827;
	wire [4-1:0] node9831;
	wire [4-1:0] node9833;
	wire [4-1:0] node9834;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9841;
	wire [4-1:0] node9845;
	wire [4-1:0] node9846;
	wire [4-1:0] node9847;
	wire [4-1:0] node9848;
	wire [4-1:0] node9850;
	wire [4-1:0] node9853;
	wire [4-1:0] node9856;
	wire [4-1:0] node9857;
	wire [4-1:0] node9860;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9866;
	wire [4-1:0] node9869;
	wire [4-1:0] node9870;
	wire [4-1:0] node9873;
	wire [4-1:0] node9874;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9881;
	wire [4-1:0] node9882;
	wire [4-1:0] node9883;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9894;
	wire [4-1:0] node9899;
	wire [4-1:0] node9901;
	wire [4-1:0] node9903;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9909;
	wire [4-1:0] node9912;
	wire [4-1:0] node9913;
	wire [4-1:0] node9915;
	wire [4-1:0] node9917;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9923;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9929;
	wire [4-1:0] node9930;
	wire [4-1:0] node9931;
	wire [4-1:0] node9934;
	wire [4-1:0] node9937;
	wire [4-1:0] node9938;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9949;
	wire [4-1:0] node9952;
	wire [4-1:0] node9953;
	wire [4-1:0] node9955;
	wire [4-1:0] node9958;
	wire [4-1:0] node9961;
	wire [4-1:0] node9962;
	wire [4-1:0] node9964;
	wire [4-1:0] node9966;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9972;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9979;
	wire [4-1:0] node9982;
	wire [4-1:0] node9983;
	wire [4-1:0] node9984;
	wire [4-1:0] node9985;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9991;
	wire [4-1:0] node9992;
	wire [4-1:0] node9993;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node10002;
	wire [4-1:0] node10003;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10011;
	wire [4-1:0] node10014;
	wire [4-1:0] node10016;
	wire [4-1:0] node10019;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10028;
	wire [4-1:0] node10029;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10034;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10044;
	wire [4-1:0] node10045;
	wire [4-1:0] node10047;
	wire [4-1:0] node10050;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10055;
	wire [4-1:0] node10059;
	wire [4-1:0] node10061;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10067;
	wire [4-1:0] node10069;
	wire [4-1:0] node10070;
	wire [4-1:0] node10073;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10080;
	wire [4-1:0] node10084;
	wire [4-1:0] node10085;
	wire [4-1:0] node10087;
	wire [4-1:0] node10090;
	wire [4-1:0] node10091;
	wire [4-1:0] node10094;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10100;
	wire [4-1:0] node10101;
	wire [4-1:0] node10102;
	wire [4-1:0] node10103;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10108;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10115;
	wire [4-1:0] node10118;
	wire [4-1:0] node10120;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10125;
	wire [4-1:0] node10129;
	wire [4-1:0] node10132;
	wire [4-1:0] node10133;
	wire [4-1:0] node10134;
	wire [4-1:0] node10135;
	wire [4-1:0] node10137;
	wire [4-1:0] node10141;
	wire [4-1:0] node10142;
	wire [4-1:0] node10145;
	wire [4-1:0] node10148;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10153;
	wire [4-1:0] node10156;
	wire [4-1:0] node10158;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10169;
	wire [4-1:0] node10172;
	wire [4-1:0] node10175;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10184;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10192;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10197;
	wire [4-1:0] node10200;
	wire [4-1:0] node10202;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10208;
	wire [4-1:0] node10211;
	wire [4-1:0] node10213;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10224;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10227;
	wire [4-1:0] node10233;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10236;
	wire [4-1:0] node10237;
	wire [4-1:0] node10241;
	wire [4-1:0] node10244;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10250;
	wire [4-1:0] node10254;
	wire [4-1:0] node10255;
	wire [4-1:0] node10256;
	wire [4-1:0] node10257;
	wire [4-1:0] node10258;
	wire [4-1:0] node10261;
	wire [4-1:0] node10262;
	wire [4-1:0] node10265;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10272;
	wire [4-1:0] node10275;
	wire [4-1:0] node10276;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10284;
	wire [4-1:0] node10285;
	wire [4-1:0] node10286;
	wire [4-1:0] node10288;
	wire [4-1:0] node10291;
	wire [4-1:0] node10293;
	wire [4-1:0] node10296;
	wire [4-1:0] node10297;
	wire [4-1:0] node10298;
	wire [4-1:0] node10299;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10308;
	wire [4-1:0] node10310;
	wire [4-1:0] node10313;
	wire [4-1:0] node10314;
	wire [4-1:0] node10315;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10321;
	wire [4-1:0] node10324;
	wire [4-1:0] node10325;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10336;
	wire [4-1:0] node10339;
	wire [4-1:0] node10340;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10347;
	wire [4-1:0] node10350;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10354;
	wire [4-1:0] node10355;
	wire [4-1:0] node10360;
	wire [4-1:0] node10361;
	wire [4-1:0] node10362;
	wire [4-1:0] node10365;
	wire [4-1:0] node10369;
	wire [4-1:0] node10370;
	wire [4-1:0] node10373;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10378;
	wire [4-1:0] node10381;
	wire [4-1:0] node10383;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10391;
	wire [4-1:0] node10395;
	wire [4-1:0] node10396;
	wire [4-1:0] node10397;
	wire [4-1:0] node10398;
	wire [4-1:0] node10400;
	wire [4-1:0] node10401;
	wire [4-1:0] node10405;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10409;
	wire [4-1:0] node10413;
	wire [4-1:0] node10415;
	wire [4-1:0] node10417;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10426;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10431;
	wire [4-1:0] node10435;
	wire [4-1:0] node10438;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10442;
	wire [4-1:0] node10445;
	wire [4-1:0] node10447;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10459;
	wire [4-1:0] node10462;
	wire [4-1:0] node10463;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10472;
	wire [4-1:0] node10473;
	wire [4-1:0] node10478;
	wire [4-1:0] node10480;
	wire [4-1:0] node10481;
	wire [4-1:0] node10484;
	wire [4-1:0] node10488;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10496;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10505;
	wire [4-1:0] node10507;
	wire [4-1:0] node10510;
	wire [4-1:0] node10511;
	wire [4-1:0] node10512;
	wire [4-1:0] node10515;
	wire [4-1:0] node10516;
	wire [4-1:0] node10520;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10534;
	wire [4-1:0] node10538;
	wire [4-1:0] node10539;
	wire [4-1:0] node10541;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10548;
	wire [4-1:0] node10549;
	wire [4-1:0] node10552;
	wire [4-1:0] node10555;
	wire [4-1:0] node10556;
	wire [4-1:0] node10557;
	wire [4-1:0] node10559;
	wire [4-1:0] node10562;
	wire [4-1:0] node10564;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10570;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10576;
	wire [4-1:0] node10577;
	wire [4-1:0] node10578;
	wire [4-1:0] node10582;
	wire [4-1:0] node10583;
	wire [4-1:0] node10585;
	wire [4-1:0] node10586;
	wire [4-1:0] node10589;
	wire [4-1:0] node10592;
	wire [4-1:0] node10594;
	wire [4-1:0] node10597;
	wire [4-1:0] node10598;
	wire [4-1:0] node10599;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10606;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10612;
	wire [4-1:0] node10614;
	wire [4-1:0] node10617;
	wire [4-1:0] node10619;
	wire [4-1:0] node10622;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10626;
	wire [4-1:0] node10627;
	wire [4-1:0] node10628;
	wire [4-1:0] node10632;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10638;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10651;
	wire [4-1:0] node10653;
	wire [4-1:0] node10655;
	wire [4-1:0] node10658;
	wire [4-1:0] node10659;
	wire [4-1:0] node10661;
	wire [4-1:0] node10664;
	wire [4-1:0] node10665;
	wire [4-1:0] node10667;
	wire [4-1:0] node10670;
	wire [4-1:0] node10671;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10679;
	wire [4-1:0] node10680;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10685;
	wire [4-1:0] node10688;
	wire [4-1:0] node10691;
	wire [4-1:0] node10692;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10703;
	wire [4-1:0] node10704;
	wire [4-1:0] node10708;
	wire [4-1:0] node10709;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10717;
	wire [4-1:0] node10718;
	wire [4-1:0] node10722;
	wire [4-1:0] node10724;
	wire [4-1:0] node10725;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10734;
	wire [4-1:0] node10737;
	wire [4-1:0] node10738;
	wire [4-1:0] node10739;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10746;
	wire [4-1:0] node10747;
	wire [4-1:0] node10751;
	wire [4-1:0] node10752;
	wire [4-1:0] node10753;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10768;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10774;
	wire [4-1:0] node10778;
	wire [4-1:0] node10779;
	wire [4-1:0] node10780;
	wire [4-1:0] node10783;
	wire [4-1:0] node10786;
	wire [4-1:0] node10787;
	wire [4-1:0] node10791;
	wire [4-1:0] node10792;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10797;
	wire [4-1:0] node10801;
	wire [4-1:0] node10804;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10811;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10816;
	wire [4-1:0] node10819;
	wire [4-1:0] node10822;
	wire [4-1:0] node10823;
	wire [4-1:0] node10824;
	wire [4-1:0] node10826;
	wire [4-1:0] node10827;
	wire [4-1:0] node10831;
	wire [4-1:0] node10832;
	wire [4-1:0] node10833;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10840;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10848;
	wire [4-1:0] node10850;
	wire [4-1:0] node10851;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10857;
	wire [4-1:0] node10858;
	wire [4-1:0] node10860;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10869;
	wire [4-1:0] node10870;
	wire [4-1:0] node10871;
	wire [4-1:0] node10872;
	wire [4-1:0] node10874;
	wire [4-1:0] node10877;
	wire [4-1:0] node10879;
	wire [4-1:0] node10882;
	wire [4-1:0] node10884;
	wire [4-1:0] node10886;
	wire [4-1:0] node10890;
	wire [4-1:0] node10891;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10896;
	wire [4-1:0] node10897;
	wire [4-1:0] node10901;
	wire [4-1:0] node10903;
	wire [4-1:0] node10906;
	wire [4-1:0] node10907;
	wire [4-1:0] node10908;
	wire [4-1:0] node10911;
	wire [4-1:0] node10914;
	wire [4-1:0] node10915;
	wire [4-1:0] node10918;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10923;
	wire [4-1:0] node10925;
	wire [4-1:0] node10928;
	wire [4-1:0] node10931;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10936;
	wire [4-1:0] node10939;
	wire [4-1:0] node10941;
	wire [4-1:0] node10944;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10949;
	wire [4-1:0] node10951;
	wire [4-1:0] node10952;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10962;
	wire [4-1:0] node10965;
	wire [4-1:0] node10967;
	wire [4-1:0] node10970;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10976;
	wire [4-1:0] node10980;
	wire [4-1:0] node10981;
	wire [4-1:0] node10984;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10989;
	wire [4-1:0] node10990;
	wire [4-1:0] node10991;
	wire [4-1:0] node10994;
	wire [4-1:0] node10998;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11002;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11009;
	wire [4-1:0] node11012;
	wire [4-1:0] node11014;
	wire [4-1:0] node11017;
	wire [4-1:0] node11018;
	wire [4-1:0] node11019;
	wire [4-1:0] node11020;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11029;
	wire [4-1:0] node11032;
	wire [4-1:0] node11033;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11044;
	wire [4-1:0] node11045;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11050;
	wire [4-1:0] node11053;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11058;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11066;
	wire [4-1:0] node11067;
	wire [4-1:0] node11069;
	wire [4-1:0] node11072;
	wire [4-1:0] node11073;
	wire [4-1:0] node11074;
	wire [4-1:0] node11076;
	wire [4-1:0] node11080;
	wire [4-1:0] node11082;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11087;
	wire [4-1:0] node11088;
	wire [4-1:0] node11090;
	wire [4-1:0] node11093;
	wire [4-1:0] node11096;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11102;
	wire [4-1:0] node11104;
	wire [4-1:0] node11107;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11114;
	wire [4-1:0] node11115;
	wire [4-1:0] node11116;
	wire [4-1:0] node11117;
	wire [4-1:0] node11118;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11124;
	wire [4-1:0] node11125;
	wire [4-1:0] node11129;
	wire [4-1:0] node11130;
	wire [4-1:0] node11134;
	wire [4-1:0] node11135;
	wire [4-1:0] node11138;
	wire [4-1:0] node11139;
	wire [4-1:0] node11143;
	wire [4-1:0] node11144;
	wire [4-1:0] node11146;
	wire [4-1:0] node11150;
	wire [4-1:0] node11151;
	wire [4-1:0] node11152;
	wire [4-1:0] node11154;
	wire [4-1:0] node11156;
	wire [4-1:0] node11160;
	wire [4-1:0] node11163;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11169;
	wire [4-1:0] node11170;
	wire [4-1:0] node11171;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11175;
	wire [4-1:0] node11179;
	wire [4-1:0] node11180;
	wire [4-1:0] node11181;
	wire [4-1:0] node11185;
	wire [4-1:0] node11186;
	wire [4-1:0] node11189;
	wire [4-1:0] node11193;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11203;
	wire [4-1:0] node11206;
	wire [4-1:0] node11209;
	wire [4-1:0] node11211;
	wire [4-1:0] node11213;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11223;
	wire [4-1:0] node11226;
	wire [4-1:0] node11227;
	wire [4-1:0] node11229;
	wire [4-1:0] node11233;
	wire [4-1:0] node11235;
	wire [4-1:0] node11236;
	wire [4-1:0] node11237;
	wire [4-1:0] node11239;
	wire [4-1:0] node11242;
	wire [4-1:0] node11244;
	wire [4-1:0] node11246;
	wire [4-1:0] node11249;
	wire [4-1:0] node11251;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11262;
	wire [4-1:0] node11266;
	wire [4-1:0] node11267;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11274;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11279;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11285;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11293;
	wire [4-1:0] node11295;
	wire [4-1:0] node11297;
	wire [4-1:0] node11300;
	wire [4-1:0] node11301;
	wire [4-1:0] node11302;
	wire [4-1:0] node11303;
	wire [4-1:0] node11304;
	wire [4-1:0] node11308;
	wire [4-1:0] node11310;
	wire [4-1:0] node11313;
	wire [4-1:0] node11314;
	wire [4-1:0] node11315;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11324;
	wire [4-1:0] node11327;
	wire [4-1:0] node11329;
	wire [4-1:0] node11332;
	wire [4-1:0] node11333;
	wire [4-1:0] node11334;
	wire [4-1:0] node11335;
	wire [4-1:0] node11338;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11344;
	wire [4-1:0] node11348;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11354;
	wire [4-1:0] node11355;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11362;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11369;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11375;
	wire [4-1:0] node11376;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11383;
	wire [4-1:0] node11384;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11392;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11398;
	wire [4-1:0] node11402;
	wire [4-1:0] node11403;
	wire [4-1:0] node11404;
	wire [4-1:0] node11408;
	wire [4-1:0] node11410;
	wire [4-1:0] node11413;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11419;
	wire [4-1:0] node11423;
	wire [4-1:0] node11424;
	wire [4-1:0] node11428;
	wire [4-1:0] node11429;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11435;
	wire [4-1:0] node11438;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11447;
	wire [4-1:0] node11449;
	wire [4-1:0] node11452;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11455;
	wire [4-1:0] node11457;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11465;
	wire [4-1:0] node11468;
	wire [4-1:0] node11469;
	wire [4-1:0] node11472;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11477;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11483;
	wire [4-1:0] node11484;
	wire [4-1:0] node11488;
	wire [4-1:0] node11489;
	wire [4-1:0] node11490;
	wire [4-1:0] node11494;
	wire [4-1:0] node11495;
	wire [4-1:0] node11499;
	wire [4-1:0] node11500;
	wire [4-1:0] node11502;
	wire [4-1:0] node11506;
	wire [4-1:0] node11507;
	wire [4-1:0] node11508;
	wire [4-1:0] node11509;
	wire [4-1:0] node11510;
	wire [4-1:0] node11513;
	wire [4-1:0] node11514;
	wire [4-1:0] node11517;
	wire [4-1:0] node11519;
	wire [4-1:0] node11522;
	wire [4-1:0] node11523;
	wire [4-1:0] node11524;
	wire [4-1:0] node11525;
	wire [4-1:0] node11529;
	wire [4-1:0] node11530;
	wire [4-1:0] node11534;
	wire [4-1:0] node11537;
	wire [4-1:0] node11538;
	wire [4-1:0] node11539;
	wire [4-1:0] node11541;
	wire [4-1:0] node11544;
	wire [4-1:0] node11545;
	wire [4-1:0] node11547;
	wire [4-1:0] node11550;
	wire [4-1:0] node11553;
	wire [4-1:0] node11554;
	wire [4-1:0] node11556;
	wire [4-1:0] node11560;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11566;
	wire [4-1:0] node11568;
	wire [4-1:0] node11570;
	wire [4-1:0] node11573;
	wire [4-1:0] node11574;
	wire [4-1:0] node11575;
	wire [4-1:0] node11576;
	wire [4-1:0] node11580;
	wire [4-1:0] node11582;
	wire [4-1:0] node11586;
	wire [4-1:0] node11587;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11601;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11607;
	wire [4-1:0] node11608;
	wire [4-1:0] node11609;
	wire [4-1:0] node11611;
	wire [4-1:0] node11612;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11619;
	wire [4-1:0] node11623;
	wire [4-1:0] node11625;
	wire [4-1:0] node11629;
	wire [4-1:0] node11630;
	wire [4-1:0] node11631;
	wire [4-1:0] node11632;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11638;
	wire [4-1:0] node11639;
	wire [4-1:0] node11643;
	wire [4-1:0] node11644;
	wire [4-1:0] node11645;
	wire [4-1:0] node11647;
	wire [4-1:0] node11651;
	wire [4-1:0] node11655;
	wire [4-1:0] node11656;
	wire [4-1:0] node11657;
	wire [4-1:0] node11658;
	wire [4-1:0] node11661;
	wire [4-1:0] node11664;
	wire [4-1:0] node11665;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11681;
	wire [4-1:0] node11686;
	wire [4-1:0] node11687;
	wire [4-1:0] node11688;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11692;
	wire [4-1:0] node11693;
	wire [4-1:0] node11694;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11697;
	wire [4-1:0] node11699;
	wire [4-1:0] node11700;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11713;
	wire [4-1:0] node11715;
	wire [4-1:0] node11718;
	wire [4-1:0] node11719;
	wire [4-1:0] node11720;
	wire [4-1:0] node11721;
	wire [4-1:0] node11725;
	wire [4-1:0] node11727;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11740;
	wire [4-1:0] node11742;
	wire [4-1:0] node11743;
	wire [4-1:0] node11747;
	wire [4-1:0] node11749;
	wire [4-1:0] node11752;
	wire [4-1:0] node11753;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11760;
	wire [4-1:0] node11761;
	wire [4-1:0] node11765;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11768;
	wire [4-1:0] node11772;
	wire [4-1:0] node11773;
	wire [4-1:0] node11775;
	wire [4-1:0] node11776;
	wire [4-1:0] node11780;
	wire [4-1:0] node11783;
	wire [4-1:0] node11784;
	wire [4-1:0] node11786;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11791;
	wire [4-1:0] node11795;
	wire [4-1:0] node11798;
	wire [4-1:0] node11799;
	wire [4-1:0] node11800;
	wire [4-1:0] node11801;
	wire [4-1:0] node11803;
	wire [4-1:0] node11805;
	wire [4-1:0] node11808;
	wire [4-1:0] node11810;
	wire [4-1:0] node11813;
	wire [4-1:0] node11814;
	wire [4-1:0] node11816;
	wire [4-1:0] node11817;
	wire [4-1:0] node11819;
	wire [4-1:0] node11822;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11827;
	wire [4-1:0] node11831;
	wire [4-1:0] node11832;
	wire [4-1:0] node11834;
	wire [4-1:0] node11837;
	wire [4-1:0] node11840;
	wire [4-1:0] node11841;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11846;
	wire [4-1:0] node11848;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11866;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11872;
	wire [4-1:0] node11876;
	wire [4-1:0] node11877;
	wire [4-1:0] node11881;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11884;
	wire [4-1:0] node11885;
	wire [4-1:0] node11886;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11893;
	wire [4-1:0] node11895;
	wire [4-1:0] node11898;
	wire [4-1:0] node11899;
	wire [4-1:0] node11900;
	wire [4-1:0] node11902;
	wire [4-1:0] node11905;
	wire [4-1:0] node11906;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11912;
	wire [4-1:0] node11914;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11925;
	wire [4-1:0] node11926;
	wire [4-1:0] node11929;
	wire [4-1:0] node11930;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11937;
	wire [4-1:0] node11940;
	wire [4-1:0] node11943;
	wire [4-1:0] node11944;
	wire [4-1:0] node11946;
	wire [4-1:0] node11948;
	wire [4-1:0] node11951;
	wire [4-1:0] node11953;
	wire [4-1:0] node11956;
	wire [4-1:0] node11957;
	wire [4-1:0] node11958;
	wire [4-1:0] node11959;
	wire [4-1:0] node11961;
	wire [4-1:0] node11962;
	wire [4-1:0] node11964;
	wire [4-1:0] node11967;
	wire [4-1:0] node11969;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11974;
	wire [4-1:0] node11978;
	wire [4-1:0] node11979;
	wire [4-1:0] node11982;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11987;
	wire [4-1:0] node11990;
	wire [4-1:0] node11992;
	wire [4-1:0] node11995;
	wire [4-1:0] node11997;
	wire [4-1:0] node12000;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12003;
	wire [4-1:0] node12006;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12013;
	wire [4-1:0] node12014;
	wire [4-1:0] node12016;
	wire [4-1:0] node12020;
	wire [4-1:0] node12021;
	wire [4-1:0] node12023;
	wire [4-1:0] node12026;
	wire [4-1:0] node12027;
	wire [4-1:0] node12029;
	wire [4-1:0] node12032;
	wire [4-1:0] node12034;
	wire [4-1:0] node12037;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12043;
	wire [4-1:0] node12047;
	wire [4-1:0] node12048;
	wire [4-1:0] node12052;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12058;
	wire [4-1:0] node12061;
	wire [4-1:0] node12062;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12069;
	wire [4-1:0] node12074;
	wire [4-1:0] node12076;
	wire [4-1:0] node12079;
	wire [4-1:0] node12080;
	wire [4-1:0] node12081;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12091;
	wire [4-1:0] node12092;
	wire [4-1:0] node12096;
	wire [4-1:0] node12097;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12103;
	wire [4-1:0] node12105;
	wire [4-1:0] node12108;
	wire [4-1:0] node12109;
	wire [4-1:0] node12113;
	wire [4-1:0] node12114;
	wire [4-1:0] node12118;
	wire [4-1:0] node12120;
	wire [4-1:0] node12121;
	wire [4-1:0] node12122;
	wire [4-1:0] node12123;
	wire [4-1:0] node12124;
	wire [4-1:0] node12125;
	wire [4-1:0] node12127;
	wire [4-1:0] node12130;
	wire [4-1:0] node12131;
	wire [4-1:0] node12134;
	wire [4-1:0] node12136;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12142;
	wire [4-1:0] node12146;
	wire [4-1:0] node12148;
	wire [4-1:0] node12151;
	wire [4-1:0] node12153;
	wire [4-1:0] node12156;
	wire [4-1:0] node12157;
	wire [4-1:0] node12158;
	wire [4-1:0] node12160;
	wire [4-1:0] node12163;
	wire [4-1:0] node12164;
	wire [4-1:0] node12166;
	wire [4-1:0] node12169;
	wire [4-1:0] node12171;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12181;
	wire [4-1:0] node12183;
	wire [4-1:0] node12186;
	wire [4-1:0] node12187;
	wire [4-1:0] node12191;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12196;
	wire [4-1:0] node12200;
	wire [4-1:0] node12201;
	wire [4-1:0] node12203;
	wire [4-1:0] node12204;
	wire [4-1:0] node12207;
	wire [4-1:0] node12210;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12217;
	wire [4-1:0] node12218;
	wire [4-1:0] node12219;
	wire [4-1:0] node12221;
	wire [4-1:0] node12224;
	wire [4-1:0] node12226;
	wire [4-1:0] node12229;
	wire [4-1:0] node12230;
	wire [4-1:0] node12232;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12245;
	wire [4-1:0] node12247;
	wire [4-1:0] node12250;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12256;
	wire [4-1:0] node12258;
	wire [4-1:0] node12261;
	wire [4-1:0] node12262;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12274;
	wire [4-1:0] node12275;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12284;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12292;
	wire [4-1:0] node12295;
	wire [4-1:0] node12296;
	wire [4-1:0] node12297;
	wire [4-1:0] node12299;
	wire [4-1:0] node12302;
	wire [4-1:0] node12304;
	wire [4-1:0] node12307;
	wire [4-1:0] node12309;
	wire [4-1:0] node12312;
	wire [4-1:0] node12313;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12318;
	wire [4-1:0] node12319;
	wire [4-1:0] node12323;
	wire [4-1:0] node12324;
	wire [4-1:0] node12328;
	wire [4-1:0] node12329;
	wire [4-1:0] node12331;
	wire [4-1:0] node12333;
	wire [4-1:0] node12336;
	wire [4-1:0] node12337;
	wire [4-1:0] node12341;
	wire [4-1:0] node12342;
	wire [4-1:0] node12343;
	wire [4-1:0] node12347;
	wire [4-1:0] node12349;
	wire [4-1:0] node12352;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12355;
	wire [4-1:0] node12357;
	wire [4-1:0] node12360;
	wire [4-1:0] node12362;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12371;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12377;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12386;
	wire [4-1:0] node12389;
	wire [4-1:0] node12392;
	wire [4-1:0] node12393;
	wire [4-1:0] node12394;
	wire [4-1:0] node12398;
	wire [4-1:0] node12399;
	wire [4-1:0] node12401;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12409;
	wire [4-1:0] node12410;
	wire [4-1:0] node12411;
	wire [4-1:0] node12412;
	wire [4-1:0] node12413;
	wire [4-1:0] node12414;
	wire [4-1:0] node12416;
	wire [4-1:0] node12419;
	wire [4-1:0] node12421;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12426;
	wire [4-1:0] node12428;
	wire [4-1:0] node12431;
	wire [4-1:0] node12433;
	wire [4-1:0] node12436;
	wire [4-1:0] node12437;
	wire [4-1:0] node12440;
	wire [4-1:0] node12443;
	wire [4-1:0] node12444;
	wire [4-1:0] node12445;
	wire [4-1:0] node12447;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12453;
	wire [4-1:0] node12454;
	wire [4-1:0] node12458;
	wire [4-1:0] node12460;
	wire [4-1:0] node12463;
	wire [4-1:0] node12464;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12475;
	wire [4-1:0] node12476;
	wire [4-1:0] node12479;
	wire [4-1:0] node12480;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12487;
	wire [4-1:0] node12488;
	wire [4-1:0] node12491;
	wire [4-1:0] node12492;
	wire [4-1:0] node12495;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12506;
	wire [4-1:0] node12509;
	wire [4-1:0] node12510;
	wire [4-1:0] node12511;
	wire [4-1:0] node12512;
	wire [4-1:0] node12515;
	wire [4-1:0] node12519;
	wire [4-1:0] node12520;
	wire [4-1:0] node12521;
	wire [4-1:0] node12524;
	wire [4-1:0] node12527;
	wire [4-1:0] node12529;
	wire [4-1:0] node12532;
	wire [4-1:0] node12533;
	wire [4-1:0] node12534;
	wire [4-1:0] node12535;
	wire [4-1:0] node12536;
	wire [4-1:0] node12540;
	wire [4-1:0] node12541;
	wire [4-1:0] node12545;
	wire [4-1:0] node12546;
	wire [4-1:0] node12547;
	wire [4-1:0] node12549;
	wire [4-1:0] node12553;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12560;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12564;
	wire [4-1:0] node12567;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12573;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12578;
	wire [4-1:0] node12582;
	wire [4-1:0] node12583;
	wire [4-1:0] node12585;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12593;
	wire [4-1:0] node12595;
	wire [4-1:0] node12596;
	wire [4-1:0] node12598;
	wire [4-1:0] node12601;
	wire [4-1:0] node12604;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12609;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12616;
	wire [4-1:0] node12619;
	wire [4-1:0] node12620;
	wire [4-1:0] node12621;
	wire [4-1:0] node12624;
	wire [4-1:0] node12626;
	wire [4-1:0] node12627;
	wire [4-1:0] node12631;
	wire [4-1:0] node12632;
	wire [4-1:0] node12633;
	wire [4-1:0] node12638;
	wire [4-1:0] node12639;
	wire [4-1:0] node12640;
	wire [4-1:0] node12641;
	wire [4-1:0] node12643;
	wire [4-1:0] node12646;
	wire [4-1:0] node12647;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12654;
	wire [4-1:0] node12657;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12667;
	wire [4-1:0] node12669;
	wire [4-1:0] node12672;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12677;
	wire [4-1:0] node12681;
	wire [4-1:0] node12682;
	wire [4-1:0] node12683;
	wire [4-1:0] node12684;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12694;
	wire [4-1:0] node12695;
	wire [4-1:0] node12699;
	wire [4-1:0] node12700;
	wire [4-1:0] node12701;
	wire [4-1:0] node12704;
	wire [4-1:0] node12707;
	wire [4-1:0] node12708;
	wire [4-1:0] node12710;
	wire [4-1:0] node12713;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12719;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12731;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12739;
	wire [4-1:0] node12740;
	wire [4-1:0] node12741;
	wire [4-1:0] node12742;
	wire [4-1:0] node12744;
	wire [4-1:0] node12745;
	wire [4-1:0] node12749;
	wire [4-1:0] node12751;
	wire [4-1:0] node12753;
	wire [4-1:0] node12756;
	wire [4-1:0] node12757;
	wire [4-1:0] node12758;
	wire [4-1:0] node12759;
	wire [4-1:0] node12763;
	wire [4-1:0] node12766;
	wire [4-1:0] node12767;
	wire [4-1:0] node12770;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12775;
	wire [4-1:0] node12777;
	wire [4-1:0] node12781;
	wire [4-1:0] node12782;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12790;
	wire [4-1:0] node12791;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12796;
	wire [4-1:0] node12797;
	wire [4-1:0] node12800;
	wire [4-1:0] node12803;
	wire [4-1:0] node12804;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12812;
	wire [4-1:0] node12815;
	wire [4-1:0] node12816;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12821;
	wire [4-1:0] node12824;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12835;
	wire [4-1:0] node12836;
	wire [4-1:0] node12838;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12846;
	wire [4-1:0] node12847;
	wire [4-1:0] node12848;
	wire [4-1:0] node12849;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12855;
	wire [4-1:0] node12859;
	wire [4-1:0] node12860;
	wire [4-1:0] node12864;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12869;
	wire [4-1:0] node12871;
	wire [4-1:0] node12874;
	wire [4-1:0] node12876;
	wire [4-1:0] node12879;
	wire [4-1:0] node12880;
	wire [4-1:0] node12881;
	wire [4-1:0] node12882;
	wire [4-1:0] node12883;
	wire [4-1:0] node12884;
	wire [4-1:0] node12887;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12899;
	wire [4-1:0] node12900;
	wire [4-1:0] node12903;
	wire [4-1:0] node12904;
	wire [4-1:0] node12907;
	wire [4-1:0] node12910;
	wire [4-1:0] node12911;
	wire [4-1:0] node12912;
	wire [4-1:0] node12913;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12923;
	wire [4-1:0] node12926;
	wire [4-1:0] node12929;
	wire [4-1:0] node12930;
	wire [4-1:0] node12931;
	wire [4-1:0] node12932;
	wire [4-1:0] node12933;
	wire [4-1:0] node12937;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12945;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12951;
	wire [4-1:0] node12952;
	wire [4-1:0] node12955;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12960;
	wire [4-1:0] node12964;
	wire [4-1:0] node12966;
	wire [4-1:0] node12969;
	wire [4-1:0] node12970;
	wire [4-1:0] node12972;
	wire [4-1:0] node12973;
	wire [4-1:0] node12977;
	wire [4-1:0] node12978;
	wire [4-1:0] node12981;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12986;
	wire [4-1:0] node12987;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12997;
	wire [4-1:0] node12999;
	wire [4-1:0] node13000;
	wire [4-1:0] node13003;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13014;
	wire [4-1:0] node13016;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13022;
	wire [4-1:0] node13025;
	wire [4-1:0] node13026;
	wire [4-1:0] node13030;
	wire [4-1:0] node13031;
	wire [4-1:0] node13033;
	wire [4-1:0] node13036;
	wire [4-1:0] node13038;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13044;
	wire [4-1:0] node13047;
	wire [4-1:0] node13049;
	wire [4-1:0] node13050;
	wire [4-1:0] node13054;
	wire [4-1:0] node13055;
	wire [4-1:0] node13056;
	wire [4-1:0] node13057;
	wire [4-1:0] node13058;
	wire [4-1:0] node13061;
	wire [4-1:0] node13064;
	wire [4-1:0] node13065;
	wire [4-1:0] node13068;
	wire [4-1:0] node13071;
	wire [4-1:0] node13072;
	wire [4-1:0] node13073;
	wire [4-1:0] node13077;
	wire [4-1:0] node13078;
	wire [4-1:0] node13081;
	wire [4-1:0] node13084;
	wire [4-1:0] node13085;
	wire [4-1:0] node13086;
	wire [4-1:0] node13088;
	wire [4-1:0] node13092;
	wire [4-1:0] node13094;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13102;
	wire [4-1:0] node13103;
	wire [4-1:0] node13104;
	wire [4-1:0] node13108;
	wire [4-1:0] node13109;
	wire [4-1:0] node13111;
	wire [4-1:0] node13114;
	wire [4-1:0] node13115;
	wire [4-1:0] node13119;
	wire [4-1:0] node13120;
	wire [4-1:0] node13121;
	wire [4-1:0] node13123;
	wire [4-1:0] node13126;
	wire [4-1:0] node13129;
	wire [4-1:0] node13130;
	wire [4-1:0] node13132;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13150;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13154;
	wire [4-1:0] node13157;
	wire [4-1:0] node13159;
	wire [4-1:0] node13162;
	wire [4-1:0] node13164;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13169;
	wire [4-1:0] node13170;
	wire [4-1:0] node13172;
	wire [4-1:0] node13175;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13181;
	wire [4-1:0] node13184;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13189;
	wire [4-1:0] node13191;
	wire [4-1:0] node13194;
	wire [4-1:0] node13196;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13201;
	wire [4-1:0] node13203;
	wire [4-1:0] node13206;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13213;
	wire [4-1:0] node13214;
	wire [4-1:0] node13216;
	wire [4-1:0] node13217;
	wire [4-1:0] node13220;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13230;
	wire [4-1:0] node13231;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13238;
	wire [4-1:0] node13241;
	wire [4-1:0] node13242;
	wire [4-1:0] node13246;
	wire [4-1:0] node13247;
	wire [4-1:0] node13248;
	wire [4-1:0] node13250;
	wire [4-1:0] node13252;
	wire [4-1:0] node13255;
	wire [4-1:0] node13257;
	wire [4-1:0] node13260;
	wire [4-1:0] node13261;
	wire [4-1:0] node13265;
	wire [4-1:0] node13267;
	wire [4-1:0] node13268;
	wire [4-1:0] node13269;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13276;
	wire [4-1:0] node13278;
	wire [4-1:0] node13281;
	wire [4-1:0] node13282;
	wire [4-1:0] node13283;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13294;
	wire [4-1:0] node13295;
	wire [4-1:0] node13296;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13300;
	wire [4-1:0] node13301;
	wire [4-1:0] node13305;
	wire [4-1:0] node13306;
	wire [4-1:0] node13309;
	wire [4-1:0] node13312;
	wire [4-1:0] node13313;
	wire [4-1:0] node13314;
	wire [4-1:0] node13318;
	wire [4-1:0] node13320;
	wire [4-1:0] node13323;
	wire [4-1:0] node13324;
	wire [4-1:0] node13325;
	wire [4-1:0] node13328;
	wire [4-1:0] node13329;
	wire [4-1:0] node13331;
	wire [4-1:0] node13335;
	wire [4-1:0] node13336;
	wire [4-1:0] node13338;
	wire [4-1:0] node13341;
	wire [4-1:0] node13343;
	wire [4-1:0] node13346;
	wire [4-1:0] node13347;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13354;
	wire [4-1:0] node13355;
	wire [4-1:0] node13359;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13366;
	wire [4-1:0] node13369;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13375;
	wire [4-1:0] node13378;
	wire [4-1:0] node13379;
	wire [4-1:0] node13384;
	wire [4-1:0] node13385;
	wire [4-1:0] node13386;
	wire [4-1:0] node13387;
	wire [4-1:0] node13388;
	wire [4-1:0] node13389;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13393;
	wire [4-1:0] node13396;
	wire [4-1:0] node13397;
	wire [4-1:0] node13399;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13407;
	wire [4-1:0] node13408;
	wire [4-1:0] node13409;
	wire [4-1:0] node13410;
	wire [4-1:0] node13415;
	wire [4-1:0] node13416;
	wire [4-1:0] node13417;
	wire [4-1:0] node13421;
	wire [4-1:0] node13423;
	wire [4-1:0] node13426;
	wire [4-1:0] node13427;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13431;
	wire [4-1:0] node13435;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13440;
	wire [4-1:0] node13444;
	wire [4-1:0] node13445;
	wire [4-1:0] node13446;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13451;
	wire [4-1:0] node13455;
	wire [4-1:0] node13456;
	wire [4-1:0] node13458;
	wire [4-1:0] node13461;
	wire [4-1:0] node13464;
	wire [4-1:0] node13466;
	wire [4-1:0] node13468;
	wire [4-1:0] node13471;
	wire [4-1:0] node13472;
	wire [4-1:0] node13473;
	wire [4-1:0] node13474;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13480;
	wire [4-1:0] node13482;
	wire [4-1:0] node13485;
	wire [4-1:0] node13486;
	wire [4-1:0] node13488;
	wire [4-1:0] node13490;
	wire [4-1:0] node13493;
	wire [4-1:0] node13495;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13503;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13513;
	wire [4-1:0] node13516;
	wire [4-1:0] node13517;
	wire [4-1:0] node13519;
	wire [4-1:0] node13522;
	wire [4-1:0] node13524;
	wire [4-1:0] node13525;
	wire [4-1:0] node13529;
	wire [4-1:0] node13530;
	wire [4-1:0] node13531;
	wire [4-1:0] node13533;
	wire [4-1:0] node13534;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13550;
	wire [4-1:0] node13551;
	wire [4-1:0] node13554;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13564;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13567;
	wire [4-1:0] node13568;
	wire [4-1:0] node13570;
	wire [4-1:0] node13573;
	wire [4-1:0] node13576;
	wire [4-1:0] node13578;
	wire [4-1:0] node13581;
	wire [4-1:0] node13582;
	wire [4-1:0] node13583;
	wire [4-1:0] node13586;
	wire [4-1:0] node13589;
	wire [4-1:0] node13591;
	wire [4-1:0] node13594;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13601;
	wire [4-1:0] node13602;
	wire [4-1:0] node13606;
	wire [4-1:0] node13607;
	wire [4-1:0] node13608;
	wire [4-1:0] node13612;
	wire [4-1:0] node13613;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13624;
	wire [4-1:0] node13627;
	wire [4-1:0] node13629;
	wire [4-1:0] node13630;
	wire [4-1:0] node13634;
	wire [4-1:0] node13635;
	wire [4-1:0] node13636;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13646;
	wire [4-1:0] node13647;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13651;
	wire [4-1:0] node13653;
	wire [4-1:0] node13654;
	wire [4-1:0] node13658;
	wire [4-1:0] node13659;
	wire [4-1:0] node13661;
	wire [4-1:0] node13664;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13670;
	wire [4-1:0] node13671;
	wire [4-1:0] node13673;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13681;
	wire [4-1:0] node13682;
	wire [4-1:0] node13683;
	wire [4-1:0] node13686;
	wire [4-1:0] node13689;
	wire [4-1:0] node13690;
	wire [4-1:0] node13694;
	wire [4-1:0] node13695;
	wire [4-1:0] node13696;
	wire [4-1:0] node13697;
	wire [4-1:0] node13698;
	wire [4-1:0] node13699;
	wire [4-1:0] node13703;
	wire [4-1:0] node13706;
	wire [4-1:0] node13708;
	wire [4-1:0] node13711;
	wire [4-1:0] node13712;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13723;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13726;
	wire [4-1:0] node13727;
	wire [4-1:0] node13729;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13737;
	wire [4-1:0] node13739;
	wire [4-1:0] node13742;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13746;
	wire [4-1:0] node13749;
	wire [4-1:0] node13750;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13766;
	wire [4-1:0] node13769;
	wire [4-1:0] node13770;
	wire [4-1:0] node13771;
	wire [4-1:0] node13772;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13779;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13788;
	wire [4-1:0] node13789;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13796;
	wire [4-1:0] node13800;
	wire [4-1:0] node13801;
	wire [4-1:0] node13802;
	wire [4-1:0] node13805;
	wire [4-1:0] node13809;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13814;
	wire [4-1:0] node13817;
	wire [4-1:0] node13820;
	wire [4-1:0] node13821;
	wire [4-1:0] node13822;
	wire [4-1:0] node13823;
	wire [4-1:0] node13824;
	wire [4-1:0] node13827;
	wire [4-1:0] node13830;
	wire [4-1:0] node13831;
	wire [4-1:0] node13832;
	wire [4-1:0] node13836;
	wire [4-1:0] node13839;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13842;
	wire [4-1:0] node13843;
	wire [4-1:0] node13846;
	wire [4-1:0] node13849;
	wire [4-1:0] node13850;
	wire [4-1:0] node13853;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13860;
	wire [4-1:0] node13863;
	wire [4-1:0] node13864;
	wire [4-1:0] node13868;
	wire [4-1:0] node13869;
	wire [4-1:0] node13870;
	wire [4-1:0] node13871;
	wire [4-1:0] node13872;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13881;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13887;
	wire [4-1:0] node13889;
	wire [4-1:0] node13892;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13898;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13903;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13914;
	wire [4-1:0] node13917;
	wire [4-1:0] node13920;
	wire [4-1:0] node13922;
	wire [4-1:0] node13923;
	wire [4-1:0] node13927;
	wire [4-1:0] node13928;
	wire [4-1:0] node13929;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13934;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13943;
	wire [4-1:0] node13945;
	wire [4-1:0] node13948;
	wire [4-1:0] node13949;
	wire [4-1:0] node13950;
	wire [4-1:0] node13951;
	wire [4-1:0] node13952;
	wire [4-1:0] node13954;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13963;
	wire [4-1:0] node13967;
	wire [4-1:0] node13968;
	wire [4-1:0] node13971;
	wire [4-1:0] node13974;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13977;
	wire [4-1:0] node13980;
	wire [4-1:0] node13983;
	wire [4-1:0] node13986;
	wire [4-1:0] node13987;
	wire [4-1:0] node13988;
	wire [4-1:0] node13989;
	wire [4-1:0] node13993;
	wire [4-1:0] node13996;
	wire [4-1:0] node13998;
	wire [4-1:0] node14001;
	wire [4-1:0] node14002;
	wire [4-1:0] node14003;
	wire [4-1:0] node14004;
	wire [4-1:0] node14006;
	wire [4-1:0] node14010;
	wire [4-1:0] node14011;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14017;
	wire [4-1:0] node14018;
	wire [4-1:0] node14021;
	wire [4-1:0] node14024;
	wire [4-1:0] node14026;
	wire [4-1:0] node14028;
	wire [4-1:0] node14031;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14038;
	wire [4-1:0] node14039;
	wire [4-1:0] node14044;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14047;
	wire [4-1:0] node14048;
	wire [4-1:0] node14049;
	wire [4-1:0] node14051;
	wire [4-1:0] node14052;
	wire [4-1:0] node14054;
	wire [4-1:0] node14057;
	wire [4-1:0] node14058;
	wire [4-1:0] node14062;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14070;
	wire [4-1:0] node14072;
	wire [4-1:0] node14075;
	wire [4-1:0] node14076;
	wire [4-1:0] node14077;
	wire [4-1:0] node14081;
	wire [4-1:0] node14084;
	wire [4-1:0] node14085;
	wire [4-1:0] node14087;
	wire [4-1:0] node14089;
	wire [4-1:0] node14092;
	wire [4-1:0] node14093;
	wire [4-1:0] node14095;
	wire [4-1:0] node14099;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14102;
	wire [4-1:0] node14103;
	wire [4-1:0] node14104;
	wire [4-1:0] node14109;
	wire [4-1:0] node14110;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14116;
	wire [4-1:0] node14117;
	wire [4-1:0] node14121;
	wire [4-1:0] node14122;
	wire [4-1:0] node14126;
	wire [4-1:0] node14127;
	wire [4-1:0] node14131;
	wire [4-1:0] node14132;
	wire [4-1:0] node14133;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14143;
	wire [4-1:0] node14145;
	wire [4-1:0] node14146;
	wire [4-1:0] node14150;
	wire [4-1:0] node14151;
	wire [4-1:0] node14152;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14155;
	wire [4-1:0] node14158;
	wire [4-1:0] node14159;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14168;
	wire [4-1:0] node14171;
	wire [4-1:0] node14174;
	wire [4-1:0] node14175;
	wire [4-1:0] node14177;
	wire [4-1:0] node14180;
	wire [4-1:0] node14183;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14188;
	wire [4-1:0] node14189;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14195;
	wire [4-1:0] node14199;
	wire [4-1:0] node14200;
	wire [4-1:0] node14202;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14209;
	wire [4-1:0] node14212;
	wire [4-1:0] node14213;
	wire [4-1:0] node14214;
	wire [4-1:0] node14215;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14222;
	wire [4-1:0] node14225;
	wire [4-1:0] node14226;
	wire [4-1:0] node14228;
	wire [4-1:0] node14230;
	wire [4-1:0] node14233;
	wire [4-1:0] node14234;
	wire [4-1:0] node14235;
	wire [4-1:0] node14240;
	wire [4-1:0] node14241;
	wire [4-1:0] node14242;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14254;
	wire [4-1:0] node14255;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14262;
	wire [4-1:0] node14265;
	wire [4-1:0] node14266;
	wire [4-1:0] node14267;
	wire [4-1:0] node14268;
	wire [4-1:0] node14269;
	wire [4-1:0] node14270;
	wire [4-1:0] node14272;
	wire [4-1:0] node14275;
	wire [4-1:0] node14276;
	wire [4-1:0] node14279;
	wire [4-1:0] node14282;
	wire [4-1:0] node14283;
	wire [4-1:0] node14285;
	wire [4-1:0] node14288;
	wire [4-1:0] node14290;
	wire [4-1:0] node14293;
	wire [4-1:0] node14294;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14308;
	wire [4-1:0] node14312;
	wire [4-1:0] node14313;
	wire [4-1:0] node14314;
	wire [4-1:0] node14315;
	wire [4-1:0] node14316;
	wire [4-1:0] node14320;
	wire [4-1:0] node14321;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14330;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14337;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14344;
	wire [4-1:0] node14347;
	wire [4-1:0] node14348;
	wire [4-1:0] node14351;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14357;
	wire [4-1:0] node14360;
	wire [4-1:0] node14361;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14367;
	wire [4-1:0] node14368;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14374;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14386;
	wire [4-1:0] node14388;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14401;
	wire [4-1:0] node14404;
	wire [4-1:0] node14406;
	wire [4-1:0] node14407;
	wire [4-1:0] node14409;
	wire [4-1:0] node14412;
	wire [4-1:0] node14414;
	wire [4-1:0] node14415;
	wire [4-1:0] node14418;
	wire [4-1:0] node14421;
	wire [4-1:0] node14422;
	wire [4-1:0] node14423;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14428;
	wire [4-1:0] node14429;
	wire [4-1:0] node14433;
	wire [4-1:0] node14435;
	wire [4-1:0] node14437;
	wire [4-1:0] node14440;
	wire [4-1:0] node14442;
	wire [4-1:0] node14443;
	wire [4-1:0] node14448;
	wire [4-1:0] node14449;
	wire [4-1:0] node14450;
	wire [4-1:0] node14451;
	wire [4-1:0] node14452;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14459;
	wire [4-1:0] node14461;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14468;
	wire [4-1:0] node14469;
	wire [4-1:0] node14471;
	wire [4-1:0] node14474;
	wire [4-1:0] node14477;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14482;
	wire [4-1:0] node14483;
	wire [4-1:0] node14484;
	wire [4-1:0] node14488;
	wire [4-1:0] node14491;
	wire [4-1:0] node14492;
	wire [4-1:0] node14495;
	wire [4-1:0] node14498;
	wire [4-1:0] node14499;
	wire [4-1:0] node14500;
	wire [4-1:0] node14501;
	wire [4-1:0] node14502;
	wire [4-1:0] node14505;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14525;
	wire [4-1:0] node14527;
	wire [4-1:0] node14530;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14535;
	wire [4-1:0] node14539;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14548;
	wire [4-1:0] node14550;
	wire [4-1:0] node14551;
	wire [4-1:0] node14554;
	wire [4-1:0] node14557;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14562;
	wire [4-1:0] node14566;
	wire [4-1:0] node14568;
	wire [4-1:0] node14571;
	wire [4-1:0] node14572;
	wire [4-1:0] node14573;
	wire [4-1:0] node14574;
	wire [4-1:0] node14579;
	wire [4-1:0] node14581;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14589;
	wire [4-1:0] node14591;
	wire [4-1:0] node14593;
	wire [4-1:0] node14596;
	wire [4-1:0] node14597;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14605;
	wire [4-1:0] node14606;
	wire [4-1:0] node14607;
	wire [4-1:0] node14608;
	wire [4-1:0] node14610;
	wire [4-1:0] node14613;
	wire [4-1:0] node14614;
	wire [4-1:0] node14617;
	wire [4-1:0] node14620;
	wire [4-1:0] node14621;
	wire [4-1:0] node14623;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14632;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14636;
	wire [4-1:0] node14637;
	wire [4-1:0] node14640;
	wire [4-1:0] node14642;
	wire [4-1:0] node14643;
	wire [4-1:0] node14647;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14658;
	wire [4-1:0] node14659;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14672;
	wire [4-1:0] node14673;
	wire [4-1:0] node14674;
	wire [4-1:0] node14675;
	wire [4-1:0] node14678;
	wire [4-1:0] node14683;
	wire [4-1:0] node14684;
	wire [4-1:0] node14685;
	wire [4-1:0] node14686;
	wire [4-1:0] node14687;
	wire [4-1:0] node14690;
	wire [4-1:0] node14691;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14697;
	wire [4-1:0] node14700;
	wire [4-1:0] node14704;
	wire [4-1:0] node14706;
	wire [4-1:0] node14707;
	wire [4-1:0] node14710;
	wire [4-1:0] node14714;
	wire [4-1:0] node14715;
	wire [4-1:0] node14716;
	wire [4-1:0] node14717;
	wire [4-1:0] node14719;
	wire [4-1:0] node14721;
	wire [4-1:0] node14722;
	wire [4-1:0] node14725;
	wire [4-1:0] node14728;
	wire [4-1:0] node14729;
	wire [4-1:0] node14730;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14738;
	wire [4-1:0] node14739;
	wire [4-1:0] node14740;
	wire [4-1:0] node14743;
	wire [4-1:0] node14749;
	wire [4-1:0] node14750;
	wire [4-1:0] node14751;
	wire [4-1:0] node14752;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14756;
	wire [4-1:0] node14757;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14760;
	wire [4-1:0] node14762;
	wire [4-1:0] node14763;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14769;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14778;
	wire [4-1:0] node14779;
	wire [4-1:0] node14781;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14787;
	wire [4-1:0] node14789;
	wire [4-1:0] node14792;
	wire [4-1:0] node14793;
	wire [4-1:0] node14797;
	wire [4-1:0] node14798;
	wire [4-1:0] node14800;
	wire [4-1:0] node14803;
	wire [4-1:0] node14804;
	wire [4-1:0] node14809;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14816;
	wire [4-1:0] node14818;
	wire [4-1:0] node14821;
	wire [4-1:0] node14823;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14832;
	wire [4-1:0] node14836;
	wire [4-1:0] node14837;
	wire [4-1:0] node14840;
	wire [4-1:0] node14843;
	wire [4-1:0] node14844;
	wire [4-1:0] node14845;
	wire [4-1:0] node14846;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14855;
	wire [4-1:0] node14856;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14867;
	wire [4-1:0] node14869;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14876;
	wire [4-1:0] node14877;
	wire [4-1:0] node14878;
	wire [4-1:0] node14879;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14887;
	wire [4-1:0] node14888;
	wire [4-1:0] node14889;
	wire [4-1:0] node14891;
	wire [4-1:0] node14894;
	wire [4-1:0] node14896;
	wire [4-1:0] node14897;
	wire [4-1:0] node14901;
	wire [4-1:0] node14903;
	wire [4-1:0] node14905;
	wire [4-1:0] node14908;
	wire [4-1:0] node14909;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14915;
	wire [4-1:0] node14917;
	wire [4-1:0] node14920;
	wire [4-1:0] node14921;
	wire [4-1:0] node14922;
	wire [4-1:0] node14923;
	wire [4-1:0] node14924;
	wire [4-1:0] node14928;
	wire [4-1:0] node14932;
	wire [4-1:0] node14933;
	wire [4-1:0] node14934;
	wire [4-1:0] node14936;
	wire [4-1:0] node14940;
	wire [4-1:0] node14941;
	wire [4-1:0] node14943;
	wire [4-1:0] node14946;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14952;
	wire [4-1:0] node14953;
	wire [4-1:0] node14955;
	wire [4-1:0] node14958;
	wire [4-1:0] node14959;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14971;
	wire [4-1:0] node14974;
	wire [4-1:0] node14975;
	wire [4-1:0] node14977;
	wire [4-1:0] node14978;
	wire [4-1:0] node14982;
	wire [4-1:0] node14983;
	wire [4-1:0] node14985;
	wire [4-1:0] node14989;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14995;
	wire [4-1:0] node14996;
	wire [4-1:0] node14998;
	wire [4-1:0] node15001;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15008;
	wire [4-1:0] node15009;
	wire [4-1:0] node15012;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15019;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15025;
	wire [4-1:0] node15027;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15033;
	wire [4-1:0] node15038;
	wire [4-1:0] node15039;
	wire [4-1:0] node15040;
	wire [4-1:0] node15041;
	wire [4-1:0] node15042;
	wire [4-1:0] node15044;
	wire [4-1:0] node15045;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15053;
	wire [4-1:0] node15055;
	wire [4-1:0] node15058;
	wire [4-1:0] node15059;
	wire [4-1:0] node15060;
	wire [4-1:0] node15061;
	wire [4-1:0] node15065;
	wire [4-1:0] node15067;
	wire [4-1:0] node15070;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15075;
	wire [4-1:0] node15078;
	wire [4-1:0] node15081;
	wire [4-1:0] node15082;
	wire [4-1:0] node15083;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15087;
	wire [4-1:0] node15090;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15095;
	wire [4-1:0] node15099;
	wire [4-1:0] node15101;
	wire [4-1:0] node15104;
	wire [4-1:0] node15105;
	wire [4-1:0] node15107;
	wire [4-1:0] node15110;
	wire [4-1:0] node15112;
	wire [4-1:0] node15115;
	wire [4-1:0] node15116;
	wire [4-1:0] node15118;
	wire [4-1:0] node15119;
	wire [4-1:0] node15122;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15127;
	wire [4-1:0] node15131;
	wire [4-1:0] node15132;
	wire [4-1:0] node15136;
	wire [4-1:0] node15137;
	wire [4-1:0] node15138;
	wire [4-1:0] node15139;
	wire [4-1:0] node15140;
	wire [4-1:0] node15144;
	wire [4-1:0] node15145;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15152;
	wire [4-1:0] node15153;
	wire [4-1:0] node15157;
	wire [4-1:0] node15159;
	wire [4-1:0] node15160;
	wire [4-1:0] node15163;
	wire [4-1:0] node15166;
	wire [4-1:0] node15167;
	wire [4-1:0] node15168;
	wire [4-1:0] node15169;
	wire [4-1:0] node15171;
	wire [4-1:0] node15174;
	wire [4-1:0] node15176;
	wire [4-1:0] node15179;
	wire [4-1:0] node15180;
	wire [4-1:0] node15181;
	wire [4-1:0] node15185;
	wire [4-1:0] node15187;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15196;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15203;
	wire [4-1:0] node15204;
	wire [4-1:0] node15205;
	wire [4-1:0] node15206;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15211;
	wire [4-1:0] node15213;
	wire [4-1:0] node15214;
	wire [4-1:0] node15217;
	wire [4-1:0] node15220;
	wire [4-1:0] node15221;
	wire [4-1:0] node15223;
	wire [4-1:0] node15227;
	wire [4-1:0] node15228;
	wire [4-1:0] node15229;
	wire [4-1:0] node15230;
	wire [4-1:0] node15234;
	wire [4-1:0] node15235;
	wire [4-1:0] node15239;
	wire [4-1:0] node15240;
	wire [4-1:0] node15241;
	wire [4-1:0] node15245;
	wire [4-1:0] node15246;
	wire [4-1:0] node15248;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15255;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15263;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15271;
	wire [4-1:0] node15273;
	wire [4-1:0] node15274;
	wire [4-1:0] node15275;
	wire [4-1:0] node15280;
	wire [4-1:0] node15281;
	wire [4-1:0] node15282;
	wire [4-1:0] node15286;
	wire [4-1:0] node15288;
	wire [4-1:0] node15291;
	wire [4-1:0] node15292;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15301;
	wire [4-1:0] node15303;
	wire [4-1:0] node15306;
	wire [4-1:0] node15307;
	wire [4-1:0] node15308;
	wire [4-1:0] node15311;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15318;
	wire [4-1:0] node15319;
	wire [4-1:0] node15321;
	wire [4-1:0] node15325;
	wire [4-1:0] node15326;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15332;
	wire [4-1:0] node15333;
	wire [4-1:0] node15334;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15339;
	wire [4-1:0] node15341;
	wire [4-1:0] node15344;
	wire [4-1:0] node15347;
	wire [4-1:0] node15349;
	wire [4-1:0] node15350;
	wire [4-1:0] node15354;
	wire [4-1:0] node15355;
	wire [4-1:0] node15356;
	wire [4-1:0] node15357;
	wire [4-1:0] node15361;
	wire [4-1:0] node15364;
	wire [4-1:0] node15365;
	wire [4-1:0] node15368;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15375;
	wire [4-1:0] node15378;
	wire [4-1:0] node15379;
	wire [4-1:0] node15380;
	wire [4-1:0] node15385;
	wire [4-1:0] node15387;
	wire [4-1:0] node15390;
	wire [4-1:0] node15391;
	wire [4-1:0] node15392;
	wire [4-1:0] node15393;
	wire [4-1:0] node15395;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15401;
	wire [4-1:0] node15405;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15408;
	wire [4-1:0] node15412;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15418;
	wire [4-1:0] node15421;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15426;
	wire [4-1:0] node15427;
	wire [4-1:0] node15431;
	wire [4-1:0] node15432;
	wire [4-1:0] node15435;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15442;
	wire [4-1:0] node15445;
	wire [4-1:0] node15446;
	wire [4-1:0] node15447;
	wire [4-1:0] node15448;
	wire [4-1:0] node15449;
	wire [4-1:0] node15450;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15457;
	wire [4-1:0] node15460;
	wire [4-1:0] node15463;
	wire [4-1:0] node15464;
	wire [4-1:0] node15466;
	wire [4-1:0] node15469;
	wire [4-1:0] node15472;
	wire [4-1:0] node15473;
	wire [4-1:0] node15474;
	wire [4-1:0] node15476;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15484;
	wire [4-1:0] node15486;
	wire [4-1:0] node15488;
	wire [4-1:0] node15491;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15495;
	wire [4-1:0] node15499;
	wire [4-1:0] node15501;
	wire [4-1:0] node15503;
	wire [4-1:0] node15506;
	wire [4-1:0] node15508;
	wire [4-1:0] node15510;
	wire [4-1:0] node15513;
	wire [4-1:0] node15514;
	wire [4-1:0] node15515;
	wire [4-1:0] node15516;
	wire [4-1:0] node15520;
	wire [4-1:0] node15523;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15534;
	wire [4-1:0] node15535;
	wire [4-1:0] node15536;
	wire [4-1:0] node15537;
	wire [4-1:0] node15538;
	wire [4-1:0] node15539;
	wire [4-1:0] node15540;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15547;
	wire [4-1:0] node15551;
	wire [4-1:0] node15553;
	wire [4-1:0] node15556;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15562;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15578;
	wire [4-1:0] node15579;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15586;
	wire [4-1:0] node15587;
	wire [4-1:0] node15590;
	wire [4-1:0] node15592;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15602;
	wire [4-1:0] node15603;
	wire [4-1:0] node15606;
	wire [4-1:0] node15609;
	wire [4-1:0] node15610;
	wire [4-1:0] node15611;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15622;
	wire [4-1:0] node15623;
	wire [4-1:0] node15624;
	wire [4-1:0] node15628;
	wire [4-1:0] node15629;
	wire [4-1:0] node15630;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15643;
	wire [4-1:0] node15644;
	wire [4-1:0] node15647;
	wire [4-1:0] node15650;
	wire [4-1:0] node15651;
	wire [4-1:0] node15653;
	wire [4-1:0] node15656;
	wire [4-1:0] node15657;
	wire [4-1:0] node15661;
	wire [4-1:0] node15662;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15668;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15675;
	wire [4-1:0] node15678;
	wire [4-1:0] node15679;
	wire [4-1:0] node15680;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15687;
	wire [4-1:0] node15688;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15695;
	wire [4-1:0] node15696;
	wire [4-1:0] node15700;
	wire [4-1:0] node15703;
	wire [4-1:0] node15705;
	wire [4-1:0] node15708;
	wire [4-1:0] node15709;
	wire [4-1:0] node15711;
	wire [4-1:0] node15712;
	wire [4-1:0] node15716;
	wire [4-1:0] node15718;
	wire [4-1:0] node15721;
	wire [4-1:0] node15722;
	wire [4-1:0] node15723;
	wire [4-1:0] node15724;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15727;
	wire [4-1:0] node15728;
	wire [4-1:0] node15732;
	wire [4-1:0] node15733;
	wire [4-1:0] node15737;
	wire [4-1:0] node15738;
	wire [4-1:0] node15741;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15747;
	wire [4-1:0] node15749;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15755;
	wire [4-1:0] node15756;
	wire [4-1:0] node15759;
	wire [4-1:0] node15760;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15767;
	wire [4-1:0] node15768;
	wire [4-1:0] node15771;
	wire [4-1:0] node15774;
	wire [4-1:0] node15776;
	wire [4-1:0] node15779;
	wire [4-1:0] node15780;
	wire [4-1:0] node15782;
	wire [4-1:0] node15785;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15791;
	wire [4-1:0] node15792;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15799;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15807;
	wire [4-1:0] node15811;
	wire [4-1:0] node15813;
	wire [4-1:0] node15816;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15819;
	wire [4-1:0] node15820;
	wire [4-1:0] node15821;
	wire [4-1:0] node15825;
	wire [4-1:0] node15827;
	wire [4-1:0] node15830;
	wire [4-1:0] node15831;
	wire [4-1:0] node15834;
	wire [4-1:0] node15837;
	wire [4-1:0] node15838;
	wire [4-1:0] node15839;
	wire [4-1:0] node15840;
	wire [4-1:0] node15844;
	wire [4-1:0] node15847;
	wire [4-1:0] node15849;
	wire [4-1:0] node15852;
	wire [4-1:0] node15853;
	wire [4-1:0] node15854;
	wire [4-1:0] node15855;
	wire [4-1:0] node15858;
	wire [4-1:0] node15862;
	wire [4-1:0] node15863;
	wire [4-1:0] node15866;
	wire [4-1:0] node15867;
	wire [4-1:0] node15870;
	wire [4-1:0] node15873;
	wire [4-1:0] node15874;
	wire [4-1:0] node15875;
	wire [4-1:0] node15876;
	wire [4-1:0] node15877;
	wire [4-1:0] node15878;
	wire [4-1:0] node15879;
	wire [4-1:0] node15883;
	wire [4-1:0] node15886;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15892;
	wire [4-1:0] node15893;
	wire [4-1:0] node15895;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15903;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15908;
	wire [4-1:0] node15909;
	wire [4-1:0] node15913;
	wire [4-1:0] node15914;
	wire [4-1:0] node15915;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15926;
	wire [4-1:0] node15927;
	wire [4-1:0] node15928;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15934;
	wire [4-1:0] node15937;
	wire [4-1:0] node15938;
	wire [4-1:0] node15939;
	wire [4-1:0] node15944;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15948;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15960;
	wire [4-1:0] node15962;
	wire [4-1:0] node15965;
	wire [4-1:0] node15966;
	wire [4-1:0] node15967;
	wire [4-1:0] node15968;
	wire [4-1:0] node15969;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15975;
	wire [4-1:0] node15978;
	wire [4-1:0] node15979;
	wire [4-1:0] node15983;
	wire [4-1:0] node15986;
	wire [4-1:0] node15987;
	wire [4-1:0] node15989;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15999;
	wire [4-1:0] node16000;
	wire [4-1:0] node16001;
	wire [4-1:0] node16003;
	wire [4-1:0] node16006;
	wire [4-1:0] node16009;
	wire [4-1:0] node16010;
	wire [4-1:0] node16014;
	wire [4-1:0] node16015;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16018;
	wire [4-1:0] node16019;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16022;
	wire [4-1:0] node16023;
	wire [4-1:0] node16027;
	wire [4-1:0] node16029;
	wire [4-1:0] node16032;
	wire [4-1:0] node16033;
	wire [4-1:0] node16037;
	wire [4-1:0] node16038;
	wire [4-1:0] node16039;
	wire [4-1:0] node16042;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16048;
	wire [4-1:0] node16051;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16056;
	wire [4-1:0] node16059;
	wire [4-1:0] node16060;
	wire [4-1:0] node16064;
	wire [4-1:0] node16065;
	wire [4-1:0] node16066;
	wire [4-1:0] node16070;
	wire [4-1:0] node16071;
	wire [4-1:0] node16074;
	wire [4-1:0] node16077;
	wire [4-1:0] node16078;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16089;
	wire [4-1:0] node16090;
	wire [4-1:0] node16091;
	wire [4-1:0] node16093;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16098;
	wire [4-1:0] node16103;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16114;
	wire [4-1:0] node16115;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16118;
	wire [4-1:0] node16119;
	wire [4-1:0] node16122;
	wire [4-1:0] node16125;
	wire [4-1:0] node16126;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16132;
	wire [4-1:0] node16133;
	wire [4-1:0] node16137;
	wire [4-1:0] node16140;
	wire [4-1:0] node16141;
	wire [4-1:0] node16143;
	wire [4-1:0] node16146;
	wire [4-1:0] node16149;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16152;
	wire [4-1:0] node16155;
	wire [4-1:0] node16156;
	wire [4-1:0] node16160;
	wire [4-1:0] node16163;
	wire [4-1:0] node16164;
	wire [4-1:0] node16165;
	wire [4-1:0] node16168;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16175;
	wire [4-1:0] node16178;
	wire [4-1:0] node16179;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16184;
	wire [4-1:0] node16186;
	wire [4-1:0] node16188;
	wire [4-1:0] node16191;
	wire [4-1:0] node16192;
	wire [4-1:0] node16193;
	wire [4-1:0] node16197;
	wire [4-1:0] node16198;
	wire [4-1:0] node16200;
	wire [4-1:0] node16203;
	wire [4-1:0] node16205;
	wire [4-1:0] node16208;
	wire [4-1:0] node16209;
	wire [4-1:0] node16210;
	wire [4-1:0] node16211;
	wire [4-1:0] node16214;
	wire [4-1:0] node16216;
	wire [4-1:0] node16219;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16225;
	wire [4-1:0] node16227;
	wire [4-1:0] node16230;
	wire [4-1:0] node16231;
	wire [4-1:0] node16232;
	wire [4-1:0] node16235;
	wire [4-1:0] node16237;
	wire [4-1:0] node16240;
	wire [4-1:0] node16243;
	wire [4-1:0] node16244;
	wire [4-1:0] node16245;
	wire [4-1:0] node16246;
	wire [4-1:0] node16247;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16257;
	wire [4-1:0] node16260;
	wire [4-1:0] node16261;
	wire [4-1:0] node16263;
	wire [4-1:0] node16266;
	wire [4-1:0] node16267;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16276;
	wire [4-1:0] node16278;
	wire [4-1:0] node16281;
	wire [4-1:0] node16282;
	wire [4-1:0] node16285;
	wire [4-1:0] node16286;
	wire [4-1:0] node16290;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16295;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16302;
	wire [4-1:0] node16305;
	wire [4-1:0] node16307;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16315;
	wire [4-1:0] node16317;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16323;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16329;
	wire [4-1:0] node16330;
	wire [4-1:0] node16332;
	wire [4-1:0] node16335;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16346;
	wire [4-1:0] node16347;
	wire [4-1:0] node16348;
	wire [4-1:0] node16350;
	wire [4-1:0] node16353;
	wire [4-1:0] node16355;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16365;
	wire [4-1:0] node16366;
	wire [4-1:0] node16367;
	wire [4-1:0] node16371;
	wire [4-1:0] node16372;
	wire [4-1:0] node16376;
	wire [4-1:0] node16377;
	wire [4-1:0] node16379;
	wire [4-1:0] node16382;
	wire [4-1:0] node16383;
	wire [4-1:0] node16386;
	wire [4-1:0] node16389;
	wire [4-1:0] node16391;
	wire [4-1:0] node16393;
	wire [4-1:0] node16396;
	wire [4-1:0] node16397;
	wire [4-1:0] node16398;
	wire [4-1:0] node16399;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16403;
	wire [4-1:0] node16404;
	wire [4-1:0] node16407;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16416;
	wire [4-1:0] node16417;
	wire [4-1:0] node16421;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16426;
	wire [4-1:0] node16430;
	wire [4-1:0] node16433;
	wire [4-1:0] node16434;
	wire [4-1:0] node16436;
	wire [4-1:0] node16439;
	wire [4-1:0] node16442;
	wire [4-1:0] node16443;
	wire [4-1:0] node16444;
	wire [4-1:0] node16446;
	wire [4-1:0] node16448;
	wire [4-1:0] node16451;
	wire [4-1:0] node16452;
	wire [4-1:0] node16453;
	wire [4-1:0] node16456;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16464;
	wire [4-1:0] node16465;
	wire [4-1:0] node16466;
	wire [4-1:0] node16468;
	wire [4-1:0] node16471;
	wire [4-1:0] node16474;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16481;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16484;
	wire [4-1:0] node16485;
	wire [4-1:0] node16486;
	wire [4-1:0] node16489;
	wire [4-1:0] node16491;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16497;
	wire [4-1:0] node16500;
	wire [4-1:0] node16503;
	wire [4-1:0] node16504;
	wire [4-1:0] node16506;
	wire [4-1:0] node16508;
	wire [4-1:0] node16511;
	wire [4-1:0] node16513;
	wire [4-1:0] node16516;
	wire [4-1:0] node16517;
	wire [4-1:0] node16519;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16527;
	wire [4-1:0] node16528;
	wire [4-1:0] node16529;
	wire [4-1:0] node16530;
	wire [4-1:0] node16533;
	wire [4-1:0] node16536;
	wire [4-1:0] node16537;
	wire [4-1:0] node16538;
	wire [4-1:0] node16540;
	wire [4-1:0] node16545;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16550;
	wire [4-1:0] node16554;
	wire [4-1:0] node16555;
	wire [4-1:0] node16556;
	wire [4-1:0] node16557;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16562;
	wire [4-1:0] node16564;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16569;
	wire [4-1:0] node16573;
	wire [4-1:0] node16574;
	wire [4-1:0] node16577;
	wire [4-1:0] node16580;
	wire [4-1:0] node16581;
	wire [4-1:0] node16582;
	wire [4-1:0] node16583;
	wire [4-1:0] node16586;
	wire [4-1:0] node16587;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16594;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16602;
	wire [4-1:0] node16603;
	wire [4-1:0] node16605;
	wire [4-1:0] node16608;
	wire [4-1:0] node16610;
	wire [4-1:0] node16613;
	wire [4-1:0] node16614;
	wire [4-1:0] node16615;
	wire [4-1:0] node16616;
	wire [4-1:0] node16617;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16625;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16636;
	wire [4-1:0] node16637;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16643;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16651;
	wire [4-1:0] node16652;
	wire [4-1:0] node16653;
	wire [4-1:0] node16656;
	wire [4-1:0] node16662;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16667;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16676;
	wire [4-1:0] node16677;
	wire [4-1:0] node16680;
	wire [4-1:0] node16683;
	wire [4-1:0] node16684;
	wire [4-1:0] node16686;
	wire [4-1:0] node16687;
	wire [4-1:0] node16690;
	wire [4-1:0] node16694;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16699;
	wire [4-1:0] node16703;
	wire [4-1:0] node16705;
	wire [4-1:0] node16706;
	wire [4-1:0] node16707;
	wire [4-1:0] node16709;
	wire [4-1:0] node16710;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16716;
	wire [4-1:0] node16717;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16724;
	wire [4-1:0] node16726;
	wire [4-1:0] node16729;
	wire [4-1:0] node16730;
	wire [4-1:0] node16731;
	wire [4-1:0] node16733;
	wire [4-1:0] node16736;
	wire [4-1:0] node16737;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16747;
	wire [4-1:0] node16748;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16757;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16761;
	wire [4-1:0] node16763;
	wire [4-1:0] node16766;
	wire [4-1:0] node16768;
	wire [4-1:0] node16770;
	wire [4-1:0] node16773;
	wire [4-1:0] node16774;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16784;
	wire [4-1:0] node16785;
	wire [4-1:0] node16787;
	wire [4-1:0] node16790;
	wire [4-1:0] node16791;
	wire [4-1:0] node16795;
	wire [4-1:0] node16796;
	wire [4-1:0] node16797;
	wire [4-1:0] node16798;
	wire [4-1:0] node16799;
	wire [4-1:0] node16803;
	wire [4-1:0] node16806;
	wire [4-1:0] node16807;
	wire [4-1:0] node16808;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16816;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16822;
	wire [4-1:0] node16825;
	wire [4-1:0] node16827;
	wire [4-1:0] node16830;
	wire [4-1:0] node16831;
	wire [4-1:0] node16832;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16835;
	wire [4-1:0] node16836;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16843;
	wire [4-1:0] node16847;
	wire [4-1:0] node16848;
	wire [4-1:0] node16849;
	wire [4-1:0] node16850;
	wire [4-1:0] node16852;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16858;
	wire [4-1:0] node16861;
	wire [4-1:0] node16865;
	wire [4-1:0] node16867;
	wire [4-1:0] node16868;
	wire [4-1:0] node16870;
	wire [4-1:0] node16873;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16878;
	wire [4-1:0] node16880;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16887;
	wire [4-1:0] node16891;
	wire [4-1:0] node16892;
	wire [4-1:0] node16894;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16901;
	wire [4-1:0] node16902;
	wire [4-1:0] node16904;
	wire [4-1:0] node16908;
	wire [4-1:0] node16909;
	wire [4-1:0] node16910;
	wire [4-1:0] node16912;
	wire [4-1:0] node16915;
	wire [4-1:0] node16916;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16923;
	wire [4-1:0] node16926;
	wire [4-1:0] node16929;
	wire [4-1:0] node16930;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16937;
	wire [4-1:0] node16938;
	wire [4-1:0] node16942;
	wire [4-1:0] node16943;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16953;
	wire [4-1:0] node16956;
	wire [4-1:0] node16957;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16965;
	wire [4-1:0] node16967;
	wire [4-1:0] node16970;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16979;
	wire [4-1:0] node16980;
	wire [4-1:0] node16984;
	wire [4-1:0] node16985;
	wire [4-1:0] node16989;
	wire [4-1:0] node16990;
	wire [4-1:0] node16991;
	wire [4-1:0] node16992;
	wire [4-1:0] node16993;
	wire [4-1:0] node16996;
	wire [4-1:0] node16999;
	wire [4-1:0] node17000;
	wire [4-1:0] node17002;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17010;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17015;
	wire [4-1:0] node17017;
	wire [4-1:0] node17019;
	wire [4-1:0] node17022;
	wire [4-1:0] node17023;
	wire [4-1:0] node17027;
	wire [4-1:0] node17028;
	wire [4-1:0] node17030;
	wire [4-1:0] node17034;
	wire [4-1:0] node17035;
	wire [4-1:0] node17036;
	wire [4-1:0] node17037;
	wire [4-1:0] node17038;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17041;
	wire [4-1:0] node17045;
	wire [4-1:0] node17048;
	wire [4-1:0] node17050;
	wire [4-1:0] node17051;
	wire [4-1:0] node17054;
	wire [4-1:0] node17057;
	wire [4-1:0] node17058;
	wire [4-1:0] node17060;
	wire [4-1:0] node17064;
	wire [4-1:0] node17065;
	wire [4-1:0] node17066;
	wire [4-1:0] node17068;
	wire [4-1:0] node17072;
	wire [4-1:0] node17073;
	wire [4-1:0] node17074;
	wire [4-1:0] node17076;
	wire [4-1:0] node17080;
	wire [4-1:0] node17082;
	wire [4-1:0] node17085;
	wire [4-1:0] node17086;
	wire [4-1:0] node17087;
	wire [4-1:0] node17088;
	wire [4-1:0] node17089;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17096;
	wire [4-1:0] node17100;
	wire [4-1:0] node17101;
	wire [4-1:0] node17102;
	wire [4-1:0] node17105;
	wire [4-1:0] node17108;
	wire [4-1:0] node17109;
	wire [4-1:0] node17112;
	wire [4-1:0] node17113;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17119;
	wire [4-1:0] node17120;
	wire [4-1:0] node17125;
	wire [4-1:0] node17127;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17134;
	wire [4-1:0] node17137;
	wire [4-1:0] node17138;
	wire [4-1:0] node17141;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17151;
	wire [4-1:0] node17152;
	wire [4-1:0] node17157;
	wire [4-1:0] node17158;
	wire [4-1:0] node17159;
	wire [4-1:0] node17161;
	wire [4-1:0] node17163;
	wire [4-1:0] node17166;
	wire [4-1:0] node17167;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17178;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17181;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17187;
	wire [4-1:0] node17190;
	wire [4-1:0] node17192;
	wire [4-1:0] node17195;
	wire [4-1:0] node17196;
	wire [4-1:0] node17197;
	wire [4-1:0] node17198;
	wire [4-1:0] node17202;
	wire [4-1:0] node17203;
	wire [4-1:0] node17209;
	wire [4-1:0] node17211;
	wire [4-1:0] node17213;
	wire [4-1:0] node17214;
	wire [4-1:0] node17215;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17224;
	wire [4-1:0] node17225;
	wire [4-1:0] node17228;
	wire [4-1:0] node17230;
	wire [4-1:0] node17233;
	wire [4-1:0] node17234;
	wire [4-1:0] node17235;
	wire [4-1:0] node17236;
	wire [4-1:0] node17240;
	wire [4-1:0] node17242;
	wire [4-1:0] node17245;
	wire [4-1:0] node17246;
	wire [4-1:0] node17249;
	wire [4-1:0] node17250;
	wire [4-1:0] node17251;
	wire [4-1:0] node17254;
	wire [4-1:0] node17257;
	wire [4-1:0] node17259;
	wire [4-1:0] node17263;
	wire [4-1:0] node17264;
	wire [4-1:0] node17265;
	wire [4-1:0] node17266;
	wire [4-1:0] node17267;
	wire [4-1:0] node17268;
	wire [4-1:0] node17269;
	wire [4-1:0] node17274;
	wire [4-1:0] node17276;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17284;
	wire [4-1:0] node17285;
	wire [4-1:0] node17286;
	wire [4-1:0] node17287;
	wire [4-1:0] node17289;
	wire [4-1:0] node17293;
	wire [4-1:0] node17294;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17303;
	wire [4-1:0] node17307;
	wire [4-1:0] node17308;
	wire [4-1:0] node17309;
	wire [4-1:0] node17310;
	wire [4-1:0] node17312;
	wire [4-1:0] node17315;
	wire [4-1:0] node17316;
	wire [4-1:0] node17318;
	wire [4-1:0] node17321;
	wire [4-1:0] node17324;
	wire [4-1:0] node17325;
	wire [4-1:0] node17326;
	wire [4-1:0] node17327;
	wire [4-1:0] node17331;
	wire [4-1:0] node17335;
	wire [4-1:0] node17336;
	wire [4-1:0] node17337;
	wire [4-1:0] node17339;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17347;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17350;
	wire [4-1:0] node17351;
	wire [4-1:0] node17352;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17359;
	wire [4-1:0] node17360;
	wire [4-1:0] node17362;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17370;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17381;
	wire [4-1:0] node17382;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17388;
	wire [4-1:0] node17392;
	wire [4-1:0] node17393;
	wire [4-1:0] node17397;
	wire [4-1:0] node17398;
	wire [4-1:0] node17399;
	wire [4-1:0] node17401;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17407;
	wire [4-1:0] node17412;
	wire [4-1:0] node17414;
	wire [4-1:0] node17416;
	wire [4-1:0] node17417;
	wire [4-1:0] node17418;
	wire [4-1:0] node17420;
	wire [4-1:0] node17423;
	wire [4-1:0] node17424;
	wire [4-1:0] node17426;
	wire [4-1:0] node17429;
	wire [4-1:0] node17432;
	wire [4-1:0] node17434;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17441;
	wire [4-1:0] node17442;
	wire [4-1:0] node17443;
	wire [4-1:0] node17444;
	wire [4-1:0] node17445;
	wire [4-1:0] node17447;
	wire [4-1:0] node17450;
	wire [4-1:0] node17452;
	wire [4-1:0] node17454;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17459;
	wire [4-1:0] node17463;
	wire [4-1:0] node17466;
	wire [4-1:0] node17467;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17473;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17479;
	wire [4-1:0] node17482;
	wire [4-1:0] node17483;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17489;
	wire [4-1:0] node17490;
	wire [4-1:0] node17494;
	wire [4-1:0] node17496;
	wire [4-1:0] node17498;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17504;
	wire [4-1:0] node17505;
	wire [4-1:0] node17507;
	wire [4-1:0] node17510;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17517;
	wire [4-1:0] node17520;
	wire [4-1:0] node17521;
	wire [4-1:0] node17523;
	wire [4-1:0] node17525;
	wire [4-1:0] node17528;
	wire [4-1:0] node17529;
	wire [4-1:0] node17530;
	wire [4-1:0] node17532;
	wire [4-1:0] node17535;
	wire [4-1:0] node17536;
	wire [4-1:0] node17541;
	wire [4-1:0] node17542;
	wire [4-1:0] node17543;
	wire [4-1:0] node17544;
	wire [4-1:0] node17547;
	wire [4-1:0] node17549;
	wire [4-1:0] node17552;
	wire [4-1:0] node17553;
	wire [4-1:0] node17555;
	wire [4-1:0] node17558;
	wire [4-1:0] node17560;
	wire [4-1:0] node17563;
	wire [4-1:0] node17564;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17570;
	wire [4-1:0] node17572;
	wire [4-1:0] node17574;
	wire [4-1:0] node17577;
	wire [4-1:0] node17578;
	wire [4-1:0] node17579;
	wire [4-1:0] node17581;
	wire [4-1:0] node17585;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17592;
	wire [4-1:0] node17593;
	wire [4-1:0] node17594;
	wire [4-1:0] node17595;
	wire [4-1:0] node17596;
	wire [4-1:0] node17597;
	wire [4-1:0] node17599;
	wire [4-1:0] node17602;
	wire [4-1:0] node17603;
	wire [4-1:0] node17604;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17612;
	wire [4-1:0] node17615;
	wire [4-1:0] node17616;
	wire [4-1:0] node17618;
	wire [4-1:0] node17622;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17628;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17637;
	wire [4-1:0] node17638;
	wire [4-1:0] node17639;
	wire [4-1:0] node17643;
	wire [4-1:0] node17645;
	wire [4-1:0] node17648;
	wire [4-1:0] node17649;
	wire [4-1:0] node17650;
	wire [4-1:0] node17654;
	wire [4-1:0] node17655;
	wire [4-1:0] node17656;
	wire [4-1:0] node17660;
	wire [4-1:0] node17662;
	wire [4-1:0] node17665;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17670;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17677;
	wire [4-1:0] node17681;
	wire [4-1:0] node17683;
	wire [4-1:0] node17684;
	wire [4-1:0] node17688;
	wire [4-1:0] node17689;
	wire [4-1:0] node17690;
	wire [4-1:0] node17691;
	wire [4-1:0] node17692;
	wire [4-1:0] node17693;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17701;
	wire [4-1:0] node17704;
	wire [4-1:0] node17705;
	wire [4-1:0] node17706;
	wire [4-1:0] node17710;
	wire [4-1:0] node17712;
	wire [4-1:0] node17713;
	wire [4-1:0] node17717;
	wire [4-1:0] node17718;
	wire [4-1:0] node17719;
	wire [4-1:0] node17723;
	wire [4-1:0] node17724;
	wire [4-1:0] node17726;
	wire [4-1:0] node17729;
	wire [4-1:0] node17731;
	wire [4-1:0] node17734;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17738;
	wire [4-1:0] node17741;
	wire [4-1:0] node17743;
	wire [4-1:0] node17746;
	wire [4-1:0] node17747;
	wire [4-1:0] node17749;
	wire [4-1:0] node17752;
	wire [4-1:0] node17754;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17760;
	wire [4-1:0] node17763;
	wire [4-1:0] node17765;
	wire [4-1:0] node17768;
	wire [4-1:0] node17769;
	wire [4-1:0] node17770;
	wire [4-1:0] node17771;
	wire [4-1:0] node17773;
	wire [4-1:0] node17777;
	wire [4-1:0] node17779;
	wire [4-1:0] node17782;
	wire [4-1:0] node17783;
	wire [4-1:0] node17785;
	wire [4-1:0] node17788;
	wire [4-1:0] node17789;
	wire [4-1:0] node17790;
	wire [4-1:0] node17794;
	wire [4-1:0] node17796;
	wire [4-1:0] node17799;
	wire [4-1:0] node17801;
	wire [4-1:0] node17802;
	wire [4-1:0] node17803;
	wire [4-1:0] node17804;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17808;
	wire [4-1:0] node17810;
	wire [4-1:0] node17812;
	wire [4-1:0] node17815;
	wire [4-1:0] node17817;
	wire [4-1:0] node17820;
	wire [4-1:0] node17822;
	wire [4-1:0] node17826;
	wire [4-1:0] node17827;
	wire [4-1:0] node17828;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17833;
	wire [4-1:0] node17834;
	wire [4-1:0] node17835;
	wire [4-1:0] node17838;
	wire [4-1:0] node17842;
	wire [4-1:0] node17843;
	wire [4-1:0] node17844;
	wire [4-1:0] node17848;
	wire [4-1:0] node17850;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17855;
	wire [4-1:0] node17857;
	wire [4-1:0] node17860;
	wire [4-1:0] node17862;
	wire [4-1:0] node17865;
	wire [4-1:0] node17866;
	wire [4-1:0] node17868;
	wire [4-1:0] node17870;
	wire [4-1:0] node17873;
	wire [4-1:0] node17876;
	wire [4-1:0] node17878;
	wire [4-1:0] node17879;
	wire [4-1:0] node17880;
	wire [4-1:0] node17883;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17892;
	wire [4-1:0] node17894;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17900;
	wire [4-1:0] node17901;
	wire [4-1:0] node17903;
	wire [4-1:0] node17906;
	wire [4-1:0] node17907;
	wire [4-1:0] node17909;
	wire [4-1:0] node17913;
	wire [4-1:0] node17914;
	wire [4-1:0] node17915;
	wire [4-1:0] node17916;
	wire [4-1:0] node17920;
	wire [4-1:0] node17922;
	wire [4-1:0] node17923;
	wire [4-1:0] node17927;
	wire [4-1:0] node17928;
	wire [4-1:0] node17930;
	wire [4-1:0] node17933;
	wire [4-1:0] node17935;
	wire [4-1:0] node17938;
	wire [4-1:0] node17939;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17943;
	wire [4-1:0] node17947;
	wire [4-1:0] node17948;
	wire [4-1:0] node17949;
	wire [4-1:0] node17953;
	wire [4-1:0] node17954;
	wire [4-1:0] node17958;
	wire [4-1:0] node17959;
	wire [4-1:0] node17961;
	wire [4-1:0] node17964;
	wire [4-1:0] node17965;
	wire [4-1:0] node17967;
	wire [4-1:0] node17970;
	wire [4-1:0] node17971;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17978;
	wire [4-1:0] node17980;
	wire [4-1:0] node17981;
	wire [4-1:0] node17984;
	wire [4-1:0] node17986;
	wire [4-1:0] node17989;
	wire [4-1:0] node17990;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17998;
	wire [4-1:0] node17999;
	wire [4-1:0] node18000;
	wire [4-1:0] node18001;
	wire [4-1:0] node18004;
	wire [4-1:0] node18006;
	wire [4-1:0] node18009;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18015;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18022;
	wire [4-1:0] node18023;
	wire [4-1:0] node18027;
	wire [4-1:0] node18028;
	wire [4-1:0] node18029;
	wire [4-1:0] node18031;
	wire [4-1:0] node18033;
	wire [4-1:0] node18035;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18044;
	wire [4-1:0] node18046;
	wire [4-1:0] node18049;
	wire [4-1:0] node18050;
	wire [4-1:0] node18051;
	wire [4-1:0] node18053;
	wire [4-1:0] node18056;
	wire [4-1:0] node18059;
	wire [4-1:0] node18060;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18069;
	wire [4-1:0] node18070;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18073;
	wire [4-1:0] node18074;
	wire [4-1:0] node18075;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18078;
	wire [4-1:0] node18081;
	wire [4-1:0] node18082;
	wire [4-1:0] node18086;
	wire [4-1:0] node18087;
	wire [4-1:0] node18088;
	wire [4-1:0] node18091;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18098;
	wire [4-1:0] node18101;
	wire [4-1:0] node18102;
	wire [4-1:0] node18103;
	wire [4-1:0] node18105;
	wire [4-1:0] node18108;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18115;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18123;
	wire [4-1:0] node18124;
	wire [4-1:0] node18125;
	wire [4-1:0] node18128;
	wire [4-1:0] node18131;
	wire [4-1:0] node18132;
	wire [4-1:0] node18136;
	wire [4-1:0] node18137;
	wire [4-1:0] node18138;
	wire [4-1:0] node18139;
	wire [4-1:0] node18140;
	wire [4-1:0] node18143;
	wire [4-1:0] node18147;
	wire [4-1:0] node18148;
	wire [4-1:0] node18149;
	wire [4-1:0] node18152;
	wire [4-1:0] node18155;
	wire [4-1:0] node18157;
	wire [4-1:0] node18160;
	wire [4-1:0] node18161;
	wire [4-1:0] node18163;
	wire [4-1:0] node18164;
	wire [4-1:0] node18166;
	wire [4-1:0] node18169;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18176;
	wire [4-1:0] node18177;
	wire [4-1:0] node18181;
	wire [4-1:0] node18182;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18185;
	wire [4-1:0] node18186;
	wire [4-1:0] node18190;
	wire [4-1:0] node18191;
	wire [4-1:0] node18195;
	wire [4-1:0] node18196;
	wire [4-1:0] node18197;
	wire [4-1:0] node18201;
	wire [4-1:0] node18202;
	wire [4-1:0] node18206;
	wire [4-1:0] node18207;
	wire [4-1:0] node18209;
	wire [4-1:0] node18212;
	wire [4-1:0] node18214;
	wire [4-1:0] node18215;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18221;
	wire [4-1:0] node18223;
	wire [4-1:0] node18226;
	wire [4-1:0] node18227;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18232;
	wire [4-1:0] node18235;
	wire [4-1:0] node18239;
	wire [4-1:0] node18240;
	wire [4-1:0] node18241;
	wire [4-1:0] node18242;
	wire [4-1:0] node18245;
	wire [4-1:0] node18246;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18257;
	wire [4-1:0] node18258;
	wire [4-1:0] node18259;
	wire [4-1:0] node18260;
	wire [4-1:0] node18265;
	wire [4-1:0] node18266;
	wire [4-1:0] node18267;
	wire [4-1:0] node18271;
	wire [4-1:0] node18273;
	wire [4-1:0] node18276;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18280;
	wire [4-1:0] node18281;
	wire [4-1:0] node18285;
	wire [4-1:0] node18286;
	wire [4-1:0] node18288;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18295;
	wire [4-1:0] node18296;
	wire [4-1:0] node18300;
	wire [4-1:0] node18303;
	wire [4-1:0] node18305;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18313;
	wire [4-1:0] node18314;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18319;
	wire [4-1:0] node18323;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18338;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18344;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18349;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18355;
	wire [4-1:0] node18357;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18363;
	wire [4-1:0] node18366;
	wire [4-1:0] node18368;
	wire [4-1:0] node18371;
	wire [4-1:0] node18372;
	wire [4-1:0] node18375;
	wire [4-1:0] node18376;
	wire [4-1:0] node18377;
	wire [4-1:0] node18381;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18387;
	wire [4-1:0] node18388;
	wire [4-1:0] node18389;
	wire [4-1:0] node18390;
	wire [4-1:0] node18392;
	wire [4-1:0] node18393;
	wire [4-1:0] node18397;
	wire [4-1:0] node18398;
	wire [4-1:0] node18401;
	wire [4-1:0] node18403;
	wire [4-1:0] node18406;
	wire [4-1:0] node18407;
	wire [4-1:0] node18409;
	wire [4-1:0] node18412;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18419;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18425;
	wire [4-1:0] node18428;
	wire [4-1:0] node18429;
	wire [4-1:0] node18433;
	wire [4-1:0] node18434;
	wire [4-1:0] node18435;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18442;
	wire [4-1:0] node18444;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18450;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18457;
	wire [4-1:0] node18458;
	wire [4-1:0] node18462;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18471;
	wire [4-1:0] node18475;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18480;
	wire [4-1:0] node18481;
	wire [4-1:0] node18482;
	wire [4-1:0] node18486;
	wire [4-1:0] node18487;
	wire [4-1:0] node18491;
	wire [4-1:0] node18492;
	wire [4-1:0] node18493;
	wire [4-1:0] node18498;
	wire [4-1:0] node18499;
	wire [4-1:0] node18500;
	wire [4-1:0] node18501;
	wire [4-1:0] node18505;
	wire [4-1:0] node18506;
	wire [4-1:0] node18509;
	wire [4-1:0] node18512;
	wire [4-1:0] node18513;
	wire [4-1:0] node18514;
	wire [4-1:0] node18518;
	wire [4-1:0] node18521;
	wire [4-1:0] node18522;
	wire [4-1:0] node18523;
	wire [4-1:0] node18524;
	wire [4-1:0] node18527;
	wire [4-1:0] node18528;
	wire [4-1:0] node18532;
	wire [4-1:0] node18533;
	wire [4-1:0] node18535;
	wire [4-1:0] node18538;
	wire [4-1:0] node18539;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18545;
	wire [4-1:0] node18549;
	wire [4-1:0] node18552;
	wire [4-1:0] node18553;
	wire [4-1:0] node18554;
	wire [4-1:0] node18555;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18560;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18567;
	wire [4-1:0] node18570;
	wire [4-1:0] node18571;
	wire [4-1:0] node18573;
	wire [4-1:0] node18575;
	wire [4-1:0] node18578;
	wire [4-1:0] node18580;
	wire [4-1:0] node18583;
	wire [4-1:0] node18584;
	wire [4-1:0] node18585;
	wire [4-1:0] node18586;
	wire [4-1:0] node18589;
	wire [4-1:0] node18593;
	wire [4-1:0] node18594;
	wire [4-1:0] node18598;
	wire [4-1:0] node18599;
	wire [4-1:0] node18600;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18606;
	wire [4-1:0] node18609;
	wire [4-1:0] node18610;
	wire [4-1:0] node18611;
	wire [4-1:0] node18615;
	wire [4-1:0] node18616;
	wire [4-1:0] node18620;
	wire [4-1:0] node18621;
	wire [4-1:0] node18622;
	wire [4-1:0] node18625;
	wire [4-1:0] node18628;
	wire [4-1:0] node18629;
	wire [4-1:0] node18631;
	wire [4-1:0] node18632;
	wire [4-1:0] node18635;
	wire [4-1:0] node18638;
	wire [4-1:0] node18640;
	wire [4-1:0] node18643;
	wire [4-1:0] node18644;
	wire [4-1:0] node18645;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18649;
	wire [4-1:0] node18652;
	wire [4-1:0] node18655;
	wire [4-1:0] node18656;
	wire [4-1:0] node18657;
	wire [4-1:0] node18659;
	wire [4-1:0] node18662;
	wire [4-1:0] node18665;
	wire [4-1:0] node18666;
	wire [4-1:0] node18669;
	wire [4-1:0] node18671;
	wire [4-1:0] node18674;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18681;
	wire [4-1:0] node18682;
	wire [4-1:0] node18684;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18691;
	wire [4-1:0] node18694;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;
	wire [4-1:0] node18701;
	wire [4-1:0] node18703;
	wire [4-1:0] node18706;
	wire [4-1:0] node18707;
	wire [4-1:0] node18708;
	wire [4-1:0] node18711;
	wire [4-1:0] node18715;
	wire [4-1:0] node18716;
	wire [4-1:0] node18717;
	wire [4-1:0] node18718;
	wire [4-1:0] node18719;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18726;
	wire [4-1:0] node18729;
	wire [4-1:0] node18730;
	wire [4-1:0] node18734;
	wire [4-1:0] node18735;
	wire [4-1:0] node18736;
	wire [4-1:0] node18740;
	wire [4-1:0] node18741;
	wire [4-1:0] node18744;
	wire [4-1:0] node18747;
	wire [4-1:0] node18748;
	wire [4-1:0] node18750;
	wire [4-1:0] node18751;
	wire [4-1:0] node18755;
	wire [4-1:0] node18756;
	wire [4-1:0] node18760;
	wire [4-1:0] node18761;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18765;
	wire [4-1:0] node18766;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18770;
	wire [4-1:0] node18773;
	wire [4-1:0] node18775;
	wire [4-1:0] node18776;
	wire [4-1:0] node18780;
	wire [4-1:0] node18782;
	wire [4-1:0] node18784;
	wire [4-1:0] node18788;
	wire [4-1:0] node18789;
	wire [4-1:0] node18790;
	wire [4-1:0] node18791;
	wire [4-1:0] node18792;
	wire [4-1:0] node18793;
	wire [4-1:0] node18794;
	wire [4-1:0] node18798;
	wire [4-1:0] node18799;
	wire [4-1:0] node18804;
	wire [4-1:0] node18805;
	wire [4-1:0] node18806;
	wire [4-1:0] node18810;
	wire [4-1:0] node18813;
	wire [4-1:0] node18814;
	wire [4-1:0] node18815;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18822;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18828;
	wire [4-1:0] node18829;
	wire [4-1:0] node18833;
	wire [4-1:0] node18834;
	wire [4-1:0] node18835;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18844;
	wire [4-1:0] node18846;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18852;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18858;
	wire [4-1:0] node18860;
	wire [4-1:0] node18862;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18875;
	wire [4-1:0] node18877;
	wire [4-1:0] node18880;
	wire [4-1:0] node18881;
	wire [4-1:0] node18882;
	wire [4-1:0] node18886;
	wire [4-1:0] node18887;
	wire [4-1:0] node18891;
	wire [4-1:0] node18892;
	wire [4-1:0] node18893;
	wire [4-1:0] node18896;
	wire [4-1:0] node18897;
	wire [4-1:0] node18901;
	wire [4-1:0] node18902;
	wire [4-1:0] node18903;
	wire [4-1:0] node18906;
	wire [4-1:0] node18908;
	wire [4-1:0] node18911;
	wire [4-1:0] node18912;
	wire [4-1:0] node18916;
	wire [4-1:0] node18917;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18921;
	wire [4-1:0] node18924;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18931;
	wire [4-1:0] node18935;
	wire [4-1:0] node18936;
	wire [4-1:0] node18940;
	wire [4-1:0] node18941;
	wire [4-1:0] node18942;
	wire [4-1:0] node18946;
	wire [4-1:0] node18947;
	wire [4-1:0] node18949;
	wire [4-1:0] node18953;
	wire [4-1:0] node18954;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18961;
	wire [4-1:0] node18962;
	wire [4-1:0] node18965;
	wire [4-1:0] node18966;
	wire [4-1:0] node18969;
	wire [4-1:0] node18970;
	wire [4-1:0] node18974;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18980;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18986;
	wire [4-1:0] node18989;
	wire [4-1:0] node18990;
	wire [4-1:0] node18991;
	wire [4-1:0] node18993;
	wire [4-1:0] node18996;
	wire [4-1:0] node18997;
	wire [4-1:0] node18999;
	wire [4-1:0] node19002;
	wire [4-1:0] node19003;
	wire [4-1:0] node19007;
	wire [4-1:0] node19008;
	wire [4-1:0] node19009;
	wire [4-1:0] node19010;
	wire [4-1:0] node19014;
	wire [4-1:0] node19016;
	wire [4-1:0] node19019;
	wire [4-1:0] node19020;
	wire [4-1:0] node19025;
	wire [4-1:0] node19026;
	wire [4-1:0] node19027;
	wire [4-1:0] node19028;
	wire [4-1:0] node19029;
	wire [4-1:0] node19030;
	wire [4-1:0] node19031;
	wire [4-1:0] node19032;
	wire [4-1:0] node19033;
	wire [4-1:0] node19034;
	wire [4-1:0] node19038;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19046;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19051;
	wire [4-1:0] node19054;
	wire [4-1:0] node19055;
	wire [4-1:0] node19057;
	wire [4-1:0] node19060;
	wire [4-1:0] node19063;
	wire [4-1:0] node19064;
	wire [4-1:0] node19065;
	wire [4-1:0] node19066;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19074;
	wire [4-1:0] node19075;
	wire [4-1:0] node19076;
	wire [4-1:0] node19080;
	wire [4-1:0] node19081;
	wire [4-1:0] node19083;
	wire [4-1:0] node19087;
	wire [4-1:0] node19088;
	wire [4-1:0] node19089;
	wire [4-1:0] node19091;
	wire [4-1:0] node19093;
	wire [4-1:0] node19096;
	wire [4-1:0] node19098;
	wire [4-1:0] node19101;
	wire [4-1:0] node19102;
	wire [4-1:0] node19105;
	wire [4-1:0] node19107;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19113;
	wire [4-1:0] node19114;
	wire [4-1:0] node19118;
	wire [4-1:0] node19119;
	wire [4-1:0] node19120;
	wire [4-1:0] node19124;
	wire [4-1:0] node19126;
	wire [4-1:0] node19129;
	wire [4-1:0] node19130;
	wire [4-1:0] node19132;
	wire [4-1:0] node19134;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19139;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19149;
	wire [4-1:0] node19150;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19153;
	wire [4-1:0] node19156;
	wire [4-1:0] node19157;
	wire [4-1:0] node19159;
	wire [4-1:0] node19162;
	wire [4-1:0] node19165;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19171;
	wire [4-1:0] node19172;
	wire [4-1:0] node19176;
	wire [4-1:0] node19177;
	wire [4-1:0] node19178;
	wire [4-1:0] node19181;
	wire [4-1:0] node19184;
	wire [4-1:0] node19187;
	wire [4-1:0] node19188;
	wire [4-1:0] node19191;
	wire [4-1:0] node19193;
	wire [4-1:0] node19196;
	wire [4-1:0] node19197;
	wire [4-1:0] node19198;
	wire [4-1:0] node19199;
	wire [4-1:0] node19202;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19207;
	wire [4-1:0] node19211;
	wire [4-1:0] node19213;
	wire [4-1:0] node19214;
	wire [4-1:0] node19217;
	wire [4-1:0] node19220;
	wire [4-1:0] node19222;
	wire [4-1:0] node19223;
	wire [4-1:0] node19224;
	wire [4-1:0] node19225;
	wire [4-1:0] node19231;
	wire [4-1:0] node19232;
	wire [4-1:0] node19233;
	wire [4-1:0] node19234;
	wire [4-1:0] node19235;
	wire [4-1:0] node19236;
	wire [4-1:0] node19237;
	wire [4-1:0] node19241;
	wire [4-1:0] node19243;
	wire [4-1:0] node19246;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19253;
	wire [4-1:0] node19254;
	wire [4-1:0] node19255;
	wire [4-1:0] node19259;
	wire [4-1:0] node19260;
	wire [4-1:0] node19261;
	wire [4-1:0] node19264;
	wire [4-1:0] node19267;
	wire [4-1:0] node19270;
	wire [4-1:0] node19271;
	wire [4-1:0] node19272;
	wire [4-1:0] node19273;
	wire [4-1:0] node19277;
	wire [4-1:0] node19278;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19285;
	wire [4-1:0] node19288;
	wire [4-1:0] node19291;
	wire [4-1:0] node19292;
	wire [4-1:0] node19293;
	wire [4-1:0] node19294;
	wire [4-1:0] node19297;
	wire [4-1:0] node19300;
	wire [4-1:0] node19301;
	wire [4-1:0] node19303;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19311;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19317;
	wire [4-1:0] node19320;
	wire [4-1:0] node19321;
	wire [4-1:0] node19322;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19327;
	wire [4-1:0] node19331;
	wire [4-1:0] node19333;
	wire [4-1:0] node19335;
	wire [4-1:0] node19338;
	wire [4-1:0] node19339;
	wire [4-1:0] node19340;
	wire [4-1:0] node19343;
	wire [4-1:0] node19347;
	wire [4-1:0] node19348;
	wire [4-1:0] node19349;
	wire [4-1:0] node19351;
	wire [4-1:0] node19354;
	wire [4-1:0] node19356;
	wire [4-1:0] node19357;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19364;
	wire [4-1:0] node19366;
	wire [4-1:0] node19370;
	wire [4-1:0] node19371;
	wire [4-1:0] node19372;
	wire [4-1:0] node19373;
	wire [4-1:0] node19374;
	wire [4-1:0] node19375;
	wire [4-1:0] node19378;
	wire [4-1:0] node19381;
	wire [4-1:0] node19383;
	wire [4-1:0] node19386;
	wire [4-1:0] node19387;
	wire [4-1:0] node19388;
	wire [4-1:0] node19391;
	wire [4-1:0] node19394;
	wire [4-1:0] node19397;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19403;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19410;
	wire [4-1:0] node19413;
	wire [4-1:0] node19416;
	wire [4-1:0] node19418;
	wire [4-1:0] node19419;
	wire [4-1:0] node19423;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19430;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19435;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19444;
	wire [4-1:0] node19446;
	wire [4-1:0] node19447;
	wire [4-1:0] node19449;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19457;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19468;
	wire [4-1:0] node19471;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19478;
	wire [4-1:0] node19481;
	wire [4-1:0] node19482;
	wire [4-1:0] node19484;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19492;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19495;
	wire [4-1:0] node19496;
	wire [4-1:0] node19497;
	wire [4-1:0] node19498;
	wire [4-1:0] node19501;
	wire [4-1:0] node19504;
	wire [4-1:0] node19505;
	wire [4-1:0] node19508;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19514;
	wire [4-1:0] node19516;
	wire [4-1:0] node19520;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19527;
	wire [4-1:0] node19529;
	wire [4-1:0] node19532;
	wire [4-1:0] node19533;
	wire [4-1:0] node19535;
	wire [4-1:0] node19538;
	wire [4-1:0] node19539;
	wire [4-1:0] node19543;
	wire [4-1:0] node19544;
	wire [4-1:0] node19545;
	wire [4-1:0] node19546;
	wire [4-1:0] node19548;
	wire [4-1:0] node19551;
	wire [4-1:0] node19552;
	wire [4-1:0] node19556;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19561;
	wire [4-1:0] node19563;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19571;
	wire [4-1:0] node19572;
	wire [4-1:0] node19573;
	wire [4-1:0] node19577;
	wire [4-1:0] node19578;
	wire [4-1:0] node19580;
	wire [4-1:0] node19583;
	wire [4-1:0] node19584;
	wire [4-1:0] node19588;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19593;
	wire [4-1:0] node19596;
	wire [4-1:0] node19599;
	wire [4-1:0] node19600;
	wire [4-1:0] node19604;
	wire [4-1:0] node19606;
	wire [4-1:0] node19607;
	wire [4-1:0] node19609;
	wire [4-1:0] node19613;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19619;
	wire [4-1:0] node19620;
	wire [4-1:0] node19624;
	wire [4-1:0] node19626;
	wire [4-1:0] node19627;
	wire [4-1:0] node19629;
	wire [4-1:0] node19632;
	wire [4-1:0] node19633;
	wire [4-1:0] node19636;
	wire [4-1:0] node19638;
	wire [4-1:0] node19639;
	wire [4-1:0] node19643;
	wire [4-1:0] node19644;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19649;
	wire [4-1:0] node19650;
	wire [4-1:0] node19652;
	wire [4-1:0] node19655;
	wire [4-1:0] node19656;
	wire [4-1:0] node19659;
	wire [4-1:0] node19662;
	wire [4-1:0] node19663;
	wire [4-1:0] node19664;
	wire [4-1:0] node19665;
	wire [4-1:0] node19670;
	wire [4-1:0] node19671;
	wire [4-1:0] node19673;
	wire [4-1:0] node19676;
	wire [4-1:0] node19678;
	wire [4-1:0] node19681;
	wire [4-1:0] node19682;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19686;
	wire [4-1:0] node19689;
	wire [4-1:0] node19691;
	wire [4-1:0] node19694;
	wire [4-1:0] node19697;
	wire [4-1:0] node19698;
	wire [4-1:0] node19699;
	wire [4-1:0] node19702;
	wire [4-1:0] node19704;
	wire [4-1:0] node19707;
	wire [4-1:0] node19708;
	wire [4-1:0] node19711;
	wire [4-1:0] node19712;
	wire [4-1:0] node19716;
	wire [4-1:0] node19717;
	wire [4-1:0] node19718;
	wire [4-1:0] node19719;
	wire [4-1:0] node19720;
	wire [4-1:0] node19724;
	wire [4-1:0] node19726;
	wire [4-1:0] node19727;
	wire [4-1:0] node19731;
	wire [4-1:0] node19733;
	wire [4-1:0] node19734;
	wire [4-1:0] node19737;
	wire [4-1:0] node19740;
	wire [4-1:0] node19741;
	wire [4-1:0] node19742;
	wire [4-1:0] node19743;
	wire [4-1:0] node19746;
	wire [4-1:0] node19749;
	wire [4-1:0] node19751;
	wire [4-1:0] node19754;
	wire [4-1:0] node19755;
	wire [4-1:0] node19756;
	wire [4-1:0] node19757;
	wire [4-1:0] node19761;
	wire [4-1:0] node19762;
	wire [4-1:0] node19766;
	wire [4-1:0] node19768;
	wire [4-1:0] node19769;
	wire [4-1:0] node19773;
	wire [4-1:0] node19774;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19781;
	wire [4-1:0] node19785;
	wire [4-1:0] node19786;
	wire [4-1:0] node19788;
	wire [4-1:0] node19791;
	wire [4-1:0] node19792;
	wire [4-1:0] node19795;
	wire [4-1:0] node19798;
	wire [4-1:0] node19799;
	wire [4-1:0] node19800;
	wire [4-1:0] node19801;
	wire [4-1:0] node19804;
	wire [4-1:0] node19806;
	wire [4-1:0] node19809;
	wire [4-1:0] node19810;
	wire [4-1:0] node19814;
	wire [4-1:0] node19815;
	wire [4-1:0] node19818;
	wire [4-1:0] node19819;
	wire [4-1:0] node19821;
	wire [4-1:0] node19825;
	wire [4-1:0] node19826;
	wire [4-1:0] node19827;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19833;
	wire [4-1:0] node19834;
	wire [4-1:0] node19835;
	wire [4-1:0] node19838;
	wire [4-1:0] node19841;
	wire [4-1:0] node19844;
	wire [4-1:0] node19845;
	wire [4-1:0] node19846;
	wire [4-1:0] node19848;
	wire [4-1:0] node19852;
	wire [4-1:0] node19854;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19859;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19865;
	wire [4-1:0] node19866;
	wire [4-1:0] node19870;
	wire [4-1:0] node19871;
	wire [4-1:0] node19874;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19881;
	wire [4-1:0] node19882;
	wire [4-1:0] node19884;
	wire [4-1:0] node19887;
	wire [4-1:0] node19890;
	wire [4-1:0] node19891;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19894;
	wire [4-1:0] node19895;
	wire [4-1:0] node19897;
	wire [4-1:0] node19900;
	wire [4-1:0] node19901;
	wire [4-1:0] node19905;
	wire [4-1:0] node19906;
	wire [4-1:0] node19908;
	wire [4-1:0] node19911;
	wire [4-1:0] node19912;
	wire [4-1:0] node19916;
	wire [4-1:0] node19917;
	wire [4-1:0] node19918;
	wire [4-1:0] node19921;
	wire [4-1:0] node19922;
	wire [4-1:0] node19927;
	wire [4-1:0] node19928;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19933;
	wire [4-1:0] node19934;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19941;
	wire [4-1:0] node19944;
	wire [4-1:0] node19946;
	wire [4-1:0] node19949;
	wire [4-1:0] node19950;
	wire [4-1:0] node19951;
	wire [4-1:0] node19953;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19960;
	wire [4-1:0] node19963;
	wire [4-1:0] node19964;
	wire [4-1:0] node19965;
	wire [4-1:0] node19967;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19976;
	wire [4-1:0] node19977;
	wire [4-1:0] node19979;
	wire [4-1:0] node19980;
	wire [4-1:0] node19981;
	wire [4-1:0] node19983;
	wire [4-1:0] node19987;
	wire [4-1:0] node19988;
	wire [4-1:0] node19990;
	wire [4-1:0] node19991;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node19999;
	wire [4-1:0] node20000;
	wire [4-1:0] node20003;
	wire [4-1:0] node20005;
	wire [4-1:0] node20009;
	wire [4-1:0] node20010;
	wire [4-1:0] node20011;
	wire [4-1:0] node20015;
	wire [4-1:0] node20016;
	wire [4-1:0] node20018;
	wire [4-1:0] node20022;
	wire [4-1:0] node20023;
	wire [4-1:0] node20024;
	wire [4-1:0] node20026;
	wire [4-1:0] node20029;
	wire [4-1:0] node20030;
	wire [4-1:0] node20035;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20040;
	wire [4-1:0] node20041;
	wire [4-1:0] node20043;
	wire [4-1:0] node20045;
	wire [4-1:0] node20048;
	wire [4-1:0] node20051;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20055;
	wire [4-1:0] node20058;
	wire [4-1:0] node20060;
	wire [4-1:0] node20063;
	wire [4-1:0] node20065;
	wire [4-1:0] node20067;
	wire [4-1:0] node20070;
	wire [4-1:0] node20071;
	wire [4-1:0] node20072;
	wire [4-1:0] node20073;
	wire [4-1:0] node20074;
	wire [4-1:0] node20077;
	wire [4-1:0] node20080;
	wire [4-1:0] node20081;
	wire [4-1:0] node20085;
	wire [4-1:0] node20086;
	wire [4-1:0] node20089;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20098;
	wire [4-1:0] node20100;
	wire [4-1:0] node20101;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20108;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20116;
	wire [4-1:0] node20117;
	wire [4-1:0] node20118;
	wire [4-1:0] node20121;
	wire [4-1:0] node20124;
	wire [4-1:0] node20126;
	wire [4-1:0] node20129;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20133;
	wire [4-1:0] node20136;
	wire [4-1:0] node20138;
	wire [4-1:0] node20141;
	wire [4-1:0] node20142;
	wire [4-1:0] node20143;
	wire [4-1:0] node20147;
	wire [4-1:0] node20149;
	wire [4-1:0] node20152;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20156;
	wire [4-1:0] node20159;
	wire [4-1:0] node20161;
	wire [4-1:0] node20164;
	wire [4-1:0] node20165;
	wire [4-1:0] node20168;
	wire [4-1:0] node20169;
	wire [4-1:0] node20170;
	wire [4-1:0] node20174;
	wire [4-1:0] node20176;
	wire [4-1:0] node20179;
	wire [4-1:0] node20180;
	wire [4-1:0] node20181;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20187;
	wire [4-1:0] node20189;
	wire [4-1:0] node20192;
	wire [4-1:0] node20193;
	wire [4-1:0] node20197;
	wire [4-1:0] node20198;
	wire [4-1:0] node20199;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20207;
	wire [4-1:0] node20209;
	wire [4-1:0] node20210;
	wire [4-1:0] node20213;
	wire [4-1:0] node20216;
	wire [4-1:0] node20217;
	wire [4-1:0] node20218;
	wire [4-1:0] node20219;
	wire [4-1:0] node20221;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20228;
	wire [4-1:0] node20231;
	wire [4-1:0] node20232;
	wire [4-1:0] node20237;
	wire [4-1:0] node20238;
	wire [4-1:0] node20239;
	wire [4-1:0] node20240;
	wire [4-1:0] node20241;
	wire [4-1:0] node20242;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20247;
	wire [4-1:0] node20251;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20257;
	wire [4-1:0] node20259;
	wire [4-1:0] node20262;
	wire [4-1:0] node20264;
	wire [4-1:0] node20265;
	wire [4-1:0] node20269;
	wire [4-1:0] node20270;
	wire [4-1:0] node20271;
	wire [4-1:0] node20273;
	wire [4-1:0] node20276;
	wire [4-1:0] node20278;
	wire [4-1:0] node20281;
	wire [4-1:0] node20282;
	wire [4-1:0] node20284;
	wire [4-1:0] node20286;
	wire [4-1:0] node20289;
	wire [4-1:0] node20292;
	wire [4-1:0] node20293;
	wire [4-1:0] node20294;
	wire [4-1:0] node20295;
	wire [4-1:0] node20296;
	wire [4-1:0] node20298;
	wire [4-1:0] node20301;
	wire [4-1:0] node20303;
	wire [4-1:0] node20306;
	wire [4-1:0] node20308;
	wire [4-1:0] node20309;
	wire [4-1:0] node20313;
	wire [4-1:0] node20314;
	wire [4-1:0] node20315;
	wire [4-1:0] node20316;
	wire [4-1:0] node20320;
	wire [4-1:0] node20323;
	wire [4-1:0] node20325;
	wire [4-1:0] node20327;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20334;
	wire [4-1:0] node20335;
	wire [4-1:0] node20337;
	wire [4-1:0] node20340;
	wire [4-1:0] node20341;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20347;
	wire [4-1:0] node20351;
	wire [4-1:0] node20353;
	wire [4-1:0] node20358;
	wire [4-1:0] node20359;
	wire [4-1:0] node20360;
	wire [4-1:0] node20361;
	wire [4-1:0] node20362;
	wire [4-1:0] node20364;
	wire [4-1:0] node20365;
	wire [4-1:0] node20366;
	wire [4-1:0] node20368;
	wire [4-1:0] node20369;
	wire [4-1:0] node20371;
	wire [4-1:0] node20374;
	wire [4-1:0] node20375;
	wire [4-1:0] node20376;
	wire [4-1:0] node20378;
	wire [4-1:0] node20381;
	wire [4-1:0] node20383;
	wire [4-1:0] node20386;
	wire [4-1:0] node20389;
	wire [4-1:0] node20390;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20394;
	wire [4-1:0] node20397;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20404;
	wire [4-1:0] node20405;
	wire [4-1:0] node20406;
	wire [4-1:0] node20408;
	wire [4-1:0] node20413;
	wire [4-1:0] node20414;
	wire [4-1:0] node20415;
	wire [4-1:0] node20419;
	wire [4-1:0] node20420;
	wire [4-1:0] node20421;
	wire [4-1:0] node20425;
	wire [4-1:0] node20428;
	wire [4-1:0] node20430;
	wire [4-1:0] node20432;
	wire [4-1:0] node20433;
	wire [4-1:0] node20434;
	wire [4-1:0] node20437;
	wire [4-1:0] node20439;
	wire [4-1:0] node20440;
	wire [4-1:0] node20443;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20449;
	wire [4-1:0] node20450;
	wire [4-1:0] node20451;
	wire [4-1:0] node20452;
	wire [4-1:0] node20453;
	wire [4-1:0] node20455;
	wire [4-1:0] node20458;
	wire [4-1:0] node20461;
	wire [4-1:0] node20462;
	wire [4-1:0] node20464;
	wire [4-1:0] node20466;
	wire [4-1:0] node20469;
	wire [4-1:0] node20470;
	wire [4-1:0] node20473;
	wire [4-1:0] node20476;
	wire [4-1:0] node20477;
	wire [4-1:0] node20478;
	wire [4-1:0] node20479;
	wire [4-1:0] node20483;
	wire [4-1:0] node20485;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20491;
	wire [4-1:0] node20492;
	wire [4-1:0] node20496;
	wire [4-1:0] node20499;
	wire [4-1:0] node20500;
	wire [4-1:0] node20501;
	wire [4-1:0] node20503;
	wire [4-1:0] node20506;
	wire [4-1:0] node20507;
	wire [4-1:0] node20509;
	wire [4-1:0] node20512;
	wire [4-1:0] node20513;
	wire [4-1:0] node20517;
	wire [4-1:0] node20518;
	wire [4-1:0] node20520;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20529;
	wire [4-1:0] node20530;
	wire [4-1:0] node20532;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20539;
	wire [4-1:0] node20541;
	wire [4-1:0] node20544;
	wire [4-1:0] node20545;
	wire [4-1:0] node20549;
	wire [4-1:0] node20550;
	wire [4-1:0] node20551;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20559;
	wire [4-1:0] node20561;
	wire [4-1:0] node20564;
	wire [4-1:0] node20565;
	wire [4-1:0] node20566;
	wire [4-1:0] node20567;
	wire [4-1:0] node20569;
	wire [4-1:0] node20572;
	wire [4-1:0] node20574;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20583;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20591;
	wire [4-1:0] node20592;
	wire [4-1:0] node20596;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20600;
	wire [4-1:0] node20603;
	wire [4-1:0] node20605;
	wire [4-1:0] node20608;
	wire [4-1:0] node20609;
	wire [4-1:0] node20612;
	wire [4-1:0] node20614;
	wire [4-1:0] node20615;
	wire [4-1:0] node20618;
	wire [4-1:0] node20621;
	wire [4-1:0] node20622;
	wire [4-1:0] node20623;
	wire [4-1:0] node20624;
	wire [4-1:0] node20625;
	wire [4-1:0] node20626;
	wire [4-1:0] node20628;
	wire [4-1:0] node20631;
	wire [4-1:0] node20633;
	wire [4-1:0] node20635;
	wire [4-1:0] node20638;
	wire [4-1:0] node20639;
	wire [4-1:0] node20640;
	wire [4-1:0] node20641;
	wire [4-1:0] node20645;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20654;
	wire [4-1:0] node20655;
	wire [4-1:0] node20656;
	wire [4-1:0] node20660;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20665;
	wire [4-1:0] node20669;
	wire [4-1:0] node20671;
	wire [4-1:0] node20674;
	wire [4-1:0] node20675;
	wire [4-1:0] node20676;
	wire [4-1:0] node20677;
	wire [4-1:0] node20679;
	wire [4-1:0] node20681;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20689;
	wire [4-1:0] node20690;
	wire [4-1:0] node20691;
	wire [4-1:0] node20692;
	wire [4-1:0] node20696;
	wire [4-1:0] node20698;
	wire [4-1:0] node20701;
	wire [4-1:0] node20702;
	wire [4-1:0] node20705;
	wire [4-1:0] node20708;
	wire [4-1:0] node20709;
	wire [4-1:0] node20710;
	wire [4-1:0] node20711;
	wire [4-1:0] node20715;
	wire [4-1:0] node20716;
	wire [4-1:0] node20720;
	wire [4-1:0] node20721;
	wire [4-1:0] node20722;
	wire [4-1:0] node20725;
	wire [4-1:0] node20728;
	wire [4-1:0] node20731;
	wire [4-1:0] node20732;
	wire [4-1:0] node20733;
	wire [4-1:0] node20734;
	wire [4-1:0] node20736;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20743;
	wire [4-1:0] node20744;
	wire [4-1:0] node20745;
	wire [4-1:0] node20749;
	wire [4-1:0] node20751;
	wire [4-1:0] node20754;
	wire [4-1:0] node20755;
	wire [4-1:0] node20757;
	wire [4-1:0] node20760;
	wire [4-1:0] node20762;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20772;
	wire [4-1:0] node20773;
	wire [4-1:0] node20777;
	wire [4-1:0] node20778;
	wire [4-1:0] node20779;
	wire [4-1:0] node20782;
	wire [4-1:0] node20783;
	wire [4-1:0] node20785;
	wire [4-1:0] node20788;
	wire [4-1:0] node20789;
	wire [4-1:0] node20792;
	wire [4-1:0] node20795;
	wire [4-1:0] node20796;
	wire [4-1:0] node20797;
	wire [4-1:0] node20800;
	wire [4-1:0] node20804;
	wire [4-1:0] node20806;
	wire [4-1:0] node20808;
	wire [4-1:0] node20809;
	wire [4-1:0] node20811;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20814;
	wire [4-1:0] node20816;
	wire [4-1:0] node20819;
	wire [4-1:0] node20822;
	wire [4-1:0] node20824;
	wire [4-1:0] node20826;
	wire [4-1:0] node20827;
	wire [4-1:0] node20832;
	wire [4-1:0] node20833;
	wire [4-1:0] node20834;
	wire [4-1:0] node20835;
	wire [4-1:0] node20836;
	wire [4-1:0] node20839;
	wire [4-1:0] node20840;
	wire [4-1:0] node20841;
	wire [4-1:0] node20845;
	wire [4-1:0] node20846;
	wire [4-1:0] node20850;
	wire [4-1:0] node20851;
	wire [4-1:0] node20853;
	wire [4-1:0] node20856;
	wire [4-1:0] node20857;
	wire [4-1:0] node20861;
	wire [4-1:0] node20862;
	wire [4-1:0] node20863;
	wire [4-1:0] node20865;
	wire [4-1:0] node20868;
	wire [4-1:0] node20871;
	wire [4-1:0] node20872;
	wire [4-1:0] node20875;
	wire [4-1:0] node20877;
	wire [4-1:0] node20880;
	wire [4-1:0] node20882;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20885;
	wire [4-1:0] node20889;
	wire [4-1:0] node20891;
	wire [4-1:0] node20894;
	wire [4-1:0] node20896;
	wire [4-1:0] node20898;
	wire [4-1:0] node20901;
	wire [4-1:0] node20902;
	wire [4-1:0] node20903;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20907;
	wire [4-1:0] node20908;
	wire [4-1:0] node20910;
	wire [4-1:0] node20913;
	wire [4-1:0] node20914;
	wire [4-1:0] node20918;
	wire [4-1:0] node20919;
	wire [4-1:0] node20923;
	wire [4-1:0] node20924;
	wire [4-1:0] node20925;
	wire [4-1:0] node20927;
	wire [4-1:0] node20928;
	wire [4-1:0] node20932;
	wire [4-1:0] node20933;
	wire [4-1:0] node20937;
	wire [4-1:0] node20938;
	wire [4-1:0] node20939;
	wire [4-1:0] node20942;
	wire [4-1:0] node20943;
	wire [4-1:0] node20947;
	wire [4-1:0] node20949;
	wire [4-1:0] node20952;
	wire [4-1:0] node20953;
	wire [4-1:0] node20954;
	wire [4-1:0] node20955;
	wire [4-1:0] node20956;
	wire [4-1:0] node20958;
	wire [4-1:0] node20961;
	wire [4-1:0] node20963;
	wire [4-1:0] node20966;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20974;
	wire [4-1:0] node20976;
	wire [4-1:0] node20979;
	wire [4-1:0] node20980;
	wire [4-1:0] node20981;
	wire [4-1:0] node20982;
	wire [4-1:0] node20987;
	wire [4-1:0] node20988;
	wire [4-1:0] node20989;
	wire [4-1:0] node20993;
	wire [4-1:0] node20994;
	wire [4-1:0] node20998;
	wire [4-1:0] node20999;
	wire [4-1:0] node21001;
	wire [4-1:0] node21002;
	wire [4-1:0] node21003;
	wire [4-1:0] node21005;
	wire [4-1:0] node21010;
	wire [4-1:0] node21011;
	wire [4-1:0] node21012;
	wire [4-1:0] node21014;
	wire [4-1:0] node21015;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21024;
	wire [4-1:0] node21025;
	wire [4-1:0] node21026;
	wire [4-1:0] node21028;
	wire [4-1:0] node21031;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21037;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21041;
	wire [4-1:0] node21044;
	wire [4-1:0] node21045;
	wire [4-1:0] node21049;
	wire [4-1:0] node21050;
	wire [4-1:0] node21052;
	wire [4-1:0] node21053;
	wire [4-1:0] node21057;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21062;
	wire [4-1:0] node21065;
	wire [4-1:0] node21068;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21076;
	wire [4-1:0] node21078;
	wire [4-1:0] node21081;
	wire [4-1:0] node21082;
	wire [4-1:0] node21084;
	wire [4-1:0] node21087;
	wire [4-1:0] node21088;
	wire [4-1:0] node21092;
	wire [4-1:0] node21093;
	wire [4-1:0] node21094;
	wire [4-1:0] node21098;
	wire [4-1:0] node21099;
	wire [4-1:0] node21101;
	wire [4-1:0] node21105;
	wire [4-1:0] node21106;
	wire [4-1:0] node21107;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21113;
	wire [4-1:0] node21114;
	wire [4-1:0] node21116;
	wire [4-1:0] node21120;
	wire [4-1:0] node21121;
	wire [4-1:0] node21122;
	wire [4-1:0] node21124;
	wire [4-1:0] node21125;
	wire [4-1:0] node21128;
	wire [4-1:0] node21131;
	wire [4-1:0] node21133;
	wire [4-1:0] node21134;
	wire [4-1:0] node21138;
	wire [4-1:0] node21139;
	wire [4-1:0] node21140;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21150;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21157;
	wire [4-1:0] node21158;
	wire [4-1:0] node21160;
	wire [4-1:0] node21163;
	wire [4-1:0] node21165;
	wire [4-1:0] node21168;
	wire [4-1:0] node21169;
	wire [4-1:0] node21171;
	wire [4-1:0] node21174;
	wire [4-1:0] node21176;
	wire [4-1:0] node21179;
	wire [4-1:0] node21180;
	wire [4-1:0] node21181;
	wire [4-1:0] node21184;
	wire [4-1:0] node21185;
	wire [4-1:0] node21189;
	wire [4-1:0] node21191;
	wire [4-1:0] node21193;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21198;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21210;
	wire [4-1:0] node21213;
	wire [4-1:0] node21214;
	wire [4-1:0] node21215;
	wire [4-1:0] node21216;
	wire [4-1:0] node21217;
	wire [4-1:0] node21220;
	wire [4-1:0] node21223;
	wire [4-1:0] node21225;
	wire [4-1:0] node21228;
	wire [4-1:0] node21229;
	wire [4-1:0] node21232;
	wire [4-1:0] node21234;
	wire [4-1:0] node21237;
	wire [4-1:0] node21238;
	wire [4-1:0] node21239;
	wire [4-1:0] node21243;
	wire [4-1:0] node21244;
	wire [4-1:0] node21246;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21253;
	wire [4-1:0] node21254;
	wire [4-1:0] node21255;
	wire [4-1:0] node21258;
	wire [4-1:0] node21262;
	wire [4-1:0] node21264;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21271;
	wire [4-1:0] node21272;
	wire [4-1:0] node21273;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21281;
	wire [4-1:0] node21284;
	wire [4-1:0] node21285;
	wire [4-1:0] node21286;
	wire [4-1:0] node21288;
	wire [4-1:0] node21291;
	wire [4-1:0] node21292;
	wire [4-1:0] node21296;
	wire [4-1:0] node21297;
	wire [4-1:0] node21298;
	wire [4-1:0] node21299;
	wire [4-1:0] node21302;
	wire [4-1:0] node21305;
	wire [4-1:0] node21308;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21313;
	wire [4-1:0] node21314;
	wire [4-1:0] node21315;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21322;
	wire [4-1:0] node21325;
	wire [4-1:0] node21326;
	wire [4-1:0] node21330;
	wire [4-1:0] node21331;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21337;
	wire [4-1:0] node21338;
	wire [4-1:0] node21340;
	wire [4-1:0] node21343;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21353;
	wire [4-1:0] node21354;
	wire [4-1:0] node21356;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21364;
	wire [4-1:0] node21365;
	wire [4-1:0] node21366;
	wire [4-1:0] node21368;
	wire [4-1:0] node21371;
	wire [4-1:0] node21372;
	wire [4-1:0] node21375;
	wire [4-1:0] node21378;
	wire [4-1:0] node21379;
	wire [4-1:0] node21382;
	wire [4-1:0] node21383;
	wire [4-1:0] node21387;
	wire [4-1:0] node21388;
	wire [4-1:0] node21389;
	wire [4-1:0] node21390;
	wire [4-1:0] node21393;
	wire [4-1:0] node21395;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21401;
	wire [4-1:0] node21405;
	wire [4-1:0] node21406;
	wire [4-1:0] node21408;
	wire [4-1:0] node21411;
	wire [4-1:0] node21413;
	wire [4-1:0] node21416;
	wire [4-1:0] node21417;
	wire [4-1:0] node21418;
	wire [4-1:0] node21419;
	wire [4-1:0] node21420;
	wire [4-1:0] node21421;
	wire [4-1:0] node21424;
	wire [4-1:0] node21427;
	wire [4-1:0] node21428;
	wire [4-1:0] node21431;
	wire [4-1:0] node21434;
	wire [4-1:0] node21435;
	wire [4-1:0] node21436;
	wire [4-1:0] node21439;
	wire [4-1:0] node21442;
	wire [4-1:0] node21443;
	wire [4-1:0] node21446;
	wire [4-1:0] node21449;
	wire [4-1:0] node21450;
	wire [4-1:0] node21451;
	wire [4-1:0] node21453;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21459;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21468;
	wire [4-1:0] node21471;
	wire [4-1:0] node21473;
	wire [4-1:0] node21476;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21480;
	wire [4-1:0] node21481;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21487;
	wire [4-1:0] node21490;
	wire [4-1:0] node21493;
	wire [4-1:0] node21494;
	wire [4-1:0] node21498;
	wire [4-1:0] node21499;
	wire [4-1:0] node21500;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21517;
	wire [4-1:0] node21518;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21521;
	wire [4-1:0] node21525;
	wire [4-1:0] node21526;
	wire [4-1:0] node21528;
	wire [4-1:0] node21531;
	wire [4-1:0] node21534;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21544;
	wire [4-1:0] node21547;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21554;
	wire [4-1:0] node21556;
	wire [4-1:0] node21557;
	wire [4-1:0] node21561;
	wire [4-1:0] node21562;
	wire [4-1:0] node21563;
	wire [4-1:0] node21566;
	wire [4-1:0] node21569;
	wire [4-1:0] node21570;
	wire [4-1:0] node21571;
	wire [4-1:0] node21575;
	wire [4-1:0] node21578;
	wire [4-1:0] node21579;
	wire [4-1:0] node21580;
	wire [4-1:0] node21581;
	wire [4-1:0] node21584;
	wire [4-1:0] node21586;
	wire [4-1:0] node21589;
	wire [4-1:0] node21590;
	wire [4-1:0] node21593;
	wire [4-1:0] node21594;
	wire [4-1:0] node21596;
	wire [4-1:0] node21600;
	wire [4-1:0] node21601;
	wire [4-1:0] node21602;
	wire [4-1:0] node21604;
	wire [4-1:0] node21605;
	wire [4-1:0] node21608;
	wire [4-1:0] node21611;
	wire [4-1:0] node21613;
	wire [4-1:0] node21615;
	wire [4-1:0] node21618;
	wire [4-1:0] node21619;
	wire [4-1:0] node21623;
	wire [4-1:0] node21624;
	wire [4-1:0] node21625;
	wire [4-1:0] node21626;
	wire [4-1:0] node21628;
	wire [4-1:0] node21631;
	wire [4-1:0] node21632;
	wire [4-1:0] node21633;
	wire [4-1:0] node21637;
	wire [4-1:0] node21639;
	wire [4-1:0] node21642;
	wire [4-1:0] node21643;
	wire [4-1:0] node21644;
	wire [4-1:0] node21645;
	wire [4-1:0] node21649;
	wire [4-1:0] node21650;
	wire [4-1:0] node21653;
	wire [4-1:0] node21656;
	wire [4-1:0] node21658;
	wire [4-1:0] node21661;
	wire [4-1:0] node21662;
	wire [4-1:0] node21663;
	wire [4-1:0] node21664;
	wire [4-1:0] node21666;
	wire [4-1:0] node21669;
	wire [4-1:0] node21671;
	wire [4-1:0] node21674;
	wire [4-1:0] node21675;
	wire [4-1:0] node21676;
	wire [4-1:0] node21680;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21685;
	wire [4-1:0] node21688;
	wire [4-1:0] node21691;
	wire [4-1:0] node21692;
	wire [4-1:0] node21693;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21700;
	wire [4-1:0] node21703;
	wire [4-1:0] node21704;
	wire [4-1:0] node21705;
	wire [4-1:0] node21706;
	wire [4-1:0] node21709;
	wire [4-1:0] node21712;
	wire [4-1:0] node21713;
	wire [4-1:0] node21716;
	wire [4-1:0] node21719;
	wire [4-1:0] node21720;
	wire [4-1:0] node21721;
	wire [4-1:0] node21726;
	wire [4-1:0] node21727;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21731;
	wire [4-1:0] node21734;
	wire [4-1:0] node21737;
	wire [4-1:0] node21738;
	wire [4-1:0] node21741;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21746;
	wire [4-1:0] node21748;
	wire [4-1:0] node21751;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21756;
	wire [4-1:0] node21759;
	wire [4-1:0] node21762;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21769;
	wire [4-1:0] node21770;
	wire [4-1:0] node21771;
	wire [4-1:0] node21772;
	wire [4-1:0] node21774;
	wire [4-1:0] node21778;
	wire [4-1:0] node21779;
	wire [4-1:0] node21781;
	wire [4-1:0] node21785;
	wire [4-1:0] node21786;
	wire [4-1:0] node21788;
	wire [4-1:0] node21789;
	wire [4-1:0] node21793;
	wire [4-1:0] node21794;
	wire [4-1:0] node21795;
	wire [4-1:0] node21799;
	wire [4-1:0] node21800;
	wire [4-1:0] node21804;
	wire [4-1:0] node21805;
	wire [4-1:0] node21806;
	wire [4-1:0] node21807;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21812;
	wire [4-1:0] node21816;
	wire [4-1:0] node21818;
	wire [4-1:0] node21819;
	wire [4-1:0] node21822;
	wire [4-1:0] node21825;
	wire [4-1:0] node21826;
	wire [4-1:0] node21828;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21835;
	wire [4-1:0] node21836;
	wire [4-1:0] node21840;
	wire [4-1:0] node21841;
	wire [4-1:0] node21842;
	wire [4-1:0] node21843;
	wire [4-1:0] node21845;
	wire [4-1:0] node21848;
	wire [4-1:0] node21851;
	wire [4-1:0] node21852;
	wire [4-1:0] node21853;
	wire [4-1:0] node21856;
	wire [4-1:0] node21859;
	wire [4-1:0] node21862;
	wire [4-1:0] node21864;
	wire [4-1:0] node21867;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21870;
	wire [4-1:0] node21871;
	wire [4-1:0] node21872;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21877;
	wire [4-1:0] node21880;
	wire [4-1:0] node21881;
	wire [4-1:0] node21885;
	wire [4-1:0] node21886;
	wire [4-1:0] node21887;
	wire [4-1:0] node21888;
	wire [4-1:0] node21892;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21898;
	wire [4-1:0] node21902;
	wire [4-1:0] node21903;
	wire [4-1:0] node21904;
	wire [4-1:0] node21905;
	wire [4-1:0] node21908;
	wire [4-1:0] node21911;
	wire [4-1:0] node21912;
	wire [4-1:0] node21914;
	wire [4-1:0] node21918;
	wire [4-1:0] node21919;
	wire [4-1:0] node21920;
	wire [4-1:0] node21923;
	wire [4-1:0] node21924;
	wire [4-1:0] node21928;
	wire [4-1:0] node21930;
	wire [4-1:0] node21933;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21940;
	wire [4-1:0] node21943;
	wire [4-1:0] node21944;
	wire [4-1:0] node21948;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21955;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21959;
	wire [4-1:0] node21960;
	wire [4-1:0] node21964;
	wire [4-1:0] node21965;
	wire [4-1:0] node21968;
	wire [4-1:0] node21971;
	wire [4-1:0] node21973;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21978;
	wire [4-1:0] node21979;
	wire [4-1:0] node21980;
	wire [4-1:0] node21981;
	wire [4-1:0] node21982;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21991;
	wire [4-1:0] node21993;
	wire [4-1:0] node21996;
	wire [4-1:0] node21998;
	wire [4-1:0] node22000;
	wire [4-1:0] node22001;
	wire [4-1:0] node22005;
	wire [4-1:0] node22006;
	wire [4-1:0] node22007;
	wire [4-1:0] node22009;
	wire [4-1:0] node22010;
	wire [4-1:0] node22013;
	wire [4-1:0] node22016;
	wire [4-1:0] node22017;
	wire [4-1:0] node22018;
	wire [4-1:0] node22023;
	wire [4-1:0] node22024;
	wire [4-1:0] node22025;
	wire [4-1:0] node22026;
	wire [4-1:0] node22029;
	wire [4-1:0] node22032;
	wire [4-1:0] node22035;
	wire [4-1:0] node22036;
	wire [4-1:0] node22040;
	wire [4-1:0] node22041;
	wire [4-1:0] node22042;
	wire [4-1:0] node22043;
	wire [4-1:0] node22044;
	wire [4-1:0] node22047;
	wire [4-1:0] node22049;
	wire [4-1:0] node22052;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22058;
	wire [4-1:0] node22061;
	wire [4-1:0] node22062;
	wire [4-1:0] node22064;
	wire [4-1:0] node22067;
	wire [4-1:0] node22069;
	wire [4-1:0] node22071;
	wire [4-1:0] node22074;
	wire [4-1:0] node22075;
	wire [4-1:0] node22076;
	wire [4-1:0] node22078;
	wire [4-1:0] node22079;
	wire [4-1:0] node22083;
	wire [4-1:0] node22084;
	wire [4-1:0] node22087;
	wire [4-1:0] node22089;
	wire [4-1:0] node22093;
	wire [4-1:0] node22094;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22097;
	wire [4-1:0] node22098;
	wire [4-1:0] node22101;
	wire [4-1:0] node22103;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22109;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22117;
	wire [4-1:0] node22118;
	wire [4-1:0] node22120;
	wire [4-1:0] node22121;
	wire [4-1:0] node22124;
	wire [4-1:0] node22127;
	wire [4-1:0] node22128;
	wire [4-1:0] node22131;
	wire [4-1:0] node22133;
	wire [4-1:0] node22136;
	wire [4-1:0] node22137;
	wire [4-1:0] node22138;
	wire [4-1:0] node22140;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22146;
	wire [4-1:0] node22149;
	wire [4-1:0] node22152;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22155;
	wire [4-1:0] node22159;
	wire [4-1:0] node22161;
	wire [4-1:0] node22165;
	wire [4-1:0] node22166;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22169;
	wire [4-1:0] node22172;
	wire [4-1:0] node22173;
	wire [4-1:0] node22177;
	wire [4-1:0] node22178;
	wire [4-1:0] node22180;
	wire [4-1:0] node22181;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22189;
	wire [4-1:0] node22191;
	wire [4-1:0] node22194;
	wire [4-1:0] node22196;
	wire [4-1:0] node22197;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22203;
	wire [4-1:0] node22204;
	wire [4-1:0] node22205;
	wire [4-1:0] node22206;
	wire [4-1:0] node22211;
	wire [4-1:0] node22213;
	wire [4-1:0] node22215;
	wire [4-1:0] node22220;
	wire [4-1:0] node22222;
	wire [4-1:0] node22223;
	wire [4-1:0] node22224;
	wire [4-1:0] node22226;
	wire [4-1:0] node22227;
	wire [4-1:0] node22228;
	wire [4-1:0] node22230;
	wire [4-1:0] node22232;
	wire [4-1:0] node22233;
	wire [4-1:0] node22235;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22241;
	wire [4-1:0] node22242;
	wire [4-1:0] node22245;
	wire [4-1:0] node22246;
	wire [4-1:0] node22250;
	wire [4-1:0] node22251;
	wire [4-1:0] node22253;
	wire [4-1:0] node22256;
	wire [4-1:0] node22258;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22263;
	wire [4-1:0] node22266;
	wire [4-1:0] node22268;
	wire [4-1:0] node22271;
	wire [4-1:0] node22272;
	wire [4-1:0] node22274;
	wire [4-1:0] node22276;
	wire [4-1:0] node22279;
	wire [4-1:0] node22281;
	wire [4-1:0] node22284;
	wire [4-1:0] node22286;
	wire [4-1:0] node22287;
	wire [4-1:0] node22289;
	wire [4-1:0] node22290;
	wire [4-1:0] node22291;
	wire [4-1:0] node22293;
	wire [4-1:0] node22299;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22303;
	wire [4-1:0] node22304;
	wire [4-1:0] node22305;
	wire [4-1:0] node22306;
	wire [4-1:0] node22310;
	wire [4-1:0] node22312;
	wire [4-1:0] node22315;
	wire [4-1:0] node22317;
	wire [4-1:0] node22320;
	wire [4-1:0] node22321;
	wire [4-1:0] node22323;
	wire [4-1:0] node22325;
	wire [4-1:0] node22328;
	wire [4-1:0] node22329;
	wire [4-1:0] node22330;
	wire [4-1:0] node22332;
	wire [4-1:0] node22335;
	wire [4-1:0] node22337;
	wire [4-1:0] node22341;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22344;
	wire [4-1:0] node22346;
	wire [4-1:0] node22348;
	wire [4-1:0] node22351;
	wire [4-1:0] node22352;
	wire [4-1:0] node22356;
	wire [4-1:0] node22357;
	wire [4-1:0] node22359;
	wire [4-1:0] node22362;
	wire [4-1:0] node22363;
	wire [4-1:0] node22367;
	wire [4-1:0] node22368;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22373;
	wire [4-1:0] node22374;
	wire [4-1:0] node22378;
	wire [4-1:0] node22380;
	wire [4-1:0] node22383;
	wire [4-1:0] node22384;
	wire [4-1:0] node22386;
	wire [4-1:0] node22389;
	wire [4-1:0] node22390;
	wire [4-1:0] node22391;
	wire [4-1:0] node22395;
	wire [4-1:0] node22397;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22402;
	wire [4-1:0] node22403;
	wire [4-1:0] node22405;
	wire [4-1:0] node22406;
	wire [4-1:0] node22409;
	wire [4-1:0] node22410;
	wire [4-1:0] node22414;
	wire [4-1:0] node22415;
	wire [4-1:0] node22418;
	wire [4-1:0] node22419;
	wire [4-1:0] node22422;
	wire [4-1:0] node22425;
	wire [4-1:0] node22426;
	wire [4-1:0] node22428;
	wire [4-1:0] node22431;
	wire [4-1:0] node22432;
	wire [4-1:0] node22433;
	wire [4-1:0] node22436;
	wire [4-1:0] node22439;
	wire [4-1:0] node22440;
	wire [4-1:0] node22444;
	wire [4-1:0] node22445;
	wire [4-1:0] node22446;
	wire [4-1:0] node22447;
	wire [4-1:0] node22448;
	wire [4-1:0] node22449;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22458;
	wire [4-1:0] node22460;
	wire [4-1:0] node22463;
	wire [4-1:0] node22464;
	wire [4-1:0] node22465;
	wire [4-1:0] node22468;
	wire [4-1:0] node22470;
	wire [4-1:0] node22474;
	wire [4-1:0] node22475;
	wire [4-1:0] node22476;
	wire [4-1:0] node22478;
	wire [4-1:0] node22481;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22487;
	wire [4-1:0] node22488;
	wire [4-1:0] node22491;
	wire [4-1:0] node22494;
	wire [4-1:0] node22495;
	wire [4-1:0] node22497;
	wire [4-1:0] node22498;
	wire [4-1:0] node22501;
	wire [4-1:0] node22505;
	wire [4-1:0] node22506;
	wire [4-1:0] node22507;
	wire [4-1:0] node22508;
	wire [4-1:0] node22509;
	wire [4-1:0] node22510;
	wire [4-1:0] node22511;
	wire [4-1:0] node22513;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22522;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22527;
	wire [4-1:0] node22529;
	wire [4-1:0] node22532;
	wire [4-1:0] node22534;
	wire [4-1:0] node22537;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22541;
	wire [4-1:0] node22544;
	wire [4-1:0] node22547;
	wire [4-1:0] node22548;
	wire [4-1:0] node22549;
	wire [4-1:0] node22551;
	wire [4-1:0] node22555;
	wire [4-1:0] node22556;
	wire [4-1:0] node22557;
	wire [4-1:0] node22561;
	wire [4-1:0] node22563;
	wire [4-1:0] node22566;
	wire [4-1:0] node22567;
	wire [4-1:0] node22568;
	wire [4-1:0] node22569;
	wire [4-1:0] node22570;
	wire [4-1:0] node22571;
	wire [4-1:0] node22574;
	wire [4-1:0] node22578;
	wire [4-1:0] node22580;
	wire [4-1:0] node22582;
	wire [4-1:0] node22585;
	wire [4-1:0] node22587;
	wire [4-1:0] node22589;
	wire [4-1:0] node22592;
	wire [4-1:0] node22593;
	wire [4-1:0] node22594;
	wire [4-1:0] node22596;
	wire [4-1:0] node22599;
	wire [4-1:0] node22601;
	wire [4-1:0] node22604;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22608;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22616;
	wire [4-1:0] node22618;
	wire [4-1:0] node22619;
	wire [4-1:0] node22622;
	wire [4-1:0] node22625;
	wire [4-1:0] node22626;
	wire [4-1:0] node22629;
	wire [4-1:0] node22632;
	wire [4-1:0] node22633;
	wire [4-1:0] node22634;
	wire [4-1:0] node22635;
	wire [4-1:0] node22638;
	wire [4-1:0] node22641;
	wire [4-1:0] node22642;
	wire [4-1:0] node22643;
	wire [4-1:0] node22646;
	wire [4-1:0] node22649;
	wire [4-1:0] node22650;
	wire [4-1:0] node22654;
	wire [4-1:0] node22656;
	wire [4-1:0] node22659;
	wire [4-1:0] node22660;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22663;
	wire [4-1:0] node22666;
	wire [4-1:0] node22670;
	wire [4-1:0] node22671;
	wire [4-1:0] node22675;
	wire [4-1:0] node22677;
	wire [4-1:0] node22678;
	wire [4-1:0] node22679;
	wire [4-1:0] node22684;
	wire [4-1:0] node22686;
	wire [4-1:0] node22688;
	wire [4-1:0] node22689;
	wire [4-1:0] node22690;
	wire [4-1:0] node22692;
	wire [4-1:0] node22694;
	wire [4-1:0] node22695;
	wire [4-1:0] node22696;
	wire [4-1:0] node22697;
	wire [4-1:0] node22701;
	wire [4-1:0] node22705;
	wire [4-1:0] node22706;
	wire [4-1:0] node22707;
	wire [4-1:0] node22708;
	wire [4-1:0] node22709;
	wire [4-1:0] node22712;
	wire [4-1:0] node22715;
	wire [4-1:0] node22716;
	wire [4-1:0] node22720;
	wire [4-1:0] node22721;
	wire [4-1:0] node22722;
	wire [4-1:0] node22726;
	wire [4-1:0] node22728;
	wire [4-1:0] node22731;
	wire [4-1:0] node22732;
	wire [4-1:0] node22733;
	wire [4-1:0] node22735;
	wire [4-1:0] node22740;
	wire [4-1:0] node22741;
	wire [4-1:0] node22743;
	wire [4-1:0] node22744;
	wire [4-1:0] node22746;
	wire [4-1:0] node22747;

	assign outp = (inp[8]) ? node11686 : node1;
		assign node1 = (inp[9]) ? node6089 : node2;
			assign node2 = (inp[6]) ? node1372 : node3;
				assign node3 = (inp[15]) ? node755 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[2]) ? node481 : node6;
							assign node6 = (inp[1]) ? node230 : node7;
								assign node7 = (inp[14]) ? node87 : node8;
									assign node8 = (inp[13]) ? node50 : node9;
										assign node9 = (inp[10]) ? node37 : node10;
											assign node10 = (inp[12]) ? node24 : node11;
												assign node11 = (inp[3]) ? node19 : node12;
													assign node12 = (inp[4]) ? 4'b0000 : node13;
														assign node13 = (inp[7]) ? node15 : 4'b0000;
															assign node15 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node19 = (inp[4]) ? 4'b0100 : node20;
														assign node20 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node24 = (inp[3]) ? node32 : node25;
													assign node25 = (inp[5]) ? node27 : 4'b1000;
														assign node27 = (inp[4]) ? node29 : 4'b1100;
															assign node29 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node32 = (inp[7]) ? 4'b1000 : node33;
														assign node33 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node37 = (inp[3]) ? node45 : node38;
												assign node38 = (inp[7]) ? node40 : 4'b0000;
													assign node40 = (inp[4]) ? 4'b0000 : node41;
														assign node41 = (inp[5]) ? 4'b0100 : 4'b1111;
												assign node45 = (inp[7]) ? node47 : 4'b0100;
													assign node47 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node50 = (inp[3]) ? node70 : node51;
											assign node51 = (inp[4]) ? node65 : node52;
												assign node52 = (inp[7]) ? node58 : node53;
													assign node53 = (inp[12]) ? node55 : 4'b1000;
														assign node55 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node58 = (inp[5]) ? node60 : 4'b1111;
														assign node60 = (inp[12]) ? node62 : 4'b1100;
															assign node62 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node65 = (inp[12]) ? node67 : 4'b1000;
													assign node67 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node70 = (inp[7]) ? node76 : node71;
												assign node71 = (inp[10]) ? 4'b1100 : node72;
													assign node72 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node76 = (inp[4]) ? node82 : node77;
													assign node77 = (inp[10]) ? 4'b1000 : node78;
														assign node78 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node82 = (inp[12]) ? node84 : 4'b1100;
														assign node84 = (inp[10]) ? 4'b1100 : 4'b0100;
									assign node87 = (inp[11]) ? node161 : node88;
										assign node88 = (inp[13]) ? node128 : node89;
											assign node89 = (inp[3]) ? node113 : node90;
												assign node90 = (inp[5]) ? node104 : node91;
													assign node91 = (inp[7]) ? 4'b1111 : node92;
														assign node92 = (inp[4]) ? node98 : node93;
															assign node93 = (inp[10]) ? node95 : 4'b1111;
																assign node95 = (inp[12]) ? 4'b1111 : 4'b0001;
															assign node98 = (inp[10]) ? node100 : 4'b1001;
																assign node100 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node104 = (inp[4]) ? node106 : 4'b1101;
														assign node106 = (inp[7]) ? node108 : 4'b1001;
															assign node108 = (inp[12]) ? 4'b1101 : node109;
																assign node109 = (inp[10]) ? 4'b0001 : 4'b1101;
												assign node113 = (inp[12]) ? node123 : node114;
													assign node114 = (inp[10]) ? node118 : node115;
														assign node115 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node118 = (inp[7]) ? node120 : 4'b0101;
															assign node120 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node123 = (inp[7]) ? 4'b1001 : node124;
														assign node124 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node128 = (inp[12]) ? node150 : node129;
												assign node129 = (inp[10]) ? node141 : node130;
													assign node130 = (inp[7]) ? node134 : node131;
														assign node131 = (inp[3]) ? 4'b0101 : 4'b0001;
														assign node134 = (inp[5]) ? node136 : 4'b1111;
															assign node136 = (inp[3]) ? node138 : 4'b0101;
																assign node138 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node141 = (inp[3]) ? node145 : node142;
														assign node142 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node145 = (inp[4]) ? 4'b1101 : node146;
															assign node146 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node150 = (inp[3]) ? node156 : node151;
													assign node151 = (inp[4]) ? 4'b0001 : node152;
														assign node152 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node156 = (inp[7]) ? node158 : 4'b0101;
														assign node158 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node161 = (inp[13]) ? node197 : node162;
											assign node162 = (inp[10]) ? node184 : node163;
												assign node163 = (inp[12]) ? node175 : node164;
													assign node164 = (inp[7]) ? node168 : node165;
														assign node165 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node168 = (inp[5]) ? node172 : node169;
															assign node169 = (inp[3]) ? 4'b0100 : 4'b1111;
															assign node172 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node175 = (inp[4]) ? node177 : 4'b1000;
														assign node177 = (inp[7]) ? node181 : node178;
															assign node178 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node181 = (inp[5]) ? 4'b1100 : 4'b1111;
												assign node184 = (inp[3]) ? node192 : node185;
													assign node185 = (inp[7]) ? node187 : 4'b0000;
														assign node187 = (inp[4]) ? 4'b0000 : node188;
															assign node188 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node192 = (inp[7]) ? node194 : 4'b0100;
														assign node194 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node197 = (inp[3]) ? node213 : node198;
												assign node198 = (inp[4]) ? node208 : node199;
													assign node199 = (inp[7]) ? node205 : node200;
														assign node200 = (inp[12]) ? node202 : 4'b1000;
															assign node202 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node205 = (inp[5]) ? 4'b1100 : 4'b1111;
													assign node208 = (inp[10]) ? 4'b1000 : node209;
														assign node209 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node213 = (inp[12]) ? node219 : node214;
													assign node214 = (inp[7]) ? node216 : 4'b1100;
														assign node216 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node219 = (inp[10]) ? node225 : node220;
														assign node220 = (inp[7]) ? node222 : 4'b0100;
															assign node222 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node225 = (inp[4]) ? 4'b1100 : node226;
															assign node226 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node230 = (inp[14]) ? node332 : node231;
									assign node231 = (inp[13]) ? node285 : node232;
										assign node232 = (inp[12]) ? node246 : node233;
											assign node233 = (inp[3]) ? node241 : node234;
												assign node234 = (inp[4]) ? 4'b0001 : node235;
													assign node235 = (inp[7]) ? node237 : 4'b0001;
														assign node237 = (inp[5]) ? 4'b0101 : 4'b1111;
												assign node241 = (inp[4]) ? 4'b0101 : node242;
													assign node242 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node246 = (inp[10]) ? node264 : node247;
												assign node247 = (inp[3]) ? node259 : node248;
													assign node248 = (inp[5]) ? node254 : node249;
														assign node249 = (inp[4]) ? node251 : 4'b1111;
															assign node251 = (inp[7]) ? 4'b1111 : 4'b1001;
														assign node254 = (inp[7]) ? 4'b1101 : node255;
															assign node255 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node259 = (inp[4]) ? node261 : 4'b1001;
														assign node261 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node264 = (inp[5]) ? node274 : node265;
													assign node265 = (inp[7]) ? node267 : 4'b0001;
														assign node267 = (inp[3]) ? node271 : node268;
															assign node268 = (inp[4]) ? 4'b0001 : 4'b1111;
															assign node271 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node274 = (inp[11]) ? node280 : node275;
														assign node275 = (inp[4]) ? node277 : 4'b0101;
															assign node277 = (inp[3]) ? 4'b0101 : 4'b0001;
														assign node280 = (inp[4]) ? 4'b0001 : node281;
															assign node281 = (inp[3]) ? 4'b0001 : 4'b0101;
										assign node285 = (inp[12]) ? node299 : node286;
											assign node286 = (inp[3]) ? node294 : node287;
												assign node287 = (inp[4]) ? 4'b1001 : node288;
													assign node288 = (inp[7]) ? node290 : 4'b1001;
														assign node290 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node294 = (inp[4]) ? 4'b1101 : node295;
													assign node295 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node299 = (inp[10]) ? node313 : node300;
												assign node300 = (inp[3]) ? node308 : node301;
													assign node301 = (inp[4]) ? 4'b0001 : node302;
														assign node302 = (inp[7]) ? node304 : 4'b0001;
															assign node304 = (inp[5]) ? 4'b0101 : 4'b1111;
													assign node308 = (inp[4]) ? 4'b0101 : node309;
														assign node309 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node313 = (inp[5]) ? node325 : node314;
													assign node314 = (inp[3]) ? node320 : node315;
														assign node315 = (inp[7]) ? node317 : 4'b1001;
															assign node317 = (inp[4]) ? 4'b1001 : 4'b1111;
														assign node320 = (inp[7]) ? node322 : 4'b1101;
															assign node322 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node325 = (inp[7]) ? node327 : 4'b1101;
														assign node327 = (inp[3]) ? node329 : 4'b1101;
															assign node329 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node332 = (inp[11]) ? node414 : node333;
										assign node333 = (inp[13]) ? node375 : node334;
											assign node334 = (inp[12]) ? node348 : node335;
												assign node335 = (inp[3]) ? node343 : node336;
													assign node336 = (inp[4]) ? 4'b0000 : node337;
														assign node337 = (inp[7]) ? node339 : 4'b0000;
															assign node339 = (inp[5]) ? 4'b0100 : 4'b1111;
													assign node343 = (inp[7]) ? node345 : 4'b0100;
														assign node345 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node348 = (inp[10]) ? node362 : node349;
													assign node349 = (inp[4]) ? node351 : 4'b1000;
														assign node351 = (inp[5]) ? node355 : node352;
															assign node352 = (inp[7]) ? 4'b1111 : 4'b1100;
															assign node355 = (inp[7]) ? node359 : node356;
																assign node356 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node359 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node362 = (inp[3]) ? node368 : node363;
														assign node363 = (inp[7]) ? node365 : 4'b0000;
															assign node365 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node368 = (inp[5]) ? 4'b0100 : node369;
															assign node369 = (inp[4]) ? 4'b0100 : node370;
																assign node370 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node375 = (inp[10]) ? node401 : node376;
												assign node376 = (inp[12]) ? node390 : node377;
													assign node377 = (inp[3]) ? node385 : node378;
														assign node378 = (inp[4]) ? 4'b1000 : node379;
															assign node379 = (inp[5]) ? node381 : 4'b1111;
																assign node381 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node385 = (inp[7]) ? node387 : 4'b1100;
															assign node387 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node390 = (inp[3]) ? node396 : node391;
														assign node391 = (inp[4]) ? 4'b0000 : node392;
															assign node392 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node396 = (inp[4]) ? 4'b0100 : node397;
															assign node397 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node401 = (inp[4]) ? node411 : node402;
													assign node402 = (inp[3]) ? node408 : node403;
														assign node403 = (inp[7]) ? node405 : 4'b1000;
															assign node405 = (inp[5]) ? 4'b1100 : 4'b1111;
														assign node408 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node411 = (inp[3]) ? 4'b1100 : 4'b1000;
										assign node414 = (inp[3]) ? node452 : node415;
											assign node415 = (inp[4]) ? node439 : node416;
												assign node416 = (inp[7]) ? node430 : node417;
													assign node417 = (inp[13]) ? node425 : node418;
														assign node418 = (inp[10]) ? 4'b0001 : node419;
															assign node419 = (inp[12]) ? node421 : 4'b0001;
																assign node421 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node425 = (inp[12]) ? node427 : 4'b1001;
															assign node427 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node430 = (inp[5]) ? node432 : 4'b1111;
														assign node432 = (inp[13]) ? node436 : node433;
															assign node433 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node436 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node439 = (inp[13]) ? node447 : node440;
													assign node440 = (inp[10]) ? 4'b0001 : node441;
														assign node441 = (inp[12]) ? node443 : 4'b0001;
															assign node443 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node447 = (inp[12]) ? node449 : 4'b1001;
														assign node449 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node452 = (inp[13]) ? node466 : node453;
												assign node453 = (inp[12]) ? node459 : node454;
													assign node454 = (inp[4]) ? 4'b0101 : node455;
														assign node455 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node459 = (inp[10]) ? 4'b0101 : node460;
														assign node460 = (inp[4]) ? node462 : 4'b1001;
															assign node462 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node466 = (inp[10]) ? node476 : node467;
													assign node467 = (inp[12]) ? node471 : node468;
														assign node468 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node471 = (inp[4]) ? 4'b0101 : node472;
															assign node472 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node476 = (inp[4]) ? 4'b1101 : node477;
														assign node477 = (inp[7]) ? 4'b1001 : 4'b1101;
							assign node481 = (inp[5]) ? node483 : 4'b1111;
								assign node483 = (inp[3]) ? node597 : node484;
									assign node484 = (inp[4]) ? node526 : node485;
										assign node485 = (inp[7]) ? 4'b1111 : node486;
											assign node486 = (inp[13]) ? node508 : node487;
												assign node487 = (inp[12]) ? node499 : node488;
													assign node488 = (inp[1]) ? node494 : node489;
														assign node489 = (inp[11]) ? 4'b0000 : node490;
															assign node490 = (inp[14]) ? 4'b1111 : 4'b0000;
														assign node494 = (inp[10]) ? 4'b0001 : node495;
															assign node495 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node499 = (inp[10]) ? node501 : 4'b1111;
														assign node501 = (inp[14]) ? node505 : node502;
															assign node502 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node505 = (inp[11]) ? 4'b0000 : 4'b1111;
												assign node508 = (inp[1]) ? node514 : node509;
													assign node509 = (inp[10]) ? 4'b1000 : node510;
														assign node510 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node514 = (inp[12]) ? node520 : node515;
														assign node515 = (inp[11]) ? 4'b1001 : node516;
															assign node516 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node520 = (inp[10]) ? node522 : 4'b0001;
															assign node522 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node526 = (inp[1]) ? node564 : node527;
											assign node527 = (inp[14]) ? node541 : node528;
												assign node528 = (inp[13]) ? node536 : node529;
													assign node529 = (inp[10]) ? 4'b0000 : node530;
														assign node530 = (inp[12]) ? node532 : 4'b0000;
															assign node532 = (inp[7]) ? 4'b1111 : 4'b1000;
													assign node536 = (inp[10]) ? 4'b1000 : node537;
														assign node537 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node541 = (inp[11]) ? node551 : node542;
													assign node542 = (inp[13]) ? 4'b0001 : node543;
														assign node543 = (inp[7]) ? 4'b1111 : node544;
															assign node544 = (inp[10]) ? node546 : 4'b1001;
																assign node546 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node551 = (inp[13]) ? node559 : node552;
														assign node552 = (inp[10]) ? 4'b0000 : node553;
															assign node553 = (inp[7]) ? 4'b1111 : node554;
																assign node554 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node559 = (inp[12]) ? node561 : 4'b1000;
															assign node561 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node564 = (inp[14]) ? node578 : node565;
												assign node565 = (inp[13]) ? node573 : node566;
													assign node566 = (inp[10]) ? 4'b0001 : node567;
														assign node567 = (inp[12]) ? node569 : 4'b0001;
															assign node569 = (inp[11]) ? 4'b1111 : 4'b1001;
													assign node573 = (inp[10]) ? 4'b1001 : node574;
														assign node574 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node578 = (inp[11]) ? node590 : node579;
													assign node579 = (inp[13]) ? node587 : node580;
														assign node580 = (inp[10]) ? 4'b0000 : node581;
															assign node581 = (inp[12]) ? node583 : 4'b0000;
																assign node583 = (inp[7]) ? 4'b1111 : 4'b1000;
														assign node587 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node590 = (inp[13]) ? 4'b1001 : node591;
														assign node591 = (inp[12]) ? node593 : 4'b0001;
															assign node593 = (inp[10]) ? 4'b0001 : 4'b1111;
									assign node597 = (inp[1]) ? node683 : node598;
										assign node598 = (inp[4]) ? node646 : node599;
											assign node599 = (inp[7]) ? node621 : node600;
												assign node600 = (inp[13]) ? node610 : node601;
													assign node601 = (inp[10]) ? 4'b0100 : node602;
														assign node602 = (inp[12]) ? 4'b1000 : node603;
															assign node603 = (inp[14]) ? node605 : 4'b0100;
																assign node605 = (inp[11]) ? 4'b0100 : 4'b1001;
													assign node610 = (inp[11]) ? node616 : node611;
														assign node611 = (inp[14]) ? node613 : 4'b1100;
															assign node613 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node616 = (inp[12]) ? node618 : 4'b1100;
															assign node618 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node621 = (inp[11]) ? node637 : node622;
													assign node622 = (inp[14]) ? node630 : node623;
														assign node623 = (inp[13]) ? 4'b1000 : node624;
															assign node624 = (inp[12]) ? node626 : 4'b0000;
																assign node626 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node630 = (inp[13]) ? 4'b0001 : node631;
															assign node631 = (inp[12]) ? 4'b1001 : node632;
																assign node632 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node637 = (inp[13]) ? node643 : node638;
														assign node638 = (inp[14]) ? 4'b0000 : node639;
															assign node639 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node643 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node646 = (inp[11]) ? node670 : node647;
												assign node647 = (inp[14]) ? node659 : node648;
													assign node648 = (inp[13]) ? node654 : node649;
														assign node649 = (inp[10]) ? 4'b0100 : node650;
															assign node650 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node654 = (inp[10]) ? 4'b1100 : node655;
															assign node655 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node659 = (inp[13]) ? node667 : node660;
														assign node660 = (inp[12]) ? node664 : node661;
															assign node661 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node664 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node667 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node670 = (inp[13]) ? node678 : node671;
													assign node671 = (inp[12]) ? node673 : 4'b0100;
														assign node673 = (inp[10]) ? 4'b0100 : node674;
															assign node674 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node678 = (inp[10]) ? 4'b1100 : node679;
														assign node679 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node683 = (inp[13]) ? node719 : node684;
											assign node684 = (inp[12]) ? node702 : node685;
												assign node685 = (inp[7]) ? node691 : node686;
													assign node686 = (inp[14]) ? node688 : 4'b0101;
														assign node688 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node691 = (inp[4]) ? node697 : node692;
														assign node692 = (inp[14]) ? node694 : 4'b0001;
															assign node694 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node697 = (inp[11]) ? 4'b0101 : node698;
															assign node698 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node702 = (inp[10]) ? node710 : node703;
													assign node703 = (inp[7]) ? node707 : node704;
														assign node704 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node707 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node710 = (inp[4]) ? node714 : node711;
														assign node711 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node714 = (inp[11]) ? 4'b0101 : node715;
															assign node715 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node719 = (inp[14]) ? node737 : node720;
												assign node720 = (inp[7]) ? node726 : node721;
													assign node721 = (inp[12]) ? node723 : 4'b1101;
														assign node723 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node726 = (inp[4]) ? node732 : node727;
														assign node727 = (inp[10]) ? 4'b1001 : node728;
															assign node728 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node732 = (inp[12]) ? node734 : 4'b1101;
															assign node734 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node737 = (inp[11]) ? node745 : node738;
													assign node738 = (inp[4]) ? 4'b1100 : node739;
														assign node739 = (inp[7]) ? 4'b1000 : node740;
															assign node740 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node745 = (inp[10]) ? node749 : node746;
														assign node746 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node749 = (inp[4]) ? 4'b1101 : node750;
															assign node750 = (inp[7]) ? 4'b1001 : 4'b1101;
					assign node755 = (inp[0]) ? 4'b1001 : node756;
						assign node756 = (inp[5]) ? node900 : node757;
							assign node757 = (inp[3]) ? node759 : 4'b1011;
								assign node759 = (inp[2]) ? 4'b1011 : node760;
									assign node760 = (inp[4]) ? node816 : node761;
										assign node761 = (inp[7]) ? 4'b1011 : node762;
											assign node762 = (inp[13]) ? node788 : node763;
												assign node763 = (inp[12]) ? node777 : node764;
													assign node764 = (inp[1]) ? node772 : node765;
														assign node765 = (inp[11]) ? 4'b0000 : node766;
															assign node766 = (inp[14]) ? node768 : 4'b0000;
																assign node768 = (inp[10]) ? 4'b0001 : 4'b1011;
														assign node772 = (inp[14]) ? node774 : 4'b0001;
															assign node774 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node777 = (inp[10]) ? node779 : 4'b1011;
														assign node779 = (inp[1]) ? node783 : node780;
															assign node780 = (inp[14]) ? 4'b1011 : 4'b0000;
															assign node783 = (inp[11]) ? 4'b0001 : node784;
																assign node784 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node788 = (inp[10]) ? node802 : node789;
													assign node789 = (inp[12]) ? node795 : node790;
														assign node790 = (inp[1]) ? 4'b1001 : node791;
															assign node791 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node795 = (inp[1]) ? 4'b0001 : node796;
															assign node796 = (inp[14]) ? node798 : 4'b0000;
																assign node798 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node802 = (inp[1]) ? node810 : node803;
														assign node803 = (inp[11]) ? 4'b1000 : node804;
															assign node804 = (inp[14]) ? node806 : 4'b1000;
																assign node806 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node810 = (inp[14]) ? node812 : 4'b1001;
															assign node812 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node816 = (inp[1]) ? node862 : node817;
											assign node817 = (inp[14]) ? node831 : node818;
												assign node818 = (inp[13]) ? node826 : node819;
													assign node819 = (inp[10]) ? 4'b0000 : node820;
														assign node820 = (inp[12]) ? node822 : 4'b0000;
															assign node822 = (inp[7]) ? 4'b1011 : 4'b1000;
													assign node826 = (inp[12]) ? node828 : 4'b1000;
														assign node828 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node831 = (inp[11]) ? node849 : node832;
													assign node832 = (inp[13]) ? node844 : node833;
														assign node833 = (inp[7]) ? node839 : node834;
															assign node834 = (inp[10]) ? node836 : 4'b1001;
																assign node836 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node839 = (inp[10]) ? node841 : 4'b1011;
																assign node841 = (inp[12]) ? 4'b1011 : 4'b0001;
														assign node844 = (inp[10]) ? node846 : 4'b0001;
															assign node846 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node849 = (inp[13]) ? node857 : node850;
														assign node850 = (inp[10]) ? 4'b0000 : node851;
															assign node851 = (inp[7]) ? 4'b1011 : node852;
																assign node852 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node857 = (inp[10]) ? 4'b1000 : node858;
															assign node858 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node862 = (inp[13]) ? node882 : node863;
												assign node863 = (inp[12]) ? node869 : node864;
													assign node864 = (inp[11]) ? 4'b0001 : node865;
														assign node865 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node869 = (inp[10]) ? node877 : node870;
														assign node870 = (inp[7]) ? 4'b1011 : node871;
															assign node871 = (inp[14]) ? node873 : 4'b1001;
																assign node873 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node877 = (inp[14]) ? node879 : 4'b0001;
															assign node879 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node882 = (inp[11]) ? node894 : node883;
													assign node883 = (inp[14]) ? node889 : node884;
														assign node884 = (inp[12]) ? node886 : 4'b1001;
															assign node886 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node889 = (inp[10]) ? 4'b1000 : node890;
															assign node890 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node894 = (inp[12]) ? node896 : 4'b1001;
														assign node896 = (inp[10]) ? 4'b1001 : 4'b0001;
							assign node900 = (inp[2]) ? node1242 : node901;
								assign node901 = (inp[1]) ? node1071 : node902;
									assign node902 = (inp[11]) ? node1012 : node903;
										assign node903 = (inp[14]) ? node961 : node904;
											assign node904 = (inp[13]) ? node932 : node905;
												assign node905 = (inp[10]) ? node921 : node906;
													assign node906 = (inp[12]) ? node914 : node907;
														assign node907 = (inp[4]) ? 4'b0000 : node908;
															assign node908 = (inp[3]) ? 4'b0100 : node909;
																assign node909 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node914 = (inp[3]) ? node916 : 4'b1000;
															assign node916 = (inp[4]) ? node918 : 4'b1100;
																assign node918 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node921 = (inp[3]) ? node927 : node922;
														assign node922 = (inp[4]) ? 4'b0100 : node923;
															assign node923 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node927 = (inp[4]) ? 4'b0000 : node928;
															assign node928 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node932 = (inp[12]) ? node944 : node933;
													assign node933 = (inp[3]) ? node939 : node934;
														assign node934 = (inp[4]) ? 4'b1100 : node935;
															assign node935 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node939 = (inp[7]) ? node941 : 4'b1000;
															assign node941 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node944 = (inp[10]) ? node952 : node945;
														assign node945 = (inp[4]) ? 4'b0100 : node946;
															assign node946 = (inp[7]) ? node948 : 4'b0000;
																assign node948 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node952 = (inp[7]) ? node956 : node953;
															assign node953 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node956 = (inp[3]) ? node958 : 4'b1000;
																assign node958 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node961 = (inp[13]) ? node989 : node962;
												assign node962 = (inp[10]) ? node972 : node963;
													assign node963 = (inp[3]) ? node967 : node964;
														assign node964 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node967 = (inp[4]) ? node969 : 4'b1101;
															assign node969 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node972 = (inp[12]) ? node980 : node973;
														assign node973 = (inp[3]) ? 4'b0001 : node974;
															assign node974 = (inp[4]) ? 4'b0101 : node975;
																assign node975 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node980 = (inp[4]) ? node982 : 4'b1101;
															assign node982 = (inp[7]) ? node986 : node983;
																assign node983 = (inp[3]) ? 4'b1001 : 4'b1101;
																assign node986 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node989 = (inp[10]) ? node1001 : node990;
													assign node990 = (inp[3]) ? node996 : node991;
														assign node991 = (inp[4]) ? 4'b0101 : node992;
															assign node992 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node996 = (inp[4]) ? 4'b0001 : node997;
															assign node997 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node1001 = (inp[12]) ? node1007 : node1002;
														assign node1002 = (inp[3]) ? 4'b1001 : node1003;
															assign node1003 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node1007 = (inp[3]) ? node1009 : 4'b0101;
															assign node1009 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node1012 = (inp[13]) ? node1046 : node1013;
											assign node1013 = (inp[10]) ? node1035 : node1014;
												assign node1014 = (inp[12]) ? node1026 : node1015;
													assign node1015 = (inp[3]) ? node1021 : node1016;
														assign node1016 = (inp[7]) ? node1018 : 4'b0100;
															assign node1018 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1021 = (inp[7]) ? node1023 : 4'b0000;
															assign node1023 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node1026 = (inp[3]) ? node1030 : node1027;
														assign node1027 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1030 = (inp[4]) ? node1032 : 4'b1100;
															assign node1032 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node1035 = (inp[3]) ? node1041 : node1036;
													assign node1036 = (inp[4]) ? 4'b0100 : node1037;
														assign node1037 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1041 = (inp[4]) ? 4'b0000 : node1042;
														assign node1042 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node1046 = (inp[3]) ? node1056 : node1047;
												assign node1047 = (inp[10]) ? node1051 : node1048;
													assign node1048 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1051 = (inp[4]) ? 4'b1100 : node1052;
														assign node1052 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node1056 = (inp[4]) ? node1066 : node1057;
													assign node1057 = (inp[7]) ? node1061 : node1058;
														assign node1058 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node1061 = (inp[10]) ? 4'b1100 : node1062;
															assign node1062 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node1066 = (inp[10]) ? 4'b1000 : node1067;
														assign node1067 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node1071 = (inp[14]) ? node1133 : node1072;
										assign node1072 = (inp[13]) ? node1102 : node1073;
											assign node1073 = (inp[10]) ? node1091 : node1074;
												assign node1074 = (inp[12]) ? node1080 : node1075;
													assign node1075 = (inp[3]) ? 4'b0001 : node1076;
														assign node1076 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1080 = (inp[3]) ? node1086 : node1081;
														assign node1081 = (inp[7]) ? 4'b1001 : node1082;
															assign node1082 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node1086 = (inp[7]) ? 4'b1101 : node1087;
															assign node1087 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node1091 = (inp[3]) ? node1097 : node1092;
													assign node1092 = (inp[4]) ? 4'b0101 : node1093;
														assign node1093 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1097 = (inp[4]) ? 4'b0001 : node1098;
														assign node1098 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node1102 = (inp[3]) ? node1120 : node1103;
												assign node1103 = (inp[10]) ? node1115 : node1104;
													assign node1104 = (inp[12]) ? node1110 : node1105;
														assign node1105 = (inp[7]) ? node1107 : 4'b1101;
															assign node1107 = (inp[11]) ? 4'b1001 : 4'b1101;
														assign node1110 = (inp[4]) ? 4'b0101 : node1111;
															assign node1111 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1115 = (inp[4]) ? 4'b1101 : node1116;
														assign node1116 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node1120 = (inp[12]) ? node1126 : node1121;
													assign node1121 = (inp[4]) ? 4'b1001 : node1122;
														assign node1122 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node1126 = (inp[10]) ? 4'b1001 : node1127;
														assign node1127 = (inp[7]) ? node1129 : 4'b0001;
															assign node1129 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node1133 = (inp[11]) ? node1185 : node1134;
											assign node1134 = (inp[13]) ? node1164 : node1135;
												assign node1135 = (inp[10]) ? node1153 : node1136;
													assign node1136 = (inp[12]) ? node1144 : node1137;
														assign node1137 = (inp[3]) ? node1139 : 4'b0100;
															assign node1139 = (inp[7]) ? node1141 : 4'b0000;
																assign node1141 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1144 = (inp[7]) ? 4'b1000 : node1145;
															assign node1145 = (inp[4]) ? node1149 : node1146;
																assign node1146 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node1149 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node1153 = (inp[3]) ? node1159 : node1154;
														assign node1154 = (inp[4]) ? 4'b0100 : node1155;
															assign node1155 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1159 = (inp[7]) ? node1161 : 4'b0000;
															assign node1161 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node1164 = (inp[10]) ? node1176 : node1165;
													assign node1165 = (inp[12]) ? node1169 : node1166;
														assign node1166 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1169 = (inp[3]) ? node1173 : node1170;
															assign node1170 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node1173 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node1176 = (inp[3]) ? node1180 : node1177;
														assign node1177 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1180 = (inp[4]) ? 4'b1000 : node1181;
															assign node1181 = (inp[12]) ? 4'b1000 : 4'b1100;
											assign node1185 = (inp[13]) ? node1213 : node1186;
												assign node1186 = (inp[10]) ? node1202 : node1187;
													assign node1187 = (inp[12]) ? node1195 : node1188;
														assign node1188 = (inp[4]) ? 4'b0101 : node1189;
															assign node1189 = (inp[7]) ? 4'b0001 : node1190;
																assign node1190 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node1195 = (inp[3]) ? node1197 : 4'b1001;
															assign node1197 = (inp[7]) ? 4'b1101 : node1198;
																assign node1198 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node1202 = (inp[3]) ? node1208 : node1203;
														assign node1203 = (inp[12]) ? node1205 : 4'b0101;
															assign node1205 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node1208 = (inp[7]) ? node1210 : 4'b0001;
															assign node1210 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node1213 = (inp[10]) ? node1231 : node1214;
													assign node1214 = (inp[12]) ? node1224 : node1215;
														assign node1215 = (inp[4]) ? 4'b1001 : node1216;
															assign node1216 = (inp[3]) ? node1220 : node1217;
																assign node1217 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node1220 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1224 = (inp[3]) ? node1226 : 4'b0101;
															assign node1226 = (inp[7]) ? node1228 : 4'b0001;
																assign node1228 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1231 = (inp[3]) ? node1237 : node1232;
														assign node1232 = (inp[7]) ? node1234 : 4'b1101;
															assign node1234 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node1237 = (inp[7]) ? node1239 : 4'b1001;
															assign node1239 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node1242 = (inp[3]) ? node1244 : 4'b1011;
									assign node1244 = (inp[4]) ? node1292 : node1245;
										assign node1245 = (inp[7]) ? 4'b1011 : node1246;
											assign node1246 = (inp[13]) ? node1272 : node1247;
												assign node1247 = (inp[12]) ? node1259 : node1248;
													assign node1248 = (inp[1]) ? node1256 : node1249;
														assign node1249 = (inp[14]) ? node1251 : 4'b0000;
															assign node1251 = (inp[11]) ? 4'b0000 : node1252;
																assign node1252 = (inp[10]) ? 4'b0001 : 4'b1011;
														assign node1256 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1259 = (inp[10]) ? node1261 : 4'b1011;
														assign node1261 = (inp[1]) ? node1267 : node1262;
															assign node1262 = (inp[11]) ? 4'b0000 : node1263;
																assign node1263 = (inp[14]) ? 4'b1011 : 4'b0000;
															assign node1267 = (inp[11]) ? 4'b0001 : node1268;
																assign node1268 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1272 = (inp[12]) ? node1280 : node1273;
													assign node1273 = (inp[1]) ? node1275 : 4'b1000;
														assign node1275 = (inp[14]) ? node1277 : 4'b1001;
															assign node1277 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node1280 = (inp[10]) ? node1286 : node1281;
														assign node1281 = (inp[14]) ? node1283 : 4'b0001;
															assign node1283 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node1286 = (inp[14]) ? node1288 : 4'b1000;
															assign node1288 = (inp[1]) ? 4'b1000 : 4'b0001;
										assign node1292 = (inp[1]) ? node1332 : node1293;
											assign node1293 = (inp[14]) ? node1307 : node1294;
												assign node1294 = (inp[13]) ? node1302 : node1295;
													assign node1295 = (inp[12]) ? node1297 : 4'b0000;
														assign node1297 = (inp[10]) ? 4'b0000 : node1298;
															assign node1298 = (inp[7]) ? 4'b1011 : 4'b1000;
													assign node1302 = (inp[10]) ? 4'b1000 : node1303;
														assign node1303 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node1307 = (inp[11]) ? node1321 : node1308;
													assign node1308 = (inp[12]) ? node1316 : node1309;
														assign node1309 = (inp[13]) ? node1313 : node1310;
															assign node1310 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node1313 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node1316 = (inp[7]) ? 4'b1011 : node1317;
															assign node1317 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node1321 = (inp[13]) ? node1327 : node1322;
														assign node1322 = (inp[12]) ? node1324 : 4'b0000;
															assign node1324 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node1327 = (inp[10]) ? 4'b1000 : node1328;
															assign node1328 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node1332 = (inp[14]) ? node1346 : node1333;
												assign node1333 = (inp[13]) ? node1341 : node1334;
													assign node1334 = (inp[12]) ? node1336 : 4'b0001;
														assign node1336 = (inp[10]) ? 4'b0001 : node1337;
															assign node1337 = (inp[7]) ? 4'b1011 : 4'b1001;
													assign node1341 = (inp[12]) ? node1343 : 4'b1001;
														assign node1343 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node1346 = (inp[11]) ? node1358 : node1347;
													assign node1347 = (inp[13]) ? node1353 : node1348;
														assign node1348 = (inp[10]) ? 4'b0000 : node1349;
															assign node1349 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node1353 = (inp[12]) ? node1355 : 4'b1000;
															assign node1355 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node1358 = (inp[10]) ? node1368 : node1359;
														assign node1359 = (inp[12]) ? node1363 : node1360;
															assign node1360 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node1363 = (inp[7]) ? 4'b1011 : node1364;
																assign node1364 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node1368 = (inp[13]) ? 4'b1001 : 4'b0001;
				assign node1372 = (inp[5]) ? node3344 : node1373;
					assign node1373 = (inp[0]) ? node2927 : node1374;
						assign node1374 = (inp[11]) ? node2320 : node1375;
							assign node1375 = (inp[10]) ? node1865 : node1376;
								assign node1376 = (inp[12]) ? node1596 : node1377;
									assign node1377 = (inp[2]) ? node1489 : node1378;
										assign node1378 = (inp[1]) ? node1438 : node1379;
											assign node1379 = (inp[14]) ? node1409 : node1380;
												assign node1380 = (inp[15]) ? node1396 : node1381;
													assign node1381 = (inp[4]) ? node1387 : node1382;
														assign node1382 = (inp[7]) ? node1384 : 4'b0000;
															assign node1384 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node1387 = (inp[3]) ? node1391 : node1388;
															assign node1388 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node1391 = (inp[13]) ? node1393 : 4'b0001;
																assign node1393 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node1396 = (inp[4]) ? node1404 : node1397;
														assign node1397 = (inp[3]) ? node1399 : 4'b1100;
															assign node1399 = (inp[13]) ? 4'b0100 : node1400;
																assign node1400 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1404 = (inp[7]) ? node1406 : 4'b0000;
															assign node1406 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node1409 = (inp[15]) ? node1421 : node1410;
													assign node1410 = (inp[4]) ? node1412 : 4'b0000;
														assign node1412 = (inp[13]) ? node1418 : node1413;
															assign node1413 = (inp[3]) ? 4'b0000 : node1414;
																assign node1414 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node1418 = (inp[3]) ? 4'b1100 : 4'b0100;
													assign node1421 = (inp[3]) ? node1429 : node1422;
														assign node1422 = (inp[4]) ? node1424 : 4'b1001;
															assign node1424 = (inp[7]) ? node1426 : 4'b0000;
																assign node1426 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node1429 = (inp[7]) ? node1433 : node1430;
															assign node1430 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node1433 = (inp[4]) ? 4'b0000 : node1434;
																assign node1434 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node1438 = (inp[13]) ? node1468 : node1439;
												assign node1439 = (inp[4]) ? node1451 : node1440;
													assign node1440 = (inp[15]) ? node1448 : node1441;
														assign node1441 = (inp[7]) ? node1443 : 4'b0000;
															assign node1443 = (inp[3]) ? 4'b0100 : node1444;
																assign node1444 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1448 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1451 = (inp[3]) ? node1461 : node1452;
														assign node1452 = (inp[15]) ? node1456 : node1453;
															assign node1453 = (inp[14]) ? 4'b0000 : 4'b0100;
															assign node1456 = (inp[7]) ? node1458 : 4'b0000;
																assign node1458 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1461 = (inp[14]) ? node1465 : node1462;
															assign node1462 = (inp[15]) ? 4'b0000 : 4'b1000;
															assign node1465 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node1468 = (inp[15]) ? node1476 : node1469;
													assign node1469 = (inp[4]) ? node1471 : 4'b0000;
														assign node1471 = (inp[3]) ? node1473 : 4'b0100;
															assign node1473 = (inp[7]) ? 4'b0100 : 4'b1101;
													assign node1476 = (inp[4]) ? node1484 : node1477;
														assign node1477 = (inp[3]) ? 4'b0100 : node1478;
															assign node1478 = (inp[14]) ? 4'b1000 : node1479;
																assign node1479 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1484 = (inp[3]) ? node1486 : 4'b0000;
															assign node1486 = (inp[7]) ? 4'b0000 : 4'b1001;
										assign node1489 = (inp[3]) ? node1555 : node1490;
											assign node1490 = (inp[13]) ? node1524 : node1491;
												assign node1491 = (inp[1]) ? node1511 : node1492;
													assign node1492 = (inp[14]) ? node1502 : node1493;
														assign node1493 = (inp[15]) ? node1497 : node1494;
															assign node1494 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node1497 = (inp[7]) ? node1499 : 4'b0100;
																assign node1499 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1502 = (inp[7]) ? 4'b1101 : node1503;
															assign node1503 = (inp[4]) ? node1507 : node1504;
																assign node1504 = (inp[15]) ? 4'b1001 : 4'b1101;
																assign node1507 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node1511 = (inp[14]) ? node1517 : node1512;
														assign node1512 = (inp[7]) ? 4'b0001 : node1513;
															assign node1513 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node1517 = (inp[7]) ? node1519 : 4'b0000;
															assign node1519 = (inp[4]) ? 4'b0100 : node1520;
																assign node1520 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node1524 = (inp[14]) ? node1542 : node1525;
													assign node1525 = (inp[1]) ? node1535 : node1526;
														assign node1526 = (inp[15]) ? node1532 : node1527;
															assign node1527 = (inp[4]) ? 4'b1000 : node1528;
																assign node1528 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1532 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1535 = (inp[15]) ? 4'b1101 : node1536;
															assign node1536 = (inp[7]) ? node1538 : 4'b1001;
																assign node1538 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node1542 = (inp[1]) ? node1552 : node1543;
														assign node1543 = (inp[15]) ? node1547 : node1544;
															assign node1544 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node1547 = (inp[4]) ? 4'b0101 : node1548;
																assign node1548 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1552 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node1555 = (inp[15]) ? node1569 : node1556;
												assign node1556 = (inp[4]) ? node1564 : node1557;
													assign node1557 = (inp[7]) ? node1559 : 4'b0000;
														assign node1559 = (inp[13]) ? 4'b0000 : node1560;
															assign node1560 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node1564 = (inp[7]) ? node1566 : 4'b0100;
														assign node1566 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node1569 = (inp[4]) ? node1585 : node1570;
													assign node1570 = (inp[7]) ? node1576 : node1571;
														assign node1571 = (inp[13]) ? node1573 : 4'b0001;
															assign node1573 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1576 = (inp[1]) ? node1582 : node1577;
															assign node1577 = (inp[14]) ? node1579 : 4'b1100;
																assign node1579 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node1582 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node1585 = (inp[13]) ? 4'b0000 : node1586;
														assign node1586 = (inp[1]) ? node1590 : node1587;
															assign node1587 = (inp[14]) ? 4'b1101 : 4'b0000;
															assign node1590 = (inp[7]) ? node1592 : 4'b0000;
																assign node1592 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node1596 = (inp[13]) ? node1724 : node1597;
										assign node1597 = (inp[1]) ? node1657 : node1598;
											assign node1598 = (inp[14]) ? node1626 : node1599;
												assign node1599 = (inp[4]) ? node1611 : node1600;
													assign node1600 = (inp[3]) ? node1602 : 4'b1100;
														assign node1602 = (inp[7]) ? 4'b1100 : node1603;
															assign node1603 = (inp[15]) ? node1607 : node1604;
																assign node1604 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node1607 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node1611 = (inp[2]) ? node1615 : node1612;
														assign node1612 = (inp[3]) ? 4'b1001 : 4'b1000;
														assign node1615 = (inp[15]) ? node1621 : node1616;
															assign node1616 = (inp[7]) ? node1618 : 4'b1000;
																assign node1618 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node1621 = (inp[7]) ? node1623 : 4'b1100;
																assign node1623 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node1626 = (inp[3]) ? node1640 : node1627;
													assign node1627 = (inp[15]) ? node1635 : node1628;
														assign node1628 = (inp[4]) ? node1630 : 4'b1101;
															assign node1630 = (inp[2]) ? node1632 : 4'b1000;
																assign node1632 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1635 = (inp[7]) ? 4'b1001 : node1636;
															assign node1636 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node1640 = (inp[2]) ? node1648 : node1641;
														assign node1641 = (inp[4]) ? node1645 : node1642;
															assign node1642 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node1645 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node1648 = (inp[15]) ? node1652 : node1649;
															assign node1649 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node1652 = (inp[7]) ? 4'b1101 : node1653;
																assign node1653 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node1657 = (inp[3]) ? node1689 : node1658;
												assign node1658 = (inp[14]) ? node1670 : node1659;
													assign node1659 = (inp[15]) ? node1663 : node1660;
														assign node1660 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1663 = (inp[2]) ? node1667 : node1664;
															assign node1664 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node1667 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node1670 = (inp[15]) ? node1684 : node1671;
														assign node1671 = (inp[2]) ? node1679 : node1672;
															assign node1672 = (inp[7]) ? node1676 : node1673;
																assign node1673 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node1676 = (inp[4]) ? 4'b0000 : 4'b1100;
															assign node1679 = (inp[4]) ? node1681 : 4'b1100;
																assign node1681 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node1684 = (inp[7]) ? 4'b1000 : node1685;
															assign node1685 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node1689 = (inp[2]) ? node1705 : node1690;
													assign node1690 = (inp[14]) ? node1696 : node1691;
														assign node1691 = (inp[7]) ? 4'b0100 : node1692;
															assign node1692 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1696 = (inp[4]) ? node1702 : node1697;
															assign node1697 = (inp[15]) ? 4'b0000 : node1698;
																assign node1698 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node1702 = (inp[15]) ? 4'b0100 : 4'b0001;
													assign node1705 = (inp[7]) ? node1715 : node1706;
														assign node1706 = (inp[14]) ? node1708 : 4'b0000;
															assign node1708 = (inp[4]) ? node1712 : node1709;
																assign node1709 = (inp[15]) ? 4'b1100 : 4'b0000;
																assign node1712 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1715 = (inp[15]) ? node1721 : node1716;
															assign node1716 = (inp[14]) ? node1718 : 4'b1001;
																assign node1718 = (inp[4]) ? 4'b0000 : 4'b1000;
															assign node1721 = (inp[4]) ? 4'b1101 : 4'b1100;
										assign node1724 = (inp[1]) ? node1792 : node1725;
											assign node1725 = (inp[2]) ? node1761 : node1726;
												assign node1726 = (inp[15]) ? node1746 : node1727;
													assign node1727 = (inp[3]) ? node1737 : node1728;
														assign node1728 = (inp[4]) ? node1734 : node1729;
															assign node1729 = (inp[7]) ? node1731 : 4'b1000;
																assign node1731 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1734 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1737 = (inp[4]) ? node1741 : node1738;
															assign node1738 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1741 = (inp[14]) ? 4'b0100 : node1742;
																assign node1742 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1746 = (inp[3]) ? node1754 : node1747;
														assign node1747 = (inp[7]) ? node1751 : node1748;
															assign node1748 = (inp[4]) ? 4'b1000 : 4'b0101;
															assign node1751 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node1754 = (inp[4]) ? node1758 : node1755;
															assign node1755 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node1758 = (inp[7]) ? 4'b1100 : 4'b0000;
												assign node1761 = (inp[14]) ? node1777 : node1762;
													assign node1762 = (inp[3]) ? node1770 : node1763;
														assign node1763 = (inp[15]) ? node1765 : 4'b0000;
															assign node1765 = (inp[4]) ? 4'b0100 : node1766;
																assign node1766 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1770 = (inp[4]) ? 4'b1000 : node1771;
															assign node1771 = (inp[15]) ? 4'b0000 : node1772;
																assign node1772 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node1777 = (inp[3]) ? node1783 : node1778;
														assign node1778 = (inp[4]) ? 4'b0001 : node1779;
															assign node1779 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node1783 = (inp[7]) ? node1787 : node1784;
															assign node1784 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node1787 = (inp[15]) ? 4'b0001 : node1788;
																assign node1788 = (inp[4]) ? 4'b1000 : 4'b0001;
											assign node1792 = (inp[14]) ? node1824 : node1793;
												assign node1793 = (inp[3]) ? node1811 : node1794;
													assign node1794 = (inp[2]) ? node1804 : node1795;
														assign node1795 = (inp[15]) ? node1799 : node1796;
															assign node1796 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node1799 = (inp[4]) ? 4'b0000 : node1800;
																assign node1800 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node1804 = (inp[15]) ? node1806 : 4'b0001;
															assign node1806 = (inp[4]) ? 4'b0101 : node1807;
																assign node1807 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1811 = (inp[2]) ? node1817 : node1812;
														assign node1812 = (inp[4]) ? 4'b1000 : node1813;
															assign node1813 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node1817 = (inp[15]) ? node1821 : node1818;
															assign node1818 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node1821 = (inp[4]) ? 4'b0000 : 4'b0001;
												assign node1824 = (inp[7]) ? node1846 : node1825;
													assign node1825 = (inp[2]) ? node1833 : node1826;
														assign node1826 = (inp[15]) ? node1830 : node1827;
															assign node1827 = (inp[3]) ? 4'b0000 : 4'b0100;
															assign node1830 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1833 = (inp[4]) ? node1839 : node1834;
															assign node1834 = (inp[15]) ? node1836 : 4'b0000;
																assign node1836 = (inp[3]) ? 4'b0000 : 4'b0100;
															assign node1839 = (inp[15]) ? node1843 : node1840;
																assign node1840 = (inp[3]) ? 4'b0100 : 4'b0000;
																assign node1843 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node1846 = (inp[2]) ? node1852 : node1847;
														assign node1847 = (inp[3]) ? node1849 : 4'b0000;
															assign node1849 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1852 = (inp[4]) ? node1858 : node1853;
															assign node1853 = (inp[3]) ? 4'b0000 : node1854;
																assign node1854 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node1858 = (inp[3]) ? node1862 : node1859;
																assign node1859 = (inp[15]) ? 4'b0100 : 4'b0000;
																assign node1862 = (inp[15]) ? 4'b0000 : 4'b0100;
								assign node1865 = (inp[13]) ? node2115 : node1866;
									assign node1866 = (inp[3]) ? node1982 : node1867;
										assign node1867 = (inp[2]) ? node1927 : node1868;
											assign node1868 = (inp[7]) ? node1892 : node1869;
												assign node1869 = (inp[4]) ? node1885 : node1870;
													assign node1870 = (inp[15]) ? node1876 : node1871;
														assign node1871 = (inp[12]) ? node1873 : 4'b1000;
															assign node1873 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node1876 = (inp[14]) ? node1880 : node1877;
															assign node1877 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node1880 = (inp[1]) ? 4'b0100 : node1881;
																assign node1881 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node1885 = (inp[15]) ? 4'b1000 : node1886;
														assign node1886 = (inp[1]) ? 4'b1100 : node1887;
															assign node1887 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node1892 = (inp[15]) ? node1904 : node1893;
													assign node1893 = (inp[4]) ? node1901 : node1894;
														assign node1894 = (inp[14]) ? node1898 : node1895;
															assign node1895 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node1898 = (inp[1]) ? 4'b0100 : 4'b1101;
														assign node1901 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node1904 = (inp[4]) ? node1912 : node1905;
														assign node1905 = (inp[14]) ? node1909 : node1906;
															assign node1906 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1909 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node1912 = (inp[12]) ? node1920 : node1913;
															assign node1913 = (inp[1]) ? node1917 : node1914;
																assign node1914 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node1917 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node1920 = (inp[14]) ? node1924 : node1921;
																assign node1921 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node1924 = (inp[1]) ? 4'b0100 : 4'b1001;
											assign node1927 = (inp[15]) ? node1953 : node1928;
												assign node1928 = (inp[4]) ? node1942 : node1929;
													assign node1929 = (inp[7]) ? node1937 : node1930;
														assign node1930 = (inp[14]) ? node1934 : node1931;
															assign node1931 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1934 = (inp[1]) ? 4'b0000 : 4'b1101;
														assign node1937 = (inp[1]) ? node1939 : 4'b0100;
															assign node1939 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1942 = (inp[12]) ? node1948 : node1943;
														assign node1943 = (inp[14]) ? node1945 : 4'b0001;
															assign node1945 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node1948 = (inp[7]) ? 4'b0000 : node1949;
															assign node1949 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node1953 = (inp[7]) ? node1965 : node1954;
													assign node1954 = (inp[12]) ? node1960 : node1955;
														assign node1955 = (inp[14]) ? node1957 : 4'b0100;
															assign node1957 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node1960 = (inp[14]) ? 4'b0100 : node1961;
															assign node1961 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node1965 = (inp[4]) ? node1975 : node1966;
														assign node1966 = (inp[14]) ? node1970 : node1967;
															assign node1967 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1970 = (inp[1]) ? 4'b0000 : node1971;
																assign node1971 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node1975 = (inp[1]) ? node1979 : node1976;
															assign node1976 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1979 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node1982 = (inp[2]) ? node2050 : node1983;
											assign node1983 = (inp[12]) ? node2017 : node1984;
												assign node1984 = (inp[1]) ? node2004 : node1985;
													assign node1985 = (inp[4]) ? node1999 : node1986;
														assign node1986 = (inp[14]) ? node1992 : node1987;
															assign node1987 = (inp[7]) ? 4'b1000 : node1988;
																assign node1988 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node1992 = (inp[15]) ? node1996 : node1993;
																assign node1993 = (inp[7]) ? 4'b1100 : 4'b1000;
																assign node1996 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1999 = (inp[15]) ? 4'b1000 : node2000;
															assign node2000 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node2004 = (inp[4]) ? node2012 : node2005;
														assign node2005 = (inp[7]) ? node2009 : node2006;
															assign node2006 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node2009 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node2012 = (inp[7]) ? 4'b1100 : node2013;
															assign node2013 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node2017 = (inp[1]) ? node2031 : node2018;
													assign node2018 = (inp[15]) ? node2024 : node2019;
														assign node2019 = (inp[4]) ? 4'b1001 : node2020;
															assign node2020 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node2024 = (inp[4]) ? node2028 : node2025;
															assign node2025 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node2028 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2031 = (inp[14]) ? node2041 : node2032;
														assign node2032 = (inp[4]) ? node2034 : 4'b1100;
															assign node2034 = (inp[15]) ? node2038 : node2035;
																assign node2035 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node2038 = (inp[7]) ? 4'b1100 : 4'b0000;
														assign node2041 = (inp[15]) ? node2045 : node2042;
															assign node2042 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node2045 = (inp[7]) ? node2047 : 4'b1000;
																assign node2047 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node2050 = (inp[15]) ? node2078 : node2051;
												assign node2051 = (inp[7]) ? node2063 : node2052;
													assign node2052 = (inp[4]) ? node2058 : node2053;
														assign node2053 = (inp[1]) ? 4'b1000 : node2054;
															assign node2054 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2058 = (inp[1]) ? 4'b1100 : node2059;
															assign node2059 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2063 = (inp[4]) ? node2073 : node2064;
														assign node2064 = (inp[1]) ? node2070 : node2065;
															assign node2065 = (inp[12]) ? 4'b1001 : node2066;
																assign node2066 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node2070 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node2073 = (inp[12]) ? node2075 : 4'b1000;
															assign node2075 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node2078 = (inp[7]) ? node2096 : node2079;
													assign node2079 = (inp[4]) ? node2091 : node2080;
														assign node2080 = (inp[12]) ? node2088 : node2081;
															assign node2081 = (inp[1]) ? node2085 : node2082;
																assign node2082 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node2085 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node2088 = (inp[1]) ? 4'b0001 : 4'b1101;
														assign node2091 = (inp[1]) ? 4'b1000 : node2092;
															assign node2092 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2096 = (inp[4]) ? node2108 : node2097;
														assign node2097 = (inp[12]) ? node2105 : node2098;
															assign node2098 = (inp[14]) ? node2102 : node2099;
																assign node2099 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node2102 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node2105 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node2108 = (inp[14]) ? node2112 : node2109;
															assign node2109 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2112 = (inp[12]) ? 4'b1101 : 4'b0001;
									assign node2115 = (inp[1]) ? node2241 : node2116;
										assign node2116 = (inp[12]) ? node2178 : node2117;
											assign node2117 = (inp[2]) ? node2143 : node2118;
												assign node2118 = (inp[3]) ? node2132 : node2119;
													assign node2119 = (inp[4]) ? node2129 : node2120;
														assign node2120 = (inp[15]) ? node2122 : 4'b1000;
															assign node2122 = (inp[7]) ? node2126 : node2123;
																assign node2123 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node2126 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node2129 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node2132 = (inp[4]) ? node2138 : node2133;
														assign node2133 = (inp[15]) ? 4'b1100 : node2134;
															assign node2134 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node2138 = (inp[14]) ? 4'b0100 : node2139;
															assign node2139 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node2143 = (inp[14]) ? node2167 : node2144;
													assign node2144 = (inp[7]) ? node2154 : node2145;
														assign node2145 = (inp[3]) ? node2149 : node2146;
															assign node2146 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node2149 = (inp[15]) ? 4'b1000 : node2150;
																assign node2150 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2154 = (inp[4]) ? node2160 : node2155;
															assign node2155 = (inp[15]) ? 4'b1100 : node2156;
																assign node2156 = (inp[3]) ? 4'b1000 : 4'b1100;
															assign node2160 = (inp[3]) ? node2164 : node2161;
																assign node2161 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node2164 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node2167 = (inp[3]) ? node2173 : node2168;
														assign node2168 = (inp[15]) ? node2170 : 4'b1001;
															assign node2170 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node2173 = (inp[7]) ? node2175 : 4'b1000;
															assign node2175 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node2178 = (inp[14]) ? node2216 : node2179;
												assign node2179 = (inp[2]) ? node2197 : node2180;
													assign node2180 = (inp[3]) ? node2190 : node2181;
														assign node2181 = (inp[4]) ? node2187 : node2182;
															assign node2182 = (inp[15]) ? node2184 : 4'b0000;
																assign node2184 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node2187 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node2190 = (inp[4]) ? 4'b0001 : node2191;
															assign node2191 = (inp[15]) ? 4'b0100 : node2192;
																assign node2192 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node2197 = (inp[3]) ? node2209 : node2198;
														assign node2198 = (inp[15]) ? node2204 : node2199;
															assign node2199 = (inp[4]) ? 4'b1000 : node2200;
																assign node2200 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node2204 = (inp[7]) ? node2206 : 4'b1100;
																assign node2206 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2209 = (inp[4]) ? node2213 : node2210;
															assign node2210 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node2213 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node2216 = (inp[2]) ? node2226 : node2217;
													assign node2217 = (inp[15]) ? node2221 : node2218;
														assign node2218 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node2221 = (inp[4]) ? 4'b0000 : node2222;
															assign node2222 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node2226 = (inp[3]) ? node2234 : node2227;
														assign node2227 = (inp[4]) ? 4'b0101 : node2228;
															assign node2228 = (inp[15]) ? node2230 : 4'b0001;
																assign node2230 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2234 = (inp[4]) ? node2238 : node2235;
															assign node2235 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node2238 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node2241 = (inp[14]) ? node2277 : node2242;
											assign node2242 = (inp[3]) ? node2266 : node2243;
												assign node2243 = (inp[2]) ? node2255 : node2244;
													assign node2244 = (inp[12]) ? node2250 : node2245;
														assign node2245 = (inp[7]) ? node2247 : 4'b1000;
															assign node2247 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node2250 = (inp[15]) ? 4'b1101 : node2251;
															assign node2251 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2255 = (inp[15]) ? node2261 : node2256;
														assign node2256 = (inp[4]) ? 4'b1001 : node2257;
															assign node2257 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node2261 = (inp[7]) ? node2263 : 4'b1101;
															assign node2263 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node2266 = (inp[15]) ? node2270 : node2267;
													assign node2267 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2270 = (inp[4]) ? 4'b1000 : node2271;
														assign node2271 = (inp[2]) ? node2273 : 4'b1100;
															assign node2273 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node2277 = (inp[3]) ? node2299 : node2278;
												assign node2278 = (inp[4]) ? node2290 : node2279;
													assign node2279 = (inp[2]) ? node2285 : node2280;
														assign node2280 = (inp[7]) ? 4'b1000 : node2281;
															assign node2281 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node2285 = (inp[15]) ? 4'b1000 : node2286;
															assign node2286 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node2290 = (inp[7]) ? 4'b1100 : node2291;
														assign node2291 = (inp[2]) ? node2295 : node2292;
															assign node2292 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node2295 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node2299 = (inp[2]) ? node2311 : node2300;
													assign node2300 = (inp[4]) ? node2304 : node2301;
														assign node2301 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node2304 = (inp[12]) ? node2308 : node2305;
															assign node2305 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node2308 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2311 = (inp[15]) ? node2315 : node2312;
														assign node2312 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2315 = (inp[4]) ? 4'b1000 : node2316;
															assign node2316 = (inp[7]) ? 4'b1100 : 4'b1000;
							assign node2320 = (inp[1]) ? node2658 : node2321;
								assign node2321 = (inp[3]) ? node2483 : node2322;
									assign node2322 = (inp[2]) ? node2428 : node2323;
										assign node2323 = (inp[15]) ? node2379 : node2324;
											assign node2324 = (inp[4]) ? node2354 : node2325;
												assign node2325 = (inp[13]) ? node2337 : node2326;
													assign node2326 = (inp[7]) ? node2334 : node2327;
														assign node2327 = (inp[12]) ? node2331 : node2328;
															assign node2328 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2331 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node2334 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node2337 = (inp[7]) ? node2347 : node2338;
														assign node2338 = (inp[14]) ? 4'b1001 : node2339;
															assign node2339 = (inp[10]) ? node2343 : node2340;
																assign node2340 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node2343 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2347 = (inp[12]) ? node2351 : node2348;
															assign node2348 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2351 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node2354 = (inp[7]) ? node2362 : node2355;
													assign node2355 = (inp[10]) ? node2359 : node2356;
														assign node2356 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node2359 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node2362 = (inp[13]) ? node2374 : node2363;
														assign node2363 = (inp[14]) ? node2369 : node2364;
															assign node2364 = (inp[12]) ? 4'b0001 : node2365;
																assign node2365 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2369 = (inp[10]) ? 4'b1001 : node2370;
																assign node2370 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2374 = (inp[12]) ? 4'b1001 : node2375;
															assign node2375 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node2379 = (inp[4]) ? node2397 : node2380;
												assign node2380 = (inp[7]) ? node2390 : node2381;
													assign node2381 = (inp[13]) ? node2385 : node2382;
														assign node2382 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node2385 = (inp[12]) ? node2387 : 4'b1100;
															assign node2387 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2390 = (inp[13]) ? 4'b1000 : node2391;
														assign node2391 = (inp[12]) ? node2393 : 4'b0000;
															assign node2393 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node2397 = (inp[13]) ? node2407 : node2398;
													assign node2398 = (inp[10]) ? node2402 : node2399;
														assign node2399 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node2402 = (inp[7]) ? 4'b0100 : node2403;
															assign node2403 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2407 = (inp[14]) ? node2419 : node2408;
														assign node2408 = (inp[7]) ? node2414 : node2409;
															assign node2409 = (inp[12]) ? 4'b1001 : node2410;
																assign node2410 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2414 = (inp[10]) ? node2416 : 4'b0001;
																assign node2416 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2419 = (inp[7]) ? node2425 : node2420;
															assign node2420 = (inp[12]) ? node2422 : 4'b0001;
																assign node2422 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node2425 = (inp[10]) ? 4'b0001 : 4'b0100;
										assign node2428 = (inp[13]) ? node2460 : node2429;
											assign node2429 = (inp[10]) ? node2449 : node2430;
												assign node2430 = (inp[12]) ? node2436 : node2431;
													assign node2431 = (inp[4]) ? node2433 : 4'b0000;
														assign node2433 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node2436 = (inp[15]) ? node2444 : node2437;
														assign node2437 = (inp[14]) ? node2439 : 4'b1100;
															assign node2439 = (inp[4]) ? node2441 : 4'b1100;
																assign node2441 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node2444 = (inp[4]) ? node2446 : 4'b1000;
															assign node2446 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node2449 = (inp[15]) ? node2455 : node2450;
													assign node2450 = (inp[7]) ? node2452 : 4'b0000;
														assign node2452 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node2455 = (inp[7]) ? node2457 : 4'b0100;
														assign node2457 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node2460 = (inp[15]) ? node2470 : node2461;
												assign node2461 = (inp[10]) ? node2465 : node2462;
													assign node2462 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2465 = (inp[7]) ? node2467 : 4'b1000;
														assign node2467 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node2470 = (inp[7]) ? node2476 : node2471;
													assign node2471 = (inp[12]) ? node2473 : 4'b1100;
														assign node2473 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2476 = (inp[4]) ? node2478 : 4'b1000;
														assign node2478 = (inp[10]) ? 4'b1100 : node2479;
															assign node2479 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node2483 = (inp[7]) ? node2563 : node2484;
										assign node2484 = (inp[2]) ? node2528 : node2485;
											assign node2485 = (inp[4]) ? node2509 : node2486;
												assign node2486 = (inp[15]) ? node2500 : node2487;
													assign node2487 = (inp[13]) ? node2495 : node2488;
														assign node2488 = (inp[12]) ? node2492 : node2489;
															assign node2489 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2492 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node2495 = (inp[10]) ? node2497 : 4'b1001;
															assign node2497 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node2500 = (inp[10]) ? node2506 : node2501;
														assign node2501 = (inp[12]) ? node2503 : 4'b0101;
															assign node2503 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node2506 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node2509 = (inp[13]) ? node2521 : node2510;
													assign node2510 = (inp[15]) ? node2514 : node2511;
														assign node2511 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node2514 = (inp[14]) ? node2516 : 4'b1101;
															assign node2516 = (inp[10]) ? node2518 : 4'b0001;
																assign node2518 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node2521 = (inp[15]) ? node2525 : node2522;
														assign node2522 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node2525 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2528 = (inp[4]) ? node2550 : node2529;
												assign node2529 = (inp[15]) ? node2539 : node2530;
													assign node2530 = (inp[10]) ? node2536 : node2531;
														assign node2531 = (inp[12]) ? node2533 : 4'b0001;
															assign node2533 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node2536 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2539 = (inp[13]) ? node2545 : node2540;
														assign node2540 = (inp[12]) ? node2542 : 4'b0000;
															assign node2542 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node2545 = (inp[10]) ? 4'b1000 : node2546;
															assign node2546 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2550 = (inp[15]) ? node2556 : node2551;
													assign node2551 = (inp[12]) ? 4'b0101 : node2552;
														assign node2552 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node2556 = (inp[10]) ? node2560 : node2557;
														assign node2557 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2560 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2563 = (inp[13]) ? node2607 : node2564;
											assign node2564 = (inp[2]) ? node2590 : node2565;
												assign node2565 = (inp[4]) ? node2579 : node2566;
													assign node2566 = (inp[15]) ? node2574 : node2567;
														assign node2567 = (inp[14]) ? node2569 : 4'b1101;
															assign node2569 = (inp[12]) ? node2571 : 4'b0101;
																assign node2571 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node2574 = (inp[10]) ? node2576 : 4'b0001;
															assign node2576 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node2579 = (inp[15]) ? node2585 : node2580;
														assign node2580 = (inp[12]) ? node2582 : 4'b0000;
															assign node2582 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node2585 = (inp[12]) ? 4'b0101 : node2586;
															assign node2586 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node2590 = (inp[15]) ? node2600 : node2591;
													assign node2591 = (inp[4]) ? node2597 : node2592;
														assign node2592 = (inp[12]) ? node2594 : 4'b0000;
															assign node2594 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node2597 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2600 = (inp[4]) ? 4'b0000 : node2601;
														assign node2601 = (inp[12]) ? node2603 : 4'b0100;
															assign node2603 = (inp[10]) ? 4'b0100 : 4'b1100;
											assign node2607 = (inp[15]) ? node2629 : node2608;
												assign node2608 = (inp[4]) ? node2616 : node2609;
													assign node2609 = (inp[10]) ? node2613 : node2610;
														assign node2610 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node2613 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2616 = (inp[2]) ? node2622 : node2617;
														assign node2617 = (inp[12]) ? 4'b0100 : node2618;
															assign node2618 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node2622 = (inp[12]) ? node2626 : node2623;
															assign node2623 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node2626 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node2629 = (inp[4]) ? node2643 : node2630;
													assign node2630 = (inp[2]) ? node2638 : node2631;
														assign node2631 = (inp[12]) ? node2635 : node2632;
															assign node2632 = (inp[14]) ? 4'b0101 : 4'b1101;
															assign node2635 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node2638 = (inp[12]) ? node2640 : 4'b1100;
															assign node2640 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2643 = (inp[10]) ? node2651 : node2644;
														assign node2644 = (inp[2]) ? node2648 : node2645;
															assign node2645 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node2648 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node2651 = (inp[12]) ? node2655 : node2652;
															assign node2652 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node2655 = (inp[2]) ? 4'b0001 : 4'b0000;
								assign node2658 = (inp[10]) ? node2820 : node2659;
									assign node2659 = (inp[3]) ? node2749 : node2660;
										assign node2660 = (inp[2]) ? node2696 : node2661;
											assign node2661 = (inp[15]) ? node2675 : node2662;
												assign node2662 = (inp[4]) ? node2670 : node2663;
													assign node2663 = (inp[7]) ? node2665 : 4'b0001;
														assign node2665 = (inp[13]) ? 4'b0001 : node2666;
															assign node2666 = (inp[14]) ? 4'b0101 : 4'b1101;
													assign node2670 = (inp[7]) ? node2672 : 4'b0101;
														assign node2672 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node2675 = (inp[4]) ? node2689 : node2676;
													assign node2676 = (inp[7]) ? node2684 : node2677;
														assign node2677 = (inp[13]) ? node2681 : node2678;
															assign node2678 = (inp[14]) ? 4'b0101 : 4'b1001;
															assign node2681 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2684 = (inp[12]) ? 4'b1001 : node2685;
															assign node2685 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node2689 = (inp[7]) ? node2691 : 4'b0001;
														assign node2691 = (inp[12]) ? 4'b1001 : node2692;
															assign node2692 = (inp[14]) ? 4'b0101 : 4'b0001;
											assign node2696 = (inp[15]) ? node2718 : node2697;
												assign node2697 = (inp[12]) ? node2711 : node2698;
													assign node2698 = (inp[13]) ? node2706 : node2699;
														assign node2699 = (inp[14]) ? 4'b0001 : node2700;
															assign node2700 = (inp[7]) ? node2702 : 4'b0001;
																assign node2702 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2706 = (inp[7]) ? node2708 : 4'b1001;
															assign node2708 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node2711 = (inp[13]) ? node2713 : 4'b1101;
														assign node2713 = (inp[7]) ? node2715 : 4'b0001;
															assign node2715 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node2718 = (inp[7]) ? node2738 : node2719;
													assign node2719 = (inp[4]) ? node2727 : node2720;
														assign node2720 = (inp[13]) ? node2724 : node2721;
															assign node2721 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node2724 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2727 = (inp[14]) ? node2733 : node2728;
															assign node2728 = (inp[13]) ? 4'b1101 : node2729;
																assign node2729 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node2733 = (inp[12]) ? node2735 : 4'b0101;
																assign node2735 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node2738 = (inp[4]) ? node2744 : node2739;
														assign node2739 = (inp[13]) ? node2741 : 4'b0001;
															assign node2741 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2744 = (inp[12]) ? 4'b1001 : node2745;
															assign node2745 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node2749 = (inp[12]) ? node2781 : node2750;
											assign node2750 = (inp[4]) ? node2770 : node2751;
												assign node2751 = (inp[15]) ? node2759 : node2752;
													assign node2752 = (inp[13]) ? 4'b0001 : node2753;
														assign node2753 = (inp[2]) ? 4'b0001 : node2754;
															assign node2754 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node2759 = (inp[13]) ? node2765 : node2760;
														assign node2760 = (inp[2]) ? node2762 : 4'b0001;
															assign node2762 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node2765 = (inp[7]) ? node2767 : 4'b1001;
															assign node2767 = (inp[14]) ? 4'b0101 : 4'b1101;
												assign node2770 = (inp[15]) ? node2776 : node2771;
													assign node2771 = (inp[13]) ? 4'b0101 : node2772;
														assign node2772 = (inp[7]) ? 4'b1001 : 4'b0101;
													assign node2776 = (inp[13]) ? 4'b0001 : node2777;
														assign node2777 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node2781 = (inp[15]) ? node2799 : node2782;
												assign node2782 = (inp[4]) ? node2788 : node2783;
													assign node2783 = (inp[13]) ? 4'b0001 : node2784;
														assign node2784 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node2788 = (inp[13]) ? node2794 : node2789;
														assign node2789 = (inp[2]) ? node2791 : 4'b0001;
															assign node2791 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2794 = (inp[2]) ? 4'b0101 : node2795;
															assign node2795 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2799 = (inp[4]) ? node2811 : node2800;
													assign node2800 = (inp[2]) ? node2806 : node2801;
														assign node2801 = (inp[7]) ? node2803 : 4'b0101;
															assign node2803 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node2806 = (inp[13]) ? node2808 : 4'b1101;
															assign node2808 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node2811 = (inp[2]) ? 4'b0001 : node2812;
														assign node2812 = (inp[7]) ? node2816 : node2813;
															assign node2813 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node2816 = (inp[14]) ? 4'b0001 : 4'b0101;
									assign node2820 = (inp[13]) ? node2878 : node2821;
										assign node2821 = (inp[3]) ? node2849 : node2822;
											assign node2822 = (inp[2]) ? node2838 : node2823;
												assign node2823 = (inp[4]) ? node2831 : node2824;
													assign node2824 = (inp[15]) ? node2828 : node2825;
														assign node2825 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node2828 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2831 = (inp[7]) ? node2835 : node2832;
														assign node2832 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node2835 = (inp[15]) ? 4'b0101 : 4'b1001;
												assign node2838 = (inp[15]) ? node2844 : node2839;
													assign node2839 = (inp[7]) ? node2841 : 4'b0001;
														assign node2841 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node2844 = (inp[4]) ? 4'b0101 : node2845;
														assign node2845 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node2849 = (inp[7]) ? node2863 : node2850;
												assign node2850 = (inp[2]) ? node2858 : node2851;
													assign node2851 = (inp[4]) ? node2855 : node2852;
														assign node2852 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node2855 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2858 = (inp[15]) ? 4'b1001 : node2859;
														assign node2859 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node2863 = (inp[2]) ? node2871 : node2864;
													assign node2864 = (inp[15]) ? node2868 : node2865;
														assign node2865 = (inp[4]) ? 4'b0001 : 4'b1101;
														assign node2868 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node2871 = (inp[15]) ? node2875 : node2872;
														assign node2872 = (inp[4]) ? 4'b1001 : 4'b0001;
														assign node2875 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node2878 = (inp[4]) ? node2916 : node2879;
											assign node2879 = (inp[15]) ? node2887 : node2880;
												assign node2880 = (inp[3]) ? 4'b1001 : node2881;
													assign node2881 = (inp[2]) ? node2883 : 4'b1001;
														assign node2883 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node2887 = (inp[2]) ? node2893 : node2888;
													assign node2888 = (inp[7]) ? node2890 : 4'b1101;
														assign node2890 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node2893 = (inp[12]) ? node2903 : node2894;
														assign node2894 = (inp[14]) ? node2896 : 4'b1101;
															assign node2896 = (inp[7]) ? node2900 : node2897;
																assign node2897 = (inp[3]) ? 4'b1001 : 4'b1101;
																assign node2900 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node2903 = (inp[14]) ? node2909 : node2904;
															assign node2904 = (inp[3]) ? node2906 : 4'b1001;
																assign node2906 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node2909 = (inp[3]) ? node2913 : node2910;
																assign node2910 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node2913 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node2916 = (inp[15]) ? node2922 : node2917;
												assign node2917 = (inp[3]) ? 4'b1101 : node2918;
													assign node2918 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node2922 = (inp[3]) ? 4'b1001 : node2923;
													assign node2923 = (inp[2]) ? 4'b1101 : 4'b1001;
						assign node2927 = (inp[15]) ? node3217 : node2928;
							assign node2928 = (inp[2]) ? 4'b1101 : node2929;
								assign node2929 = (inp[1]) ? node3063 : node2930;
									assign node2930 = (inp[14]) ? node2988 : node2931;
										assign node2931 = (inp[3]) ? node2957 : node2932;
											assign node2932 = (inp[4]) ? node2944 : node2933;
												assign node2933 = (inp[7]) ? 4'b1101 : node2934;
													assign node2934 = (inp[12]) ? node2938 : node2935;
														assign node2935 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node2938 = (inp[10]) ? 4'b0000 : node2939;
															assign node2939 = (inp[13]) ? 4'b0000 : 4'b1101;
												assign node2944 = (inp[13]) ? node2952 : node2945;
													assign node2945 = (inp[12]) ? node2947 : 4'b0000;
														assign node2947 = (inp[10]) ? 4'b0000 : node2948;
															assign node2948 = (inp[7]) ? 4'b1101 : 4'b1000;
													assign node2952 = (inp[10]) ? 4'b1000 : node2953;
														assign node2953 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2957 = (inp[13]) ? node2971 : node2958;
												assign node2958 = (inp[12]) ? node2964 : node2959;
													assign node2959 = (inp[7]) ? node2961 : 4'b0100;
														assign node2961 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2964 = (inp[10]) ? node2966 : 4'b1000;
														assign node2966 = (inp[7]) ? node2968 : 4'b0100;
															assign node2968 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node2971 = (inp[10]) ? node2983 : node2972;
													assign node2972 = (inp[12]) ? node2978 : node2973;
														assign node2973 = (inp[4]) ? 4'b1100 : node2974;
															assign node2974 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node2978 = (inp[4]) ? 4'b0100 : node2979;
															assign node2979 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node2983 = (inp[7]) ? node2985 : 4'b1100;
														assign node2985 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node2988 = (inp[11]) ? node3034 : node2989;
											assign node2989 = (inp[13]) ? node3013 : node2990;
												assign node2990 = (inp[12]) ? node3002 : node2991;
													assign node2991 = (inp[10]) ? node2995 : node2992;
														assign node2992 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node2995 = (inp[4]) ? 4'b0101 : node2996;
															assign node2996 = (inp[7]) ? node2998 : 4'b0001;
																assign node2998 = (inp[3]) ? 4'b0001 : 4'b1101;
													assign node3002 = (inp[3]) ? node3008 : node3003;
														assign node3003 = (inp[7]) ? 4'b1101 : node3004;
															assign node3004 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node3008 = (inp[4]) ? node3010 : 4'b1001;
															assign node3010 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node3013 = (inp[10]) ? node3023 : node3014;
													assign node3014 = (inp[3]) ? node3018 : node3015;
														assign node3015 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node3018 = (inp[7]) ? node3020 : 4'b0101;
															assign node3020 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node3023 = (inp[12]) ? node3029 : node3024;
														assign node3024 = (inp[3]) ? node3026 : 4'b1001;
															assign node3026 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node3029 = (inp[3]) ? node3031 : 4'b1101;
															assign node3031 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node3034 = (inp[13]) ? node3050 : node3035;
												assign node3035 = (inp[3]) ? node3041 : node3036;
													assign node3036 = (inp[7]) ? node3038 : 4'b0000;
														assign node3038 = (inp[4]) ? 4'b0000 : 4'b1101;
													assign node3041 = (inp[7]) ? node3047 : node3042;
														assign node3042 = (inp[10]) ? 4'b0100 : node3043;
															assign node3043 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node3047 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node3050 = (inp[3]) ? node3058 : node3051;
													assign node3051 = (inp[7]) ? node3055 : node3052;
														assign node3052 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3055 = (inp[4]) ? 4'b1000 : 4'b1101;
													assign node3058 = (inp[7]) ? node3060 : 4'b1100;
														assign node3060 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node3063 = (inp[14]) ? node3123 : node3064;
										assign node3064 = (inp[13]) ? node3100 : node3065;
											assign node3065 = (inp[12]) ? node3077 : node3066;
												assign node3066 = (inp[3]) ? node3072 : node3067;
													assign node3067 = (inp[4]) ? 4'b0001 : node3068;
														assign node3068 = (inp[7]) ? 4'b1101 : 4'b0001;
													assign node3072 = (inp[4]) ? 4'b0101 : node3073;
														assign node3073 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node3077 = (inp[10]) ? node3089 : node3078;
													assign node3078 = (inp[3]) ? node3084 : node3079;
														assign node3079 = (inp[7]) ? 4'b1101 : node3080;
															assign node3080 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node3084 = (inp[4]) ? node3086 : 4'b1001;
															assign node3086 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3089 = (inp[3]) ? node3095 : node3090;
														assign node3090 = (inp[7]) ? node3092 : 4'b0001;
															assign node3092 = (inp[4]) ? 4'b0001 : 4'b1101;
														assign node3095 = (inp[4]) ? 4'b0101 : node3096;
															assign node3096 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node3100 = (inp[3]) ? node3114 : node3101;
												assign node3101 = (inp[7]) ? node3107 : node3102;
													assign node3102 = (inp[10]) ? 4'b1001 : node3103;
														assign node3103 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3107 = (inp[4]) ? node3109 : 4'b1101;
														assign node3109 = (inp[10]) ? 4'b1001 : node3110;
															assign node3110 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node3114 = (inp[4]) ? node3118 : node3115;
													assign node3115 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3118 = (inp[12]) ? node3120 : 4'b1101;
														assign node3120 = (inp[10]) ? 4'b1101 : 4'b0101;
										assign node3123 = (inp[11]) ? node3173 : node3124;
											assign node3124 = (inp[3]) ? node3146 : node3125;
												assign node3125 = (inp[7]) ? node3137 : node3126;
													assign node3126 = (inp[10]) ? node3134 : node3127;
														assign node3127 = (inp[13]) ? node3131 : node3128;
															assign node3128 = (inp[4]) ? 4'b1000 : 4'b1101;
															assign node3131 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3134 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node3137 = (inp[4]) ? node3139 : 4'b1101;
														assign node3139 = (inp[13]) ? node3143 : node3140;
															assign node3140 = (inp[10]) ? 4'b0000 : 4'b1101;
															assign node3143 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3146 = (inp[4]) ? node3160 : node3147;
													assign node3147 = (inp[7]) ? node3153 : node3148;
														assign node3148 = (inp[13]) ? 4'b1100 : node3149;
															assign node3149 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node3153 = (inp[13]) ? 4'b1000 : node3154;
															assign node3154 = (inp[10]) ? 4'b0000 : node3155;
																assign node3155 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node3160 = (inp[13]) ? node3168 : node3161;
														assign node3161 = (inp[10]) ? 4'b0100 : node3162;
															assign node3162 = (inp[12]) ? node3164 : 4'b0100;
																assign node3164 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node3168 = (inp[12]) ? node3170 : 4'b1100;
															assign node3170 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node3173 = (inp[3]) ? node3195 : node3174;
												assign node3174 = (inp[4]) ? node3186 : node3175;
													assign node3175 = (inp[7]) ? 4'b1101 : node3176;
														assign node3176 = (inp[13]) ? node3180 : node3177;
															assign node3177 = (inp[10]) ? 4'b0001 : 4'b1101;
															assign node3180 = (inp[12]) ? node3182 : 4'b1001;
																assign node3182 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3186 = (inp[13]) ? node3190 : node3187;
														assign node3187 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node3190 = (inp[10]) ? 4'b1001 : node3191;
															assign node3191 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node3195 = (inp[13]) ? node3207 : node3196;
													assign node3196 = (inp[10]) ? 4'b0101 : node3197;
														assign node3197 = (inp[12]) ? node3201 : node3198;
															assign node3198 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node3201 = (inp[7]) ? 4'b1001 : node3202;
																assign node3202 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node3207 = (inp[12]) ? node3213 : node3208;
														assign node3208 = (inp[7]) ? node3210 : 4'b1101;
															assign node3210 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node3213 = (inp[10]) ? 4'b1101 : 4'b0101;
							assign node3217 = (inp[2]) ? 4'b1001 : node3218;
								assign node3218 = (inp[3]) ? node3220 : 4'b1001;
									assign node3220 = (inp[4]) ? node3276 : node3221;
										assign node3221 = (inp[7]) ? 4'b1001 : node3222;
											assign node3222 = (inp[13]) ? node3246 : node3223;
												assign node3223 = (inp[12]) ? node3237 : node3224;
													assign node3224 = (inp[14]) ? node3228 : node3225;
														assign node3225 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node3228 = (inp[10]) ? node3234 : node3229;
															assign node3229 = (inp[11]) ? node3231 : 4'b0000;
																assign node3231 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node3234 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node3237 = (inp[10]) ? node3239 : 4'b1001;
														assign node3239 = (inp[1]) ? 4'b0001 : node3240;
															assign node3240 = (inp[14]) ? node3242 : 4'b0000;
																assign node3242 = (inp[11]) ? 4'b0000 : 4'b1001;
												assign node3246 = (inp[12]) ? node3258 : node3247;
													assign node3247 = (inp[14]) ? node3249 : 4'b1001;
														assign node3249 = (inp[10]) ? node3251 : 4'b1001;
															assign node3251 = (inp[1]) ? node3255 : node3252;
																assign node3252 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node3255 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node3258 = (inp[10]) ? node3266 : node3259;
														assign node3259 = (inp[1]) ? node3261 : 4'b0000;
															assign node3261 = (inp[14]) ? node3263 : 4'b0001;
																assign node3263 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node3266 = (inp[1]) ? node3270 : node3267;
															assign node3267 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node3270 = (inp[14]) ? node3272 : 4'b1001;
																assign node3272 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node3276 = (inp[1]) ? node3310 : node3277;
											assign node3277 = (inp[14]) ? node3289 : node3278;
												assign node3278 = (inp[13]) ? node3284 : node3279;
													assign node3279 = (inp[10]) ? 4'b0000 : node3280;
														assign node3280 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node3284 = (inp[10]) ? 4'b1000 : node3285;
														assign node3285 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3289 = (inp[11]) ? node3301 : node3290;
													assign node3290 = (inp[13]) ? node3296 : node3291;
														assign node3291 = (inp[10]) ? node3293 : 4'b1001;
															assign node3293 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3296 = (inp[10]) ? node3298 : 4'b0001;
															assign node3298 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3301 = (inp[13]) ? node3305 : node3302;
														assign node3302 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node3305 = (inp[10]) ? 4'b1000 : node3306;
															assign node3306 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node3310 = (inp[14]) ? node3322 : node3311;
												assign node3311 = (inp[13]) ? node3317 : node3312;
													assign node3312 = (inp[10]) ? 4'b0001 : node3313;
														assign node3313 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node3317 = (inp[12]) ? node3319 : 4'b1001;
														assign node3319 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3322 = (inp[11]) ? node3336 : node3323;
													assign node3323 = (inp[13]) ? node3331 : node3324;
														assign node3324 = (inp[12]) ? node3326 : 4'b0000;
															assign node3326 = (inp[10]) ? 4'b0000 : node3327;
																assign node3327 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node3331 = (inp[12]) ? node3333 : 4'b1000;
															assign node3333 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3336 = (inp[13]) ? 4'b1001 : node3337;
														assign node3337 = (inp[12]) ? node3339 : 4'b0001;
															assign node3339 = (inp[10]) ? 4'b0001 : 4'b1001;
					assign node3344 = (inp[3]) ? node4680 : node3345;
						assign node3345 = (inp[1]) ? node4069 : node3346;
							assign node3346 = (inp[2]) ? node3774 : node3347;
								assign node3347 = (inp[0]) ? node3537 : node3348;
									assign node3348 = (inp[4]) ? node3442 : node3349;
										assign node3349 = (inp[11]) ? node3411 : node3350;
											assign node3350 = (inp[12]) ? node3382 : node3351;
												assign node3351 = (inp[14]) ? node3365 : node3352;
													assign node3352 = (inp[15]) ? node3358 : node3353;
														assign node3353 = (inp[10]) ? 4'b0001 : node3354;
															assign node3354 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node3358 = (inp[10]) ? node3362 : node3359;
															assign node3359 = (inp[13]) ? 4'b1101 : 4'b0001;
															assign node3362 = (inp[13]) ? 4'b0001 : 4'b1101;
													assign node3365 = (inp[13]) ? node3373 : node3366;
														assign node3366 = (inp[15]) ? node3370 : node3367;
															assign node3367 = (inp[10]) ? 4'b0001 : 4'b0100;
															assign node3370 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node3373 = (inp[10]) ? node3379 : node3374;
															assign node3374 = (inp[15]) ? 4'b1100 : node3375;
																assign node3375 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node3379 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node3382 = (inp[14]) ? node3402 : node3383;
													assign node3383 = (inp[15]) ? node3393 : node3384;
														assign node3384 = (inp[10]) ? node3388 : node3385;
															assign node3385 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node3388 = (inp[7]) ? 4'b1001 : node3389;
																assign node3389 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node3393 = (inp[13]) ? node3397 : node3394;
															assign node3394 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node3397 = (inp[7]) ? 4'b0101 : node3398;
																assign node3398 = (inp[10]) ? 4'b1001 : 4'b0101;
													assign node3402 = (inp[15]) ? node3408 : node3403;
														assign node3403 = (inp[13]) ? node3405 : 4'b1100;
															assign node3405 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node3408 = (inp[13]) ? 4'b0100 : 4'b1000;
											assign node3411 = (inp[10]) ? node3427 : node3412;
												assign node3412 = (inp[15]) ? node3420 : node3413;
													assign node3413 = (inp[13]) ? node3417 : node3414;
														assign node3414 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node3417 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3420 = (inp[13]) ? node3424 : node3421;
														assign node3421 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node3424 = (inp[7]) ? 4'b1100 : 4'b0001;
												assign node3427 = (inp[7]) ? node3435 : node3428;
													assign node3428 = (inp[15]) ? node3432 : node3429;
														assign node3429 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node3432 = (inp[13]) ? 4'b0001 : 4'b1100;
													assign node3435 = (inp[13]) ? node3439 : node3436;
														assign node3436 = (inp[15]) ? 4'b0100 : 4'b0001;
														assign node3439 = (inp[15]) ? 4'b0001 : 4'b0101;
										assign node3442 = (inp[15]) ? node3494 : node3443;
											assign node3443 = (inp[11]) ? node3471 : node3444;
												assign node3444 = (inp[10]) ? node3452 : node3445;
													assign node3445 = (inp[14]) ? node3447 : 4'b0000;
														assign node3447 = (inp[13]) ? 4'b0000 : node3448;
															assign node3448 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node3452 = (inp[12]) ? node3462 : node3453;
														assign node3453 = (inp[14]) ? node3459 : node3454;
															assign node3454 = (inp[7]) ? 4'b1000 : node3455;
																assign node3455 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node3459 = (inp[13]) ? 4'b1000 : 4'b0001;
														assign node3462 = (inp[13]) ? node3466 : node3463;
															assign node3463 = (inp[14]) ? 4'b0001 : 4'b0100;
															assign node3466 = (inp[7]) ? 4'b1000 : node3467;
																assign node3467 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3471 = (inp[13]) ? node3485 : node3472;
													assign node3472 = (inp[7]) ? node3480 : node3473;
														assign node3473 = (inp[12]) ? node3477 : node3474;
															assign node3474 = (inp[14]) ? 4'b1000 : 4'b0001;
															assign node3477 = (inp[10]) ? 4'b1100 : 4'b0000;
														assign node3480 = (inp[10]) ? 4'b1000 : node3481;
															assign node3481 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node3485 = (inp[10]) ? node3489 : node3486;
														assign node3486 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3489 = (inp[12]) ? node3491 : 4'b0000;
															assign node3491 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node3494 = (inp[13]) ? node3518 : node3495;
												assign node3495 = (inp[12]) ? node3505 : node3496;
													assign node3496 = (inp[10]) ? node3500 : node3497;
														assign node3497 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node3500 = (inp[7]) ? 4'b0101 : node3501;
															assign node3501 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node3505 = (inp[7]) ? node3513 : node3506;
														assign node3506 = (inp[10]) ? node3508 : 4'b0101;
															assign node3508 = (inp[11]) ? 4'b1000 : node3509;
																assign node3509 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node3513 = (inp[11]) ? node3515 : 4'b1001;
															assign node3515 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node3518 = (inp[11]) ? node3526 : node3519;
													assign node3519 = (inp[14]) ? node3521 : 4'b1000;
														assign node3521 = (inp[7]) ? 4'b1001 : node3522;
															assign node3522 = (inp[12]) ? 4'b0001 : 4'b1000;
													assign node3526 = (inp[10]) ? node3532 : node3527;
														assign node3527 = (inp[12]) ? 4'b1000 : node3528;
															assign node3528 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node3532 = (inp[12]) ? node3534 : 4'b0001;
															assign node3534 = (inp[7]) ? 4'b0100 : 4'b1001;
									assign node3537 = (inp[7]) ? node3643 : node3538;
										assign node3538 = (inp[15]) ? node3600 : node3539;
											assign node3539 = (inp[11]) ? node3573 : node3540;
												assign node3540 = (inp[13]) ? node3556 : node3541;
													assign node3541 = (inp[4]) ? node3549 : node3542;
														assign node3542 = (inp[10]) ? node3546 : node3543;
															assign node3543 = (inp[12]) ? 4'b1101 : 4'b0000;
															assign node3546 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3549 = (inp[12]) ? node3553 : node3550;
															assign node3550 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node3553 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node3556 = (inp[12]) ? node3568 : node3557;
														assign node3557 = (inp[14]) ? node3561 : node3558;
															assign node3558 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node3561 = (inp[10]) ? node3565 : node3562;
																assign node3562 = (inp[4]) ? 4'b1000 : 4'b0000;
																assign node3565 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node3568 = (inp[10]) ? 4'b0000 : node3569;
															assign node3569 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node3573 = (inp[13]) ? node3587 : node3574;
													assign node3574 = (inp[12]) ? node3582 : node3575;
														assign node3575 = (inp[10]) ? node3579 : node3576;
															assign node3576 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node3579 = (inp[4]) ? 4'b0000 : 4'b1001;
														assign node3582 = (inp[4]) ? node3584 : 4'b1100;
															assign node3584 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node3587 = (inp[4]) ? node3595 : node3588;
														assign node3588 = (inp[12]) ? node3592 : node3589;
															assign node3589 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node3592 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node3595 = (inp[10]) ? node3597 : 4'b1000;
															assign node3597 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node3600 = (inp[4]) ? node3626 : node3601;
												assign node3601 = (inp[11]) ? node3617 : node3602;
													assign node3602 = (inp[14]) ? node3606 : node3603;
														assign node3603 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node3606 = (inp[13]) ? node3612 : node3607;
															assign node3607 = (inp[10]) ? node3609 : 4'b1001;
																assign node3609 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node3612 = (inp[10]) ? node3614 : 4'b0101;
																assign node3614 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node3617 = (inp[13]) ? node3621 : node3618;
														assign node3618 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node3621 = (inp[10]) ? 4'b1100 : node3622;
															assign node3622 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node3626 = (inp[11]) ? node3636 : node3627;
													assign node3627 = (inp[12]) ? node3631 : node3628;
														assign node3628 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3631 = (inp[13]) ? 4'b1000 : node3632;
															assign node3632 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node3636 = (inp[10]) ? node3640 : node3637;
														assign node3637 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node3640 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node3643 = (inp[14]) ? node3705 : node3644;
											assign node3644 = (inp[13]) ? node3672 : node3645;
												assign node3645 = (inp[12]) ? node3657 : node3646;
													assign node3646 = (inp[15]) ? node3654 : node3647;
														assign node3647 = (inp[4]) ? node3649 : 4'b0100;
															assign node3649 = (inp[11]) ? node3651 : 4'b0000;
																assign node3651 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node3654 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node3657 = (inp[10]) ? node3665 : node3658;
														assign node3658 = (inp[4]) ? node3662 : node3659;
															assign node3659 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node3662 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node3665 = (inp[15]) ? node3669 : node3666;
															assign node3666 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node3669 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node3672 = (inp[12]) ? node3686 : node3673;
													assign node3673 = (inp[10]) ? node3681 : node3674;
														assign node3674 = (inp[15]) ? node3678 : node3675;
															assign node3675 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3678 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node3681 = (inp[15]) ? node3683 : 4'b1001;
															assign node3683 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node3686 = (inp[10]) ? node3694 : node3687;
														assign node3687 = (inp[4]) ? node3691 : node3688;
															assign node3688 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3691 = (inp[15]) ? 4'b0100 : 4'b1000;
														assign node3694 = (inp[4]) ? node3698 : node3695;
															assign node3695 = (inp[15]) ? 4'b1000 : 4'b0000;
															assign node3698 = (inp[11]) ? node3702 : node3699;
																assign node3699 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node3702 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node3705 = (inp[11]) ? node3741 : node3706;
												assign node3706 = (inp[15]) ? node3726 : node3707;
													assign node3707 = (inp[4]) ? node3719 : node3708;
														assign node3708 = (inp[13]) ? node3714 : node3709;
															assign node3709 = (inp[10]) ? node3711 : 4'b1101;
																assign node3711 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node3714 = (inp[12]) ? 4'b0000 : node3715;
																assign node3715 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3719 = (inp[12]) ? node3723 : node3720;
															assign node3720 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node3723 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node3726 = (inp[13]) ? node3732 : node3727;
														assign node3727 = (inp[12]) ? 4'b1001 : node3728;
															assign node3728 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node3732 = (inp[10]) ? node3738 : node3733;
															assign node3733 = (inp[12]) ? node3735 : 4'b0000;
																assign node3735 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node3738 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node3741 = (inp[4]) ? node3759 : node3742;
													assign node3742 = (inp[15]) ? node3750 : node3743;
														assign node3743 = (inp[12]) ? 4'b0100 : node3744;
															assign node3744 = (inp[13]) ? node3746 : 4'b0100;
																assign node3746 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node3750 = (inp[10]) ? node3756 : node3751;
															assign node3751 = (inp[13]) ? node3753 : 4'b1000;
																assign node3753 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node3756 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node3759 = (inp[15]) ? node3769 : node3760;
														assign node3760 = (inp[10]) ? node3764 : node3761;
															assign node3761 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3764 = (inp[13]) ? node3766 : 4'b0001;
																assign node3766 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3769 = (inp[13]) ? node3771 : 4'b0100;
															assign node3771 = (inp[10]) ? 4'b0001 : 4'b0100;
								assign node3774 = (inp[0]) ? node4008 : node3775;
									assign node3775 = (inp[4]) ? node3905 : node3776;
										assign node3776 = (inp[11]) ? node3856 : node3777;
											assign node3777 = (inp[14]) ? node3815 : node3778;
												assign node3778 = (inp[15]) ? node3794 : node3779;
													assign node3779 = (inp[13]) ? node3789 : node3780;
														assign node3780 = (inp[7]) ? node3786 : node3781;
															assign node3781 = (inp[12]) ? 4'b1100 : node3782;
																assign node3782 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node3786 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node3789 = (inp[12]) ? 4'b0001 : node3790;
															assign node3790 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node3794 = (inp[12]) ? node3806 : node3795;
														assign node3795 = (inp[10]) ? node3801 : node3796;
															assign node3796 = (inp[7]) ? node3798 : 4'b0100;
																assign node3798 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node3801 = (inp[7]) ? 4'b1100 : node3802;
																assign node3802 = (inp[13]) ? 4'b0001 : 4'b1100;
														assign node3806 = (inp[10]) ? node3812 : node3807;
															assign node3807 = (inp[13]) ? node3809 : 4'b1000;
																assign node3809 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node3812 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node3815 = (inp[13]) ? node3841 : node3816;
													assign node3816 = (inp[15]) ? node3828 : node3817;
														assign node3817 = (inp[7]) ? node3821 : node3818;
															assign node3818 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node3821 = (inp[12]) ? node3825 : node3822;
																assign node3822 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node3825 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node3828 = (inp[7]) ? node3834 : node3829;
															assign node3829 = (inp[12]) ? 4'b1000 : node3830;
																assign node3830 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node3834 = (inp[12]) ? node3838 : node3835;
																assign node3835 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node3838 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node3841 = (inp[10]) ? node3847 : node3842;
														assign node3842 = (inp[7]) ? 4'b1000 : node3843;
															assign node3843 = (inp[15]) ? 4'b0100 : 4'b1000;
														assign node3847 = (inp[15]) ? node3851 : node3848;
															assign node3848 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node3851 = (inp[7]) ? node3853 : 4'b0000;
																assign node3853 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node3856 = (inp[15]) ? node3880 : node3857;
												assign node3857 = (inp[13]) ? node3871 : node3858;
													assign node3858 = (inp[7]) ? node3864 : node3859;
														assign node3859 = (inp[10]) ? node3861 : 4'b0000;
															assign node3861 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node3864 = (inp[10]) ? node3868 : node3865;
															assign node3865 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node3868 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node3871 = (inp[10]) ? node3873 : 4'b1000;
														assign node3873 = (inp[12]) ? node3877 : node3874;
															assign node3874 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node3877 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node3880 = (inp[7]) ? node3894 : node3881;
													assign node3881 = (inp[10]) ? node3887 : node3882;
														assign node3882 = (inp[12]) ? node3884 : 4'b0101;
															assign node3884 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node3887 = (inp[13]) ? node3891 : node3888;
															assign node3888 = (inp[14]) ? 4'b0101 : 4'b1101;
															assign node3891 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node3894 = (inp[13]) ? node3900 : node3895;
														assign node3895 = (inp[10]) ? node3897 : 4'b0001;
															assign node3897 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3900 = (inp[10]) ? 4'b0101 : node3901;
															assign node3901 = (inp[12]) ? 4'b1001 : 4'b0101;
										assign node3905 = (inp[11]) ? node3973 : node3906;
											assign node3906 = (inp[12]) ? node3940 : node3907;
												assign node3907 = (inp[15]) ? node3925 : node3908;
													assign node3908 = (inp[13]) ? node3914 : node3909;
														assign node3909 = (inp[7]) ? node3911 : 4'b0001;
															assign node3911 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node3914 = (inp[14]) ? node3920 : node3915;
															assign node3915 = (inp[10]) ? 4'b0000 : node3916;
																assign node3916 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node3920 = (inp[7]) ? node3922 : 4'b0101;
																assign node3922 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node3925 = (inp[14]) ? node3935 : node3926;
														assign node3926 = (inp[10]) ? node3932 : node3927;
															assign node3927 = (inp[7]) ? node3929 : 4'b0001;
																assign node3929 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node3932 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node3935 = (inp[13]) ? 4'b0001 : node3936;
															assign node3936 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node3940 = (inp[15]) ? node3954 : node3941;
													assign node3941 = (inp[13]) ? node3947 : node3942;
														assign node3942 = (inp[14]) ? 4'b1000 : node3943;
															assign node3943 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node3947 = (inp[14]) ? 4'b1001 : node3948;
															assign node3948 = (inp[10]) ? node3950 : 4'b1001;
																assign node3950 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3954 = (inp[14]) ? node3964 : node3955;
														assign node3955 = (inp[13]) ? node3957 : 4'b1001;
															assign node3957 = (inp[7]) ? node3961 : node3958;
																assign node3958 = (inp[10]) ? 4'b1001 : 4'b0101;
																assign node3961 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node3964 = (inp[13]) ? node3968 : node3965;
															assign node3965 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node3968 = (inp[7]) ? 4'b0100 : node3969;
																assign node3969 = (inp[10]) ? 4'b1001 : 4'b0100;
											assign node3973 = (inp[15]) ? node3993 : node3974;
												assign node3974 = (inp[10]) ? node3990 : node3975;
													assign node3975 = (inp[12]) ? node3983 : node3976;
														assign node3976 = (inp[13]) ? node3980 : node3977;
															assign node3977 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node3980 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node3983 = (inp[13]) ? node3987 : node3984;
															assign node3984 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node3987 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3990 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node3993 = (inp[13]) ? node4003 : node3994;
													assign node3994 = (inp[12]) ? node4000 : node3995;
														assign node3995 = (inp[10]) ? node3997 : 4'b0000;
															assign node3997 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4000 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node4003 = (inp[7]) ? node4005 : 4'b0001;
														assign node4005 = (inp[10]) ? 4'b0001 : 4'b1000;
									assign node4008 = (inp[15]) ? 4'b1001 : node4009;
										assign node4009 = (inp[4]) ? node4031 : node4010;
											assign node4010 = (inp[7]) ? 4'b1101 : node4011;
												assign node4011 = (inp[11]) ? node4023 : node4012;
													assign node4012 = (inp[14]) ? node4018 : node4013;
														assign node4013 = (inp[13]) ? 4'b1000 : node4014;
															assign node4014 = (inp[12]) ? 4'b1101 : 4'b0000;
														assign node4018 = (inp[13]) ? 4'b0001 : node4019;
															assign node4019 = (inp[10]) ? 4'b0001 : 4'b1101;
													assign node4023 = (inp[13]) ? node4025 : 4'b0000;
														assign node4025 = (inp[10]) ? 4'b1000 : node4026;
															assign node4026 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node4031 = (inp[14]) ? node4045 : node4032;
												assign node4032 = (inp[13]) ? node4040 : node4033;
													assign node4033 = (inp[10]) ? 4'b0000 : node4034;
														assign node4034 = (inp[12]) ? node4036 : 4'b0000;
															assign node4036 = (inp[7]) ? 4'b1101 : 4'b1000;
													assign node4040 = (inp[10]) ? 4'b1000 : node4041;
														assign node4041 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4045 = (inp[11]) ? node4057 : node4046;
													assign node4046 = (inp[13]) ? node4052 : node4047;
														assign node4047 = (inp[12]) ? node4049 : 4'b0001;
															assign node4049 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node4052 = (inp[12]) ? 4'b0001 : node4053;
															assign node4053 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node4057 = (inp[13]) ? node4063 : node4058;
														assign node4058 = (inp[12]) ? node4060 : 4'b0000;
															assign node4060 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node4063 = (inp[12]) ? node4065 : 4'b1000;
															assign node4065 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node4069 = (inp[11]) ? node4423 : node4070;
								assign node4070 = (inp[2]) ? node4288 : node4071;
									assign node4071 = (inp[4]) ? node4195 : node4072;
										assign node4072 = (inp[0]) ? node4140 : node4073;
											assign node4073 = (inp[12]) ? node4103 : node4074;
												assign node4074 = (inp[14]) ? node4094 : node4075;
													assign node4075 = (inp[13]) ? node4085 : node4076;
														assign node4076 = (inp[10]) ? 4'b0100 : node4077;
															assign node4077 = (inp[7]) ? node4081 : node4078;
																assign node4078 = (inp[15]) ? 4'b1100 : 4'b1001;
																assign node4081 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node4085 = (inp[7]) ? node4087 : 4'b1001;
															assign node4087 = (inp[10]) ? node4091 : node4088;
																assign node4088 = (inp[15]) ? 4'b0100 : 4'b1001;
																assign node4091 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node4094 = (inp[13]) ? node4098 : node4095;
														assign node4095 = (inp[15]) ? 4'b0101 : 4'b1001;
														assign node4098 = (inp[7]) ? 4'b1101 : node4099;
															assign node4099 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node4103 = (inp[14]) ? node4121 : node4104;
													assign node4104 = (inp[15]) ? node4112 : node4105;
														assign node4105 = (inp[7]) ? node4107 : 4'b0001;
															assign node4107 = (inp[13]) ? 4'b0001 : node4108;
																assign node4108 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node4112 = (inp[13]) ? node4118 : node4113;
															assign node4113 = (inp[10]) ? 4'b0100 : node4114;
																assign node4114 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node4118 = (inp[7]) ? 4'b1100 : 4'b0001;
													assign node4121 = (inp[10]) ? node4131 : node4122;
														assign node4122 = (inp[15]) ? node4124 : 4'b0101;
															assign node4124 = (inp[7]) ? node4128 : node4125;
																assign node4125 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node4128 = (inp[13]) ? 4'b1101 : 4'b0001;
														assign node4131 = (inp[15]) ? node4135 : node4132;
															assign node4132 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node4135 = (inp[13]) ? 4'b0001 : node4136;
																assign node4136 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node4140 = (inp[14]) ? node4168 : node4141;
												assign node4141 = (inp[15]) ? node4151 : node4142;
													assign node4142 = (inp[10]) ? node4146 : node4143;
														assign node4143 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node4146 = (inp[7]) ? node4148 : 4'b1000;
															assign node4148 = (inp[13]) ? 4'b1000 : 4'b0101;
													assign node4151 = (inp[7]) ? node4159 : node4152;
														assign node4152 = (inp[13]) ? 4'b1101 : node4153;
															assign node4153 = (inp[10]) ? 4'b0101 : node4154;
																assign node4154 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node4159 = (inp[13]) ? node4165 : node4160;
															assign node4160 = (inp[12]) ? node4162 : 4'b0001;
																assign node4162 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node4165 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4168 = (inp[7]) ? node4180 : node4169;
													assign node4169 = (inp[15]) ? node4173 : node4170;
														assign node4170 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node4173 = (inp[13]) ? node4175 : 4'b0100;
															assign node4175 = (inp[10]) ? 4'b1100 : node4176;
																assign node4176 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node4180 = (inp[13]) ? node4188 : node4181;
														assign node4181 = (inp[10]) ? node4185 : node4182;
															assign node4182 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node4185 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node4188 = (inp[10]) ? 4'b1000 : node4189;
															assign node4189 = (inp[15]) ? node4191 : 4'b0000;
																assign node4191 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node4195 = (inp[10]) ? node4239 : node4196;
											assign node4196 = (inp[15]) ? node4216 : node4197;
												assign node4197 = (inp[0]) ? node4207 : node4198;
													assign node4198 = (inp[13]) ? node4202 : node4199;
														assign node4199 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node4202 = (inp[12]) ? 4'b1000 : node4203;
															assign node4203 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node4207 = (inp[14]) ? node4211 : node4208;
														assign node4208 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4211 = (inp[12]) ? 4'b0100 : node4212;
															assign node4212 = (inp[13]) ? 4'b1001 : 4'b0100;
												assign node4216 = (inp[7]) ? node4224 : node4217;
													assign node4217 = (inp[0]) ? 4'b0000 : node4218;
														assign node4218 = (inp[12]) ? node4220 : 4'b0000;
															assign node4220 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4224 = (inp[13]) ? node4234 : node4225;
														assign node4225 = (inp[0]) ? node4229 : node4226;
															assign node4226 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node4229 = (inp[12]) ? 4'b1001 : node4230;
																assign node4230 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node4234 = (inp[14]) ? 4'b0000 : node4235;
															assign node4235 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node4239 = (inp[0]) ? node4271 : node4240;
												assign node4240 = (inp[7]) ? node4256 : node4241;
													assign node4241 = (inp[12]) ? node4247 : node4242;
														assign node4242 = (inp[15]) ? node4244 : 4'b1000;
															assign node4244 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node4247 = (inp[15]) ? node4251 : node4248;
															assign node4248 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node4251 = (inp[13]) ? 4'b0000 : node4252;
																assign node4252 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node4256 = (inp[13]) ? node4266 : node4257;
														assign node4257 = (inp[14]) ? node4263 : node4258;
															assign node4258 = (inp[12]) ? node4260 : 4'b0101;
																assign node4260 = (inp[15]) ? 4'b0101 : 4'b1001;
															assign node4263 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node4266 = (inp[15]) ? node4268 : 4'b0001;
															assign node4268 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4271 = (inp[15]) ? node4283 : node4272;
													assign node4272 = (inp[7]) ? 4'b1000 : node4273;
														assign node4273 = (inp[14]) ? node4277 : node4274;
															assign node4274 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node4277 = (inp[12]) ? 4'b0001 : node4278;
																assign node4278 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node4283 = (inp[7]) ? node4285 : 4'b1000;
														assign node4285 = (inp[13]) ? 4'b1000 : 4'b0101;
									assign node4288 = (inp[0]) ? node4384 : node4289;
										assign node4289 = (inp[4]) ? node4327 : node4290;
											assign node4290 = (inp[10]) ? node4306 : node4291;
												assign node4291 = (inp[15]) ? node4301 : node4292;
													assign node4292 = (inp[13]) ? node4298 : node4293;
														assign node4293 = (inp[7]) ? 4'b0100 : node4294;
															assign node4294 = (inp[12]) ? 4'b0001 : 4'b1000;
														assign node4298 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node4301 = (inp[7]) ? node4303 : 4'b0100;
														assign node4303 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node4306 = (inp[15]) ? node4320 : node4307;
													assign node4307 = (inp[14]) ? node4311 : node4308;
														assign node4308 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node4311 = (inp[13]) ? node4315 : node4312;
															assign node4312 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node4315 = (inp[12]) ? node4317 : 4'b1101;
																assign node4317 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4320 = (inp[13]) ? node4324 : node4321;
														assign node4321 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node4324 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node4327 = (inp[12]) ? node4359 : node4328;
												assign node4328 = (inp[10]) ? node4348 : node4329;
													assign node4329 = (inp[7]) ? node4339 : node4330;
														assign node4330 = (inp[13]) ? node4334 : node4331;
															assign node4331 = (inp[14]) ? 4'b0001 : 4'b1001;
															assign node4334 = (inp[15]) ? 4'b1001 : node4335;
																assign node4335 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4339 = (inp[14]) ? 4'b0101 : node4340;
															assign node4340 = (inp[13]) ? node4344 : node4341;
																assign node4341 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node4344 = (inp[15]) ? 4'b0100 : 4'b1001;
													assign node4348 = (inp[13]) ? node4354 : node4349;
														assign node4349 = (inp[15]) ? node4351 : 4'b1001;
															assign node4351 = (inp[14]) ? 4'b0101 : 4'b0000;
														assign node4354 = (inp[14]) ? node4356 : 4'b1001;
															assign node4356 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node4359 = (inp[15]) ? node4363 : node4360;
													assign node4360 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node4363 = (inp[14]) ? node4373 : node4364;
														assign node4364 = (inp[13]) ? node4368 : node4365;
															assign node4365 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node4368 = (inp[7]) ? node4370 : 4'b0001;
																assign node4370 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node4373 = (inp[7]) ? node4379 : node4374;
															assign node4374 = (inp[10]) ? node4376 : 4'b0001;
																assign node4376 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node4379 = (inp[13]) ? 4'b1001 : node4380;
																assign node4380 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node4384 = (inp[15]) ? 4'b1001 : node4385;
											assign node4385 = (inp[4]) ? node4401 : node4386;
												assign node4386 = (inp[7]) ? 4'b1101 : node4387;
													assign node4387 = (inp[14]) ? node4391 : node4388;
														assign node4388 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node4391 = (inp[13]) ? node4395 : node4392;
															assign node4392 = (inp[12]) ? 4'b1101 : 4'b0000;
															assign node4395 = (inp[10]) ? 4'b1000 : node4396;
																assign node4396 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4401 = (inp[14]) ? node4413 : node4402;
													assign node4402 = (inp[13]) ? node4408 : node4403;
														assign node4403 = (inp[12]) ? node4405 : 4'b0001;
															assign node4405 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node4408 = (inp[10]) ? 4'b1001 : node4409;
															assign node4409 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4413 = (inp[13]) ? node4417 : node4414;
														assign node4414 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node4417 = (inp[10]) ? 4'b1000 : node4418;
															assign node4418 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node4423 = (inp[13]) ? node4585 : node4424;
									assign node4424 = (inp[2]) ? node4526 : node4425;
										assign node4425 = (inp[0]) ? node4463 : node4426;
											assign node4426 = (inp[15]) ? node4446 : node4427;
												assign node4427 = (inp[7]) ? node4435 : node4428;
													assign node4428 = (inp[4]) ? node4430 : 4'b1001;
														assign node4430 = (inp[10]) ? 4'b1001 : node4431;
															assign node4431 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node4435 = (inp[4]) ? node4441 : node4436;
														assign node4436 = (inp[10]) ? 4'b1001 : node4437;
															assign node4437 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4441 = (inp[10]) ? 4'b0101 : node4442;
															assign node4442 = (inp[14]) ? 4'b0001 : 4'b1001;
												assign node4446 = (inp[10]) ? node4460 : node4447;
													assign node4447 = (inp[7]) ? node4455 : node4448;
														assign node4448 = (inp[4]) ? node4452 : node4449;
															assign node4449 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node4452 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node4455 = (inp[12]) ? node4457 : 4'b1001;
															assign node4457 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node4460 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node4463 = (inp[12]) ? node4501 : node4464;
												assign node4464 = (inp[15]) ? node4488 : node4465;
													assign node4465 = (inp[10]) ? node4479 : node4466;
														assign node4466 = (inp[14]) ? node4474 : node4467;
															assign node4467 = (inp[7]) ? node4471 : node4468;
																assign node4468 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node4471 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node4474 = (inp[7]) ? 4'b0001 : node4475;
																assign node4475 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node4479 = (inp[14]) ? node4483 : node4480;
															assign node4480 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node4483 = (inp[4]) ? node4485 : 4'b1001;
																assign node4485 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node4488 = (inp[10]) ? node4496 : node4489;
														assign node4489 = (inp[7]) ? node4493 : node4490;
															assign node4490 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node4493 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node4496 = (inp[7]) ? node4498 : 4'b0101;
															assign node4498 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node4501 = (inp[15]) ? node4517 : node4502;
													assign node4502 = (inp[4]) ? node4510 : node4503;
														assign node4503 = (inp[7]) ? node4507 : node4504;
															assign node4504 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4507 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node4510 = (inp[10]) ? node4514 : node4511;
															assign node4511 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node4514 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node4517 = (inp[10]) ? node4519 : 4'b1001;
														assign node4519 = (inp[4]) ? node4523 : node4520;
															assign node4520 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node4523 = (inp[7]) ? 4'b0101 : 4'b1001;
										assign node4526 = (inp[15]) ? node4560 : node4527;
											assign node4527 = (inp[7]) ? node4541 : node4528;
												assign node4528 = (inp[0]) ? node4536 : node4529;
													assign node4529 = (inp[4]) ? 4'b1001 : node4530;
														assign node4530 = (inp[10]) ? 4'b0001 : node4531;
															assign node4531 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4536 = (inp[10]) ? 4'b0001 : node4537;
														assign node4537 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node4541 = (inp[10]) ? node4553 : node4542;
													assign node4542 = (inp[0]) ? node4548 : node4543;
														assign node4543 = (inp[4]) ? node4545 : 4'b0101;
															assign node4545 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4548 = (inp[12]) ? 4'b1101 : node4549;
															assign node4549 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node4553 = (inp[4]) ? node4557 : node4554;
														assign node4554 = (inp[0]) ? 4'b1101 : 4'b0001;
														assign node4557 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node4560 = (inp[0]) ? 4'b1001 : node4561;
												assign node4561 = (inp[7]) ? node4571 : node4562;
													assign node4562 = (inp[4]) ? node4566 : node4563;
														assign node4563 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node4566 = (inp[10]) ? 4'b0101 : node4567;
															assign node4567 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4571 = (inp[12]) ? node4579 : node4572;
														assign node4572 = (inp[10]) ? node4576 : node4573;
															assign node4573 = (inp[4]) ? 4'b1001 : 4'b0001;
															assign node4576 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node4579 = (inp[4]) ? 4'b0001 : node4580;
															assign node4580 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node4585 = (inp[10]) ? node4657 : node4586;
										assign node4586 = (inp[4]) ? node4620 : node4587;
											assign node4587 = (inp[0]) ? node4607 : node4588;
												assign node4588 = (inp[2]) ? node4598 : node4589;
													assign node4589 = (inp[15]) ? node4593 : node4590;
														assign node4590 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node4593 = (inp[7]) ? node4595 : 4'b1001;
															assign node4595 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node4598 = (inp[15]) ? node4602 : node4599;
														assign node4599 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node4602 = (inp[7]) ? 4'b0101 : node4603;
															assign node4603 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node4607 = (inp[2]) ? node4615 : node4608;
													assign node4608 = (inp[15]) ? node4610 : 4'b0001;
														assign node4610 = (inp[12]) ? node4612 : 4'b1001;
															assign node4612 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node4615 = (inp[15]) ? 4'b1001 : node4616;
														assign node4616 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node4620 = (inp[2]) ? node4638 : node4621;
												assign node4621 = (inp[15]) ? node4631 : node4622;
													assign node4622 = (inp[12]) ? node4624 : 4'b0001;
														assign node4624 = (inp[0]) ? node4628 : node4625;
															assign node4625 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node4628 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node4631 = (inp[12]) ? 4'b0001 : node4632;
														assign node4632 = (inp[7]) ? node4634 : 4'b0001;
															assign node4634 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node4638 = (inp[7]) ? node4644 : node4639;
													assign node4639 = (inp[12]) ? node4641 : 4'b1001;
														assign node4641 = (inp[15]) ? 4'b1001 : 4'b0001;
													assign node4644 = (inp[12]) ? node4652 : node4645;
														assign node4645 = (inp[14]) ? 4'b0101 : node4646;
															assign node4646 = (inp[0]) ? 4'b1001 : node4647;
																assign node4647 = (inp[15]) ? 4'b0101 : 4'b1001;
														assign node4652 = (inp[0]) ? node4654 : 4'b1001;
															assign node4654 = (inp[15]) ? 4'b1001 : 4'b0001;
										assign node4657 = (inp[4]) ? 4'b1001 : node4658;
											assign node4658 = (inp[7]) ? node4666 : node4659;
												assign node4659 = (inp[2]) ? node4661 : 4'b1001;
													assign node4661 = (inp[15]) ? 4'b1001 : node4662;
														assign node4662 = (inp[0]) ? 4'b1001 : 4'b1101;
												assign node4666 = (inp[15]) ? node4674 : node4667;
													assign node4667 = (inp[2]) ? node4671 : node4668;
														assign node4668 = (inp[0]) ? 4'b1001 : 4'b1101;
														assign node4671 = (inp[0]) ? 4'b1101 : 4'b1001;
													assign node4674 = (inp[2]) ? node4676 : 4'b1001;
														assign node4676 = (inp[0]) ? 4'b1001 : 4'b1101;
						assign node4680 = (inp[4]) ? node5460 : node4681;
							assign node4681 = (inp[1]) ? node5103 : node4682;
								assign node4682 = (inp[15]) ? node4920 : node4683;
									assign node4683 = (inp[2]) ? node4791 : node4684;
										assign node4684 = (inp[13]) ? node4736 : node4685;
											assign node4685 = (inp[7]) ? node4705 : node4686;
												assign node4686 = (inp[0]) ? node4698 : node4687;
													assign node4687 = (inp[10]) ? node4691 : node4688;
														assign node4688 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node4691 = (inp[11]) ? 4'b0000 : node4692;
															assign node4692 = (inp[14]) ? node4694 : 4'b1000;
																assign node4694 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4698 = (inp[11]) ? 4'b0001 : node4699;
														assign node4699 = (inp[12]) ? node4701 : 4'b0001;
															assign node4701 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node4705 = (inp[14]) ? node4719 : node4706;
													assign node4706 = (inp[11]) ? node4712 : node4707;
														assign node4707 = (inp[12]) ? node4709 : 4'b0001;
															assign node4709 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node4712 = (inp[10]) ? node4716 : node4713;
															assign node4713 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node4716 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4719 = (inp[10]) ? node4729 : node4720;
														assign node4720 = (inp[11]) ? node4726 : node4721;
															assign node4721 = (inp[12]) ? node4723 : 4'b0000;
																assign node4723 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node4726 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node4729 = (inp[0]) ? node4733 : node4730;
															assign node4730 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node4733 = (inp[11]) ? 4'b0001 : 4'b1000;
											assign node4736 = (inp[7]) ? node4766 : node4737;
												assign node4737 = (inp[0]) ? node4753 : node4738;
													assign node4738 = (inp[10]) ? node4742 : node4739;
														assign node4739 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node4742 = (inp[12]) ? node4748 : node4743;
															assign node4743 = (inp[11]) ? 4'b0001 : node4744;
																assign node4744 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node4748 = (inp[11]) ? 4'b0000 : node4749;
																assign node4749 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node4753 = (inp[12]) ? node4757 : node4754;
														assign node4754 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node4757 = (inp[10]) ? node4763 : node4758;
															assign node4758 = (inp[11]) ? 4'b1000 : node4759;
																assign node4759 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node4763 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4766 = (inp[11]) ? node4780 : node4767;
													assign node4767 = (inp[0]) ? node4775 : node4768;
														assign node4768 = (inp[10]) ? node4772 : node4769;
															assign node4769 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node4772 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4775 = (inp[12]) ? 4'b1001 : node4776;
															assign node4776 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4780 = (inp[12]) ? node4786 : node4781;
														assign node4781 = (inp[10]) ? 4'b0000 : node4782;
															assign node4782 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4786 = (inp[10]) ? 4'b0000 : node4787;
															assign node4787 = (inp[0]) ? 4'b0001 : 4'b1001;
										assign node4791 = (inp[11]) ? node4867 : node4792;
											assign node4792 = (inp[14]) ? node4830 : node4793;
												assign node4793 = (inp[12]) ? node4811 : node4794;
													assign node4794 = (inp[7]) ? node4806 : node4795;
														assign node4795 = (inp[10]) ? node4801 : node4796;
															assign node4796 = (inp[13]) ? node4798 : 4'b0000;
																assign node4798 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4801 = (inp[13]) ? node4803 : 4'b0001;
																assign node4803 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node4806 = (inp[13]) ? 4'b0000 : node4807;
															assign node4807 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node4811 = (inp[13]) ? node4825 : node4812;
														assign node4812 = (inp[7]) ? node4820 : node4813;
															assign node4813 = (inp[0]) ? node4817 : node4814;
																assign node4814 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node4817 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node4820 = (inp[0]) ? node4822 : 4'b1000;
																assign node4822 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node4825 = (inp[10]) ? 4'b0000 : node4826;
															assign node4826 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node4830 = (inp[7]) ? node4848 : node4831;
													assign node4831 = (inp[13]) ? node4841 : node4832;
														assign node4832 = (inp[10]) ? node4834 : 4'b0000;
															assign node4834 = (inp[12]) ? node4838 : node4835;
																assign node4835 = (inp[0]) ? 4'b1000 : 4'b0000;
																assign node4838 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node4841 = (inp[0]) ? node4845 : node4842;
															assign node4842 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4845 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4848 = (inp[13]) ? node4858 : node4849;
														assign node4849 = (inp[10]) ? node4855 : node4850;
															assign node4850 = (inp[12]) ? 4'b1001 : node4851;
																assign node4851 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node4855 = (inp[0]) ? 4'b0001 : 4'b1000;
														assign node4858 = (inp[12]) ? node4864 : node4859;
															assign node4859 = (inp[0]) ? node4861 : 4'b1000;
																assign node4861 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node4864 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node4867 = (inp[7]) ? node4897 : node4868;
												assign node4868 = (inp[10]) ? node4878 : node4869;
													assign node4869 = (inp[12]) ? node4873 : node4870;
														assign node4870 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node4873 = (inp[13]) ? 4'b1001 : node4874;
															assign node4874 = (inp[0]) ? 4'b1000 : 4'b0001;
													assign node4878 = (inp[12]) ? node4892 : node4879;
														assign node4879 = (inp[14]) ? node4885 : node4880;
															assign node4880 = (inp[13]) ? 4'b1000 : node4881;
																assign node4881 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node4885 = (inp[0]) ? node4889 : node4886;
																assign node4886 = (inp[13]) ? 4'b1001 : 4'b1000;
																assign node4889 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node4892 = (inp[0]) ? node4894 : 4'b0000;
															assign node4894 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node4897 = (inp[10]) ? node4909 : node4898;
													assign node4898 = (inp[13]) ? node4904 : node4899;
														assign node4899 = (inp[12]) ? 4'b1000 : node4900;
															assign node4900 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node4904 = (inp[0]) ? node4906 : 4'b0000;
															assign node4906 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4909 = (inp[0]) ? node4915 : node4910;
														assign node4910 = (inp[13]) ? 4'b1000 : node4911;
															assign node4911 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4915 = (inp[13]) ? node4917 : 4'b0000;
															assign node4917 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node4920 = (inp[2]) ? node5024 : node4921;
										assign node4921 = (inp[7]) ? node4971 : node4922;
											assign node4922 = (inp[11]) ? node4952 : node4923;
												assign node4923 = (inp[12]) ? node4935 : node4924;
													assign node4924 = (inp[14]) ? node4930 : node4925;
														assign node4925 = (inp[13]) ? 4'b0000 : node4926;
															assign node4926 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node4930 = (inp[0]) ? 4'b0001 : node4931;
															assign node4931 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node4935 = (inp[10]) ? node4947 : node4936;
														assign node4936 = (inp[14]) ? node4942 : node4937;
															assign node4937 = (inp[0]) ? 4'b0001 : node4938;
																assign node4938 = (inp[13]) ? 4'b1000 : 4'b0001;
															assign node4942 = (inp[0]) ? node4944 : 4'b1001;
																assign node4944 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node4947 = (inp[0]) ? 4'b1001 : node4948;
															assign node4948 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node4952 = (inp[13]) ? node4962 : node4953;
													assign node4953 = (inp[0]) ? node4957 : node4954;
														assign node4954 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node4957 = (inp[10]) ? node4959 : 4'b0000;
															assign node4959 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node4962 = (inp[0]) ? node4968 : node4963;
														assign node4963 = (inp[10]) ? 4'b0001 : node4964;
															assign node4964 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node4968 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node4971 = (inp[12]) ? node4995 : node4972;
												assign node4972 = (inp[11]) ? node4984 : node4973;
													assign node4973 = (inp[0]) ? node4975 : 4'b0000;
														assign node4975 = (inp[14]) ? node4979 : node4976;
															assign node4976 = (inp[13]) ? 4'b0001 : 4'b1000;
															assign node4979 = (inp[10]) ? 4'b1000 : node4980;
																assign node4980 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node4984 = (inp[0]) ? node4990 : node4985;
														assign node4985 = (inp[10]) ? 4'b1000 : node4986;
															assign node4986 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node4990 = (inp[10]) ? node4992 : 4'b1000;
															assign node4992 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node4995 = (inp[0]) ? node5011 : node4996;
													assign node4996 = (inp[10]) ? node5004 : node4997;
														assign node4997 = (inp[14]) ? node4999 : 4'b0000;
															assign node4999 = (inp[13]) ? 4'b0001 : node5000;
																assign node5000 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node5004 = (inp[11]) ? 4'b0000 : node5005;
															assign node5005 = (inp[13]) ? 4'b1000 : node5006;
																assign node5006 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node5011 = (inp[10]) ? node5019 : node5012;
														assign node5012 = (inp[11]) ? 4'b1000 : node5013;
															assign node5013 = (inp[13]) ? node5015 : 4'b1000;
																assign node5015 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5019 = (inp[11]) ? 4'b0001 : node5020;
															assign node5020 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node5024 = (inp[7]) ? node5082 : node5025;
											assign node5025 = (inp[14]) ? node5047 : node5026;
												assign node5026 = (inp[11]) ? node5038 : node5027;
													assign node5027 = (inp[0]) ? node5033 : node5028;
														assign node5028 = (inp[13]) ? node5030 : 4'b0000;
															assign node5030 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node5033 = (inp[13]) ? node5035 : 4'b0000;
															assign node5035 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5038 = (inp[0]) ? node5040 : 4'b1001;
														assign node5040 = (inp[13]) ? 4'b1000 : node5041;
															assign node5041 = (inp[10]) ? 4'b0000 : node5042;
																assign node5042 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node5047 = (inp[11]) ? node5063 : node5048;
													assign node5048 = (inp[13]) ? node5054 : node5049;
														assign node5049 = (inp[0]) ? 4'b1001 : node5050;
															assign node5050 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node5054 = (inp[10]) ? node5058 : node5055;
															assign node5055 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5058 = (inp[12]) ? 4'b0001 : node5059;
																assign node5059 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node5063 = (inp[0]) ? node5073 : node5064;
														assign node5064 = (inp[13]) ? 4'b1001 : node5065;
															assign node5065 = (inp[12]) ? node5069 : node5066;
																assign node5066 = (inp[10]) ? 4'b0001 : 4'b1000;
																assign node5069 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node5073 = (inp[12]) ? node5075 : 4'b0000;
															assign node5075 = (inp[10]) ? node5079 : node5076;
																assign node5076 = (inp[13]) ? 4'b0000 : 4'b1001;
																assign node5079 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node5082 = (inp[0]) ? 4'b1001 : node5083;
												assign node5083 = (inp[11]) ? node5097 : node5084;
													assign node5084 = (inp[13]) ? node5092 : node5085;
														assign node5085 = (inp[10]) ? node5089 : node5086;
															assign node5086 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5089 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5092 = (inp[14]) ? 4'b0000 : node5093;
															assign node5093 = (inp[10]) ? 4'b1001 : 4'b0000;
													assign node5097 = (inp[10]) ? 4'b1000 : node5098;
														assign node5098 = (inp[13]) ? 4'b1001 : 4'b0001;
								assign node5103 = (inp[11]) ? node5321 : node5104;
									assign node5104 = (inp[15]) ? node5206 : node5105;
										assign node5105 = (inp[10]) ? node5157 : node5106;
											assign node5106 = (inp[2]) ? node5136 : node5107;
												assign node5107 = (inp[13]) ? node5117 : node5108;
													assign node5108 = (inp[0]) ? node5110 : 4'b0001;
														assign node5110 = (inp[7]) ? node5112 : 4'b0001;
															assign node5112 = (inp[14]) ? 4'b0001 : node5113;
																assign node5113 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5117 = (inp[12]) ? node5127 : node5118;
														assign node5118 = (inp[0]) ? node5122 : node5119;
															assign node5119 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node5122 = (inp[14]) ? 4'b0000 : node5123;
																assign node5123 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node5127 = (inp[7]) ? node5129 : 4'b0001;
															assign node5129 = (inp[14]) ? node5133 : node5130;
																assign node5130 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node5133 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node5136 = (inp[12]) ? node5150 : node5137;
													assign node5137 = (inp[14]) ? 4'b0000 : node5138;
														assign node5138 = (inp[7]) ? node5144 : node5139;
															assign node5139 = (inp[13]) ? node5141 : 4'b0000;
																assign node5141 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5144 = (inp[0]) ? node5146 : 4'b0000;
																assign node5146 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node5150 = (inp[13]) ? 4'b0001 : node5151;
														assign node5151 = (inp[0]) ? node5153 : 4'b1000;
															assign node5153 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node5157 = (inp[13]) ? node5183 : node5158;
												assign node5158 = (inp[2]) ? node5170 : node5159;
													assign node5159 = (inp[7]) ? node5163 : node5160;
														assign node5160 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node5163 = (inp[0]) ? node5167 : node5164;
															assign node5164 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5167 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5170 = (inp[14]) ? node5178 : node5171;
														assign node5171 = (inp[0]) ? 4'b1000 : node5172;
															assign node5172 = (inp[7]) ? 4'b0000 : node5173;
																assign node5173 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5178 = (inp[0]) ? 4'b1000 : node5179;
															assign node5179 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node5183 = (inp[2]) ? node5203 : node5184;
													assign node5184 = (inp[0]) ? node5192 : node5185;
														assign node5185 = (inp[12]) ? node5187 : 4'b0000;
															assign node5187 = (inp[14]) ? 4'b1000 : node5188;
																assign node5188 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node5192 = (inp[12]) ? node5198 : node5193;
															assign node5193 = (inp[7]) ? 4'b1000 : node5194;
																assign node5194 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node5198 = (inp[14]) ? node5200 : 4'b0000;
																assign node5200 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node5203 = (inp[0]) ? 4'b1000 : 4'b0000;
										assign node5206 = (inp[2]) ? node5274 : node5207;
											assign node5207 = (inp[13]) ? node5231 : node5208;
												assign node5208 = (inp[14]) ? node5220 : node5209;
													assign node5209 = (inp[0]) ? node5213 : node5210;
														assign node5210 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node5213 = (inp[12]) ? 4'b0000 : node5214;
															assign node5214 = (inp[10]) ? 4'b0000 : node5215;
																assign node5215 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node5220 = (inp[7]) ? node5226 : node5221;
														assign node5221 = (inp[12]) ? node5223 : 4'b0001;
															assign node5223 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node5226 = (inp[10]) ? 4'b0001 : node5227;
															assign node5227 = (inp[0]) ? 4'b0000 : 4'b1000;
												assign node5231 = (inp[10]) ? node5247 : node5232;
													assign node5232 = (inp[0]) ? node5240 : node5233;
														assign node5233 = (inp[12]) ? node5235 : 4'b0001;
															assign node5235 = (inp[14]) ? 4'b1000 : node5236;
																assign node5236 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node5240 = (inp[7]) ? node5244 : node5241;
															assign node5241 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node5244 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node5247 = (inp[7]) ? node5259 : node5248;
														assign node5248 = (inp[14]) ? node5254 : node5249;
															assign node5249 = (inp[12]) ? node5251 : 4'b1001;
																assign node5251 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node5254 = (inp[12]) ? node5256 : 4'b0000;
																assign node5256 = (inp[0]) ? 4'b0000 : 4'b1001;
														assign node5259 = (inp[14]) ? node5267 : node5260;
															assign node5260 = (inp[0]) ? node5264 : node5261;
																assign node5261 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node5264 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node5267 = (inp[12]) ? node5271 : node5268;
																assign node5268 = (inp[0]) ? 4'b1001 : 4'b0001;
																assign node5271 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node5274 = (inp[7]) ? node5304 : node5275;
												assign node5275 = (inp[14]) ? node5289 : node5276;
													assign node5276 = (inp[0]) ? node5284 : node5277;
														assign node5277 = (inp[10]) ? node5281 : node5278;
															assign node5278 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node5281 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5284 = (inp[13]) ? node5286 : 4'b0001;
															assign node5286 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5289 = (inp[10]) ? 4'b0000 : node5290;
														assign node5290 = (inp[0]) ? node5296 : node5291;
															assign node5291 = (inp[13]) ? node5293 : 4'b1000;
																assign node5293 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node5296 = (inp[13]) ? node5300 : node5297;
																assign node5297 = (inp[12]) ? 4'b1001 : 4'b0000;
																assign node5300 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5304 = (inp[0]) ? 4'b1001 : node5305;
													assign node5305 = (inp[10]) ? node5311 : node5306;
														assign node5306 = (inp[13]) ? 4'b1000 : node5307;
															assign node5307 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5311 = (inp[13]) ? 4'b0001 : node5312;
															assign node5312 = (inp[12]) ? node5316 : node5313;
																assign node5313 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node5316 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node5321 = (inp[13]) ? node5401 : node5322;
										assign node5322 = (inp[2]) ? node5360 : node5323;
											assign node5323 = (inp[15]) ? node5347 : node5324;
												assign node5324 = (inp[7]) ? node5336 : node5325;
													assign node5325 = (inp[12]) ? node5333 : node5326;
														assign node5326 = (inp[10]) ? node5330 : node5327;
															assign node5327 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node5330 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node5333 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node5336 = (inp[14]) ? 4'b1001 : node5337;
														assign node5337 = (inp[12]) ? node5339 : 4'b1001;
															assign node5339 = (inp[0]) ? node5343 : node5340;
																assign node5340 = (inp[10]) ? 4'b0001 : 4'b1001;
																assign node5343 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node5347 = (inp[12]) ? 4'b0001 : node5348;
													assign node5348 = (inp[0]) ? node5354 : node5349;
														assign node5349 = (inp[10]) ? node5351 : 4'b1001;
															assign node5351 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node5354 = (inp[7]) ? 4'b0001 : node5355;
															assign node5355 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node5360 = (inp[12]) ? node5376 : node5361;
												assign node5361 = (inp[15]) ? node5367 : node5362;
													assign node5362 = (inp[0]) ? node5364 : 4'b0001;
														assign node5364 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node5367 = (inp[0]) ? node5373 : node5368;
														assign node5368 = (inp[7]) ? 4'b0001 : node5369;
															assign node5369 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node5373 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node5376 = (inp[15]) ? node5392 : node5377;
													assign node5377 = (inp[0]) ? node5379 : 4'b0001;
														assign node5379 = (inp[14]) ? node5387 : node5380;
															assign node5380 = (inp[10]) ? node5384 : node5381;
																assign node5381 = (inp[7]) ? 4'b1001 : 4'b0001;
																assign node5384 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node5387 = (inp[10]) ? node5389 : 4'b1001;
																assign node5389 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node5392 = (inp[10]) ? node5394 : 4'b1001;
														assign node5394 = (inp[7]) ? node5398 : node5395;
															assign node5395 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node5398 = (inp[0]) ? 4'b1001 : 4'b0001;
										assign node5401 = (inp[10]) ? 4'b1001 : node5402;
											assign node5402 = (inp[14]) ? node5430 : node5403;
												assign node5403 = (inp[2]) ? node5425 : node5404;
													assign node5404 = (inp[7]) ? node5418 : node5405;
														assign node5405 = (inp[12]) ? node5413 : node5406;
															assign node5406 = (inp[15]) ? node5410 : node5407;
																assign node5407 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node5410 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node5413 = (inp[0]) ? node5415 : 4'b1001;
																assign node5415 = (inp[15]) ? 4'b1001 : 4'b0001;
														assign node5418 = (inp[0]) ? node5420 : 4'b0001;
															assign node5420 = (inp[15]) ? 4'b0001 : node5421;
																assign node5421 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5425 = (inp[12]) ? 4'b0001 : node5426;
														assign node5426 = (inp[15]) ? 4'b0001 : 4'b1001;
												assign node5430 = (inp[12]) ? node5446 : node5431;
													assign node5431 = (inp[0]) ? node5439 : node5432;
														assign node5432 = (inp[15]) ? 4'b0001 : node5433;
															assign node5433 = (inp[2]) ? 4'b1001 : node5434;
																assign node5434 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node5439 = (inp[2]) ? 4'b1001 : node5440;
															assign node5440 = (inp[15]) ? node5442 : 4'b1001;
																assign node5442 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node5446 = (inp[0]) ? node5454 : node5447;
														assign node5447 = (inp[15]) ? node5449 : 4'b1001;
															assign node5449 = (inp[7]) ? 4'b0001 : node5450;
																assign node5450 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node5454 = (inp[15]) ? node5456 : 4'b0001;
															assign node5456 = (inp[2]) ? 4'b0001 : 4'b1001;
							assign node5460 = (inp[13]) ? node5860 : node5461;
								assign node5461 = (inp[1]) ? node5673 : node5462;
									assign node5462 = (inp[10]) ? node5576 : node5463;
										assign node5463 = (inp[2]) ? node5519 : node5464;
											assign node5464 = (inp[0]) ? node5488 : node5465;
												assign node5465 = (inp[7]) ? node5477 : node5466;
													assign node5466 = (inp[15]) ? 4'b1000 : node5467;
														assign node5467 = (inp[14]) ? node5473 : node5468;
															assign node5468 = (inp[12]) ? node5470 : 4'b0000;
																assign node5470 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node5473 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node5477 = (inp[12]) ? node5485 : node5478;
														assign node5478 = (inp[11]) ? 4'b1001 : node5479;
															assign node5479 = (inp[14]) ? 4'b1000 : node5480;
																assign node5480 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node5485 = (inp[15]) ? 4'b0001 : 4'b1001;
												assign node5488 = (inp[11]) ? node5506 : node5489;
													assign node5489 = (inp[12]) ? node5501 : node5490;
														assign node5490 = (inp[15]) ? node5496 : node5491;
															assign node5491 = (inp[7]) ? node5493 : 4'b0001;
																assign node5493 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node5496 = (inp[7]) ? node5498 : 4'b0000;
																assign node5498 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5501 = (inp[15]) ? 4'b1001 : node5502;
															assign node5502 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node5506 = (inp[7]) ? node5514 : node5507;
														assign node5507 = (inp[12]) ? node5511 : node5508;
															assign node5508 = (inp[15]) ? 4'b1001 : 4'b0000;
															assign node5511 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node5514 = (inp[15]) ? node5516 : 4'b1000;
															assign node5516 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node5519 = (inp[15]) ? node5545 : node5520;
												assign node5520 = (inp[14]) ? node5530 : node5521;
													assign node5521 = (inp[0]) ? node5525 : node5522;
														assign node5522 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5525 = (inp[12]) ? node5527 : 4'b0001;
															assign node5527 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node5530 = (inp[12]) ? node5536 : node5531;
														assign node5531 = (inp[0]) ? node5533 : 4'b1000;
															assign node5533 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node5536 = (inp[0]) ? 4'b0000 : node5537;
															assign node5537 = (inp[11]) ? node5541 : node5538;
																assign node5538 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node5541 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node5545 = (inp[7]) ? node5559 : node5546;
													assign node5546 = (inp[11]) ? node5556 : node5547;
														assign node5547 = (inp[12]) ? node5551 : node5548;
															assign node5548 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node5551 = (inp[0]) ? node5553 : 4'b0000;
																assign node5553 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node5556 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node5559 = (inp[14]) ? node5569 : node5560;
														assign node5560 = (inp[11]) ? node5566 : node5561;
															assign node5561 = (inp[12]) ? 4'b0000 : node5562;
																assign node5562 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node5566 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5569 = (inp[0]) ? 4'b1001 : node5570;
															assign node5570 = (inp[12]) ? node5572 : 4'b0001;
																assign node5572 = (inp[11]) ? 4'b1000 : 4'b0001;
										assign node5576 = (inp[11]) ? node5634 : node5577;
											assign node5577 = (inp[14]) ? node5599 : node5578;
												assign node5578 = (inp[7]) ? node5584 : node5579;
													assign node5579 = (inp[2]) ? node5581 : 4'b0001;
														assign node5581 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5584 = (inp[2]) ? node5596 : node5585;
														assign node5585 = (inp[15]) ? node5591 : node5586;
															assign node5586 = (inp[12]) ? node5588 : 4'b0000;
																assign node5588 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node5591 = (inp[12]) ? node5593 : 4'b1000;
																assign node5593 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node5596 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node5599 = (inp[2]) ? node5617 : node5600;
													assign node5600 = (inp[0]) ? node5610 : node5601;
														assign node5601 = (inp[12]) ? node5607 : node5602;
															assign node5602 = (inp[15]) ? node5604 : 4'b0001;
																assign node5604 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node5607 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node5610 = (inp[12]) ? node5612 : 4'b0000;
															assign node5612 = (inp[15]) ? 4'b0001 : node5613;
																assign node5613 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node5617 = (inp[12]) ? node5625 : node5618;
														assign node5618 = (inp[7]) ? node5622 : node5619;
															assign node5619 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node5622 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node5625 = (inp[7]) ? node5629 : node5626;
															assign node5626 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node5629 = (inp[15]) ? node5631 : 4'b1000;
																assign node5631 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node5634 = (inp[2]) ? node5654 : node5635;
												assign node5635 = (inp[15]) ? node5647 : node5636;
													assign node5636 = (inp[0]) ? node5642 : node5637;
														assign node5637 = (inp[12]) ? 4'b0000 : node5638;
															assign node5638 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node5642 = (inp[12]) ? 4'b0001 : node5643;
															assign node5643 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node5647 = (inp[7]) ? 4'b1000 : node5648;
														assign node5648 = (inp[0]) ? 4'b0000 : node5649;
															assign node5649 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node5654 = (inp[7]) ? node5668 : node5655;
													assign node5655 = (inp[12]) ? node5663 : node5656;
														assign node5656 = (inp[15]) ? node5660 : node5657;
															assign node5657 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5660 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node5663 = (inp[0]) ? node5665 : 4'b0001;
															assign node5665 = (inp[15]) ? 4'b0001 : 4'b1000;
													assign node5668 = (inp[0]) ? 4'b0000 : node5669;
														assign node5669 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node5673 = (inp[11]) ? node5811 : node5674;
										assign node5674 = (inp[10]) ? node5734 : node5675;
											assign node5675 = (inp[15]) ? node5703 : node5676;
												assign node5676 = (inp[0]) ? node5692 : node5677;
													assign node5677 = (inp[7]) ? node5687 : node5678;
														assign node5678 = (inp[12]) ? node5684 : node5679;
															assign node5679 = (inp[2]) ? 4'b1000 : node5680;
																assign node5680 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node5684 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node5687 = (inp[2]) ? node5689 : 4'b0000;
															assign node5689 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5692 = (inp[12]) ? node5696 : node5693;
														assign node5693 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node5696 = (inp[2]) ? node5698 : 4'b0001;
															assign node5698 = (inp[7]) ? node5700 : 4'b0001;
																assign node5700 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node5703 = (inp[12]) ? node5719 : node5704;
													assign node5704 = (inp[0]) ? node5714 : node5705;
														assign node5705 = (inp[7]) ? node5711 : node5706;
															assign node5706 = (inp[2]) ? 4'b0001 : node5707;
																assign node5707 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node5711 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node5714 = (inp[2]) ? 4'b0000 : node5715;
															assign node5715 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node5719 = (inp[2]) ? node5727 : node5720;
														assign node5720 = (inp[0]) ? node5724 : node5721;
															assign node5721 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node5724 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5727 = (inp[7]) ? node5731 : node5728;
															assign node5728 = (inp[0]) ? 4'b0000 : 4'b1001;
															assign node5731 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node5734 = (inp[14]) ? node5778 : node5735;
												assign node5735 = (inp[15]) ? node5757 : node5736;
													assign node5736 = (inp[2]) ? node5750 : node5737;
														assign node5737 = (inp[12]) ? node5743 : node5738;
															assign node5738 = (inp[7]) ? 4'b0001 : node5739;
																assign node5739 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5743 = (inp[0]) ? node5747 : node5744;
																assign node5744 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node5747 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node5750 = (inp[7]) ? node5754 : node5751;
															assign node5751 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5754 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node5757 = (inp[12]) ? node5763 : node5758;
														assign node5758 = (inp[0]) ? 4'b0000 : node5759;
															assign node5759 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node5763 = (inp[2]) ? node5771 : node5764;
															assign node5764 = (inp[0]) ? node5768 : node5765;
																assign node5765 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node5768 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node5771 = (inp[7]) ? node5775 : node5772;
																assign node5772 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node5775 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node5778 = (inp[2]) ? node5790 : node5779;
													assign node5779 = (inp[7]) ? node5783 : node5780;
														assign node5780 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node5783 = (inp[0]) ? 4'b0001 : node5784;
															assign node5784 = (inp[15]) ? node5786 : 4'b0000;
																assign node5786 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5790 = (inp[0]) ? node5800 : node5791;
														assign node5791 = (inp[12]) ? node5795 : node5792;
															assign node5792 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node5795 = (inp[7]) ? node5797 : 4'b0001;
																assign node5797 = (inp[15]) ? 4'b0001 : 4'b1000;
														assign node5800 = (inp[7]) ? node5806 : node5801;
															assign node5801 = (inp[12]) ? 4'b1000 : node5802;
																assign node5802 = (inp[15]) ? 4'b0001 : 4'b1000;
															assign node5806 = (inp[15]) ? 4'b0000 : node5807;
																assign node5807 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node5811 = (inp[10]) ? 4'b0001 : node5812;
											assign node5812 = (inp[15]) ? node5846 : node5813;
												assign node5813 = (inp[14]) ? node5835 : node5814;
													assign node5814 = (inp[7]) ? node5824 : node5815;
														assign node5815 = (inp[2]) ? node5817 : 4'b0001;
															assign node5817 = (inp[12]) ? node5821 : node5818;
																assign node5818 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node5821 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node5824 = (inp[0]) ? node5830 : node5825;
															assign node5825 = (inp[2]) ? 4'b0001 : node5826;
																assign node5826 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node5830 = (inp[2]) ? node5832 : 4'b1001;
																assign node5832 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5835 = (inp[7]) ? 4'b0001 : node5836;
														assign node5836 = (inp[0]) ? 4'b0001 : node5837;
															assign node5837 = (inp[12]) ? node5841 : node5838;
																assign node5838 = (inp[2]) ? 4'b1001 : 4'b0001;
																assign node5841 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node5846 = (inp[2]) ? 4'b0001 : node5847;
													assign node5847 = (inp[7]) ? node5853 : node5848;
														assign node5848 = (inp[12]) ? 4'b0001 : node5849;
															assign node5849 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node5853 = (inp[0]) ? 4'b0001 : node5854;
															assign node5854 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node5860 = (inp[10]) ? node6016 : node5861;
									assign node5861 = (inp[1]) ? node5975 : node5862;
										assign node5862 = (inp[11]) ? node5920 : node5863;
											assign node5863 = (inp[0]) ? node5889 : node5864;
												assign node5864 = (inp[7]) ? node5880 : node5865;
													assign node5865 = (inp[14]) ? node5873 : node5866;
														assign node5866 = (inp[2]) ? node5868 : 4'b0001;
															assign node5868 = (inp[12]) ? 4'b0000 : node5869;
																assign node5869 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node5873 = (inp[12]) ? 4'b0000 : node5874;
															assign node5874 = (inp[2]) ? 4'b0000 : node5875;
																assign node5875 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node5880 = (inp[2]) ? 4'b0001 : node5881;
														assign node5881 = (inp[14]) ? node5883 : 4'b0000;
															assign node5883 = (inp[15]) ? 4'b0001 : node5884;
																assign node5884 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node5889 = (inp[7]) ? node5909 : node5890;
													assign node5890 = (inp[14]) ? node5898 : node5891;
														assign node5891 = (inp[2]) ? node5893 : 4'b0000;
															assign node5893 = (inp[15]) ? 4'b0001 : node5894;
																assign node5894 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node5898 = (inp[12]) ? node5904 : node5899;
															assign node5899 = (inp[2]) ? 4'b0001 : node5900;
																assign node5900 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node5904 = (inp[15]) ? node5906 : 4'b0001;
																assign node5906 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node5909 = (inp[12]) ? node5911 : 4'b0000;
														assign node5911 = (inp[15]) ? node5917 : node5912;
															assign node5912 = (inp[14]) ? 4'b0000 : node5913;
																assign node5913 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node5917 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node5920 = (inp[15]) ? node5950 : node5921;
												assign node5921 = (inp[14]) ? node5935 : node5922;
													assign node5922 = (inp[0]) ? 4'b0000 : node5923;
														assign node5923 = (inp[2]) ? node5929 : node5924;
															assign node5924 = (inp[12]) ? 4'b0000 : node5925;
																assign node5925 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node5929 = (inp[7]) ? node5931 : 4'b0000;
																assign node5931 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node5935 = (inp[2]) ? node5945 : node5936;
														assign node5936 = (inp[0]) ? node5938 : 4'b0000;
															assign node5938 = (inp[12]) ? node5942 : node5939;
																assign node5939 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node5942 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node5945 = (inp[12]) ? node5947 : 4'b0001;
															assign node5947 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node5950 = (inp[2]) ? node5962 : node5951;
													assign node5951 = (inp[7]) ? node5957 : node5952;
														assign node5952 = (inp[0]) ? 4'b0000 : node5953;
															assign node5953 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node5957 = (inp[12]) ? node5959 : 4'b0001;
															assign node5959 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node5962 = (inp[7]) ? node5970 : node5963;
														assign node5963 = (inp[0]) ? node5967 : node5964;
															assign node5964 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node5967 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node5970 = (inp[12]) ? 4'b0000 : node5971;
															assign node5971 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node5975 = (inp[11]) ? 4'b0001 : node5976;
											assign node5976 = (inp[0]) ? node5998 : node5977;
												assign node5977 = (inp[15]) ? node5989 : node5978;
													assign node5978 = (inp[14]) ? node5984 : node5979;
														assign node5979 = (inp[2]) ? node5981 : 4'b0000;
															assign node5981 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node5984 = (inp[7]) ? node5986 : 4'b0000;
															assign node5986 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node5989 = (inp[7]) ? 4'b0001 : node5990;
														assign node5990 = (inp[14]) ? node5992 : 4'b0000;
															assign node5992 = (inp[2]) ? node5994 : 4'b0001;
																assign node5994 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node5998 = (inp[15]) ? 4'b0000 : node5999;
													assign node5999 = (inp[12]) ? node6007 : node6000;
														assign node6000 = (inp[7]) ? 4'b0000 : node6001;
															assign node6001 = (inp[2]) ? 4'b0001 : node6002;
																assign node6002 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6007 = (inp[7]) ? node6011 : node6008;
															assign node6008 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6011 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node6016 = (inp[11]) ? 4'b0000 : node6017;
										assign node6017 = (inp[1]) ? 4'b0000 : node6018;
											assign node6018 = (inp[2]) ? node6060 : node6019;
												assign node6019 = (inp[12]) ? node6039 : node6020;
													assign node6020 = (inp[0]) ? node6034 : node6021;
														assign node6021 = (inp[15]) ? node6029 : node6022;
															assign node6022 = (inp[7]) ? node6026 : node6023;
																assign node6023 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node6026 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6029 = (inp[14]) ? node6031 : 4'b0000;
																assign node6031 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6034 = (inp[14]) ? 4'b0000 : node6035;
															assign node6035 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node6039 = (inp[15]) ? node6051 : node6040;
														assign node6040 = (inp[7]) ? node6046 : node6041;
															assign node6041 = (inp[14]) ? 4'b0001 : node6042;
																assign node6042 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6046 = (inp[0]) ? node6048 : 4'b0000;
																assign node6048 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6051 = (inp[14]) ? node6055 : node6052;
															assign node6052 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6055 = (inp[0]) ? 4'b0001 : node6056;
																assign node6056 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node6060 = (inp[15]) ? node6072 : node6061;
													assign node6061 = (inp[14]) ? 4'b0000 : node6062;
														assign node6062 = (inp[7]) ? 4'b0000 : node6063;
															assign node6063 = (inp[0]) ? node6067 : node6064;
																assign node6064 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node6067 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node6072 = (inp[0]) ? node6080 : node6073;
														assign node6073 = (inp[14]) ? 4'b0000 : node6074;
															assign node6074 = (inp[7]) ? 4'b0000 : node6075;
																assign node6075 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node6080 = (inp[14]) ? 4'b0001 : node6081;
															assign node6081 = (inp[7]) ? node6083 : 4'b0000;
																assign node6083 = (inp[12]) ? 4'b0001 : 4'b0000;
			assign node6089 = (inp[15]) ? node9189 : node6090;
				assign node6090 = (inp[6]) ? node6828 : node6091;
					assign node6091 = (inp[0]) ? 4'b0101 : node6092;
						assign node6092 = (inp[2]) ? node6560 : node6093;
							assign node6093 = (inp[1]) ? node6331 : node6094;
								assign node6094 = (inp[11]) ? node6242 : node6095;
									assign node6095 = (inp[14]) ? node6169 : node6096;
										assign node6096 = (inp[3]) ? node6138 : node6097;
											assign node6097 = (inp[5]) ? node6119 : node6098;
												assign node6098 = (inp[13]) ? node6104 : node6099;
													assign node6099 = (inp[7]) ? 4'b0111 : node6100;
														assign node6100 = (inp[4]) ? 4'b1000 : 4'b0111;
													assign node6104 = (inp[7]) ? node6114 : node6105;
														assign node6105 = (inp[4]) ? node6111 : node6106;
															assign node6106 = (inp[10]) ? 4'b0000 : node6107;
																assign node6107 = (inp[12]) ? 4'b0111 : 4'b0000;
															assign node6111 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node6114 = (inp[4]) ? node6116 : 4'b0111;
															assign node6116 = (inp[12]) ? 4'b0111 : 4'b0000;
												assign node6119 = (inp[13]) ? node6129 : node6120;
													assign node6120 = (inp[10]) ? node6124 : node6121;
														assign node6121 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node6124 = (inp[4]) ? node6126 : 4'b1100;
															assign node6126 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node6129 = (inp[12]) ? node6135 : node6130;
														assign node6130 = (inp[7]) ? node6132 : 4'b0000;
															assign node6132 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node6135 = (inp[10]) ? 4'b0100 : 4'b1100;
											assign node6138 = (inp[13]) ? node6152 : node6139;
												assign node6139 = (inp[12]) ? node6141 : 4'b1000;
													assign node6141 = (inp[10]) ? node6147 : node6142;
														assign node6142 = (inp[7]) ? 4'b0000 : node6143;
															assign node6143 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node6147 = (inp[7]) ? 4'b1000 : node6148;
															assign node6148 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6152 = (inp[7]) ? node6158 : node6153;
													assign node6153 = (inp[12]) ? node6155 : 4'b0100;
														assign node6155 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node6158 = (inp[4]) ? node6164 : node6159;
														assign node6159 = (inp[10]) ? 4'b0000 : node6160;
															assign node6160 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node6164 = (inp[12]) ? node6166 : 4'b0100;
															assign node6166 = (inp[10]) ? 4'b0100 : 4'b1000;
										assign node6169 = (inp[3]) ? node6205 : node6170;
											assign node6170 = (inp[5]) ? node6184 : node6171;
												assign node6171 = (inp[4]) ? node6173 : 4'b0111;
													assign node6173 = (inp[7]) ? 4'b0111 : node6174;
														assign node6174 = (inp[13]) ? node6180 : node6175;
															assign node6175 = (inp[12]) ? 4'b0001 : node6176;
																assign node6176 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node6180 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node6184 = (inp[4]) ? node6198 : node6185;
													assign node6185 = (inp[13]) ? node6191 : node6186;
														assign node6186 = (inp[12]) ? 4'b0101 : node6187;
															assign node6187 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node6191 = (inp[10]) ? node6193 : 4'b1101;
															assign node6193 = (inp[7]) ? node6195 : 4'b0001;
																assign node6195 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node6198 = (inp[7]) ? node6202 : node6199;
														assign node6199 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6202 = (inp[13]) ? 4'b0001 : 4'b0101;
											assign node6205 = (inp[7]) ? node6229 : node6206;
												assign node6206 = (inp[4]) ? node6218 : node6207;
													assign node6207 = (inp[13]) ? node6213 : node6208;
														assign node6208 = (inp[12]) ? 4'b0001 : node6209;
															assign node6209 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6213 = (inp[10]) ? node6215 : 4'b1001;
															assign node6215 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node6218 = (inp[13]) ? node6224 : node6219;
														assign node6219 = (inp[12]) ? 4'b0101 : node6220;
															assign node6220 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node6224 = (inp[12]) ? 4'b1101 : node6225;
															assign node6225 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node6229 = (inp[13]) ? node6235 : node6230;
													assign node6230 = (inp[10]) ? node6232 : 4'b0001;
														assign node6232 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6235 = (inp[10]) ? node6237 : 4'b1001;
														assign node6237 = (inp[12]) ? 4'b1001 : node6238;
															assign node6238 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node6242 = (inp[13]) ? node6286 : node6243;
										assign node6243 = (inp[3]) ? node6269 : node6244;
											assign node6244 = (inp[5]) ? node6254 : node6245;
												assign node6245 = (inp[7]) ? 4'b0111 : node6246;
													assign node6246 = (inp[4]) ? node6248 : 4'b0111;
														assign node6248 = (inp[12]) ? node6250 : 4'b1000;
															assign node6250 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node6254 = (inp[12]) ? node6260 : node6255;
													assign node6255 = (inp[7]) ? 4'b1100 : node6256;
														assign node6256 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node6260 = (inp[10]) ? node6266 : node6261;
														assign node6261 = (inp[4]) ? node6263 : 4'b0100;
															assign node6263 = (inp[14]) ? 4'b0000 : 4'b0100;
														assign node6266 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node6269 = (inp[10]) ? node6281 : node6270;
												assign node6270 = (inp[12]) ? node6276 : node6271;
													assign node6271 = (inp[7]) ? 4'b1000 : node6272;
														assign node6272 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node6276 = (inp[4]) ? node6278 : 4'b0000;
														assign node6278 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node6281 = (inp[7]) ? 4'b1000 : node6282;
													assign node6282 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node6286 = (inp[10]) ? node6318 : node6287;
											assign node6287 = (inp[12]) ? node6301 : node6288;
												assign node6288 = (inp[3]) ? node6296 : node6289;
													assign node6289 = (inp[4]) ? 4'b0000 : node6290;
														assign node6290 = (inp[7]) ? node6292 : 4'b0000;
															assign node6292 = (inp[14]) ? 4'b0100 : 4'b0111;
													assign node6296 = (inp[4]) ? 4'b0100 : node6297;
														assign node6297 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node6301 = (inp[3]) ? node6313 : node6302;
													assign node6302 = (inp[5]) ? node6308 : node6303;
														assign node6303 = (inp[14]) ? 4'b0111 : node6304;
															assign node6304 = (inp[4]) ? 4'b1000 : 4'b0111;
														assign node6308 = (inp[7]) ? 4'b1100 : node6309;
															assign node6309 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node6313 = (inp[7]) ? 4'b1000 : node6314;
														assign node6314 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node6318 = (inp[3]) ? node6326 : node6319;
												assign node6319 = (inp[7]) ? node6321 : 4'b0000;
													assign node6321 = (inp[4]) ? 4'b0000 : node6322;
														assign node6322 = (inp[5]) ? 4'b0100 : 4'b0111;
												assign node6326 = (inp[4]) ? 4'b0100 : node6327;
													assign node6327 = (inp[7]) ? 4'b0000 : 4'b0100;
								assign node6331 = (inp[14]) ? node6417 : node6332;
									assign node6332 = (inp[13]) ? node6374 : node6333;
										assign node6333 = (inp[3]) ? node6361 : node6334;
											assign node6334 = (inp[5]) ? node6344 : node6335;
												assign node6335 = (inp[7]) ? 4'b0111 : node6336;
													assign node6336 = (inp[4]) ? node6338 : 4'b0111;
														assign node6338 = (inp[12]) ? node6340 : 4'b1001;
															assign node6340 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node6344 = (inp[7]) ? node6356 : node6345;
													assign node6345 = (inp[4]) ? node6351 : node6346;
														assign node6346 = (inp[10]) ? 4'b1101 : node6347;
															assign node6347 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node6351 = (inp[12]) ? node6353 : 4'b1001;
															assign node6353 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6356 = (inp[12]) ? node6358 : 4'b1101;
														assign node6358 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node6361 = (inp[10]) ? node6369 : node6362;
												assign node6362 = (inp[12]) ? node6364 : 4'b1001;
													assign node6364 = (inp[7]) ? 4'b0001 : node6365;
														assign node6365 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node6369 = (inp[7]) ? 4'b1001 : node6370;
													assign node6370 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node6374 = (inp[10]) ? node6404 : node6375;
											assign node6375 = (inp[12]) ? node6389 : node6376;
												assign node6376 = (inp[3]) ? node6384 : node6377;
													assign node6377 = (inp[4]) ? 4'b0001 : node6378;
														assign node6378 = (inp[7]) ? node6380 : 4'b0001;
															assign node6380 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node6384 = (inp[4]) ? 4'b0101 : node6385;
														assign node6385 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node6389 = (inp[3]) ? node6399 : node6390;
													assign node6390 = (inp[5]) ? node6394 : node6391;
														assign node6391 = (inp[7]) ? 4'b0111 : 4'b1001;
														assign node6394 = (inp[4]) ? node6396 : 4'b1101;
															assign node6396 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node6399 = (inp[4]) ? node6401 : 4'b1001;
														assign node6401 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node6404 = (inp[3]) ? node6412 : node6405;
												assign node6405 = (inp[4]) ? 4'b0001 : node6406;
													assign node6406 = (inp[7]) ? node6408 : 4'b0001;
														assign node6408 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node6412 = (inp[7]) ? node6414 : 4'b0101;
													assign node6414 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node6417 = (inp[11]) ? node6491 : node6418;
										assign node6418 = (inp[13]) ? node6458 : node6419;
											assign node6419 = (inp[3]) ? node6441 : node6420;
												assign node6420 = (inp[5]) ? node6426 : node6421;
													assign node6421 = (inp[7]) ? 4'b0111 : node6422;
														assign node6422 = (inp[4]) ? 4'b1000 : 4'b0111;
													assign node6426 = (inp[12]) ? node6432 : node6427;
														assign node6427 = (inp[7]) ? 4'b1100 : node6428;
															assign node6428 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node6432 = (inp[10]) ? node6438 : node6433;
															assign node6433 = (inp[4]) ? node6435 : 4'b0100;
																assign node6435 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node6438 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node6441 = (inp[7]) ? node6453 : node6442;
													assign node6442 = (inp[4]) ? node6448 : node6443;
														assign node6443 = (inp[12]) ? node6445 : 4'b1000;
															assign node6445 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6448 = (inp[10]) ? 4'b1100 : node6449;
															assign node6449 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node6453 = (inp[12]) ? node6455 : 4'b1000;
														assign node6455 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node6458 = (inp[12]) ? node6472 : node6459;
												assign node6459 = (inp[3]) ? node6467 : node6460;
													assign node6460 = (inp[4]) ? 4'b0000 : node6461;
														assign node6461 = (inp[7]) ? node6463 : 4'b0000;
															assign node6463 = (inp[5]) ? 4'b0100 : 4'b0111;
													assign node6467 = (inp[4]) ? 4'b0100 : node6468;
														assign node6468 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node6472 = (inp[10]) ? node6480 : node6473;
													assign node6473 = (inp[3]) ? 4'b1000 : node6474;
														assign node6474 = (inp[7]) ? 4'b0111 : node6475;
															assign node6475 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node6480 = (inp[4]) ? 4'b0000 : node6481;
														assign node6481 = (inp[5]) ? node6483 : 4'b0100;
															assign node6483 = (inp[3]) ? node6487 : node6484;
																assign node6484 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node6487 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node6491 = (inp[13]) ? node6523 : node6492;
											assign node6492 = (inp[3]) ? node6508 : node6493;
												assign node6493 = (inp[5]) ? node6499 : node6494;
													assign node6494 = (inp[7]) ? 4'b0111 : node6495;
														assign node6495 = (inp[4]) ? 4'b1001 : 4'b0111;
													assign node6499 = (inp[10]) ? node6503 : node6500;
														assign node6500 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node6503 = (inp[4]) ? node6505 : 4'b1101;
															assign node6505 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node6508 = (inp[7]) ? node6518 : node6509;
													assign node6509 = (inp[4]) ? node6513 : node6510;
														assign node6510 = (inp[5]) ? 4'b1001 : 4'b0001;
														assign node6513 = (inp[12]) ? node6515 : 4'b1101;
															assign node6515 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node6518 = (inp[10]) ? 4'b1001 : node6519;
														assign node6519 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6523 = (inp[10]) ? node6549 : node6524;
												assign node6524 = (inp[12]) ? node6538 : node6525;
													assign node6525 = (inp[3]) ? node6533 : node6526;
														assign node6526 = (inp[4]) ? 4'b0001 : node6527;
															assign node6527 = (inp[5]) ? node6529 : 4'b0111;
																assign node6529 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node6533 = (inp[7]) ? node6535 : 4'b0101;
															assign node6535 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node6538 = (inp[7]) ? node6546 : node6539;
														assign node6539 = (inp[3]) ? node6543 : node6540;
															assign node6540 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node6543 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node6546 = (inp[3]) ? 4'b1001 : 4'b0111;
												assign node6549 = (inp[3]) ? node6555 : node6550;
													assign node6550 = (inp[7]) ? node6552 : 4'b0001;
														assign node6552 = (inp[4]) ? 4'b0001 : 4'b0111;
													assign node6555 = (inp[4]) ? 4'b0101 : node6556;
														assign node6556 = (inp[7]) ? 4'b0001 : 4'b0101;
							assign node6560 = (inp[5]) ? node6562 : 4'b0111;
								assign node6562 = (inp[3]) ? node6658 : node6563;
									assign node6563 = (inp[4]) ? node6581 : node6564;
										assign node6564 = (inp[7]) ? 4'b0111 : node6565;
											assign node6565 = (inp[13]) ? node6567 : 4'b0111;
												assign node6567 = (inp[12]) ? node6575 : node6568;
													assign node6568 = (inp[1]) ? 4'b0001 : node6569;
														assign node6569 = (inp[14]) ? node6571 : 4'b0000;
															assign node6571 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node6575 = (inp[10]) ? node6577 : 4'b0111;
														assign node6577 = (inp[14]) ? 4'b0111 : 4'b0000;
										assign node6581 = (inp[7]) ? node6633 : node6582;
											assign node6582 = (inp[13]) ? node6612 : node6583;
												assign node6583 = (inp[10]) ? node6601 : node6584;
													assign node6584 = (inp[12]) ? node6592 : node6585;
														assign node6585 = (inp[14]) ? node6589 : node6586;
															assign node6586 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node6589 = (inp[1]) ? 4'b1000 : 4'b0001;
														assign node6592 = (inp[14]) ? node6594 : 4'b0000;
															assign node6594 = (inp[1]) ? node6598 : node6595;
																assign node6595 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node6598 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node6601 = (inp[1]) ? node6607 : node6602;
														assign node6602 = (inp[12]) ? node6604 : 4'b1000;
															assign node6604 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node6607 = (inp[14]) ? node6609 : 4'b1001;
															assign node6609 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node6612 = (inp[1]) ? node6620 : node6613;
													assign node6613 = (inp[12]) ? node6617 : node6614;
														assign node6614 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node6617 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node6620 = (inp[10]) ? node6628 : node6621;
														assign node6621 = (inp[12]) ? 4'b1001 : node6622;
															assign node6622 = (inp[11]) ? 4'b0001 : node6623;
																assign node6623 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6628 = (inp[11]) ? 4'b0001 : node6629;
															assign node6629 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node6633 = (inp[13]) ? node6635 : 4'b0111;
												assign node6635 = (inp[10]) ? node6647 : node6636;
													assign node6636 = (inp[12]) ? 4'b0111 : node6637;
														assign node6637 = (inp[11]) ? node6643 : node6638;
															assign node6638 = (inp[1]) ? node6640 : 4'b0111;
																assign node6640 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6643 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node6647 = (inp[1]) ? node6653 : node6648;
														assign node6648 = (inp[11]) ? 4'b0000 : node6649;
															assign node6649 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6653 = (inp[11]) ? 4'b0001 : node6654;
															assign node6654 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node6658 = (inp[1]) ? node6742 : node6659;
										assign node6659 = (inp[14]) ? node6693 : node6660;
											assign node6660 = (inp[13]) ? node6676 : node6661;
												assign node6661 = (inp[10]) ? node6671 : node6662;
													assign node6662 = (inp[12]) ? node6666 : node6663;
														assign node6663 = (inp[11]) ? 4'b1100 : 4'b1000;
														assign node6666 = (inp[7]) ? 4'b0000 : node6667;
															assign node6667 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node6671 = (inp[7]) ? 4'b1000 : node6672;
														assign node6672 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6676 = (inp[4]) ? node6688 : node6677;
													assign node6677 = (inp[7]) ? node6683 : node6678;
														assign node6678 = (inp[12]) ? node6680 : 4'b0100;
															assign node6680 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node6683 = (inp[12]) ? node6685 : 4'b0000;
															assign node6685 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node6688 = (inp[10]) ? 4'b0100 : node6689;
														assign node6689 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node6693 = (inp[11]) ? node6723 : node6694;
												assign node6694 = (inp[4]) ? node6706 : node6695;
													assign node6695 = (inp[13]) ? node6701 : node6696;
														assign node6696 = (inp[12]) ? 4'b0001 : node6697;
															assign node6697 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node6701 = (inp[10]) ? node6703 : 4'b1001;
															assign node6703 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node6706 = (inp[7]) ? node6716 : node6707;
														assign node6707 = (inp[12]) ? 4'b0101 : node6708;
															assign node6708 = (inp[13]) ? node6712 : node6709;
																assign node6709 = (inp[10]) ? 4'b1101 : 4'b0101;
																assign node6712 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node6716 = (inp[12]) ? node6720 : node6717;
															assign node6717 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node6720 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node6723 = (inp[13]) ? node6733 : node6724;
													assign node6724 = (inp[4]) ? node6730 : node6725;
														assign node6725 = (inp[12]) ? node6727 : 4'b1000;
															assign node6727 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node6730 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node6733 = (inp[7]) ? node6735 : 4'b0100;
														assign node6735 = (inp[12]) ? node6739 : node6736;
															assign node6736 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node6739 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node6742 = (inp[13]) ? node6784 : node6743;
											assign node6743 = (inp[11]) ? node6773 : node6744;
												assign node6744 = (inp[14]) ? node6756 : node6745;
													assign node6745 = (inp[7]) ? 4'b1001 : node6746;
														assign node6746 = (inp[4]) ? node6752 : node6747;
															assign node6747 = (inp[10]) ? 4'b1001 : node6748;
																assign node6748 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node6752 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node6756 = (inp[10]) ? node6768 : node6757;
														assign node6757 = (inp[12]) ? node6763 : node6758;
															assign node6758 = (inp[7]) ? 4'b1000 : node6759;
																assign node6759 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node6763 = (inp[4]) ? node6765 : 4'b0000;
																assign node6765 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node6768 = (inp[7]) ? 4'b1000 : node6769;
															assign node6769 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node6773 = (inp[7]) ? node6779 : node6774;
													assign node6774 = (inp[4]) ? 4'b1101 : node6775;
														assign node6775 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node6779 = (inp[10]) ? 4'b1001 : node6780;
														assign node6780 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node6784 = (inp[12]) ? node6798 : node6785;
												assign node6785 = (inp[7]) ? node6791 : node6786;
													assign node6786 = (inp[14]) ? node6788 : 4'b0101;
														assign node6788 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node6791 = (inp[4]) ? node6793 : 4'b0001;
														assign node6793 = (inp[11]) ? 4'b0101 : node6794;
															assign node6794 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node6798 = (inp[10]) ? node6814 : node6799;
													assign node6799 = (inp[11]) ? node6809 : node6800;
														assign node6800 = (inp[14]) ? node6804 : node6801;
															assign node6801 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node6804 = (inp[4]) ? node6806 : 4'b1000;
																assign node6806 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node6809 = (inp[7]) ? 4'b1001 : node6810;
															assign node6810 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node6814 = (inp[4]) ? node6822 : node6815;
														assign node6815 = (inp[7]) ? node6817 : 4'b0101;
															assign node6817 = (inp[14]) ? node6819 : 4'b0001;
																assign node6819 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node6822 = (inp[11]) ? 4'b0101 : node6823;
															assign node6823 = (inp[7]) ? 4'b0100 : 4'b0101;
					assign node6828 = (inp[5]) ? node7850 : node6829;
						assign node6829 = (inp[0]) ? node7555 : node6830;
							assign node6830 = (inp[11]) ? node7246 : node6831;
								assign node6831 = (inp[10]) ? node7049 : node6832;
									assign node6832 = (inp[3]) ? node6954 : node6833;
										assign node6833 = (inp[4]) ? node6897 : node6834;
											assign node6834 = (inp[7]) ? node6864 : node6835;
												assign node6835 = (inp[13]) ? node6845 : node6836;
													assign node6836 = (inp[12]) ? node6840 : node6837;
														assign node6837 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node6840 = (inp[14]) ? 4'b0100 : node6841;
															assign node6841 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node6845 = (inp[2]) ? node6851 : node6846;
														assign node6846 = (inp[1]) ? 4'b1000 : node6847;
															assign node6847 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node6851 = (inp[12]) ? node6859 : node6852;
															assign node6852 = (inp[1]) ? node6856 : node6853;
																assign node6853 = (inp[14]) ? 4'b1101 : 4'b0000;
																assign node6856 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6859 = (inp[1]) ? node6861 : 4'b1100;
																assign node6861 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node6864 = (inp[13]) ? node6882 : node6865;
													assign node6865 = (inp[12]) ? node6873 : node6866;
														assign node6866 = (inp[2]) ? 4'b0101 : node6867;
															assign node6867 = (inp[14]) ? 4'b1100 : node6868;
																assign node6868 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node6873 = (inp[2]) ? 4'b0101 : node6874;
															assign node6874 = (inp[1]) ? node6878 : node6875;
																assign node6875 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node6878 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node6882 = (inp[12]) ? node6890 : node6883;
														assign node6883 = (inp[14]) ? node6887 : node6884;
															assign node6884 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node6887 = (inp[1]) ? 4'b0100 : 4'b1101;
														assign node6890 = (inp[14]) ? node6894 : node6891;
															assign node6891 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node6894 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node6897 = (inp[2]) ? node6915 : node6898;
												assign node6898 = (inp[13]) ? node6904 : node6899;
													assign node6899 = (inp[12]) ? node6901 : 4'b1000;
														assign node6901 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node6904 = (inp[7]) ? node6910 : node6905;
														assign node6905 = (inp[12]) ? node6907 : 4'b1100;
															assign node6907 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node6910 = (inp[14]) ? 4'b1000 : node6911;
															assign node6911 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node6915 = (inp[7]) ? node6935 : node6916;
													assign node6916 = (inp[13]) ? node6926 : node6917;
														assign node6917 = (inp[12]) ? node6921 : node6918;
															assign node6918 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node6921 = (inp[1]) ? 4'b0000 : node6922;
																assign node6922 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6926 = (inp[12]) ? node6928 : 4'b0000;
															assign node6928 = (inp[14]) ? node6932 : node6929;
																assign node6929 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node6932 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node6935 = (inp[13]) ? node6943 : node6936;
														assign node6936 = (inp[1]) ? node6940 : node6937;
															assign node6937 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node6940 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node6943 = (inp[12]) ? node6949 : node6944;
															assign node6944 = (inp[14]) ? 4'b1101 : node6945;
																assign node6945 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node6949 = (inp[1]) ? node6951 : 4'b1101;
																assign node6951 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node6954 = (inp[2]) ? node7006 : node6955;
											assign node6955 = (inp[4]) ? node6969 : node6956;
												assign node6956 = (inp[7]) ? node6964 : node6957;
													assign node6957 = (inp[13]) ? node6959 : 4'b1100;
														assign node6959 = (inp[12]) ? node6961 : 4'b1000;
															assign node6961 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node6964 = (inp[1]) ? 4'b1100 : node6965;
														assign node6965 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node6969 = (inp[13]) ? node6987 : node6970;
													assign node6970 = (inp[7]) ? node6980 : node6971;
														assign node6971 = (inp[12]) ? node6977 : node6972;
															assign node6972 = (inp[14]) ? node6974 : 4'b0000;
																assign node6974 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node6977 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6980 = (inp[14]) ? node6984 : node6981;
															assign node6981 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node6984 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6987 = (inp[7]) ? node6997 : node6988;
														assign node6988 = (inp[12]) ? 4'b0100 : node6989;
															assign node6989 = (inp[1]) ? node6993 : node6990;
																assign node6990 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node6993 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node6997 = (inp[1]) ? node7003 : node6998;
															assign node6998 = (inp[12]) ? 4'b1001 : node6999;
																assign node6999 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node7003 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node7006 = (inp[4]) ? node7036 : node7007;
												assign node7007 = (inp[13]) ? node7019 : node7008;
													assign node7008 = (inp[12]) ? node7016 : node7009;
														assign node7009 = (inp[14]) ? node7013 : node7010;
															assign node7010 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node7013 = (inp[1]) ? 4'b1000 : 4'b0001;
														assign node7016 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node7019 = (inp[1]) ? node7027 : node7020;
														assign node7020 = (inp[12]) ? node7024 : node7021;
															assign node7021 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node7024 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node7027 = (inp[14]) ? node7033 : node7028;
															assign node7028 = (inp[7]) ? node7030 : 4'b1000;
																assign node7030 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node7033 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node7036 = (inp[13]) ? node7042 : node7037;
													assign node7037 = (inp[12]) ? node7039 : 4'b1000;
														assign node7039 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node7042 = (inp[7]) ? 4'b1000 : node7043;
														assign node7043 = (inp[1]) ? 4'b1100 : node7044;
															assign node7044 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node7049 = (inp[12]) ? node7141 : node7050;
										assign node7050 = (inp[13]) ? node7100 : node7051;
											assign node7051 = (inp[3]) ? node7075 : node7052;
												assign node7052 = (inp[2]) ? node7064 : node7053;
													assign node7053 = (inp[7]) ? node7057 : node7054;
														assign node7054 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7057 = (inp[4]) ? 4'b0000 : node7058;
															assign node7058 = (inp[14]) ? node7060 : 4'b1101;
																assign node7060 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node7064 = (inp[1]) ? node7068 : node7065;
														assign node7065 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node7068 = (inp[14]) ? node7070 : 4'b1101;
															assign node7070 = (inp[4]) ? node7072 : 4'b1100;
																assign node7072 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node7075 = (inp[7]) ? node7083 : node7076;
													assign node7076 = (inp[4]) ? node7078 : 4'b0000;
														assign node7078 = (inp[2]) ? 4'b0100 : node7079;
															assign node7079 = (inp[1]) ? 4'b1000 : 4'b0001;
													assign node7083 = (inp[4]) ? node7091 : node7084;
														assign node7084 = (inp[2]) ? node7086 : 4'b0100;
															assign node7086 = (inp[14]) ? node7088 : 4'b1000;
																assign node7088 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7091 = (inp[2]) ? 4'b0000 : node7092;
															assign node7092 = (inp[1]) ? node7096 : node7093;
																assign node7093 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node7096 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node7100 = (inp[4]) ? node7122 : node7101;
												assign node7101 = (inp[3]) ? node7115 : node7102;
													assign node7102 = (inp[2]) ? node7104 : 4'b0000;
														assign node7104 = (inp[7]) ? node7110 : node7105;
															assign node7105 = (inp[14]) ? node7107 : 4'b0000;
																assign node7107 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node7110 = (inp[14]) ? 4'b0100 : node7111;
																assign node7111 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node7115 = (inp[2]) ? 4'b0000 : node7116;
														assign node7116 = (inp[7]) ? 4'b0000 : node7117;
															assign node7117 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node7122 = (inp[2]) ? node7132 : node7123;
													assign node7123 = (inp[3]) ? node7125 : 4'b0100;
														assign node7125 = (inp[1]) ? node7129 : node7126;
															assign node7126 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node7129 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node7132 = (inp[3]) ? 4'b0100 : node7133;
														assign node7133 = (inp[7]) ? 4'b0001 : node7134;
															assign node7134 = (inp[14]) ? node7136 : 4'b0001;
																assign node7136 = (inp[1]) ? 4'b0000 : 4'b0001;
										assign node7141 = (inp[1]) ? node7197 : node7142;
											assign node7142 = (inp[4]) ? node7164 : node7143;
												assign node7143 = (inp[14]) ? node7153 : node7144;
													assign node7144 = (inp[13]) ? node7150 : node7145;
														assign node7145 = (inp[3]) ? node7147 : 4'b1100;
															assign node7147 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node7150 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node7153 = (inp[3]) ? node7157 : node7154;
														assign node7154 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node7157 = (inp[2]) ? node7159 : 4'b1100;
															assign node7159 = (inp[13]) ? node7161 : 4'b0001;
																assign node7161 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node7164 = (inp[13]) ? node7174 : node7165;
													assign node7165 = (inp[14]) ? node7167 : 4'b1000;
														assign node7167 = (inp[2]) ? node7171 : node7168;
															assign node7168 = (inp[3]) ? 4'b0000 : 4'b1000;
															assign node7171 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node7174 = (inp[7]) ? node7184 : node7175;
														assign node7175 = (inp[2]) ? node7181 : node7176;
															assign node7176 = (inp[14]) ? 4'b1100 : node7177;
																assign node7177 = (inp[3]) ? 4'b1101 : 4'b1100;
															assign node7181 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node7184 = (inp[3]) ? node7192 : node7185;
															assign node7185 = (inp[14]) ? node7189 : node7186;
																assign node7186 = (inp[2]) ? 4'b0000 : 4'b1000;
																assign node7189 = (inp[2]) ? 4'b1101 : 4'b1000;
															assign node7192 = (inp[2]) ? 4'b1000 : node7193;
																assign node7193 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node7197 = (inp[13]) ? node7223 : node7198;
												assign node7198 = (inp[2]) ? node7208 : node7199;
													assign node7199 = (inp[7]) ? node7203 : node7200;
														assign node7200 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7203 = (inp[4]) ? node7205 : 4'b1101;
															assign node7205 = (inp[3]) ? 4'b0001 : 4'b0000;
													assign node7208 = (inp[3]) ? node7214 : node7209;
														assign node7209 = (inp[7]) ? 4'b1100 : node7210;
															assign node7210 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node7214 = (inp[4]) ? node7220 : node7215;
															assign node7215 = (inp[14]) ? node7217 : 4'b1001;
																assign node7217 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node7220 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7223 = (inp[4]) ? node7235 : node7224;
													assign node7224 = (inp[3]) ? 4'b0000 : node7225;
														assign node7225 = (inp[14]) ? node7231 : node7226;
															assign node7226 = (inp[2]) ? node7228 : 4'b0000;
																assign node7228 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node7231 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node7235 = (inp[2]) ? node7241 : node7236;
														assign node7236 = (inp[3]) ? node7238 : 4'b0100;
															assign node7238 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node7241 = (inp[3]) ? 4'b0100 : node7242;
															assign node7242 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node7246 = (inp[1]) ? node7440 : node7247;
									assign node7247 = (inp[3]) ? node7341 : node7248;
										assign node7248 = (inp[2]) ? node7302 : node7249;
											assign node7249 = (inp[4]) ? node7281 : node7250;
												assign node7250 = (inp[7]) ? node7264 : node7251;
													assign node7251 = (inp[13]) ? node7253 : 4'b1100;
														assign node7253 = (inp[14]) ? node7259 : node7254;
															assign node7254 = (inp[10]) ? node7256 : 4'b1001;
																assign node7256 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node7259 = (inp[12]) ? node7261 : 4'b0001;
																assign node7261 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7264 = (inp[13]) ? node7270 : node7265;
														assign node7265 = (inp[10]) ? 4'b1100 : node7266;
															assign node7266 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7270 = (inp[14]) ? node7276 : node7271;
															assign node7271 = (inp[10]) ? 4'b0100 : node7272;
																assign node7272 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node7276 = (inp[12]) ? 4'b0100 : node7277;
																assign node7277 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node7281 = (inp[13]) ? node7289 : node7282;
													assign node7282 = (inp[12]) ? node7286 : node7283;
														assign node7283 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node7286 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7289 = (inp[7]) ? node7295 : node7290;
														assign node7290 = (inp[12]) ? node7292 : 4'b0101;
															assign node7292 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node7295 = (inp[14]) ? node7297 : 4'b1001;
															assign node7297 = (inp[12]) ? node7299 : 4'b0101;
																assign node7299 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node7302 = (inp[4]) ? node7320 : node7303;
												assign node7303 = (inp[13]) ? node7309 : node7304;
													assign node7304 = (inp[10]) ? 4'b1100 : node7305;
														assign node7305 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node7309 = (inp[7]) ? node7315 : node7310;
														assign node7310 = (inp[12]) ? node7312 : 4'b0000;
															assign node7312 = (inp[14]) ? 4'b1100 : 4'b0000;
														assign node7315 = (inp[10]) ? 4'b0100 : node7316;
															assign node7316 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node7320 = (inp[7]) ? node7334 : node7321;
													assign node7321 = (inp[10]) ? node7331 : node7322;
														assign node7322 = (inp[14]) ? node7328 : node7323;
															assign node7323 = (inp[12]) ? 4'b0000 : node7324;
																assign node7324 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node7328 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node7331 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node7334 = (inp[10]) ? 4'b0000 : node7335;
														assign node7335 = (inp[12]) ? node7337 : 4'b0000;
															assign node7337 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node7341 = (inp[2]) ? node7385 : node7342;
											assign node7342 = (inp[4]) ? node7364 : node7343;
												assign node7343 = (inp[10]) ? node7355 : node7344;
													assign node7344 = (inp[12]) ? node7350 : node7345;
														assign node7345 = (inp[7]) ? 4'b1101 : node7346;
															assign node7346 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node7350 = (inp[7]) ? 4'b0101 : node7351;
															assign node7351 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node7355 = (inp[12]) ? node7361 : node7356;
														assign node7356 = (inp[13]) ? node7358 : 4'b0001;
															assign node7358 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node7361 = (inp[13]) ? 4'b1001 : 4'b1101;
												assign node7364 = (inp[13]) ? node7374 : node7365;
													assign node7365 = (inp[12]) ? node7369 : node7366;
														assign node7366 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node7369 = (inp[10]) ? 4'b0000 : node7370;
															assign node7370 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node7374 = (inp[12]) ? node7380 : node7375;
														assign node7375 = (inp[10]) ? 4'b0100 : node7376;
															assign node7376 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7380 = (inp[10]) ? node7382 : 4'b0000;
															assign node7382 = (inp[14]) ? 4'b1000 : 4'b1100;
											assign node7385 = (inp[4]) ? node7411 : node7386;
												assign node7386 = (inp[7]) ? node7400 : node7387;
													assign node7387 = (inp[13]) ? node7393 : node7388;
														assign node7388 = (inp[12]) ? node7390 : 4'b0001;
															assign node7390 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7393 = (inp[12]) ? node7397 : node7394;
															assign node7394 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node7397 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7400 = (inp[13]) ? node7406 : node7401;
														assign node7401 = (inp[12]) ? node7403 : 4'b1000;
															assign node7403 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node7406 = (inp[12]) ? 4'b1000 : node7407;
															assign node7407 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node7411 = (inp[7]) ? node7425 : node7412;
													assign node7412 = (inp[13]) ? node7420 : node7413;
														assign node7413 = (inp[10]) ? node7417 : node7414;
															assign node7414 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7417 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node7420 = (inp[14]) ? 4'b1101 : node7421;
															assign node7421 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node7425 = (inp[14]) ? node7435 : node7426;
														assign node7426 = (inp[10]) ? node7430 : node7427;
															assign node7427 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7430 = (inp[13]) ? 4'b0101 : node7431;
																assign node7431 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7435 = (inp[10]) ? 4'b1001 : node7436;
															assign node7436 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node7440 = (inp[10]) ? node7516 : node7441;
										assign node7441 = (inp[4]) ? node7477 : node7442;
											assign node7442 = (inp[3]) ? node7458 : node7443;
												assign node7443 = (inp[13]) ? node7447 : node7444;
													assign node7444 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node7447 = (inp[12]) ? node7453 : node7448;
														assign node7448 = (inp[7]) ? 4'b0101 : node7449;
															assign node7449 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node7453 = (inp[14]) ? node7455 : 4'b1101;
															assign node7455 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node7458 = (inp[2]) ? node7464 : node7459;
													assign node7459 = (inp[7]) ? 4'b1101 : node7460;
														assign node7460 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node7464 = (inp[14]) ? node7472 : node7465;
														assign node7465 = (inp[13]) ? node7469 : node7466;
															assign node7466 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7469 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7472 = (inp[13]) ? node7474 : 4'b0001;
															assign node7474 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node7477 = (inp[3]) ? node7499 : node7478;
												assign node7478 = (inp[2]) ? node7484 : node7479;
													assign node7479 = (inp[13]) ? node7481 : 4'b1001;
														assign node7481 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7484 = (inp[7]) ? node7492 : node7485;
														assign node7485 = (inp[12]) ? node7489 : node7486;
															assign node7486 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node7489 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node7492 = (inp[13]) ? node7496 : node7493;
															assign node7493 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7496 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node7499 = (inp[2]) ? node7511 : node7500;
													assign node7500 = (inp[13]) ? node7504 : node7501;
														assign node7501 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7504 = (inp[7]) ? node7508 : node7505;
															assign node7505 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7508 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7511 = (inp[13]) ? node7513 : 4'b1001;
														assign node7513 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node7516 = (inp[13]) ? node7542 : node7517;
											assign node7517 = (inp[3]) ? node7531 : node7518;
												assign node7518 = (inp[2]) ? node7526 : node7519;
													assign node7519 = (inp[4]) ? node7523 : node7520;
														assign node7520 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node7523 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node7526 = (inp[7]) ? 4'b1101 : node7527;
														assign node7527 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node7531 = (inp[4]) ? node7537 : node7532;
													assign node7532 = (inp[7]) ? node7534 : 4'b0001;
														assign node7534 = (inp[2]) ? 4'b1001 : 4'b0101;
													assign node7537 = (inp[2]) ? node7539 : 4'b1001;
														assign node7539 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node7542 = (inp[4]) ? node7550 : node7543;
												assign node7543 = (inp[7]) ? node7545 : 4'b0001;
													assign node7545 = (inp[3]) ? 4'b0001 : node7546;
														assign node7546 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node7550 = (inp[2]) ? node7552 : 4'b0101;
													assign node7552 = (inp[3]) ? 4'b0101 : 4'b0001;
							assign node7555 = (inp[2]) ? 4'b0101 : node7556;
								assign node7556 = (inp[3]) ? node7654 : node7557;
									assign node7557 = (inp[4]) ? node7579 : node7558;
										assign node7558 = (inp[13]) ? node7560 : 4'b0101;
											assign node7560 = (inp[7]) ? 4'b0101 : node7561;
												assign node7561 = (inp[1]) ? node7573 : node7562;
													assign node7562 = (inp[11]) ? node7568 : node7563;
														assign node7563 = (inp[14]) ? 4'b0101 : node7564;
															assign node7564 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node7568 = (inp[12]) ? node7570 : 4'b0000;
															assign node7570 = (inp[10]) ? 4'b0000 : 4'b0101;
													assign node7573 = (inp[12]) ? node7575 : 4'b0001;
														assign node7575 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node7579 = (inp[7]) ? node7635 : node7580;
											assign node7580 = (inp[1]) ? node7608 : node7581;
												assign node7581 = (inp[14]) ? node7593 : node7582;
													assign node7582 = (inp[13]) ? node7588 : node7583;
														assign node7583 = (inp[10]) ? 4'b1000 : node7584;
															assign node7584 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7588 = (inp[12]) ? node7590 : 4'b0000;
															assign node7590 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node7593 = (inp[11]) ? node7603 : node7594;
														assign node7594 = (inp[12]) ? 4'b1001 : node7595;
															assign node7595 = (inp[13]) ? node7599 : node7596;
																assign node7596 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node7599 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node7603 = (inp[13]) ? 4'b0000 : node7604;
															assign node7604 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node7608 = (inp[14]) ? node7620 : node7609;
													assign node7609 = (inp[13]) ? node7615 : node7610;
														assign node7610 = (inp[10]) ? 4'b1001 : node7611;
															assign node7611 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7615 = (inp[12]) ? node7617 : 4'b0001;
															assign node7617 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node7620 = (inp[11]) ? node7630 : node7621;
														assign node7621 = (inp[10]) ? node7627 : node7622;
															assign node7622 = (inp[12]) ? node7624 : 4'b1000;
																assign node7624 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node7627 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node7630 = (inp[13]) ? 4'b0001 : node7631;
															assign node7631 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node7635 = (inp[13]) ? node7637 : 4'b0101;
												assign node7637 = (inp[10]) ? node7645 : node7638;
													assign node7638 = (inp[12]) ? 4'b0101 : node7639;
														assign node7639 = (inp[14]) ? 4'b0101 : node7640;
															assign node7640 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node7645 = (inp[1]) ? node7649 : node7646;
														assign node7646 = (inp[11]) ? 4'b0000 : 4'b0101;
														assign node7649 = (inp[11]) ? 4'b0001 : node7650;
															assign node7650 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node7654 = (inp[4]) ? node7728 : node7655;
										assign node7655 = (inp[1]) ? node7689 : node7656;
											assign node7656 = (inp[11]) ? node7672 : node7657;
												assign node7657 = (inp[14]) ? node7665 : node7658;
													assign node7658 = (inp[13]) ? node7660 : 4'b1000;
														assign node7660 = (inp[7]) ? node7662 : 4'b0100;
															assign node7662 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node7665 = (inp[13]) ? 4'b1001 : node7666;
														assign node7666 = (inp[10]) ? node7668 : 4'b0001;
															assign node7668 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node7672 = (inp[13]) ? node7678 : node7673;
													assign node7673 = (inp[12]) ? node7675 : 4'b1000;
														assign node7675 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node7678 = (inp[7]) ? node7684 : node7679;
														assign node7679 = (inp[12]) ? node7681 : 4'b0100;
															assign node7681 = (inp[14]) ? 4'b0100 : 4'b1000;
														assign node7684 = (inp[10]) ? 4'b0000 : node7685;
															assign node7685 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node7689 = (inp[13]) ? node7705 : node7690;
												assign node7690 = (inp[11]) ? node7700 : node7691;
													assign node7691 = (inp[14]) ? node7695 : node7692;
														assign node7692 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7695 = (inp[10]) ? 4'b1000 : node7696;
															assign node7696 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7700 = (inp[10]) ? 4'b1001 : node7701;
														assign node7701 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node7705 = (inp[7]) ? node7715 : node7706;
													assign node7706 = (inp[12]) ? node7712 : node7707;
														assign node7707 = (inp[11]) ? 4'b0101 : node7708;
															assign node7708 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node7712 = (inp[11]) ? 4'b1001 : 4'b0100;
													assign node7715 = (inp[11]) ? node7723 : node7716;
														assign node7716 = (inp[14]) ? node7718 : 4'b0001;
															assign node7718 = (inp[10]) ? 4'b0000 : node7719;
																assign node7719 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node7723 = (inp[12]) ? node7725 : 4'b0001;
															assign node7725 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node7728 = (inp[7]) ? node7790 : node7729;
											assign node7729 = (inp[1]) ? node7757 : node7730;
												assign node7730 = (inp[14]) ? node7744 : node7731;
													assign node7731 = (inp[10]) ? 4'b1100 : node7732;
														assign node7732 = (inp[11]) ? node7738 : node7733;
															assign node7733 = (inp[12]) ? node7735 : 4'b1100;
																assign node7735 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node7738 = (inp[12]) ? 4'b0100 : node7739;
																assign node7739 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node7744 = (inp[11]) ? node7752 : node7745;
														assign node7745 = (inp[13]) ? node7749 : node7746;
															assign node7746 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node7749 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node7752 = (inp[13]) ? 4'b0100 : node7753;
															assign node7753 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node7757 = (inp[11]) ? node7777 : node7758;
													assign node7758 = (inp[14]) ? node7768 : node7759;
														assign node7759 = (inp[10]) ? 4'b1101 : node7760;
															assign node7760 = (inp[12]) ? node7764 : node7761;
																assign node7761 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node7764 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node7768 = (inp[12]) ? node7770 : 4'b0100;
															assign node7770 = (inp[13]) ? node7774 : node7771;
																assign node7771 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node7774 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node7777 = (inp[13]) ? node7783 : node7778;
														assign node7778 = (inp[10]) ? 4'b1101 : node7779;
															assign node7779 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7783 = (inp[14]) ? 4'b0101 : node7784;
															assign node7784 = (inp[10]) ? 4'b0101 : node7785;
																assign node7785 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node7790 = (inp[13]) ? node7818 : node7791;
												assign node7791 = (inp[12]) ? node7803 : node7792;
													assign node7792 = (inp[1]) ? node7798 : node7793;
														assign node7793 = (inp[10]) ? 4'b1000 : node7794;
															assign node7794 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node7798 = (inp[11]) ? 4'b1001 : node7799;
															assign node7799 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7803 = (inp[10]) ? node7811 : node7804;
														assign node7804 = (inp[11]) ? 4'b0001 : node7805;
															assign node7805 = (inp[14]) ? node7807 : 4'b0001;
																assign node7807 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node7811 = (inp[11]) ? 4'b1000 : node7812;
															assign node7812 = (inp[14]) ? 4'b0001 : node7813;
																assign node7813 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node7818 = (inp[10]) ? node7836 : node7819;
													assign node7819 = (inp[12]) ? node7829 : node7820;
														assign node7820 = (inp[1]) ? node7824 : node7821;
															assign node7821 = (inp[14]) ? 4'b1001 : 4'b0100;
															assign node7824 = (inp[11]) ? 4'b0101 : node7825;
																assign node7825 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node7829 = (inp[1]) ? 4'b1001 : node7830;
															assign node7830 = (inp[14]) ? node7832 : 4'b1000;
																assign node7832 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node7836 = (inp[1]) ? node7844 : node7837;
														assign node7837 = (inp[14]) ? node7839 : 4'b0100;
															assign node7839 = (inp[12]) ? 4'b1001 : node7840;
																assign node7840 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node7844 = (inp[11]) ? 4'b0101 : node7845;
															assign node7845 = (inp[14]) ? 4'b0100 : 4'b0101;
						assign node7850 = (inp[3]) ? node8504 : node7851;
							assign node7851 = (inp[4]) ? node8143 : node7852;
								assign node7852 = (inp[13]) ? node8006 : node7853;
									assign node7853 = (inp[0]) ? node7943 : node7854;
										assign node7854 = (inp[7]) ? node7898 : node7855;
											assign node7855 = (inp[10]) ? node7877 : node7856;
												assign node7856 = (inp[12]) ? node7866 : node7857;
													assign node7857 = (inp[1]) ? node7859 : 4'b1100;
														assign node7859 = (inp[11]) ? 4'b0001 : node7860;
															assign node7860 = (inp[14]) ? 4'b1100 : node7861;
																assign node7861 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node7866 = (inp[1]) ? node7872 : node7867;
														assign node7867 = (inp[11]) ? node7869 : 4'b0100;
															assign node7869 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node7872 = (inp[11]) ? 4'b1101 : node7873;
															assign node7873 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node7877 = (inp[2]) ? node7885 : node7878;
													assign node7878 = (inp[1]) ? 4'b0001 : node7879;
														assign node7879 = (inp[12]) ? node7881 : 4'b1001;
															assign node7881 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node7885 = (inp[1]) ? node7893 : node7886;
														assign node7886 = (inp[11]) ? node7890 : node7887;
															assign node7887 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node7890 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7893 = (inp[11]) ? 4'b1001 : node7894;
															assign node7894 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node7898 = (inp[10]) ? node7920 : node7899;
												assign node7899 = (inp[11]) ? node7909 : node7900;
													assign node7900 = (inp[2]) ? 4'b1100 : node7901;
														assign node7901 = (inp[1]) ? 4'b1101 : node7902;
															assign node7902 = (inp[12]) ? 4'b0100 : node7903;
																assign node7903 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7909 = (inp[2]) ? node7915 : node7910;
														assign node7910 = (inp[1]) ? node7912 : 4'b1100;
															assign node7912 = (inp[14]) ? 4'b1101 : 4'b0101;
														assign node7915 = (inp[12]) ? node7917 : 4'b1101;
															assign node7917 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node7920 = (inp[1]) ? node7934 : node7921;
													assign node7921 = (inp[11]) ? node7927 : node7922;
														assign node7922 = (inp[2]) ? node7924 : 4'b0101;
															assign node7924 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node7927 = (inp[2]) ? node7931 : node7928;
															assign node7928 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node7931 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node7934 = (inp[2]) ? node7940 : node7935;
														assign node7935 = (inp[12]) ? node7937 : 4'b0001;
															assign node7937 = (inp[11]) ? 4'b0001 : 4'b1100;
														assign node7940 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node7943 = (inp[2]) ? 4'b0101 : node7944;
											assign node7944 = (inp[7]) ? node7978 : node7945;
												assign node7945 = (inp[10]) ? node7967 : node7946;
													assign node7946 = (inp[12]) ? node7958 : node7947;
														assign node7947 = (inp[1]) ? node7953 : node7948;
															assign node7948 = (inp[14]) ? node7950 : 4'b1100;
																assign node7950 = (inp[11]) ? 4'b1100 : 4'b0101;
															assign node7953 = (inp[14]) ? node7955 : 4'b1101;
																assign node7955 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node7958 = (inp[11]) ? 4'b0101 : node7959;
															assign node7959 = (inp[14]) ? node7963 : node7960;
																assign node7960 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node7963 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node7967 = (inp[11]) ? node7973 : node7968;
														assign node7968 = (inp[12]) ? node7970 : 4'b0000;
															assign node7970 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node7973 = (inp[12]) ? node7975 : 4'b0001;
															assign node7975 = (inp[1]) ? 4'b0001 : 4'b1100;
												assign node7978 = (inp[1]) ? node7990 : node7979;
													assign node7979 = (inp[11]) ? 4'b1100 : node7980;
														assign node7980 = (inp[14]) ? node7986 : node7981;
															assign node7981 = (inp[12]) ? node7983 : 4'b1100;
																assign node7983 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node7986 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node7990 = (inp[10]) ? node8000 : node7991;
														assign node7991 = (inp[12]) ? node7995 : node7992;
															assign node7992 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node7995 = (inp[11]) ? 4'b0101 : node7996;
																assign node7996 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node8000 = (inp[11]) ? 4'b1101 : node8001;
															assign node8001 = (inp[14]) ? 4'b1100 : 4'b1101;
									assign node8006 = (inp[0]) ? node8088 : node8007;
										assign node8007 = (inp[2]) ? node8051 : node8008;
											assign node8008 = (inp[1]) ? node8024 : node8009;
												assign node8009 = (inp[7]) ? node8019 : node8010;
													assign node8010 = (inp[10]) ? node8014 : node8011;
														assign node8011 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node8014 = (inp[11]) ? 4'b1101 : node8015;
															assign node8015 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node8019 = (inp[12]) ? node8021 : 4'b1001;
														assign node8021 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node8024 = (inp[12]) ? node8040 : node8025;
													assign node8025 = (inp[11]) ? 4'b0001 : node8026;
														assign node8026 = (inp[14]) ? node8032 : node8027;
															assign node8027 = (inp[7]) ? 4'b0101 : node8028;
																assign node8028 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node8032 = (inp[7]) ? node8036 : node8033;
																assign node8033 = (inp[10]) ? 4'b0000 : 4'b0101;
																assign node8036 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node8040 = (inp[11]) ? node8046 : node8041;
														assign node8041 = (inp[7]) ? 4'b1001 : node8042;
															assign node8042 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node8046 = (inp[14]) ? 4'b0001 : node8047;
															assign node8047 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node8051 = (inp[1]) ? node8063 : node8052;
												assign node8052 = (inp[11]) ? node8058 : node8053;
													assign node8053 = (inp[14]) ? 4'b1000 : node8054;
														assign node8054 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8058 = (inp[10]) ? node8060 : 4'b0000;
														assign node8060 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8063 = (inp[10]) ? node8077 : node8064;
													assign node8064 = (inp[14]) ? node8072 : node8065;
														assign node8065 = (inp[12]) ? node8069 : node8066;
															assign node8066 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node8069 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node8072 = (inp[11]) ? node8074 : 4'b0001;
															assign node8074 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8077 = (inp[7]) ? node8083 : node8078;
														assign node8078 = (inp[11]) ? 4'b0101 : node8079;
															assign node8079 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node8083 = (inp[11]) ? 4'b0001 : node8084;
															assign node8084 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node8088 = (inp[2]) ? node8122 : node8089;
											assign node8089 = (inp[10]) ? node8109 : node8090;
												assign node8090 = (inp[7]) ? node8100 : node8091;
													assign node8091 = (inp[11]) ? node8095 : node8092;
														assign node8092 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8095 = (inp[1]) ? 4'b1001 : node8096;
															assign node8096 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8100 = (inp[12]) ? node8106 : node8101;
														assign node8101 = (inp[1]) ? node8103 : 4'b0100;
															assign node8103 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node8106 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node8109 = (inp[11]) ? node8117 : node8110;
													assign node8110 = (inp[1]) ? 4'b0000 : node8111;
														assign node8111 = (inp[12]) ? node8113 : 4'b0000;
															assign node8113 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node8117 = (inp[1]) ? 4'b0001 : node8118;
														assign node8118 = (inp[12]) ? 4'b0100 : 4'b0001;
											assign node8122 = (inp[7]) ? 4'b0101 : node8123;
												assign node8123 = (inp[12]) ? node8133 : node8124;
													assign node8124 = (inp[1]) ? node8130 : node8125;
														assign node8125 = (inp[14]) ? node8127 : 4'b0000;
															assign node8127 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node8130 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8133 = (inp[10]) ? node8135 : 4'b0101;
														assign node8135 = (inp[14]) ? node8139 : node8136;
															assign node8136 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node8139 = (inp[1]) ? 4'b0000 : 4'b0101;
								assign node8143 = (inp[1]) ? node8353 : node8144;
									assign node8144 = (inp[7]) ? node8246 : node8145;
										assign node8145 = (inp[0]) ? node8187 : node8146;
											assign node8146 = (inp[2]) ? node8164 : node8147;
												assign node8147 = (inp[10]) ? node8157 : node8148;
													assign node8148 = (inp[13]) ? node8154 : node8149;
														assign node8149 = (inp[11]) ? node8151 : 4'b1000;
															assign node8151 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node8154 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8157 = (inp[11]) ? 4'b0100 : node8158;
														assign node8158 = (inp[13]) ? node8160 : 4'b1001;
															assign node8160 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node8164 = (inp[11]) ? node8180 : node8165;
													assign node8165 = (inp[12]) ? node8173 : node8166;
														assign node8166 = (inp[13]) ? node8170 : node8167;
															assign node8167 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node8170 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8173 = (inp[13]) ? node8177 : node8174;
															assign node8174 = (inp[10]) ? 4'b0001 : 4'b0100;
															assign node8177 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node8180 = (inp[14]) ? 4'b1001 : node8181;
														assign node8181 = (inp[13]) ? node8183 : 4'b1100;
															assign node8183 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node8187 = (inp[13]) ? node8223 : node8188;
												assign node8188 = (inp[12]) ? node8204 : node8189;
													assign node8189 = (inp[2]) ? node8197 : node8190;
														assign node8190 = (inp[10]) ? node8194 : node8191;
															assign node8191 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node8194 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node8197 = (inp[10]) ? node8199 : 4'b1000;
															assign node8199 = (inp[11]) ? 4'b1000 : node8200;
																assign node8200 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8204 = (inp[10]) ? node8216 : node8205;
														assign node8205 = (inp[14]) ? node8211 : node8206;
															assign node8206 = (inp[2]) ? 4'b0000 : node8207;
																assign node8207 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node8211 = (inp[11]) ? node8213 : 4'b0001;
																assign node8213 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node8216 = (inp[11]) ? node8220 : node8217;
															assign node8217 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node8220 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node8223 = (inp[11]) ? node8237 : node8224;
													assign node8224 = (inp[14]) ? node8232 : node8225;
														assign node8225 = (inp[2]) ? node8227 : 4'b1001;
															assign node8227 = (inp[12]) ? node8229 : 4'b0000;
																assign node8229 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node8232 = (inp[2]) ? 4'b1001 : node8233;
															assign node8233 = (inp[12]) ? 4'b0100 : 4'b1000;
													assign node8237 = (inp[12]) ? node8239 : 4'b0000;
														assign node8239 = (inp[10]) ? node8243 : node8240;
															assign node8240 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node8243 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node8246 = (inp[2]) ? node8314 : node8247;
											assign node8247 = (inp[11]) ? node8283 : node8248;
												assign node8248 = (inp[0]) ? node8260 : node8249;
													assign node8249 = (inp[14]) ? node8253 : node8250;
														assign node8250 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node8253 = (inp[10]) ? 4'b1001 : node8254;
															assign node8254 = (inp[13]) ? 4'b1001 : node8255;
																assign node8255 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node8260 = (inp[13]) ? node8276 : node8261;
														assign node8261 = (inp[14]) ? node8269 : node8262;
															assign node8262 = (inp[10]) ? node8266 : node8263;
																assign node8263 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node8266 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node8269 = (inp[10]) ? node8273 : node8270;
																assign node8270 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node8273 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node8276 = (inp[10]) ? node8280 : node8277;
															assign node8277 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node8280 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node8283 = (inp[0]) ? node8293 : node8284;
													assign node8284 = (inp[10]) ? node8290 : node8285;
														assign node8285 = (inp[12]) ? node8287 : 4'b0000;
															assign node8287 = (inp[13]) ? 4'b0100 : 4'b1101;
														assign node8290 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node8293 = (inp[13]) ? node8305 : node8294;
														assign node8294 = (inp[14]) ? node8300 : node8295;
															assign node8295 = (inp[12]) ? node8297 : 4'b0001;
																assign node8297 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node8300 = (inp[12]) ? 4'b0001 : node8301;
																assign node8301 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8305 = (inp[14]) ? 4'b0000 : node8306;
															assign node8306 = (inp[10]) ? node8310 : node8307;
																assign node8307 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node8310 = (inp[12]) ? 4'b1001 : 4'b0000;
											assign node8314 = (inp[0]) ? node8340 : node8315;
												assign node8315 = (inp[13]) ? node8335 : node8316;
													assign node8316 = (inp[10]) ? node8328 : node8317;
														assign node8317 = (inp[14]) ? node8323 : node8318;
															assign node8318 = (inp[11]) ? 4'b1000 : node8319;
																assign node8319 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8323 = (inp[11]) ? 4'b1000 : node8324;
																assign node8324 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8328 = (inp[11]) ? node8332 : node8329;
															assign node8329 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8332 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node8335 = (inp[11]) ? 4'b1001 : node8336;
														assign node8336 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8340 = (inp[13]) ? node8342 : 4'b0101;
													assign node8342 = (inp[10]) ? node8346 : node8343;
														assign node8343 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node8346 = (inp[14]) ? node8348 : 4'b0000;
															assign node8348 = (inp[11]) ? 4'b0000 : node8349;
																assign node8349 = (inp[12]) ? 4'b0101 : 4'b0001;
									assign node8353 = (inp[11]) ? node8451 : node8354;
										assign node8354 = (inp[2]) ? node8398 : node8355;
											assign node8355 = (inp[10]) ? node8369 : node8356;
												assign node8356 = (inp[0]) ? node8364 : node8357;
													assign node8357 = (inp[13]) ? node8361 : node8358;
														assign node8358 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8361 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8364 = (inp[7]) ? 4'b1000 : node8365;
														assign node8365 = (inp[13]) ? 4'b0001 : 4'b1000;
												assign node8369 = (inp[0]) ? node8387 : node8370;
													assign node8370 = (inp[14]) ? node8378 : node8371;
														assign node8371 = (inp[7]) ? node8375 : node8372;
															assign node8372 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node8375 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8378 = (inp[7]) ? node8380 : 4'b0100;
															assign node8380 = (inp[12]) ? node8384 : node8381;
																assign node8381 = (inp[13]) ? 4'b0100 : 4'b1000;
																assign node8384 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8387 = (inp[14]) ? node8393 : node8388;
														assign node8388 = (inp[7]) ? 4'b0000 : node8389;
															assign node8389 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node8393 = (inp[12]) ? 4'b0100 : node8394;
															assign node8394 = (inp[13]) ? 4'b0001 : 4'b0100;
											assign node8398 = (inp[12]) ? node8416 : node8399;
												assign node8399 = (inp[0]) ? node8409 : node8400;
													assign node8400 = (inp[10]) ? 4'b0001 : node8401;
														assign node8401 = (inp[7]) ? node8403 : 4'b0101;
															assign node8403 = (inp[13]) ? 4'b0001 : node8404;
																assign node8404 = (inp[14]) ? 4'b1001 : 4'b0100;
													assign node8409 = (inp[14]) ? node8413 : node8410;
														assign node8410 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node8413 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node8416 = (inp[0]) ? node8436 : node8417;
													assign node8417 = (inp[13]) ? node8429 : node8418;
														assign node8418 = (inp[14]) ? node8426 : node8419;
															assign node8419 = (inp[10]) ? node8423 : node8420;
																assign node8420 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node8423 = (inp[7]) ? 4'b1100 : 4'b1001;
															assign node8426 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node8429 = (inp[10]) ? node8431 : 4'b1001;
															assign node8431 = (inp[7]) ? 4'b1001 : node8432;
																assign node8432 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node8436 = (inp[7]) ? node8444 : node8437;
														assign node8437 = (inp[14]) ? node8441 : node8438;
															assign node8438 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node8441 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node8444 = (inp[10]) ? node8446 : 4'b0101;
															assign node8446 = (inp[13]) ? node8448 : 4'b0101;
																assign node8448 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node8451 = (inp[10]) ? node8489 : node8452;
											assign node8452 = (inp[2]) ? node8468 : node8453;
												assign node8453 = (inp[12]) ? node8455 : 4'b1001;
													assign node8455 = (inp[7]) ? node8463 : node8456;
														assign node8456 = (inp[13]) ? node8460 : node8457;
															assign node8457 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node8460 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node8463 = (inp[0]) ? 4'b1001 : node8464;
															assign node8464 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node8468 = (inp[7]) ? node8482 : node8469;
													assign node8469 = (inp[0]) ? node8475 : node8470;
														assign node8470 = (inp[12]) ? node8472 : 4'b0001;
															assign node8472 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node8475 = (inp[12]) ? node8479 : node8476;
															assign node8476 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node8479 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node8482 = (inp[13]) ? 4'b0001 : node8483;
														assign node8483 = (inp[12]) ? node8485 : 4'b0101;
															assign node8485 = (inp[14]) ? 4'b1001 : 4'b0101;
											assign node8489 = (inp[13]) ? 4'b0001 : node8490;
												assign node8490 = (inp[0]) ? node8496 : node8491;
													assign node8491 = (inp[7]) ? node8493 : 4'b0001;
														assign node8493 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node8496 = (inp[2]) ? node8500 : node8497;
														assign node8497 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node8500 = (inp[7]) ? 4'b0101 : 4'b1001;
							assign node8504 = (inp[4]) ? node8922 : node8505;
								assign node8505 = (inp[11]) ? node8777 : node8506;
									assign node8506 = (inp[7]) ? node8628 : node8507;
										assign node8507 = (inp[13]) ? node8581 : node8508;
											assign node8508 = (inp[2]) ? node8544 : node8509;
												assign node8509 = (inp[10]) ? node8527 : node8510;
													assign node8510 = (inp[1]) ? node8518 : node8511;
														assign node8511 = (inp[14]) ? node8513 : 4'b1001;
															assign node8513 = (inp[0]) ? node8515 : 4'b1000;
																assign node8515 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8518 = (inp[12]) ? node8522 : node8519;
															assign node8519 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node8522 = (inp[0]) ? node8524 : 4'b1001;
																assign node8524 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8527 = (inp[0]) ? node8535 : node8528;
														assign node8528 = (inp[1]) ? node8532 : node8529;
															assign node8529 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node8532 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8535 = (inp[14]) ? 4'b1001 : node8536;
															assign node8536 = (inp[12]) ? node8540 : node8537;
																assign node8537 = (inp[1]) ? 4'b0001 : 4'b1001;
																assign node8540 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node8544 = (inp[12]) ? node8566 : node8545;
													assign node8545 = (inp[10]) ? node8555 : node8546;
														assign node8546 = (inp[0]) ? node8548 : 4'b1000;
															assign node8548 = (inp[1]) ? node8552 : node8549;
																assign node8549 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node8552 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8555 = (inp[14]) ? node8561 : node8556;
															assign node8556 = (inp[1]) ? node8558 : 4'b0000;
																assign node8558 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node8561 = (inp[0]) ? 4'b0000 : node8562;
																assign node8562 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node8566 = (inp[14]) ? node8578 : node8567;
														assign node8567 = (inp[0]) ? node8573 : node8568;
															assign node8568 = (inp[10]) ? 4'b0000 : node8569;
																assign node8569 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node8573 = (inp[10]) ? 4'b0000 : node8574;
																assign node8574 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node8578 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node8581 = (inp[1]) ? node8607 : node8582;
												assign node8582 = (inp[10]) ? node8596 : node8583;
													assign node8583 = (inp[12]) ? node8593 : node8584;
														assign node8584 = (inp[0]) ? node8590 : node8585;
															assign node8585 = (inp[2]) ? node8587 : 4'b0000;
																assign node8587 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8590 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node8593 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node8596 = (inp[0]) ? node8602 : node8597;
														assign node8597 = (inp[14]) ? node8599 : 4'b1000;
															assign node8599 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8602 = (inp[12]) ? node8604 : 4'b0000;
															assign node8604 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node8607 = (inp[10]) ? node8617 : node8608;
													assign node8608 = (inp[2]) ? node8614 : node8609;
														assign node8609 = (inp[14]) ? 4'b1000 : node8610;
															assign node8610 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node8614 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node8617 = (inp[0]) ? node8623 : node8618;
														assign node8618 = (inp[2]) ? 4'b1000 : node8619;
															assign node8619 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8623 = (inp[2]) ? 4'b0000 : node8624;
															assign node8624 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node8628 = (inp[1]) ? node8708 : node8629;
											assign node8629 = (inp[12]) ? node8673 : node8630;
												assign node8630 = (inp[13]) ? node8654 : node8631;
													assign node8631 = (inp[10]) ? node8643 : node8632;
														assign node8632 = (inp[0]) ? node8640 : node8633;
															assign node8633 = (inp[14]) ? node8637 : node8634;
																assign node8634 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node8637 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node8640 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node8643 = (inp[2]) ? node8649 : node8644;
															assign node8644 = (inp[0]) ? node8646 : 4'b1001;
																assign node8646 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8649 = (inp[0]) ? node8651 : 4'b0000;
																assign node8651 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8654 = (inp[0]) ? node8664 : node8655;
														assign node8655 = (inp[10]) ? node8661 : node8656;
															assign node8656 = (inp[2]) ? node8658 : 4'b0000;
																assign node8658 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8661 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node8664 = (inp[14]) ? node8670 : node8665;
															assign node8665 = (inp[2]) ? 4'b0000 : node8666;
																assign node8666 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node8670 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node8673 = (inp[0]) ? node8693 : node8674;
													assign node8674 = (inp[13]) ? node8686 : node8675;
														assign node8675 = (inp[2]) ? node8681 : node8676;
															assign node8676 = (inp[10]) ? 4'b1001 : node8677;
																assign node8677 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node8681 = (inp[14]) ? node8683 : 4'b1000;
																assign node8683 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8686 = (inp[14]) ? 4'b0000 : node8687;
															assign node8687 = (inp[10]) ? 4'b1001 : node8688;
																assign node8688 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node8693 = (inp[13]) ? node8705 : node8694;
														assign node8694 = (inp[10]) ? node8700 : node8695;
															assign node8695 = (inp[14]) ? 4'b0000 : node8696;
																assign node8696 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node8700 = (inp[14]) ? node8702 : 4'b0001;
																assign node8702 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node8705 = (inp[2]) ? 4'b1001 : 4'b0001;
											assign node8708 = (inp[13]) ? node8744 : node8709;
												assign node8709 = (inp[0]) ? node8723 : node8710;
													assign node8710 = (inp[2]) ? node8718 : node8711;
														assign node8711 = (inp[10]) ? node8715 : node8712;
															assign node8712 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node8715 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node8718 = (inp[14]) ? 4'b0000 : node8719;
															assign node8719 = (inp[10]) ? 4'b1000 : 4'b0001;
													assign node8723 = (inp[12]) ? node8733 : node8724;
														assign node8724 = (inp[2]) ? node8730 : node8725;
															assign node8725 = (inp[14]) ? node8727 : 4'b0000;
																assign node8727 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8730 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8733 = (inp[2]) ? node8739 : node8734;
															assign node8734 = (inp[14]) ? node8736 : 4'b1000;
																assign node8736 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8739 = (inp[10]) ? 4'b1001 : node8740;
																assign node8740 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node8744 = (inp[12]) ? node8758 : node8745;
													assign node8745 = (inp[10]) ? node8755 : node8746;
														assign node8746 = (inp[0]) ? node8752 : node8747;
															assign node8747 = (inp[2]) ? node8749 : 4'b0000;
																assign node8749 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node8752 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8755 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node8758 = (inp[10]) ? node8768 : node8759;
														assign node8759 = (inp[0]) ? node8763 : node8760;
															assign node8760 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node8763 = (inp[14]) ? node8765 : 4'b1001;
																assign node8765 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node8768 = (inp[14]) ? node8772 : node8769;
															assign node8769 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node8772 = (inp[0]) ? 4'b0000 : node8773;
																assign node8773 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node8777 = (inp[1]) ? node8875 : node8778;
										assign node8778 = (inp[2]) ? node8828 : node8779;
											assign node8779 = (inp[0]) ? node8797 : node8780;
												assign node8780 = (inp[10]) ? node8792 : node8781;
													assign node8781 = (inp[14]) ? node8783 : 4'b0000;
														assign node8783 = (inp[7]) ? node8787 : node8784;
															assign node8784 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node8787 = (inp[13]) ? node8789 : 4'b0000;
																assign node8789 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8792 = (inp[7]) ? node8794 : 4'b1000;
														assign node8794 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node8797 = (inp[14]) ? node8809 : node8798;
													assign node8798 = (inp[13]) ? node8804 : node8799;
														assign node8799 = (inp[7]) ? 4'b1000 : node8800;
															assign node8800 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node8804 = (inp[10]) ? node8806 : 4'b1001;
															assign node8806 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node8809 = (inp[12]) ? node8817 : node8810;
														assign node8810 = (inp[7]) ? node8812 : 4'b1000;
															assign node8812 = (inp[13]) ? node8814 : 4'b1000;
																assign node8814 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node8817 = (inp[13]) ? node8821 : node8818;
															assign node8818 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8821 = (inp[7]) ? node8825 : node8822;
																assign node8822 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node8825 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node8828 = (inp[7]) ? node8854 : node8829;
												assign node8829 = (inp[13]) ? node8841 : node8830;
													assign node8830 = (inp[12]) ? node8836 : node8831;
														assign node8831 = (inp[0]) ? 4'b0001 : node8832;
															assign node8832 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8836 = (inp[0]) ? node8838 : 4'b1000;
															assign node8838 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node8841 = (inp[0]) ? node8847 : node8842;
														assign node8842 = (inp[12]) ? node8844 : 4'b0001;
															assign node8844 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node8847 = (inp[10]) ? node8851 : node8848;
															assign node8848 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8851 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node8854 = (inp[10]) ? node8866 : node8855;
													assign node8855 = (inp[12]) ? node8861 : node8856;
														assign node8856 = (inp[13]) ? node8858 : 4'b0000;
															assign node8858 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node8861 = (inp[13]) ? 4'b1000 : node8862;
															assign node8862 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node8866 = (inp[13]) ? node8872 : node8867;
														assign node8867 = (inp[0]) ? 4'b1000 : node8868;
															assign node8868 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8872 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node8875 = (inp[2]) ? node8895 : node8876;
											assign node8876 = (inp[7]) ? node8886 : node8877;
												assign node8877 = (inp[10]) ? 4'b0001 : node8878;
													assign node8878 = (inp[13]) ? node8880 : 4'b0001;
														assign node8880 = (inp[0]) ? node8882 : 4'b0001;
															assign node8882 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node8886 = (inp[0]) ? 4'b0001 : node8887;
													assign node8887 = (inp[10]) ? node8891 : node8888;
														assign node8888 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node8891 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node8895 = (inp[13]) ? node8913 : node8896;
												assign node8896 = (inp[12]) ? node8906 : node8897;
													assign node8897 = (inp[10]) ? node8899 : 4'b1001;
														assign node8899 = (inp[0]) ? node8903 : node8900;
															assign node8900 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node8903 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node8906 = (inp[10]) ? node8908 : 4'b0001;
														assign node8908 = (inp[0]) ? 4'b1001 : node8909;
															assign node8909 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node8913 = (inp[0]) ? node8915 : 4'b0001;
													assign node8915 = (inp[10]) ? 4'b0001 : node8916;
														assign node8916 = (inp[7]) ? node8918 : 4'b1001;
															assign node8918 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node8922 = (inp[13]) ? node9102 : node8923;
									assign node8923 = (inp[1]) ? node9023 : node8924;
										assign node8924 = (inp[0]) ? node8968 : node8925;
											assign node8925 = (inp[2]) ? node8949 : node8926;
												assign node8926 = (inp[12]) ? node8936 : node8927;
													assign node8927 = (inp[10]) ? 4'b0000 : node8928;
														assign node8928 = (inp[14]) ? node8930 : 4'b1000;
															assign node8930 = (inp[7]) ? node8932 : 4'b0001;
																assign node8932 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node8936 = (inp[10]) ? 4'b0001 : node8937;
														assign node8937 = (inp[14]) ? node8943 : node8938;
															assign node8938 = (inp[11]) ? node8940 : 4'b0001;
																assign node8940 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node8943 = (inp[11]) ? node8945 : 4'b0000;
																assign node8945 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node8949 = (inp[12]) ? node8957 : node8950;
													assign node8950 = (inp[10]) ? 4'b0001 : node8951;
														assign node8951 = (inp[7]) ? 4'b1000 : node8952;
															assign node8952 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node8957 = (inp[10]) ? node8961 : node8958;
														assign node8958 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node8961 = (inp[11]) ? node8965 : node8962;
															assign node8962 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node8965 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node8968 = (inp[12]) ? node8998 : node8969;
												assign node8969 = (inp[2]) ? node8981 : node8970;
													assign node8970 = (inp[11]) ? node8978 : node8971;
														assign node8971 = (inp[7]) ? node8973 : 4'b1000;
															assign node8973 = (inp[10]) ? node8975 : 4'b1000;
																assign node8975 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node8978 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node8981 = (inp[10]) ? node8995 : node8982;
														assign node8982 = (inp[14]) ? node8990 : node8983;
															assign node8983 = (inp[11]) ? node8987 : node8984;
																assign node8984 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node8987 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node8990 = (inp[11]) ? node8992 : 4'b1000;
																assign node8992 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node8995 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node8998 = (inp[2]) ? node9010 : node8999;
													assign node8999 = (inp[11]) ? node9005 : node9000;
														assign node9000 = (inp[10]) ? 4'b1001 : node9001;
															assign node9001 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9005 = (inp[10]) ? 4'b1000 : node9006;
															assign node9006 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9010 = (inp[14]) ? node9018 : node9011;
														assign node9011 = (inp[11]) ? node9015 : node9012;
															assign node9012 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node9015 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node9018 = (inp[11]) ? node9020 : 4'b0000;
															assign node9020 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node9023 = (inp[11]) ? node9081 : node9024;
											assign node9024 = (inp[10]) ? node9052 : node9025;
												assign node9025 = (inp[12]) ? node9035 : node9026;
													assign node9026 = (inp[7]) ? node9030 : node9027;
														assign node9027 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node9030 = (inp[2]) ? 4'b0000 : node9031;
															assign node9031 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9035 = (inp[7]) ? node9045 : node9036;
														assign node9036 = (inp[2]) ? node9038 : 4'b1000;
															assign node9038 = (inp[14]) ? node9042 : node9039;
																assign node9039 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node9042 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node9045 = (inp[0]) ? node9049 : node9046;
															assign node9046 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9049 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node9052 = (inp[7]) ? node9068 : node9053;
													assign node9053 = (inp[2]) ? node9061 : node9054;
														assign node9054 = (inp[0]) ? 4'b0001 : node9055;
															assign node9055 = (inp[12]) ? node9057 : 4'b0001;
																assign node9057 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node9061 = (inp[0]) ? node9063 : 4'b0001;
															assign node9063 = (inp[14]) ? 4'b0000 : node9064;
																assign node9064 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node9068 = (inp[0]) ? node9074 : node9069;
														assign node9069 = (inp[14]) ? 4'b0000 : node9070;
															assign node9070 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node9074 = (inp[14]) ? 4'b0001 : node9075;
															assign node9075 = (inp[2]) ? node9077 : 4'b0000;
																assign node9077 = (inp[12]) ? 4'b1000 : 4'b0001;
											assign node9081 = (inp[10]) ? 4'b0001 : node9082;
												assign node9082 = (inp[0]) ? node9094 : node9083;
													assign node9083 = (inp[12]) ? node9089 : node9084;
														assign node9084 = (inp[7]) ? node9086 : 4'b0001;
															assign node9086 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node9089 = (inp[7]) ? node9091 : 4'b1001;
															assign node9091 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node9094 = (inp[12]) ? 4'b0001 : node9095;
														assign node9095 = (inp[7]) ? 4'b0001 : node9096;
															assign node9096 = (inp[14]) ? 4'b0001 : 4'b1001;
									assign node9102 = (inp[10]) ? node9168 : node9103;
										assign node9103 = (inp[1]) ? node9149 : node9104;
											assign node9104 = (inp[0]) ? node9130 : node9105;
												assign node9105 = (inp[7]) ? node9119 : node9106;
													assign node9106 = (inp[14]) ? node9108 : 4'b0000;
														assign node9108 = (inp[11]) ? node9114 : node9109;
															assign node9109 = (inp[12]) ? node9111 : 4'b0000;
																assign node9111 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node9114 = (inp[12]) ? node9116 : 4'b0001;
																assign node9116 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node9119 = (inp[11]) ? node9125 : node9120;
														assign node9120 = (inp[2]) ? 4'b0001 : node9121;
															assign node9121 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node9125 = (inp[2]) ? 4'b0000 : node9126;
															assign node9126 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node9130 = (inp[11]) ? node9136 : node9131;
													assign node9131 = (inp[7]) ? node9133 : 4'b0001;
														assign node9133 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node9136 = (inp[2]) ? node9142 : node9137;
														assign node9137 = (inp[12]) ? node9139 : 4'b0000;
															assign node9139 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node9142 = (inp[12]) ? node9146 : node9143;
															assign node9143 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node9146 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node9149 = (inp[11]) ? 4'b0001 : node9150;
												assign node9150 = (inp[0]) ? node9160 : node9151;
													assign node9151 = (inp[14]) ? node9157 : node9152;
														assign node9152 = (inp[2]) ? node9154 : 4'b0001;
															assign node9154 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node9157 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node9160 = (inp[14]) ? node9162 : 4'b0000;
														assign node9162 = (inp[12]) ? node9164 : 4'b0001;
															assign node9164 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node9168 = (inp[11]) ? 4'b0000 : node9169;
											assign node9169 = (inp[1]) ? 4'b0000 : node9170;
												assign node9170 = (inp[14]) ? node9182 : node9171;
													assign node9171 = (inp[12]) ? node9177 : node9172;
														assign node9172 = (inp[2]) ? 4'b0000 : node9173;
															assign node9173 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node9177 = (inp[0]) ? node9179 : 4'b0001;
															assign node9179 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node9182 = (inp[7]) ? 4'b0000 : node9183;
														assign node9183 = (inp[2]) ? 4'b0001 : 4'b0000;
				assign node9189 = (inp[0]) ? node11163 : node9190;
					assign node9190 = (inp[6]) ? node9692 : node9191;
						assign node9191 = (inp[2]) ? node9595 : node9192;
							assign node9192 = (inp[5]) ? node9282 : node9193;
								assign node9193 = (inp[3]) ? node9195 : 4'b0011;
									assign node9195 = (inp[7]) ? node9257 : node9196;
										assign node9196 = (inp[4]) ? node9222 : node9197;
											assign node9197 = (inp[13]) ? node9199 : 4'b0011;
												assign node9199 = (inp[12]) ? node9211 : node9200;
													assign node9200 = (inp[1]) ? node9206 : node9201;
														assign node9201 = (inp[14]) ? node9203 : 4'b0000;
															assign node9203 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node9206 = (inp[11]) ? 4'b0001 : node9207;
															assign node9207 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9211 = (inp[10]) ? node9213 : 4'b0011;
														assign node9213 = (inp[1]) ? node9217 : node9214;
															assign node9214 = (inp[11]) ? 4'b0000 : 4'b0011;
															assign node9217 = (inp[14]) ? node9219 : 4'b0001;
																assign node9219 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node9222 = (inp[1]) ? node9242 : node9223;
												assign node9223 = (inp[14]) ? node9231 : node9224;
													assign node9224 = (inp[13]) ? node9226 : 4'b1000;
														assign node9226 = (inp[10]) ? 4'b0000 : node9227;
															assign node9227 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node9231 = (inp[11]) ? node9237 : node9232;
														assign node9232 = (inp[13]) ? node9234 : 4'b0001;
															assign node9234 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node9237 = (inp[10]) ? node9239 : 4'b0000;
															assign node9239 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node9242 = (inp[14]) ? node9254 : node9243;
													assign node9243 = (inp[13]) ? node9249 : node9244;
														assign node9244 = (inp[10]) ? 4'b1001 : node9245;
															assign node9245 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9249 = (inp[10]) ? 4'b0001 : node9250;
															assign node9250 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node9254 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node9257 = (inp[4]) ? node9259 : 4'b0011;
											assign node9259 = (inp[13]) ? node9261 : 4'b0011;
												assign node9261 = (inp[12]) ? node9275 : node9262;
													assign node9262 = (inp[1]) ? node9270 : node9263;
														assign node9263 = (inp[14]) ? node9265 : 4'b0000;
															assign node9265 = (inp[11]) ? 4'b0000 : node9266;
																assign node9266 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node9270 = (inp[14]) ? node9272 : 4'b0001;
															assign node9272 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node9275 = (inp[10]) ? node9277 : 4'b0011;
														assign node9277 = (inp[1]) ? 4'b0001 : node9278;
															assign node9278 = (inp[14]) ? 4'b0011 : 4'b0000;
								assign node9282 = (inp[1]) ? node9446 : node9283;
									assign node9283 = (inp[14]) ? node9349 : node9284;
										assign node9284 = (inp[13]) ? node9320 : node9285;
											assign node9285 = (inp[10]) ? node9309 : node9286;
												assign node9286 = (inp[12]) ? node9298 : node9287;
													assign node9287 = (inp[3]) ? node9293 : node9288;
														assign node9288 = (inp[7]) ? 4'b1000 : node9289;
															assign node9289 = (inp[11]) ? 4'b1000 : 4'b1100;
														assign node9293 = (inp[4]) ? node9295 : 4'b1100;
															assign node9295 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node9298 = (inp[3]) ? node9304 : node9299;
														assign node9299 = (inp[7]) ? 4'b0000 : node9300;
															assign node9300 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9304 = (inp[11]) ? node9306 : 4'b0100;
															assign node9306 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node9309 = (inp[3]) ? node9315 : node9310;
													assign node9310 = (inp[4]) ? node9312 : 4'b1000;
														assign node9312 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node9315 = (inp[7]) ? 4'b1100 : node9316;
														assign node9316 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node9320 = (inp[12]) ? node9332 : node9321;
												assign node9321 = (inp[3]) ? node9327 : node9322;
													assign node9322 = (inp[7]) ? node9324 : 4'b0100;
														assign node9324 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node9327 = (inp[4]) ? 4'b0000 : node9328;
														assign node9328 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node9332 = (inp[10]) ? node9342 : node9333;
													assign node9333 = (inp[3]) ? node9339 : node9334;
														assign node9334 = (inp[7]) ? 4'b1000 : node9335;
															assign node9335 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9339 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node9342 = (inp[3]) ? 4'b0000 : node9343;
														assign node9343 = (inp[7]) ? node9345 : 4'b0100;
															assign node9345 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node9349 = (inp[11]) ? node9401 : node9350;
											assign node9350 = (inp[13]) ? node9378 : node9351;
												assign node9351 = (inp[10]) ? node9363 : node9352;
													assign node9352 = (inp[3]) ? node9358 : node9353;
														assign node9353 = (inp[7]) ? 4'b0001 : node9354;
															assign node9354 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node9358 = (inp[7]) ? 4'b0101 : node9359;
															assign node9359 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9363 = (inp[12]) ? node9371 : node9364;
														assign node9364 = (inp[7]) ? 4'b1101 : node9365;
															assign node9365 = (inp[3]) ? node9367 : 4'b1001;
																assign node9367 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node9371 = (inp[7]) ? 4'b0101 : node9372;
															assign node9372 = (inp[4]) ? node9374 : 4'b0001;
																assign node9374 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node9378 = (inp[12]) ? node9392 : node9379;
													assign node9379 = (inp[10]) ? node9383 : node9380;
														assign node9380 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node9383 = (inp[3]) ? node9387 : node9384;
															assign node9384 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node9387 = (inp[7]) ? node9389 : 4'b0001;
																assign node9389 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9392 = (inp[7]) ? 4'b1101 : node9393;
														assign node9393 = (inp[4]) ? node9397 : node9394;
															assign node9394 = (inp[3]) ? 4'b1101 : 4'b1001;
															assign node9397 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node9401 = (inp[13]) ? node9423 : node9402;
												assign node9402 = (inp[10]) ? node9414 : node9403;
													assign node9403 = (inp[12]) ? node9409 : node9404;
														assign node9404 = (inp[3]) ? 4'b1100 : node9405;
															assign node9405 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node9409 = (inp[3]) ? 4'b0100 : node9410;
															assign node9410 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node9414 = (inp[3]) ? node9420 : node9415;
														assign node9415 = (inp[4]) ? node9417 : 4'b1000;
															assign node9417 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node9420 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node9423 = (inp[10]) ? node9435 : node9424;
													assign node9424 = (inp[12]) ? node9432 : node9425;
														assign node9425 = (inp[7]) ? node9427 : 4'b0000;
															assign node9427 = (inp[4]) ? 4'b0100 : node9428;
																assign node9428 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node9432 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node9435 = (inp[3]) ? node9441 : node9436;
														assign node9436 = (inp[12]) ? 4'b0100 : node9437;
															assign node9437 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9441 = (inp[4]) ? 4'b0000 : node9442;
															assign node9442 = (inp[7]) ? 4'b0100 : 4'b0000;
									assign node9446 = (inp[14]) ? node9504 : node9447;
										assign node9447 = (inp[13]) ? node9473 : node9448;
											assign node9448 = (inp[3]) ? node9460 : node9449;
												assign node9449 = (inp[10]) ? 4'b1001 : node9450;
													assign node9450 = (inp[12]) ? node9456 : node9451;
														assign node9451 = (inp[7]) ? 4'b1001 : node9452;
															assign node9452 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9456 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node9460 = (inp[4]) ? node9466 : node9461;
													assign node9461 = (inp[10]) ? 4'b1101 : node9462;
														assign node9462 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node9466 = (inp[7]) ? node9470 : node9467;
														assign node9467 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9470 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node9473 = (inp[10]) ? node9493 : node9474;
												assign node9474 = (inp[12]) ? node9482 : node9475;
													assign node9475 = (inp[3]) ? 4'b0001 : node9476;
														assign node9476 = (inp[11]) ? 4'b0101 : node9477;
															assign node9477 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node9482 = (inp[3]) ? node9488 : node9483;
														assign node9483 = (inp[4]) ? node9485 : 4'b1001;
															assign node9485 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node9488 = (inp[4]) ? node9490 : 4'b1101;
															assign node9490 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node9493 = (inp[3]) ? node9499 : node9494;
													assign node9494 = (inp[4]) ? 4'b0101 : node9495;
														assign node9495 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9499 = (inp[4]) ? 4'b0001 : node9500;
														assign node9500 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node9504 = (inp[11]) ? node9552 : node9505;
											assign node9505 = (inp[13]) ? node9527 : node9506;
												assign node9506 = (inp[3]) ? node9518 : node9507;
													assign node9507 = (inp[10]) ? node9513 : node9508;
														assign node9508 = (inp[12]) ? node9510 : 4'b1000;
															assign node9510 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9513 = (inp[7]) ? 4'b1000 : node9514;
															assign node9514 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9518 = (inp[10]) ? node9522 : node9519;
														assign node9519 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node9522 = (inp[7]) ? 4'b1100 : node9523;
															assign node9523 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node9527 = (inp[12]) ? node9535 : node9528;
													assign node9528 = (inp[3]) ? node9530 : 4'b0100;
														assign node9530 = (inp[7]) ? node9532 : 4'b0000;
															assign node9532 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node9535 = (inp[10]) ? node9545 : node9536;
														assign node9536 = (inp[3]) ? node9540 : node9537;
															assign node9537 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node9540 = (inp[4]) ? node9542 : 4'b1100;
																assign node9542 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node9545 = (inp[4]) ? 4'b0000 : node9546;
															assign node9546 = (inp[3]) ? 4'b0100 : node9547;
																assign node9547 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node9552 = (inp[13]) ? node9572 : node9553;
												assign node9553 = (inp[3]) ? node9563 : node9554;
													assign node9554 = (inp[10]) ? node9558 : node9555;
														assign node9555 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9558 = (inp[4]) ? node9560 : 4'b1001;
															assign node9560 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node9563 = (inp[7]) ? node9567 : node9564;
														assign node9564 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node9567 = (inp[10]) ? 4'b1101 : node9568;
															assign node9568 = (inp[4]) ? 4'b1101 : 4'b0101;
												assign node9572 = (inp[12]) ? node9584 : node9573;
													assign node9573 = (inp[3]) ? node9579 : node9574;
														assign node9574 = (inp[4]) ? 4'b0101 : node9575;
															assign node9575 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node9579 = (inp[7]) ? node9581 : 4'b0001;
															assign node9581 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node9584 = (inp[10]) ? node9588 : node9585;
														assign node9585 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node9588 = (inp[3]) ? 4'b0001 : node9589;
															assign node9589 = (inp[4]) ? 4'b0101 : node9590;
																assign node9590 = (inp[7]) ? 4'b0001 : 4'b0101;
							assign node9595 = (inp[5]) ? node9597 : 4'b0011;
								assign node9597 = (inp[3]) ? node9599 : 4'b0011;
									assign node9599 = (inp[4]) ? node9621 : node9600;
										assign node9600 = (inp[7]) ? 4'b0011 : node9601;
											assign node9601 = (inp[13]) ? node9603 : 4'b0011;
												assign node9603 = (inp[10]) ? node9609 : node9604;
													assign node9604 = (inp[12]) ? 4'b0011 : node9605;
														assign node9605 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9609 = (inp[1]) ? node9617 : node9610;
														assign node9610 = (inp[14]) ? node9612 : 4'b0000;
															assign node9612 = (inp[11]) ? 4'b0000 : node9613;
																assign node9613 = (inp[12]) ? 4'b0011 : 4'b0001;
														assign node9617 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node9621 = (inp[7]) ? node9671 : node9622;
											assign node9622 = (inp[1]) ? node9652 : node9623;
												assign node9623 = (inp[14]) ? node9635 : node9624;
													assign node9624 = (inp[11]) ? 4'b1000 : node9625;
														assign node9625 = (inp[10]) ? node9631 : node9626;
															assign node9626 = (inp[13]) ? node9628 : 4'b0000;
																assign node9628 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node9631 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node9635 = (inp[11]) ? node9643 : node9636;
														assign node9636 = (inp[13]) ? 4'b1001 : node9637;
															assign node9637 = (inp[12]) ? 4'b0001 : node9638;
																assign node9638 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9643 = (inp[10]) ? 4'b0000 : node9644;
															assign node9644 = (inp[13]) ? node9648 : node9645;
																assign node9645 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node9648 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node9652 = (inp[13]) ? node9658 : node9653;
													assign node9653 = (inp[11]) ? 4'b1001 : node9654;
														assign node9654 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node9658 = (inp[12]) ? node9664 : node9659;
														assign node9659 = (inp[14]) ? node9661 : 4'b0001;
															assign node9661 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node9664 = (inp[10]) ? 4'b0001 : node9665;
															assign node9665 = (inp[11]) ? 4'b1001 : node9666;
																assign node9666 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node9671 = (inp[13]) ? node9673 : 4'b0011;
												assign node9673 = (inp[12]) ? node9683 : node9674;
													assign node9674 = (inp[1]) ? node9680 : node9675;
														assign node9675 = (inp[11]) ? 4'b0000 : node9676;
															assign node9676 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node9680 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node9683 = (inp[10]) ? node9685 : 4'b0011;
														assign node9685 = (inp[1]) ? node9687 : 4'b0000;
															assign node9687 = (inp[11]) ? 4'b0001 : node9688;
																assign node9688 = (inp[14]) ? 4'b0000 : 4'b0001;
						assign node9692 = (inp[1]) ? node10488 : node9693;
							assign node9693 = (inp[5]) ? node10097 : node9694;
								assign node9694 = (inp[14]) ? node9878 : node9695;
									assign node9695 = (inp[13]) ? node9773 : node9696;
										assign node9696 = (inp[3]) ? node9718 : node9697;
											assign node9697 = (inp[10]) ? node9709 : node9698;
												assign node9698 = (inp[12]) ? node9704 : node9699;
													assign node9699 = (inp[7]) ? 4'b1000 : node9700;
														assign node9700 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node9704 = (inp[4]) ? node9706 : 4'b0000;
														assign node9706 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9709 = (inp[7]) ? 4'b1000 : node9710;
													assign node9710 = (inp[4]) ? node9712 : 4'b1000;
														assign node9712 = (inp[12]) ? 4'b1100 : node9713;
															assign node9713 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node9718 = (inp[11]) ? node9746 : node9719;
												assign node9719 = (inp[4]) ? node9729 : node9720;
													assign node9720 = (inp[2]) ? 4'b1100 : node9721;
														assign node9721 = (inp[12]) ? 4'b1000 : node9722;
															assign node9722 = (inp[10]) ? node9724 : 4'b1000;
																assign node9724 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node9729 = (inp[7]) ? node9739 : node9730;
														assign node9730 = (inp[2]) ? 4'b0000 : node9731;
															assign node9731 = (inp[12]) ? node9735 : node9732;
																assign node9732 = (inp[10]) ? 4'b0000 : 4'b1100;
																assign node9735 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node9739 = (inp[10]) ? node9741 : 4'b0100;
															assign node9741 = (inp[2]) ? 4'b1100 : node9742;
																assign node9742 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node9746 = (inp[2]) ? node9760 : node9747;
													assign node9747 = (inp[4]) ? node9755 : node9748;
														assign node9748 = (inp[10]) ? node9752 : node9749;
															assign node9749 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node9752 = (inp[7]) ? 4'b1001 : 4'b0101;
														assign node9755 = (inp[10]) ? node9757 : 4'b1101;
															assign node9757 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node9760 = (inp[7]) ? node9768 : node9761;
														assign node9761 = (inp[4]) ? node9763 : 4'b1100;
															assign node9763 = (inp[10]) ? 4'b0001 : node9764;
																assign node9764 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9768 = (inp[12]) ? node9770 : 4'b1100;
															assign node9770 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node9773 = (inp[12]) ? node9821 : node9774;
											assign node9774 = (inp[2]) ? node9802 : node9775;
												assign node9775 = (inp[10]) ? node9789 : node9776;
													assign node9776 = (inp[3]) ? node9782 : node9777;
														assign node9777 = (inp[7]) ? node9779 : 4'b1001;
															assign node9779 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9782 = (inp[4]) ? 4'b0001 : node9783;
															assign node9783 = (inp[7]) ? node9785 : 4'b1100;
																assign node9785 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9789 = (inp[4]) ? node9797 : node9790;
														assign node9790 = (inp[3]) ? node9794 : node9791;
															assign node9791 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node9794 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node9797 = (inp[3]) ? 4'b0000 : node9798;
															assign node9798 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node9802 = (inp[3]) ? node9808 : node9803;
													assign node9803 = (inp[4]) ? 4'b0100 : node9804;
														assign node9804 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node9808 = (inp[7]) ? node9818 : node9809;
														assign node9809 = (inp[4]) ? node9811 : 4'b0000;
															assign node9811 = (inp[11]) ? node9815 : node9812;
																assign node9812 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node9815 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node9818 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node9821 = (inp[10]) ? node9845 : node9822;
												assign node9822 = (inp[2]) ? node9838 : node9823;
													assign node9823 = (inp[11]) ? node9831 : node9824;
														assign node9824 = (inp[3]) ? 4'b0000 : node9825;
															assign node9825 = (inp[4]) ? node9827 : 4'b1000;
																assign node9827 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node9831 = (inp[4]) ? node9833 : 4'b0101;
															assign node9833 = (inp[7]) ? 4'b0101 : node9834;
																assign node9834 = (inp[3]) ? 4'b0000 : 4'b0001;
													assign node9838 = (inp[3]) ? 4'b1100 : node9839;
														assign node9839 = (inp[4]) ? node9841 : 4'b1000;
															assign node9841 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node9845 = (inp[2]) ? node9863 : node9846;
													assign node9846 = (inp[3]) ? node9856 : node9847;
														assign node9847 = (inp[7]) ? node9853 : node9848;
															assign node9848 = (inp[4]) ? node9850 : 4'b0100;
																assign node9850 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node9853 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9856 = (inp[4]) ? node9860 : node9857;
															assign node9857 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node9860 = (inp[11]) ? 4'b1000 : 4'b1100;
													assign node9863 = (inp[3]) ? node9869 : node9864;
														assign node9864 = (inp[7]) ? node9866 : 4'b0100;
															assign node9866 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node9869 = (inp[4]) ? node9873 : node9870;
															assign node9870 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node9873 = (inp[7]) ? 4'b0000 : node9874;
																assign node9874 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node9878 = (inp[11]) ? node9982 : node9879;
										assign node9879 = (inp[3]) ? node9921 : node9880;
											assign node9880 = (inp[7]) ? node9906 : node9881;
												assign node9881 = (inp[4]) ? node9891 : node9882;
													assign node9882 = (inp[13]) ? node9888 : node9883;
														assign node9883 = (inp[2]) ? node9885 : 4'b0001;
															assign node9885 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9888 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node9891 = (inp[2]) ? node9899 : node9892;
														assign node9892 = (inp[13]) ? 4'b0000 : node9893;
															assign node9893 = (inp[12]) ? 4'b0101 : node9894;
																assign node9894 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node9899 = (inp[10]) ? node9901 : 4'b0101;
															assign node9901 = (inp[13]) ? node9903 : 4'b1101;
																assign node9903 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node9906 = (inp[13]) ? node9912 : node9907;
													assign node9907 = (inp[10]) ? node9909 : 4'b0001;
														assign node9909 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node9912 = (inp[12]) ? 4'b1001 : node9913;
														assign node9913 = (inp[10]) ? node9915 : 4'b1001;
															assign node9915 = (inp[2]) ? node9917 : 4'b0000;
																assign node9917 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node9921 = (inp[2]) ? node9961 : node9922;
												assign node9922 = (inp[4]) ? node9942 : node9923;
													assign node9923 = (inp[13]) ? node9929 : node9924;
														assign node9924 = (inp[10]) ? 4'b1000 : node9925;
															assign node9925 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9929 = (inp[7]) ? node9937 : node9930;
															assign node9930 = (inp[10]) ? node9934 : node9931;
																assign node9931 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node9934 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node9937 = (inp[12]) ? 4'b1000 : node9938;
																assign node9938 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node9942 = (inp[7]) ? node9952 : node9943;
														assign node9943 = (inp[13]) ? node9949 : node9944;
															assign node9944 = (inp[10]) ? 4'b0000 : node9945;
																assign node9945 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node9949 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node9952 = (inp[12]) ? node9958 : node9953;
															assign node9953 = (inp[10]) ? node9955 : 4'b1100;
																assign node9955 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node9958 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node9961 = (inp[13]) ? node9969 : node9962;
													assign node9962 = (inp[4]) ? node9964 : 4'b0101;
														assign node9964 = (inp[7]) ? node9966 : 4'b0001;
															assign node9966 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node9969 = (inp[4]) ? node9975 : node9970;
														assign node9970 = (inp[10]) ? node9972 : 4'b1101;
															assign node9972 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node9975 = (inp[7]) ? node9979 : node9976;
															assign node9976 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node9979 = (inp[12]) ? 4'b1101 : 4'b0000;
										assign node9982 = (inp[3]) ? node10028 : node9983;
											assign node9983 = (inp[13]) ? node10007 : node9984;
												assign node9984 = (inp[7]) ? node10002 : node9985;
													assign node9985 = (inp[4]) ? node9991 : node9986;
														assign node9986 = (inp[10]) ? 4'b1000 : node9987;
															assign node9987 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9991 = (inp[2]) ? node9997 : node9992;
															assign node9992 = (inp[10]) ? 4'b0001 : node9993;
																assign node9993 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node9997 = (inp[10]) ? 4'b1100 : node9998;
																assign node9998 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node10002 = (inp[10]) ? 4'b1000 : node10003;
														assign node10003 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10007 = (inp[10]) ? node10019 : node10008;
													assign node10008 = (inp[12]) ? node10014 : node10009;
														assign node10009 = (inp[7]) ? node10011 : 4'b0100;
															assign node10011 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10014 = (inp[4]) ? node10016 : 4'b1000;
															assign node10016 = (inp[2]) ? 4'b1100 : 4'b0001;
													assign node10019 = (inp[2]) ? 4'b0100 : node10020;
														assign node10020 = (inp[7]) ? node10024 : node10021;
															assign node10021 = (inp[4]) ? 4'b0001 : 4'b0100;
															assign node10024 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node10028 = (inp[2]) ? node10064 : node10029;
												assign node10029 = (inp[4]) ? node10053 : node10030;
													assign node10030 = (inp[7]) ? node10044 : node10031;
														assign node10031 = (inp[13]) ? node10037 : node10032;
															assign node10032 = (inp[12]) ? node10034 : 4'b0101;
																assign node10034 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node10037 = (inp[12]) ? node10041 : node10038;
																assign node10038 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node10041 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node10044 = (inp[12]) ? node10050 : node10045;
															assign node10045 = (inp[10]) ? node10047 : 4'b1001;
																assign node10047 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node10050 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node10053 = (inp[13]) ? node10059 : node10054;
														assign node10054 = (inp[12]) ? 4'b0101 : node10055;
															assign node10055 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node10059 = (inp[7]) ? node10061 : 4'b0000;
															assign node10061 = (inp[12]) ? 4'b1101 : 4'b0000;
												assign node10064 = (inp[4]) ? node10076 : node10065;
													assign node10065 = (inp[7]) ? node10067 : 4'b1100;
														assign node10067 = (inp[12]) ? node10069 : 4'b0100;
															assign node10069 = (inp[13]) ? node10073 : node10070;
																assign node10070 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node10073 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node10076 = (inp[13]) ? node10084 : node10077;
														assign node10077 = (inp[7]) ? 4'b1100 : node10078;
															assign node10078 = (inp[12]) ? node10080 : 4'b1000;
																assign node10080 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10084 = (inp[7]) ? node10090 : node10085;
															assign node10085 = (inp[12]) ? node10087 : 4'b1001;
																assign node10087 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node10090 = (inp[10]) ? node10094 : node10091;
																assign node10091 = (inp[12]) ? 4'b1100 : 4'b0000;
																assign node10094 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node10097 = (inp[3]) ? node10313 : node10098;
									assign node10098 = (inp[4]) ? node10216 : node10099;
										assign node10099 = (inp[13]) ? node10163 : node10100;
											assign node10100 = (inp[10]) ? node10132 : node10101;
												assign node10101 = (inp[12]) ? node10123 : node10102;
													assign node10102 = (inp[14]) ? node10118 : node10103;
														assign node10103 = (inp[7]) ? node10111 : node10104;
															assign node10104 = (inp[2]) ? node10108 : node10105;
																assign node10105 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node10108 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10111 = (inp[11]) ? node10115 : node10112;
																assign node10112 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node10115 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node10118 = (inp[11]) ? node10120 : 4'b1000;
															assign node10120 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node10123 = (inp[11]) ? node10129 : node10124;
														assign node10124 = (inp[2]) ? 4'b0000 : node10125;
															assign node10125 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10129 = (inp[2]) ? 4'b0001 : 4'b1000;
												assign node10132 = (inp[7]) ? node10148 : node10133;
													assign node10133 = (inp[2]) ? node10141 : node10134;
														assign node10134 = (inp[14]) ? 4'b0100 : node10135;
															assign node10135 = (inp[11]) ? node10137 : 4'b0101;
																assign node10137 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10141 = (inp[12]) ? node10145 : node10142;
															assign node10142 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node10145 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node10148 = (inp[14]) ? node10156 : node10149;
														assign node10149 = (inp[11]) ? node10153 : node10150;
															assign node10150 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node10153 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10156 = (inp[11]) ? node10158 : 4'b1000;
															assign node10158 = (inp[2]) ? node10160 : 4'b1000;
																assign node10160 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node10163 = (inp[10]) ? node10195 : node10164;
												assign node10164 = (inp[7]) ? node10178 : node10165;
													assign node10165 = (inp[11]) ? node10175 : node10166;
														assign node10166 = (inp[2]) ? node10172 : node10167;
															assign node10167 = (inp[14]) ? node10169 : 4'b1101;
																assign node10169 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node10172 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node10175 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node10178 = (inp[2]) ? node10188 : node10179;
														assign node10179 = (inp[11]) ? 4'b0100 : node10180;
															assign node10180 = (inp[12]) ? node10184 : node10181;
																assign node10181 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node10184 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10188 = (inp[12]) ? node10192 : node10189;
															assign node10189 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10192 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node10195 = (inp[12]) ? node10205 : node10196;
													assign node10196 = (inp[2]) ? node10200 : node10197;
														assign node10197 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node10200 = (inp[11]) ? node10202 : 4'b0100;
															assign node10202 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node10205 = (inp[7]) ? node10211 : node10206;
														assign node10206 = (inp[2]) ? node10208 : 4'b0001;
															assign node10208 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node10211 = (inp[2]) ? node10213 : 4'b1100;
															assign node10213 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node10216 = (inp[13]) ? node10254 : node10217;
											assign node10217 = (inp[2]) ? node10233 : node10218;
												assign node10218 = (inp[10]) ? node10224 : node10219;
													assign node10219 = (inp[11]) ? 4'b1001 : node10220;
														assign node10220 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10224 = (inp[7]) ? 4'b1001 : node10225;
														assign node10225 = (inp[11]) ? 4'b0000 : node10226;
															assign node10226 = (inp[12]) ? 4'b0101 : node10227;
																assign node10227 = (inp[14]) ? 4'b1101 : 4'b0000;
												assign node10233 = (inp[10]) ? node10247 : node10234;
													assign node10234 = (inp[7]) ? node10244 : node10235;
														assign node10235 = (inp[12]) ? node10241 : node10236;
															assign node10236 = (inp[14]) ? 4'b1000 : node10237;
																assign node10237 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node10241 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10244 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node10247 = (inp[14]) ? 4'b0000 : node10248;
														assign node10248 = (inp[11]) ? node10250 : 4'b0001;
															assign node10250 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node10254 = (inp[10]) ? node10284 : node10255;
												assign node10255 = (inp[11]) ? node10275 : node10256;
													assign node10256 = (inp[12]) ? node10268 : node10257;
														assign node10257 = (inp[7]) ? node10261 : node10258;
															assign node10258 = (inp[14]) ? 4'b0100 : 4'b0000;
															assign node10261 = (inp[14]) ? node10265 : node10262;
																assign node10262 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node10265 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node10268 = (inp[2]) ? node10272 : node10269;
															assign node10269 = (inp[14]) ? 4'b0101 : 4'b0000;
															assign node10272 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node10275 = (inp[7]) ? node10279 : node10276;
														assign node10276 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node10279 = (inp[2]) ? 4'b0000 : node10280;
															assign node10280 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10284 = (inp[7]) ? node10296 : node10285;
													assign node10285 = (inp[11]) ? node10291 : node10286;
														assign node10286 = (inp[2]) ? node10288 : 4'b0000;
															assign node10288 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10291 = (inp[12]) ? node10293 : 4'b1001;
															assign node10293 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node10296 = (inp[11]) ? node10308 : node10297;
														assign node10297 = (inp[12]) ? node10303 : node10298;
															assign node10298 = (inp[14]) ? 4'b1000 : node10299;
																assign node10299 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node10303 = (inp[2]) ? 4'b1001 : node10304;
																assign node10304 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node10308 = (inp[2]) ? node10310 : 4'b1000;
															assign node10310 = (inp[12]) ? 4'b1000 : 4'b0100;
									assign node10313 = (inp[4]) ? node10395 : node10314;
										assign node10314 = (inp[10]) ? node10350 : node10315;
											assign node10315 = (inp[13]) ? node10329 : node10316;
												assign node10316 = (inp[12]) ? node10324 : node10317;
													assign node10317 = (inp[11]) ? node10321 : node10318;
														assign node10318 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node10321 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node10324 = (inp[11]) ? 4'b1001 : node10325;
														assign node10325 = (inp[2]) ? 4'b0001 : 4'b1000;
												assign node10329 = (inp[11]) ? node10339 : node10330;
													assign node10330 = (inp[2]) ? node10336 : node10331;
														assign node10331 = (inp[7]) ? 4'b1001 : node10332;
															assign node10332 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node10336 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node10339 = (inp[2]) ? node10343 : node10340;
														assign node10340 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node10343 = (inp[7]) ? node10347 : node10344;
															assign node10344 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node10347 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node10350 = (inp[7]) ? node10376 : node10351;
												assign node10351 = (inp[11]) ? node10369 : node10352;
													assign node10352 = (inp[2]) ? node10360 : node10353;
														assign node10353 = (inp[14]) ? 4'b0000 : node10354;
															assign node10354 = (inp[13]) ? 4'b0001 : node10355;
																assign node10355 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10360 = (inp[14]) ? 4'b1001 : node10361;
															assign node10361 = (inp[12]) ? node10365 : node10362;
																assign node10362 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node10365 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node10369 = (inp[13]) ? node10373 : node10370;
														assign node10370 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node10373 = (inp[2]) ? 4'b0001 : 4'b1000;
												assign node10376 = (inp[2]) ? node10386 : node10377;
													assign node10377 = (inp[11]) ? node10381 : node10378;
														assign node10378 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10381 = (inp[12]) ? node10383 : 4'b0000;
															assign node10383 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node10386 = (inp[11]) ? 4'b0000 : node10387;
														assign node10387 = (inp[13]) ? node10391 : node10388;
															assign node10388 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10391 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node10395 = (inp[13]) ? node10455 : node10396;
											assign node10396 = (inp[2]) ? node10420 : node10397;
												assign node10397 = (inp[7]) ? node10405 : node10398;
													assign node10398 = (inp[10]) ? node10400 : 4'b0000;
														assign node10400 = (inp[14]) ? 4'b0000 : node10401;
															assign node10401 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node10405 = (inp[14]) ? node10413 : node10406;
														assign node10406 = (inp[11]) ? 4'b1000 : node10407;
															assign node10407 = (inp[10]) ? node10409 : 4'b0000;
																assign node10409 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node10413 = (inp[12]) ? node10415 : 4'b0001;
															assign node10415 = (inp[11]) ? node10417 : 4'b1001;
																assign node10417 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node10420 = (inp[10]) ? node10438 : node10421;
													assign node10421 = (inp[7]) ? node10429 : node10422;
														assign node10422 = (inp[11]) ? node10426 : node10423;
															assign node10423 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node10426 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10429 = (inp[11]) ? node10435 : node10430;
															assign node10430 = (inp[14]) ? 4'b1001 : node10431;
																assign node10431 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node10435 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10438 = (inp[11]) ? node10450 : node10439;
														assign node10439 = (inp[14]) ? node10445 : node10440;
															assign node10440 = (inp[7]) ? node10442 : 4'b1000;
																assign node10442 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node10445 = (inp[7]) ? node10447 : 4'b0001;
																assign node10447 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node10450 = (inp[7]) ? 4'b0000 : node10451;
															assign node10451 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node10455 = (inp[10]) ? node10469 : node10456;
												assign node10456 = (inp[7]) ? node10462 : node10457;
													assign node10457 = (inp[2]) ? node10459 : 4'b0000;
														assign node10459 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node10462 = (inp[2]) ? node10466 : node10463;
														assign node10463 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node10466 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node10469 = (inp[11]) ? 4'b0000 : node10470;
													assign node10470 = (inp[7]) ? node10478 : node10471;
														assign node10471 = (inp[14]) ? 4'b0000 : node10472;
															assign node10472 = (inp[12]) ? 4'b0000 : node10473;
																assign node10473 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node10478 = (inp[12]) ? node10480 : 4'b0000;
															assign node10480 = (inp[2]) ? node10484 : node10481;
																assign node10481 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node10484 = (inp[14]) ? 4'b0000 : 4'b0001;
							assign node10488 = (inp[11]) ? node10890 : node10489;
								assign node10489 = (inp[5]) ? node10675 : node10490;
									assign node10490 = (inp[14]) ? node10574 : node10491;
										assign node10491 = (inp[3]) ? node10527 : node10492;
											assign node10492 = (inp[13]) ? node10510 : node10493;
												assign node10493 = (inp[12]) ? node10499 : node10494;
													assign node10494 = (inp[4]) ? node10496 : 4'b1001;
														assign node10496 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node10499 = (inp[10]) ? node10505 : node10500;
														assign node10500 = (inp[7]) ? 4'b0001 : node10501;
															assign node10501 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node10505 = (inp[4]) ? node10507 : 4'b1001;
															assign node10507 = (inp[7]) ? 4'b1001 : 4'b0000;
												assign node10510 = (inp[2]) ? node10520 : node10511;
													assign node10511 = (inp[10]) ? node10515 : node10512;
														assign node10512 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node10515 = (inp[4]) ? 4'b0000 : node10516;
															assign node10516 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node10520 = (inp[4]) ? 4'b0101 : node10521;
														assign node10521 = (inp[12]) ? 4'b1001 : node10522;
															assign node10522 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node10527 = (inp[10]) ? node10555 : node10528;
												assign node10528 = (inp[2]) ? node10538 : node10529;
													assign node10529 = (inp[4]) ? node10531 : 4'b1000;
														assign node10531 = (inp[7]) ? 4'b1100 : node10532;
															assign node10532 = (inp[13]) ? node10534 : 4'b1100;
																assign node10534 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10538 = (inp[4]) ? node10544 : node10539;
														assign node10539 = (inp[13]) ? node10541 : 4'b1101;
															assign node10541 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node10544 = (inp[7]) ? node10548 : node10545;
															assign node10545 = (inp[13]) ? 4'b1000 : 4'b0001;
															assign node10548 = (inp[12]) ? node10552 : node10549;
																assign node10549 = (inp[13]) ? 4'b0001 : 4'b1101;
																assign node10552 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node10555 = (inp[4]) ? node10567 : node10556;
													assign node10556 = (inp[2]) ? node10562 : node10557;
														assign node10557 = (inp[7]) ? node10559 : 4'b0100;
															assign node10559 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node10562 = (inp[13]) ? node10564 : 4'b1101;
															assign node10564 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node10567 = (inp[13]) ? 4'b0000 : node10568;
														assign node10568 = (inp[7]) ? node10570 : 4'b0000;
															assign node10570 = (inp[2]) ? 4'b1101 : 4'b0100;
										assign node10574 = (inp[13]) ? node10622 : node10575;
											assign node10575 = (inp[3]) ? node10597 : node10576;
												assign node10576 = (inp[4]) ? node10582 : node10577;
													assign node10577 = (inp[10]) ? 4'b1000 : node10578;
														assign node10578 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10582 = (inp[7]) ? node10592 : node10583;
														assign node10583 = (inp[12]) ? node10585 : 4'b1100;
															assign node10585 = (inp[2]) ? node10589 : node10586;
																assign node10586 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node10589 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node10592 = (inp[12]) ? node10594 : 4'b1000;
															assign node10594 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node10597 = (inp[2]) ? node10609 : node10598;
													assign node10598 = (inp[10]) ? node10602 : node10599;
														assign node10599 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node10602 = (inp[7]) ? node10606 : node10603;
															assign node10603 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node10606 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node10609 = (inp[10]) ? node10617 : node10610;
														assign node10610 = (inp[12]) ? node10612 : 4'b1100;
															assign node10612 = (inp[4]) ? node10614 : 4'b0100;
																assign node10614 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node10617 = (inp[4]) ? node10619 : 4'b1100;
															assign node10619 = (inp[7]) ? 4'b1100 : 4'b0000;
											assign node10622 = (inp[10]) ? node10648 : node10623;
												assign node10623 = (inp[12]) ? node10635 : node10624;
													assign node10624 = (inp[4]) ? node10626 : 4'b0000;
														assign node10626 = (inp[7]) ? node10632 : node10627;
															assign node10627 = (inp[2]) ? 4'b0100 : node10628;
																assign node10628 = (inp[3]) ? 4'b0001 : 4'b1000;
															assign node10632 = (inp[3]) ? 4'b1100 : 4'b0100;
													assign node10635 = (inp[2]) ? node10641 : node10636;
														assign node10636 = (inp[4]) ? node10638 : 4'b1000;
															assign node10638 = (inp[3]) ? 4'b0001 : 4'b1000;
														assign node10641 = (inp[3]) ? 4'b1100 : node10642;
															assign node10642 = (inp[7]) ? 4'b1000 : node10643;
																assign node10643 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node10648 = (inp[12]) ? node10658 : node10649;
													assign node10649 = (inp[7]) ? node10651 : 4'b0100;
														assign node10651 = (inp[2]) ? node10653 : 4'b0000;
															assign node10653 = (inp[3]) ? node10655 : 4'b0100;
																assign node10655 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node10658 = (inp[2]) ? node10664 : node10659;
														assign node10659 = (inp[3]) ? node10661 : 4'b0000;
															assign node10661 = (inp[4]) ? 4'b1001 : 4'b0100;
														assign node10664 = (inp[3]) ? node10670 : node10665;
															assign node10665 = (inp[7]) ? node10667 : 4'b0100;
																assign node10667 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node10670 = (inp[4]) ? 4'b0000 : node10671;
																assign node10671 = (inp[7]) ? 4'b0100 : 4'b0000;
									assign node10675 = (inp[3]) ? node10791 : node10676;
										assign node10676 = (inp[2]) ? node10744 : node10677;
											assign node10677 = (inp[12]) ? node10713 : node10678;
												assign node10678 = (inp[13]) ? node10700 : node10679;
													assign node10679 = (inp[14]) ? node10691 : node10680;
														assign node10680 = (inp[4]) ? node10688 : node10681;
															assign node10681 = (inp[10]) ? node10685 : node10682;
																assign node10682 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node10685 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node10688 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node10691 = (inp[4]) ? node10697 : node10692;
															assign node10692 = (inp[10]) ? node10694 : 4'b1001;
																assign node10694 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node10697 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node10700 = (inp[4]) ? node10708 : node10701;
														assign node10701 = (inp[7]) ? node10703 : 4'b0001;
															assign node10703 = (inp[10]) ? 4'b0001 : node10704;
																assign node10704 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node10708 = (inp[10]) ? 4'b0000 : node10709;
															assign node10709 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node10713 = (inp[4]) ? node10731 : node10714;
													assign node10714 = (inp[14]) ? node10722 : node10715;
														assign node10715 = (inp[10]) ? node10717 : 4'b0100;
															assign node10717 = (inp[13]) ? 4'b1001 : node10718;
																assign node10718 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node10722 = (inp[10]) ? node10724 : 4'b1001;
															assign node10724 = (inp[13]) ? node10728 : node10725;
																assign node10725 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node10728 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node10731 = (inp[13]) ? node10737 : node10732;
														assign node10732 = (inp[10]) ? node10734 : 4'b1001;
															assign node10734 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node10737 = (inp[14]) ? 4'b1000 : node10738;
															assign node10738 = (inp[7]) ? 4'b1001 : node10739;
																assign node10739 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node10744 = (inp[10]) ? node10766 : node10745;
												assign node10745 = (inp[4]) ? node10751 : node10746;
													assign node10746 = (inp[7]) ? 4'b1000 : node10747;
														assign node10747 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node10751 = (inp[14]) ? node10761 : node10752;
														assign node10752 = (inp[12]) ? node10756 : node10753;
															assign node10753 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node10756 = (inp[13]) ? 4'b0100 : node10757;
																assign node10757 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node10761 = (inp[13]) ? 4'b0001 : node10762;
															assign node10762 = (inp[7]) ? 4'b1100 : 4'b1001;
												assign node10766 = (inp[4]) ? node10778 : node10767;
													assign node10767 = (inp[13]) ? node10771 : node10768;
														assign node10768 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node10771 = (inp[7]) ? 4'b0100 : node10772;
															assign node10772 = (inp[14]) ? node10774 : 4'b0000;
																assign node10774 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node10778 = (inp[7]) ? node10786 : node10779;
														assign node10779 = (inp[13]) ? node10783 : node10780;
															assign node10780 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node10783 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node10786 = (inp[14]) ? 4'b0001 : node10787;
															assign node10787 = (inp[12]) ? 4'b0100 : 4'b0001;
										assign node10791 = (inp[4]) ? node10855 : node10792;
											assign node10792 = (inp[10]) ? node10822 : node10793;
												assign node10793 = (inp[12]) ? node10811 : node10794;
													assign node10794 = (inp[7]) ? node10804 : node10795;
														assign node10795 = (inp[13]) ? node10801 : node10796;
															assign node10796 = (inp[2]) ? 4'b0000 : node10797;
																assign node10797 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node10801 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node10804 = (inp[2]) ? 4'b1000 : node10805;
															assign node10805 = (inp[14]) ? 4'b1000 : node10806;
																assign node10806 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node10811 = (inp[7]) ? node10813 : 4'b0000;
														assign node10813 = (inp[2]) ? node10819 : node10814;
															assign node10814 = (inp[13]) ? node10816 : 4'b0000;
																assign node10816 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10819 = (inp[13]) ? 4'b0000 : 4'b1001;
												assign node10822 = (inp[13]) ? node10844 : node10823;
													assign node10823 = (inp[2]) ? node10831 : node10824;
														assign node10824 = (inp[7]) ? node10826 : 4'b1001;
															assign node10826 = (inp[14]) ? 4'b0001 : node10827;
																assign node10827 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10831 = (inp[14]) ? node10839 : node10832;
															assign node10832 = (inp[7]) ? node10836 : node10833;
																assign node10833 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node10836 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10839 = (inp[12]) ? 4'b0000 : node10840;
																assign node10840 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node10844 = (inp[2]) ? node10848 : node10845;
														assign node10845 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10848 = (inp[7]) ? node10850 : 4'b1001;
															assign node10850 = (inp[14]) ? 4'b1001 : node10851;
																assign node10851 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node10855 = (inp[7]) ? node10869 : node10856;
												assign node10856 = (inp[13]) ? node10864 : node10857;
													assign node10857 = (inp[14]) ? 4'b0001 : node10858;
														assign node10858 = (inp[2]) ? node10860 : 4'b1000;
															assign node10860 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node10864 = (inp[10]) ? 4'b0000 : node10865;
														assign node10865 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node10869 = (inp[13]) ? 4'b0000 : node10870;
													assign node10870 = (inp[2]) ? node10882 : node10871;
														assign node10871 = (inp[10]) ? node10877 : node10872;
															assign node10872 = (inp[12]) ? node10874 : 4'b0001;
																assign node10874 = (inp[14]) ? 4'b1000 : 4'b0000;
															assign node10877 = (inp[12]) ? node10879 : 4'b0000;
																assign node10879 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10882 = (inp[10]) ? node10884 : 4'b0000;
															assign node10884 = (inp[14]) ? node10886 : 4'b0000;
																assign node10886 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node10890 = (inp[5]) ? node11042 : node10891;
									assign node10891 = (inp[10]) ? node10987 : node10892;
										assign node10892 = (inp[3]) ? node10944 : node10893;
											assign node10893 = (inp[7]) ? node10921 : node10894;
												assign node10894 = (inp[2]) ? node10906 : node10895;
													assign node10895 = (inp[14]) ? node10901 : node10896;
														assign node10896 = (inp[13]) ? 4'b1001 : node10897;
															assign node10897 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10901 = (inp[4]) ? node10903 : 4'b0101;
															assign node10903 = (inp[13]) ? 4'b1001 : 4'b0101;
													assign node10906 = (inp[4]) ? node10914 : node10907;
														assign node10907 = (inp[13]) ? node10911 : node10908;
															assign node10908 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10911 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node10914 = (inp[13]) ? node10918 : node10915;
															assign node10915 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node10918 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node10921 = (inp[2]) ? node10931 : node10922;
													assign node10922 = (inp[12]) ? node10928 : node10923;
														assign node10923 = (inp[13]) ? node10925 : 4'b1001;
															assign node10925 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node10928 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node10931 = (inp[4]) ? node10939 : node10932;
														assign node10932 = (inp[12]) ? node10936 : node10933;
															assign node10933 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node10936 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node10939 = (inp[12]) ? node10941 : 4'b1001;
															assign node10941 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node10944 = (inp[2]) ? node10956 : node10945;
												assign node10945 = (inp[4]) ? node10949 : node10946;
													assign node10946 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node10949 = (inp[13]) ? node10951 : 4'b1101;
														assign node10951 = (inp[7]) ? 4'b1101 : node10952;
															assign node10952 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node10956 = (inp[7]) ? node10970 : node10957;
													assign node10957 = (inp[4]) ? node10965 : node10958;
														assign node10958 = (inp[12]) ? node10962 : node10959;
															assign node10959 = (inp[13]) ? 4'b0001 : 4'b1101;
															assign node10962 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node10965 = (inp[12]) ? node10967 : 4'b1001;
															assign node10967 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node10970 = (inp[4]) ? node10980 : node10971;
														assign node10971 = (inp[14]) ? 4'b1101 : node10972;
															assign node10972 = (inp[13]) ? node10976 : node10973;
																assign node10973 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node10976 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node10980 = (inp[13]) ? node10984 : node10981;
															assign node10981 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node10984 = (inp[12]) ? 4'b1101 : 4'b0001;
										assign node10987 = (inp[13]) ? node11017 : node10988;
											assign node10988 = (inp[3]) ? node10998 : node10989;
												assign node10989 = (inp[7]) ? 4'b1001 : node10990;
													assign node10990 = (inp[2]) ? node10994 : node10991;
														assign node10991 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node10994 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node10998 = (inp[2]) ? node11012 : node10999;
													assign node10999 = (inp[14]) ? node11005 : node11000;
														assign node11000 = (inp[7]) ? node11002 : 4'b0101;
															assign node11002 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node11005 = (inp[7]) ? node11009 : node11006;
															assign node11006 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node11009 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node11012 = (inp[4]) ? node11014 : 4'b1101;
														assign node11014 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node11017 = (inp[4]) ? node11037 : node11018;
												assign node11018 = (inp[2]) ? node11024 : node11019;
													assign node11019 = (inp[3]) ? 4'b0101 : node11020;
														assign node11020 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node11024 = (inp[12]) ? node11032 : node11025;
														assign node11025 = (inp[3]) ? node11029 : node11026;
															assign node11026 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node11029 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node11032 = (inp[3]) ? 4'b0001 : node11033;
															assign node11033 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node11037 = (inp[3]) ? 4'b0001 : node11038;
													assign node11038 = (inp[2]) ? 4'b0101 : 4'b0001;
									assign node11042 = (inp[3]) ? node11114 : node11043;
										assign node11043 = (inp[13]) ? node11085 : node11044;
											assign node11044 = (inp[12]) ? node11066 : node11045;
												assign node11045 = (inp[10]) ? node11053 : node11046;
													assign node11046 = (inp[2]) ? node11050 : node11047;
														assign node11047 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11050 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node11053 = (inp[2]) ? node11061 : node11054;
														assign node11054 = (inp[4]) ? node11058 : node11055;
															assign node11055 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node11058 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node11061 = (inp[4]) ? 4'b1001 : node11062;
															assign node11062 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node11066 = (inp[10]) ? node11072 : node11067;
													assign node11067 = (inp[4]) ? node11069 : 4'b1001;
														assign node11069 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node11072 = (inp[14]) ? node11080 : node11073;
														assign node11073 = (inp[2]) ? 4'b0101 : node11074;
															assign node11074 = (inp[4]) ? node11076 : 4'b1001;
																assign node11076 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node11080 = (inp[7]) ? node11082 : 4'b1001;
															assign node11082 = (inp[4]) ? 4'b0101 : 4'b1001;
											assign node11085 = (inp[10]) ? node11107 : node11086;
												assign node11086 = (inp[4]) ? node11096 : node11087;
													assign node11087 = (inp[2]) ? node11093 : node11088;
														assign node11088 = (inp[7]) ? node11090 : 4'b0001;
															assign node11090 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node11093 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node11096 = (inp[2]) ? node11102 : node11097;
														assign node11097 = (inp[12]) ? 4'b1001 : node11098;
															assign node11098 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11102 = (inp[7]) ? node11104 : 4'b0001;
															assign node11104 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node11107 = (inp[7]) ? node11109 : 4'b0001;
													assign node11109 = (inp[4]) ? 4'b0001 : node11110;
														assign node11110 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node11114 = (inp[4]) ? node11150 : node11115;
											assign node11115 = (inp[10]) ? node11143 : node11116;
												assign node11116 = (inp[13]) ? node11134 : node11117;
													assign node11117 = (inp[7]) ? node11129 : node11118;
														assign node11118 = (inp[14]) ? node11124 : node11119;
															assign node11119 = (inp[2]) ? 4'b1001 : node11120;
																assign node11120 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node11124 = (inp[12]) ? 4'b0001 : node11125;
																assign node11125 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node11129 = (inp[2]) ? 4'b0001 : node11130;
															assign node11130 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11134 = (inp[12]) ? node11138 : node11135;
														assign node11135 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node11138 = (inp[7]) ? 4'b1001 : node11139;
															assign node11139 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node11143 = (inp[13]) ? 4'b0001 : node11144;
													assign node11144 = (inp[2]) ? node11146 : 4'b0001;
														assign node11146 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node11150 = (inp[13]) ? node11160 : node11151;
												assign node11151 = (inp[10]) ? 4'b0001 : node11152;
													assign node11152 = (inp[7]) ? node11154 : 4'b0001;
														assign node11154 = (inp[2]) ? node11156 : 4'b0001;
															assign node11156 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node11160 = (inp[10]) ? 4'b0000 : 4'b0001;
					assign node11163 = (inp[6]) ? node11165 : 4'b0001;
						assign node11165 = (inp[5]) ? node11255 : node11166;
							assign node11166 = (inp[2]) ? 4'b0001 : node11167;
								assign node11167 = (inp[3]) ? node11169 : 4'b0001;
									assign node11169 = (inp[4]) ? node11193 : node11170;
										assign node11170 = (inp[7]) ? 4'b0001 : node11171;
											assign node11171 = (inp[13]) ? node11173 : 4'b0001;
												assign node11173 = (inp[14]) ? node11179 : node11174;
													assign node11174 = (inp[1]) ? 4'b0001 : node11175;
														assign node11175 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node11179 = (inp[10]) ? node11185 : node11180;
														assign node11180 = (inp[11]) ? 4'b0001 : node11181;
															assign node11181 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node11185 = (inp[1]) ? node11189 : node11186;
															assign node11186 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node11189 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node11193 = (inp[7]) ? node11233 : node11194;
											assign node11194 = (inp[1]) ? node11216 : node11195;
												assign node11195 = (inp[11]) ? node11209 : node11196;
													assign node11196 = (inp[14]) ? node11206 : node11197;
														assign node11197 = (inp[12]) ? node11199 : 4'b0000;
															assign node11199 = (inp[13]) ? node11203 : node11200;
																assign node11200 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node11203 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node11206 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node11209 = (inp[13]) ? node11211 : 4'b1000;
														assign node11211 = (inp[12]) ? node11213 : 4'b0000;
															assign node11213 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node11216 = (inp[13]) ? node11226 : node11217;
													assign node11217 = (inp[12]) ? node11219 : 4'b1001;
														assign node11219 = (inp[10]) ? node11223 : node11220;
															assign node11220 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11223 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11226 = (inp[10]) ? 4'b0001 : node11227;
														assign node11227 = (inp[12]) ? node11229 : 4'b0001;
															assign node11229 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node11233 = (inp[13]) ? node11235 : 4'b0001;
												assign node11235 = (inp[1]) ? node11249 : node11236;
													assign node11236 = (inp[12]) ? node11242 : node11237;
														assign node11237 = (inp[10]) ? node11239 : 4'b0000;
															assign node11239 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11242 = (inp[10]) ? node11244 : 4'b0001;
															assign node11244 = (inp[14]) ? node11246 : 4'b0000;
																assign node11246 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node11249 = (inp[14]) ? node11251 : 4'b0001;
														assign node11251 = (inp[11]) ? 4'b0001 : 4'b0000;
							assign node11255 = (inp[2]) ? node11601 : node11256;
								assign node11256 = (inp[3]) ? node11428 : node11257;
									assign node11257 = (inp[1]) ? node11351 : node11258;
										assign node11258 = (inp[14]) ? node11300 : node11259;
											assign node11259 = (inp[13]) ? node11277 : node11260;
												assign node11260 = (inp[4]) ? node11266 : node11261;
													assign node11261 = (inp[10]) ? 4'b1000 : node11262;
														assign node11262 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11266 = (inp[7]) ? node11274 : node11267;
														assign node11267 = (inp[10]) ? node11269 : 4'b1100;
															assign node11269 = (inp[12]) ? 4'b1100 : node11270;
																assign node11270 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node11274 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node11277 = (inp[7]) ? node11293 : node11278;
													assign node11278 = (inp[4]) ? node11282 : node11279;
														assign node11279 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node11282 = (inp[11]) ? node11288 : node11283;
															assign node11283 = (inp[10]) ? node11285 : 4'b1000;
																assign node11285 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node11288 = (inp[12]) ? 4'b1001 : node11289;
																assign node11289 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node11293 = (inp[4]) ? node11295 : 4'b0000;
														assign node11295 = (inp[11]) ? node11297 : 4'b0100;
															assign node11297 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node11300 = (inp[11]) ? node11332 : node11301;
												assign node11301 = (inp[13]) ? node11313 : node11302;
													assign node11302 = (inp[4]) ? node11308 : node11303;
														assign node11303 = (inp[12]) ? 4'b0001 : node11304;
															assign node11304 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11308 = (inp[7]) ? node11310 : 4'b0101;
															assign node11310 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node11313 = (inp[4]) ? node11319 : node11314;
														assign node11314 = (inp[12]) ? 4'b1001 : node11315;
															assign node11315 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node11319 = (inp[7]) ? node11327 : node11320;
															assign node11320 = (inp[10]) ? node11324 : node11321;
																assign node11321 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node11324 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node11327 = (inp[10]) ? node11329 : 4'b1001;
																assign node11329 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node11332 = (inp[13]) ? node11342 : node11333;
													assign node11333 = (inp[10]) ? 4'b1000 : node11334;
														assign node11334 = (inp[12]) ? node11338 : node11335;
															assign node11335 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node11338 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node11342 = (inp[4]) ? node11348 : node11343;
														assign node11343 = (inp[7]) ? 4'b0000 : node11344;
															assign node11344 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node11348 = (inp[12]) ? 4'b0100 : 4'b0001;
										assign node11351 = (inp[11]) ? node11395 : node11352;
											assign node11352 = (inp[14]) ? node11374 : node11353;
												assign node11353 = (inp[4]) ? node11365 : node11354;
													assign node11354 = (inp[13]) ? node11358 : node11355;
														assign node11355 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node11358 = (inp[10]) ? node11362 : node11359;
															assign node11359 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node11362 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node11365 = (inp[7]) ? node11369 : node11366;
														assign node11366 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node11369 = (inp[13]) ? node11371 : 4'b1001;
															assign node11371 = (inp[10]) ? 4'b0000 : 4'b0101;
												assign node11374 = (inp[7]) ? node11388 : node11375;
													assign node11375 = (inp[10]) ? node11383 : node11376;
														assign node11376 = (inp[13]) ? node11378 : 4'b0100;
															assign node11378 = (inp[4]) ? 4'b1000 : node11379;
																assign node11379 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node11383 = (inp[4]) ? 4'b0000 : node11384;
															assign node11384 = (inp[13]) ? 4'b0100 : 4'b1000;
													assign node11388 = (inp[13]) ? node11392 : node11389;
														assign node11389 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node11392 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node11395 = (inp[13]) ? node11413 : node11396;
												assign node11396 = (inp[12]) ? node11402 : node11397;
													assign node11397 = (inp[7]) ? 4'b1001 : node11398;
														assign node11398 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node11402 = (inp[10]) ? node11408 : node11403;
														assign node11403 = (inp[7]) ? 4'b0001 : node11404;
															assign node11404 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node11408 = (inp[4]) ? node11410 : 4'b1001;
															assign node11410 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node11413 = (inp[10]) ? node11423 : node11414;
													assign node11414 = (inp[12]) ? 4'b1001 : node11415;
														assign node11415 = (inp[4]) ? node11419 : node11416;
															assign node11416 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node11419 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node11423 = (inp[4]) ? 4'b0001 : node11424;
														assign node11424 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node11428 = (inp[4]) ? node11506 : node11429;
										assign node11429 = (inp[11]) ? node11475 : node11430;
											assign node11430 = (inp[13]) ? node11452 : node11431;
												assign node11431 = (inp[10]) ? node11441 : node11432;
													assign node11432 = (inp[12]) ? node11438 : node11433;
														assign node11433 = (inp[1]) ? node11435 : 4'b1000;
															assign node11435 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node11438 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node11441 = (inp[7]) ? node11447 : node11442;
														assign node11442 = (inp[1]) ? 4'b1000 : node11443;
															assign node11443 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11447 = (inp[12]) ? node11449 : 4'b0000;
															assign node11449 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node11452 = (inp[1]) ? node11462 : node11453;
													assign node11453 = (inp[14]) ? 4'b1000 : node11454;
														assign node11454 = (inp[10]) ? 4'b1001 : node11455;
															assign node11455 = (inp[12]) ? node11457 : 4'b0001;
																assign node11457 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node11462 = (inp[12]) ? node11468 : node11463;
														assign node11463 = (inp[14]) ? node11465 : 4'b0001;
															assign node11465 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node11468 = (inp[10]) ? node11472 : node11469;
															assign node11469 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node11472 = (inp[7]) ? 4'b0000 : 4'b1001;
											assign node11475 = (inp[13]) ? node11499 : node11476;
												assign node11476 = (inp[7]) ? node11488 : node11477;
													assign node11477 = (inp[10]) ? node11483 : node11478;
														assign node11478 = (inp[12]) ? 4'b0001 : node11479;
															assign node11479 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node11483 = (inp[1]) ? 4'b1001 : node11484;
															assign node11484 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11488 = (inp[10]) ? node11494 : node11489;
														assign node11489 = (inp[1]) ? 4'b1001 : node11490;
															assign node11490 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node11494 = (inp[1]) ? 4'b0001 : node11495;
															assign node11495 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node11499 = (inp[1]) ? 4'b0001 : node11500;
													assign node11500 = (inp[10]) ? node11502 : 4'b0000;
														assign node11502 = (inp[7]) ? 4'b0000 : 4'b1001;
										assign node11506 = (inp[13]) ? node11560 : node11507;
											assign node11507 = (inp[10]) ? node11537 : node11508;
												assign node11508 = (inp[7]) ? node11522 : node11509;
													assign node11509 = (inp[14]) ? node11513 : node11510;
														assign node11510 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node11513 = (inp[11]) ? node11517 : node11514;
															assign node11514 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node11517 = (inp[1]) ? node11519 : 4'b1000;
																assign node11519 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node11522 = (inp[14]) ? node11534 : node11523;
														assign node11523 = (inp[11]) ? node11529 : node11524;
															assign node11524 = (inp[12]) ? 4'b0001 : node11525;
																assign node11525 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node11529 = (inp[12]) ? 4'b1001 : node11530;
																assign node11530 = (inp[1]) ? 4'b1001 : 4'b0000;
														assign node11534 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node11537 = (inp[11]) ? node11553 : node11538;
													assign node11538 = (inp[1]) ? node11544 : node11539;
														assign node11539 = (inp[14]) ? node11541 : 4'b0000;
															assign node11541 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11544 = (inp[14]) ? node11550 : node11545;
															assign node11545 = (inp[7]) ? node11547 : 4'b0001;
																assign node11547 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11550 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node11553 = (inp[12]) ? 4'b0001 : node11554;
														assign node11554 = (inp[7]) ? node11556 : 4'b0001;
															assign node11556 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node11560 = (inp[10]) ? node11586 : node11561;
												assign node11561 = (inp[1]) ? node11573 : node11562;
													assign node11562 = (inp[7]) ? node11566 : node11563;
														assign node11563 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node11566 = (inp[12]) ? node11568 : 4'b0000;
															assign node11568 = (inp[14]) ? node11570 : 4'b0000;
																assign node11570 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node11573 = (inp[11]) ? 4'b0001 : node11574;
														assign node11574 = (inp[12]) ? node11580 : node11575;
															assign node11575 = (inp[14]) ? 4'b0000 : node11576;
																assign node11576 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node11580 = (inp[7]) ? node11582 : 4'b0001;
																assign node11582 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node11586 = (inp[1]) ? 4'b0000 : node11587;
													assign node11587 = (inp[11]) ? 4'b0000 : node11588;
														assign node11588 = (inp[12]) ? node11594 : node11589;
															assign node11589 = (inp[14]) ? 4'b0001 : node11590;
																assign node11590 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11594 = (inp[14]) ? 4'b0000 : node11595;
																assign node11595 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node11601 = (inp[3]) ? node11603 : 4'b0001;
									assign node11603 = (inp[4]) ? node11629 : node11604;
										assign node11604 = (inp[7]) ? 4'b0001 : node11605;
											assign node11605 = (inp[13]) ? node11607 : 4'b0001;
												assign node11607 = (inp[10]) ? node11617 : node11608;
													assign node11608 = (inp[12]) ? 4'b0001 : node11609;
														assign node11609 = (inp[14]) ? node11611 : 4'b0001;
															assign node11611 = (inp[1]) ? 4'b0000 : node11612;
																assign node11612 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node11617 = (inp[1]) ? node11623 : node11618;
														assign node11618 = (inp[11]) ? 4'b0000 : node11619;
															assign node11619 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11623 = (inp[14]) ? node11625 : 4'b0001;
															assign node11625 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node11629 = (inp[13]) ? node11655 : node11630;
											assign node11630 = (inp[7]) ? 4'b0001 : node11631;
												assign node11631 = (inp[1]) ? node11643 : node11632;
													assign node11632 = (inp[11]) ? node11638 : node11633;
														assign node11633 = (inp[10]) ? 4'b0000 : node11634;
															assign node11634 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node11638 = (inp[10]) ? 4'b1000 : node11639;
															assign node11639 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node11643 = (inp[10]) ? node11651 : node11644;
														assign node11644 = (inp[12]) ? 4'b0001 : node11645;
															assign node11645 = (inp[14]) ? node11647 : 4'b1001;
																assign node11647 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11651 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node11655 = (inp[10]) ? node11673 : node11656;
												assign node11656 = (inp[1]) ? node11664 : node11657;
													assign node11657 = (inp[7]) ? node11661 : node11658;
														assign node11658 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11661 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node11664 = (inp[11]) ? 4'b0001 : node11665;
														assign node11665 = (inp[12]) ? node11667 : 4'b0000;
															assign node11667 = (inp[14]) ? 4'b0001 : node11668;
																assign node11668 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node11673 = (inp[1]) ? 4'b0000 : node11674;
													assign node11674 = (inp[11]) ? 4'b0000 : node11675;
														assign node11675 = (inp[12]) ? node11681 : node11676;
															assign node11676 = (inp[7]) ? 4'b0000 : node11677;
																assign node11677 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11681 = (inp[7]) ? 4'b0001 : 4'b0000;
		assign node11686 = (inp[9]) ? node17344 : node11687;
			assign node11687 = (inp[15]) ? node14749 : node11688;
				assign node11688 = (inp[6]) ? node12406 : node11689;
					assign node11689 = (inp[0]) ? 4'b1100 : node11690;
						assign node11690 = (inp[2]) ? node12118 : node11691;
							assign node11691 = (inp[1]) ? node11881 : node11692;
								assign node11692 = (inp[13]) ? node11798 : node11693;
									assign node11693 = (inp[10]) ? node11735 : node11694;
										assign node11694 = (inp[3]) ? node11718 : node11695;
											assign node11695 = (inp[5]) ? node11705 : node11696;
												assign node11696 = (inp[7]) ? 4'b1110 : node11697;
													assign node11697 = (inp[4]) ? node11699 : 4'b1110;
														assign node11699 = (inp[11]) ? 4'b1001 : node11700;
															assign node11700 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node11705 = (inp[7]) ? node11713 : node11706;
													assign node11706 = (inp[4]) ? node11708 : 4'b1101;
														assign node11708 = (inp[11]) ? 4'b1001 : node11709;
															assign node11709 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node11713 = (inp[14]) ? node11715 : 4'b1101;
														assign node11715 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node11718 = (inp[11]) ? node11730 : node11719;
												assign node11719 = (inp[14]) ? node11725 : node11720;
													assign node11720 = (inp[7]) ? 4'b1001 : node11721;
														assign node11721 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node11725 = (inp[4]) ? node11727 : 4'b1000;
														assign node11727 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node11730 = (inp[7]) ? 4'b1001 : node11731;
													assign node11731 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node11735 = (inp[12]) ? node11765 : node11736;
											assign node11736 = (inp[3]) ? node11752 : node11737;
												assign node11737 = (inp[4]) ? node11747 : node11738;
													assign node11738 = (inp[7]) ? node11740 : 4'b0001;
														assign node11740 = (inp[5]) ? node11742 : 4'b1110;
															assign node11742 = (inp[11]) ? 4'b0101 : node11743;
																assign node11743 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node11747 = (inp[14]) ? node11749 : 4'b0001;
														assign node11749 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node11752 = (inp[4]) ? node11760 : node11753;
													assign node11753 = (inp[7]) ? node11755 : 4'b0101;
														assign node11755 = (inp[11]) ? 4'b0001 : node11756;
															assign node11756 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11760 = (inp[11]) ? 4'b0101 : node11761;
														assign node11761 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node11765 = (inp[3]) ? node11783 : node11766;
												assign node11766 = (inp[5]) ? node11772 : node11767;
													assign node11767 = (inp[7]) ? 4'b1110 : node11768;
														assign node11768 = (inp[4]) ? 4'b1001 : 4'b1110;
													assign node11772 = (inp[11]) ? node11780 : node11773;
														assign node11773 = (inp[14]) ? node11775 : 4'b1101;
															assign node11775 = (inp[7]) ? 4'b1100 : node11776;
																assign node11776 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node11780 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node11783 = (inp[4]) ? node11789 : node11784;
													assign node11784 = (inp[14]) ? node11786 : 4'b1001;
														assign node11786 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11789 = (inp[7]) ? node11795 : node11790;
														assign node11790 = (inp[11]) ? 4'b1101 : node11791;
															assign node11791 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node11795 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node11798 = (inp[3]) ? node11840 : node11799;
										assign node11799 = (inp[7]) ? node11813 : node11800;
											assign node11800 = (inp[11]) ? node11808 : node11801;
												assign node11801 = (inp[14]) ? node11803 : 4'b0001;
													assign node11803 = (inp[10]) ? node11805 : 4'b0000;
														assign node11805 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node11808 = (inp[10]) ? node11810 : 4'b0001;
													assign node11810 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node11813 = (inp[4]) ? node11825 : node11814;
												assign node11814 = (inp[5]) ? node11816 : 4'b1110;
													assign node11816 = (inp[10]) ? node11822 : node11817;
														assign node11817 = (inp[14]) ? node11819 : 4'b0101;
															assign node11819 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node11822 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node11825 = (inp[14]) ? node11831 : node11826;
													assign node11826 = (inp[12]) ? 4'b0001 : node11827;
														assign node11827 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node11831 = (inp[11]) ? node11837 : node11832;
														assign node11832 = (inp[10]) ? node11834 : 4'b0000;
															assign node11834 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11837 = (inp[5]) ? 4'b0001 : 4'b1001;
										assign node11840 = (inp[12]) ? node11864 : node11841;
											assign node11841 = (inp[10]) ? node11851 : node11842;
												assign node11842 = (inp[11]) ? node11846 : node11843;
													assign node11843 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node11846 = (inp[7]) ? node11848 : 4'b0101;
														assign node11848 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node11851 = (inp[11]) ? node11859 : node11852;
													assign node11852 = (inp[14]) ? node11854 : 4'b1101;
														assign node11854 = (inp[4]) ? 4'b1100 : node11855;
															assign node11855 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node11859 = (inp[4]) ? 4'b1101 : node11860;
														assign node11860 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node11864 = (inp[7]) ? node11870 : node11865;
												assign node11865 = (inp[11]) ? 4'b0101 : node11866;
													assign node11866 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node11870 = (inp[4]) ? node11876 : node11871;
													assign node11871 = (inp[11]) ? 4'b0001 : node11872;
														assign node11872 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11876 = (inp[11]) ? 4'b0101 : node11877;
														assign node11877 = (inp[14]) ? 4'b0100 : 4'b0101;
								assign node11881 = (inp[11]) ? node12037 : node11882;
									assign node11882 = (inp[14]) ? node11956 : node11883;
										assign node11883 = (inp[13]) ? node11923 : node11884;
											assign node11884 = (inp[12]) ? node11898 : node11885;
												assign node11885 = (inp[3]) ? node11893 : node11886;
													assign node11886 = (inp[7]) ? node11888 : 4'b0000;
														assign node11888 = (inp[4]) ? 4'b0000 : node11889;
															assign node11889 = (inp[10]) ? 4'b1110 : 4'b0100;
													assign node11893 = (inp[7]) ? node11895 : 4'b0100;
														assign node11895 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node11898 = (inp[10]) ? node11910 : node11899;
													assign node11899 = (inp[3]) ? node11905 : node11900;
														assign node11900 = (inp[5]) ? node11902 : 4'b1110;
															assign node11902 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node11905 = (inp[7]) ? 4'b1000 : node11906;
															assign node11906 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node11910 = (inp[3]) ? node11918 : node11911;
														assign node11911 = (inp[4]) ? 4'b0000 : node11912;
															assign node11912 = (inp[5]) ? node11914 : 4'b1110;
																assign node11914 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node11918 = (inp[4]) ? 4'b0100 : node11919;
															assign node11919 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node11923 = (inp[10]) ? node11943 : node11924;
												assign node11924 = (inp[12]) ? node11934 : node11925;
													assign node11925 = (inp[3]) ? node11929 : node11926;
														assign node11926 = (inp[5]) ? 4'b1000 : 4'b1110;
														assign node11929 = (inp[4]) ? 4'b1100 : node11930;
															assign node11930 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node11934 = (inp[3]) ? node11940 : node11935;
														assign node11935 = (inp[7]) ? node11937 : 4'b0000;
															assign node11937 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node11940 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node11943 = (inp[3]) ? node11951 : node11944;
													assign node11944 = (inp[7]) ? node11946 : 4'b1000;
														assign node11946 = (inp[5]) ? node11948 : 4'b1110;
															assign node11948 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node11951 = (inp[7]) ? node11953 : 4'b1100;
														assign node11953 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node11956 = (inp[13]) ? node12000 : node11957;
											assign node11957 = (inp[3]) ? node11985 : node11958;
												assign node11958 = (inp[5]) ? node11972 : node11959;
													assign node11959 = (inp[4]) ? node11961 : 4'b1110;
														assign node11961 = (inp[7]) ? node11967 : node11962;
															assign node11962 = (inp[10]) ? node11964 : 4'b1001;
																assign node11964 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node11967 = (inp[10]) ? node11969 : 4'b1110;
																assign node11969 = (inp[12]) ? 4'b1110 : 4'b0001;
													assign node11972 = (inp[4]) ? node11978 : node11973;
														assign node11973 = (inp[12]) ? 4'b1101 : node11974;
															assign node11974 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node11978 = (inp[12]) ? node11982 : node11979;
															assign node11979 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node11982 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node11985 = (inp[12]) ? node11995 : node11986;
													assign node11986 = (inp[10]) ? node11990 : node11987;
														assign node11987 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node11990 = (inp[7]) ? node11992 : 4'b0101;
															assign node11992 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node11995 = (inp[4]) ? node11997 : 4'b1001;
														assign node11997 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node12000 = (inp[3]) ? node12020 : node12001;
												assign node12001 = (inp[12]) ? node12013 : node12002;
													assign node12002 = (inp[10]) ? node12006 : node12003;
														assign node12003 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node12006 = (inp[7]) ? node12008 : 4'b1001;
															assign node12008 = (inp[4]) ? 4'b1001 : node12009;
																assign node12009 = (inp[5]) ? 4'b1101 : 4'b1110;
													assign node12013 = (inp[4]) ? 4'b0001 : node12014;
														assign node12014 = (inp[7]) ? node12016 : 4'b0001;
															assign node12016 = (inp[5]) ? 4'b0101 : 4'b1110;
												assign node12020 = (inp[7]) ? node12026 : node12021;
													assign node12021 = (inp[10]) ? node12023 : 4'b0101;
														assign node12023 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node12026 = (inp[4]) ? node12032 : node12027;
														assign node12027 = (inp[10]) ? node12029 : 4'b0001;
															assign node12029 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12032 = (inp[10]) ? node12034 : 4'b0101;
															assign node12034 = (inp[12]) ? 4'b0101 : 4'b1101;
									assign node12037 = (inp[13]) ? node12079 : node12038;
										assign node12038 = (inp[12]) ? node12052 : node12039;
											assign node12039 = (inp[3]) ? node12047 : node12040;
												assign node12040 = (inp[4]) ? 4'b0000 : node12041;
													assign node12041 = (inp[7]) ? node12043 : 4'b0000;
														assign node12043 = (inp[5]) ? 4'b0100 : 4'b1110;
												assign node12047 = (inp[4]) ? 4'b0100 : node12048;
													assign node12048 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node12052 = (inp[10]) ? node12066 : node12053;
												assign node12053 = (inp[3]) ? node12061 : node12054;
													assign node12054 = (inp[7]) ? node12058 : node12055;
														assign node12055 = (inp[4]) ? 4'b1000 : 4'b1110;
														assign node12058 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node12061 = (inp[7]) ? 4'b1000 : node12062;
														assign node12062 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node12066 = (inp[3]) ? node12074 : node12067;
													assign node12067 = (inp[4]) ? 4'b0000 : node12068;
														assign node12068 = (inp[5]) ? 4'b0100 : node12069;
															assign node12069 = (inp[7]) ? 4'b1110 : 4'b0000;
													assign node12074 = (inp[7]) ? node12076 : 4'b0100;
														assign node12076 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node12079 = (inp[3]) ? node12101 : node12080;
											assign node12080 = (inp[12]) ? node12088 : node12081;
												assign node12081 = (inp[7]) ? node12083 : 4'b1000;
													assign node12083 = (inp[4]) ? 4'b1000 : node12084;
														assign node12084 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node12088 = (inp[10]) ? node12096 : node12089;
													assign node12089 = (inp[7]) ? node12091 : 4'b0000;
														assign node12091 = (inp[4]) ? 4'b0000 : node12092;
															assign node12092 = (inp[5]) ? 4'b0100 : 4'b1110;
													assign node12096 = (inp[4]) ? 4'b1000 : node12097;
														assign node12097 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node12101 = (inp[4]) ? node12113 : node12102;
												assign node12102 = (inp[7]) ? node12108 : node12103;
													assign node12103 = (inp[12]) ? node12105 : 4'b1100;
														assign node12105 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node12108 = (inp[10]) ? 4'b1000 : node12109;
														assign node12109 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node12113 = (inp[10]) ? 4'b1100 : node12114;
													assign node12114 = (inp[12]) ? 4'b0100 : 4'b1100;
							assign node12118 = (inp[5]) ? node12120 : 4'b1110;
								assign node12120 = (inp[3]) ? node12240 : node12121;
									assign node12121 = (inp[7]) ? node12191 : node12122;
										assign node12122 = (inp[1]) ? node12156 : node12123;
											assign node12123 = (inp[13]) ? node12139 : node12124;
												assign node12124 = (inp[4]) ? node12130 : node12125;
													assign node12125 = (inp[10]) ? node12127 : 4'b1110;
														assign node12127 = (inp[12]) ? 4'b1110 : 4'b0001;
													assign node12130 = (inp[12]) ? node12134 : node12131;
														assign node12131 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node12134 = (inp[14]) ? node12136 : 4'b1001;
															assign node12136 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node12139 = (inp[12]) ? node12151 : node12140;
													assign node12140 = (inp[10]) ? node12146 : node12141;
														assign node12141 = (inp[11]) ? 4'b0001 : node12142;
															assign node12142 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node12146 = (inp[14]) ? node12148 : 4'b1001;
															assign node12148 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12151 = (inp[14]) ? node12153 : 4'b0001;
														assign node12153 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node12156 = (inp[13]) ? node12174 : node12157;
												assign node12157 = (inp[12]) ? node12163 : node12158;
													assign node12158 = (inp[14]) ? node12160 : 4'b0000;
														assign node12160 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node12163 = (inp[10]) ? node12169 : node12164;
														assign node12164 = (inp[4]) ? node12166 : 4'b1110;
															assign node12166 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node12169 = (inp[14]) ? node12171 : 4'b0000;
															assign node12171 = (inp[11]) ? 4'b0000 : 4'b1110;
												assign node12174 = (inp[11]) ? node12186 : node12175;
													assign node12175 = (inp[14]) ? node12181 : node12176;
														assign node12176 = (inp[10]) ? 4'b1000 : node12177;
															assign node12177 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node12181 = (inp[10]) ? node12183 : 4'b0001;
															assign node12183 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node12186 = (inp[10]) ? 4'b1000 : node12187;
														assign node12187 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node12191 = (inp[4]) ? node12193 : 4'b1110;
											assign node12193 = (inp[13]) ? node12217 : node12194;
												assign node12194 = (inp[10]) ? node12200 : node12195;
													assign node12195 = (inp[12]) ? 4'b1110 : node12196;
														assign node12196 = (inp[1]) ? 4'b0000 : 4'b1110;
													assign node12200 = (inp[12]) ? node12210 : node12201;
														assign node12201 = (inp[14]) ? node12203 : 4'b0001;
															assign node12203 = (inp[1]) ? node12207 : node12204;
																assign node12204 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node12207 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node12210 = (inp[1]) ? node12212 : 4'b1110;
															assign node12212 = (inp[11]) ? 4'b0000 : node12213;
																assign node12213 = (inp[14]) ? 4'b1110 : 4'b0000;
												assign node12217 = (inp[1]) ? node12229 : node12218;
													assign node12218 = (inp[14]) ? node12224 : node12219;
														assign node12219 = (inp[10]) ? node12221 : 4'b0001;
															assign node12221 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12224 = (inp[12]) ? node12226 : 4'b1000;
															assign node12226 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node12229 = (inp[14]) ? node12235 : node12230;
														assign node12230 = (inp[12]) ? node12232 : 4'b1000;
															assign node12232 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12235 = (inp[10]) ? 4'b1001 : node12236;
															assign node12236 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node12240 = (inp[1]) ? node12312 : node12241;
										assign node12241 = (inp[13]) ? node12279 : node12242;
											assign node12242 = (inp[7]) ? node12266 : node12243;
												assign node12243 = (inp[4]) ? node12253 : node12244;
													assign node12244 = (inp[10]) ? node12250 : node12245;
														assign node12245 = (inp[14]) ? node12247 : 4'b1001;
															assign node12247 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12250 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node12253 = (inp[12]) ? node12261 : node12254;
														assign node12254 = (inp[10]) ? node12256 : 4'b1101;
															assign node12256 = (inp[14]) ? node12258 : 4'b0101;
																assign node12258 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node12261 = (inp[11]) ? 4'b1101 : node12262;
															assign node12262 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node12266 = (inp[11]) ? node12274 : node12267;
													assign node12267 = (inp[14]) ? 4'b1000 : node12268;
														assign node12268 = (inp[12]) ? 4'b1001 : node12269;
															assign node12269 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node12274 = (inp[12]) ? 4'b1001 : node12275;
														assign node12275 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node12279 = (inp[11]) ? node12295 : node12280;
												assign node12280 = (inp[14]) ? node12288 : node12281;
													assign node12281 = (inp[4]) ? 4'b0101 : node12282;
														assign node12282 = (inp[7]) ? node12284 : 4'b1101;
															assign node12284 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node12288 = (inp[12]) ? node12292 : node12289;
														assign node12289 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node12292 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node12295 = (inp[12]) ? node12307 : node12296;
													assign node12296 = (inp[10]) ? node12302 : node12297;
														assign node12297 = (inp[7]) ? node12299 : 4'b0101;
															assign node12299 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node12302 = (inp[7]) ? node12304 : 4'b1101;
															assign node12304 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node12307 = (inp[7]) ? node12309 : 4'b0101;
														assign node12309 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node12312 = (inp[7]) ? node12352 : node12313;
											assign node12313 = (inp[11]) ? node12341 : node12314;
												assign node12314 = (inp[14]) ? node12328 : node12315;
													assign node12315 = (inp[13]) ? node12323 : node12316;
														assign node12316 = (inp[12]) ? node12318 : 4'b0100;
															assign node12318 = (inp[10]) ? 4'b0100 : node12319;
																assign node12319 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12323 = (inp[10]) ? 4'b1100 : node12324;
															assign node12324 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node12328 = (inp[13]) ? node12336 : node12329;
														assign node12329 = (inp[4]) ? node12331 : 4'b1001;
															assign node12331 = (inp[10]) ? node12333 : 4'b1101;
																assign node12333 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node12336 = (inp[12]) ? 4'b0101 : node12337;
															assign node12337 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node12341 = (inp[13]) ? node12347 : node12342;
													assign node12342 = (inp[10]) ? 4'b0100 : node12343;
														assign node12343 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node12347 = (inp[12]) ? node12349 : 4'b1100;
														assign node12349 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node12352 = (inp[4]) ? node12380 : node12353;
												assign node12353 = (inp[14]) ? node12365 : node12354;
													assign node12354 = (inp[13]) ? node12360 : node12355;
														assign node12355 = (inp[12]) ? node12357 : 4'b0000;
															assign node12357 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node12360 = (inp[12]) ? node12362 : 4'b1000;
															assign node12362 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12365 = (inp[11]) ? node12371 : node12366;
														assign node12366 = (inp[13]) ? 4'b0001 : node12367;
															assign node12367 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node12371 = (inp[12]) ? node12373 : 4'b1000;
															assign node12373 = (inp[10]) ? node12377 : node12374;
																assign node12374 = (inp[13]) ? 4'b0000 : 4'b1000;
																assign node12377 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node12380 = (inp[14]) ? node12392 : node12381;
													assign node12381 = (inp[10]) ? node12389 : node12382;
														assign node12382 = (inp[13]) ? node12386 : node12383;
															assign node12383 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node12386 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node12389 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node12392 = (inp[11]) ? node12398 : node12393;
														assign node12393 = (inp[13]) ? 4'b0101 : node12394;
															assign node12394 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node12398 = (inp[10]) ? 4'b1100 : node12399;
															assign node12399 = (inp[12]) ? node12401 : 4'b0100;
																assign node12401 = (inp[13]) ? 4'b0100 : 4'b1000;
					assign node12406 = (inp[5]) ? node13384 : node12407;
						assign node12407 = (inp[0]) ? node13097 : node12408;
							assign node12408 = (inp[11]) ? node12790 : node12409;
								assign node12409 = (inp[10]) ? node12589 : node12410;
									assign node12410 = (inp[1]) ? node12484 : node12411;
										assign node12411 = (inp[13]) ? node12443 : node12412;
											assign node12412 = (inp[4]) ? node12424 : node12413;
												assign node12413 = (inp[14]) ? node12419 : node12414;
													assign node12414 = (inp[3]) ? node12416 : 4'b1101;
														assign node12416 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node12419 = (inp[3]) ? node12421 : 4'b1100;
														assign node12421 = (inp[2]) ? 4'b1000 : 4'b1101;
												assign node12424 = (inp[7]) ? node12436 : node12425;
													assign node12425 = (inp[14]) ? node12431 : node12426;
														assign node12426 = (inp[3]) ? node12428 : 4'b1001;
															assign node12428 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12431 = (inp[2]) ? node12433 : 4'b1001;
															assign node12433 = (inp[3]) ? 4'b1001 : 4'b1000;
													assign node12436 = (inp[3]) ? node12440 : node12437;
														assign node12437 = (inp[12]) ? 4'b1100 : 4'b1101;
														assign node12440 = (inp[2]) ? 4'b1001 : 4'b0000;
											assign node12443 = (inp[2]) ? node12463 : node12444;
												assign node12444 = (inp[4]) ? node12450 : node12445;
													assign node12445 = (inp[7]) ? node12447 : 4'b1001;
														assign node12447 = (inp[3]) ? 4'b1101 : 4'b0100;
													assign node12450 = (inp[7]) ? node12458 : node12451;
														assign node12451 = (inp[3]) ? node12453 : 4'b1101;
															assign node12453 = (inp[14]) ? 4'b0101 : node12454;
																assign node12454 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node12458 = (inp[3]) ? node12460 : 4'b1001;
															assign node12460 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node12463 = (inp[3]) ? node12475 : node12464;
													assign node12464 = (inp[14]) ? node12470 : node12465;
														assign node12465 = (inp[4]) ? 4'b0001 : node12466;
															assign node12466 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12470 = (inp[4]) ? 4'b0000 : node12471;
															assign node12471 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node12475 = (inp[7]) ? node12479 : node12476;
														assign node12476 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node12479 = (inp[4]) ? 4'b1001 : node12480;
															assign node12480 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node12484 = (inp[12]) ? node12532 : node12485;
											assign node12485 = (inp[3]) ? node12509 : node12486;
												assign node12486 = (inp[14]) ? node12498 : node12487;
													assign node12487 = (inp[2]) ? node12491 : node12488;
														assign node12488 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node12491 = (inp[13]) ? node12495 : node12492;
															assign node12492 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node12495 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node12498 = (inp[13]) ? node12506 : node12499;
														assign node12499 = (inp[2]) ? 4'b1101 : node12500;
															assign node12500 = (inp[7]) ? 4'b0001 : node12501;
																assign node12501 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node12506 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node12509 = (inp[4]) ? node12519 : node12510;
													assign node12510 = (inp[13]) ? 4'b0001 : node12511;
														assign node12511 = (inp[2]) ? node12515 : node12512;
															assign node12512 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node12515 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node12519 = (inp[2]) ? node12527 : node12520;
														assign node12520 = (inp[13]) ? node12524 : node12521;
															assign node12521 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12524 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node12527 = (inp[7]) ? node12529 : 4'b0101;
															assign node12529 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node12532 = (inp[14]) ? node12560 : node12533;
												assign node12533 = (inp[2]) ? node12545 : node12534;
													assign node12534 = (inp[4]) ? node12540 : node12535;
														assign node12535 = (inp[13]) ? 4'b1001 : node12536;
															assign node12536 = (inp[3]) ? 4'b1101 : 4'b1100;
														assign node12540 = (inp[13]) ? 4'b1101 : node12541;
															assign node12541 = (inp[3]) ? 4'b0001 : 4'b1001;
													assign node12545 = (inp[13]) ? node12553 : node12546;
														assign node12546 = (inp[3]) ? 4'b1000 : node12547;
															assign node12547 = (inp[4]) ? node12549 : 4'b1100;
																assign node12549 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node12553 = (inp[7]) ? node12555 : 4'b1001;
															assign node12555 = (inp[4]) ? 4'b0000 : node12556;
																assign node12556 = (inp[3]) ? 4'b0000 : 4'b0100;
												assign node12560 = (inp[4]) ? node12576 : node12561;
													assign node12561 = (inp[13]) ? node12567 : node12562;
														assign node12562 = (inp[3]) ? node12564 : 4'b1101;
															assign node12564 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node12567 = (inp[3]) ? node12571 : node12568;
															assign node12568 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node12571 = (inp[7]) ? node12573 : 4'b1001;
																assign node12573 = (inp[2]) ? 4'b0001 : 4'b1101;
													assign node12576 = (inp[7]) ? node12582 : node12577;
														assign node12577 = (inp[2]) ? 4'b0001 : node12578;
															assign node12578 = (inp[3]) ? 4'b1100 : 4'b1101;
														assign node12582 = (inp[2]) ? 4'b1001 : node12583;
															assign node12583 = (inp[3]) ? node12585 : 4'b1001;
																assign node12585 = (inp[13]) ? 4'b1000 : 4'b0000;
									assign node12589 = (inp[1]) ? node12681 : node12590;
										assign node12590 = (inp[4]) ? node12638 : node12591;
											assign node12591 = (inp[3]) ? node12619 : node12592;
												assign node12592 = (inp[7]) ? node12604 : node12593;
													assign node12593 = (inp[2]) ? node12595 : 4'b0001;
														assign node12595 = (inp[14]) ? node12601 : node12596;
															assign node12596 = (inp[13]) ? node12598 : 4'b1101;
																assign node12598 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node12601 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node12604 = (inp[14]) ? node12612 : node12605;
														assign node12605 = (inp[12]) ? node12609 : node12606;
															assign node12606 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node12609 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node12612 = (inp[13]) ? node12616 : node12613;
															assign node12613 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node12616 = (inp[2]) ? 4'b0100 : 4'b0001;
												assign node12619 = (inp[13]) ? node12631 : node12620;
													assign node12620 = (inp[2]) ? node12624 : node12621;
														assign node12621 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12624 = (inp[7]) ? node12626 : 4'b0001;
															assign node12626 = (inp[14]) ? 4'b1000 : node12627;
																assign node12627 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12631 = (inp[2]) ? 4'b0001 : node12632;
														assign node12632 = (inp[14]) ? 4'b0001 : node12633;
															assign node12633 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node12638 = (inp[13]) ? node12664 : node12639;
												assign node12639 = (inp[7]) ? node12651 : node12640;
													assign node12640 = (inp[2]) ? node12646 : node12641;
														assign node12641 = (inp[3]) ? node12643 : 4'b0101;
															assign node12643 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node12646 = (inp[3]) ? 4'b0101 : node12647;
															assign node12647 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node12651 = (inp[14]) ? node12657 : node12652;
														assign node12652 = (inp[3]) ? node12654 : 4'b0001;
															assign node12654 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node12657 = (inp[2]) ? node12659 : 4'b0001;
															assign node12659 = (inp[12]) ? 4'b1100 : node12660;
																assign node12660 = (inp[3]) ? 4'b0001 : 4'b0000;
												assign node12664 = (inp[2]) ? node12672 : node12665;
													assign node12665 = (inp[3]) ? node12667 : 4'b0101;
														assign node12667 = (inp[14]) ? node12669 : 4'b0100;
															assign node12669 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node12672 = (inp[3]) ? 4'b0101 : node12673;
														assign node12673 = (inp[14]) ? node12677 : node12674;
															assign node12674 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node12677 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node12681 = (inp[12]) ? node12739 : node12682;
											assign node12682 = (inp[13]) ? node12716 : node12683;
												assign node12683 = (inp[2]) ? node12699 : node12684;
													assign node12684 = (inp[3]) ? node12690 : node12685;
														assign node12685 = (inp[4]) ? 4'b1001 : node12686;
															assign node12686 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node12690 = (inp[4]) ? node12694 : node12691;
															assign node12691 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node12694 = (inp[7]) ? 4'b0001 : node12695;
																assign node12695 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node12699 = (inp[3]) ? node12707 : node12700;
														assign node12700 = (inp[14]) ? node12704 : node12701;
															assign node12701 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node12704 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12707 = (inp[4]) ? node12713 : node12708;
															assign node12708 = (inp[7]) ? node12710 : 4'b1001;
																assign node12710 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node12713 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node12716 = (inp[4]) ? node12728 : node12717;
													assign node12717 = (inp[3]) ? 4'b1001 : node12718;
														assign node12718 = (inp[14]) ? node12724 : node12719;
															assign node12719 = (inp[2]) ? node12721 : 4'b1001;
																assign node12721 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node12724 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node12728 = (inp[2]) ? node12734 : node12729;
														assign node12729 = (inp[14]) ? node12731 : 4'b1101;
															assign node12731 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node12734 = (inp[3]) ? 4'b1101 : node12735;
															assign node12735 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node12739 = (inp[13]) ? node12773 : node12740;
												assign node12740 = (inp[14]) ? node12756 : node12741;
													assign node12741 = (inp[2]) ? node12749 : node12742;
														assign node12742 = (inp[3]) ? node12744 : 4'b0101;
															assign node12744 = (inp[4]) ? 4'b1001 : node12745;
																assign node12745 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12749 = (inp[3]) ? node12751 : 4'b0000;
															assign node12751 = (inp[7]) ? node12753 : 4'b0101;
																assign node12753 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node12756 = (inp[2]) ? node12766 : node12757;
														assign node12757 = (inp[3]) ? node12763 : node12758;
															assign node12758 = (inp[7]) ? 4'b0001 : node12759;
																assign node12759 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node12763 = (inp[4]) ? 4'b1000 : 4'b0101;
														assign node12766 = (inp[4]) ? node12770 : node12767;
															assign node12767 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node12770 = (inp[7]) ? 4'b0001 : 4'b1001;
												assign node12773 = (inp[4]) ? node12781 : node12774;
													assign node12774 = (inp[3]) ? 4'b0001 : node12775;
														assign node12775 = (inp[7]) ? node12777 : 4'b0001;
															assign node12777 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node12781 = (inp[2]) ? node12785 : node12782;
														assign node12782 = (inp[3]) ? 4'b0100 : 4'b0101;
														assign node12785 = (inp[3]) ? 4'b0101 : node12786;
															assign node12786 = (inp[14]) ? 4'b0001 : 4'b1000;
								assign node12790 = (inp[1]) ? node12984 : node12791;
									assign node12791 = (inp[3]) ? node12879 : node12792;
										assign node12792 = (inp[2]) ? node12846 : node12793;
											assign node12793 = (inp[4]) ? node12815 : node12794;
												assign node12794 = (inp[13]) ? node12808 : node12795;
													assign node12795 = (inp[7]) ? node12803 : node12796;
														assign node12796 = (inp[10]) ? node12800 : node12797;
															assign node12797 = (inp[12]) ? 4'b1101 : 4'b0000;
															assign node12800 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node12803 = (inp[12]) ? 4'b1101 : node12804;
															assign node12804 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node12808 = (inp[12]) ? node12812 : node12809;
														assign node12809 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12812 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node12815 = (inp[13]) ? node12835 : node12816;
													assign node12816 = (inp[7]) ? node12824 : node12817;
														assign node12817 = (inp[10]) ? node12821 : node12818;
															assign node12818 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node12821 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node12824 = (inp[14]) ? node12830 : node12825;
															assign node12825 = (inp[12]) ? 4'b1000 : node12826;
																assign node12826 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node12830 = (inp[12]) ? 4'b0000 : node12831;
																assign node12831 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node12835 = (inp[14]) ? node12841 : node12836;
														assign node12836 = (inp[10]) ? node12838 : 4'b1000;
															assign node12838 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node12841 = (inp[7]) ? 4'b0100 : node12842;
															assign node12842 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node12846 = (inp[13]) ? node12864 : node12847;
												assign node12847 = (inp[10]) ? node12853 : node12848;
													assign node12848 = (inp[7]) ? 4'b1101 : node12849;
														assign node12849 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node12853 = (inp[12]) ? node12859 : node12854;
														assign node12854 = (inp[4]) ? 4'b0001 : node12855;
															assign node12855 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12859 = (inp[7]) ? 4'b1101 : node12860;
															assign node12860 = (inp[14]) ? 4'b1001 : 4'b1101;
												assign node12864 = (inp[4]) ? node12874 : node12865;
													assign node12865 = (inp[7]) ? node12869 : node12866;
														assign node12866 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node12869 = (inp[10]) ? node12871 : 4'b0101;
															assign node12871 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node12874 = (inp[10]) ? node12876 : 4'b0001;
														assign node12876 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node12879 = (inp[4]) ? node12929 : node12880;
											assign node12880 = (inp[2]) ? node12910 : node12881;
												assign node12881 = (inp[13]) ? node12899 : node12882;
													assign node12882 = (inp[7]) ? node12890 : node12883;
														assign node12883 = (inp[12]) ? node12887 : node12884;
															assign node12884 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node12887 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node12890 = (inp[14]) ? 4'b1100 : node12891;
															assign node12891 = (inp[12]) ? node12895 : node12892;
																assign node12892 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node12895 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node12899 = (inp[7]) ? node12903 : node12900;
														assign node12900 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node12903 = (inp[10]) ? node12907 : node12904;
															assign node12904 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node12907 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node12910 = (inp[13]) ? node12920 : node12911;
													assign node12911 = (inp[7]) ? node12917 : node12912;
														assign node12912 = (inp[12]) ? 4'b1001 : node12913;
															assign node12913 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12917 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node12920 = (inp[10]) ? node12926 : node12921;
														assign node12921 = (inp[12]) ? node12923 : 4'b0000;
															assign node12923 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node12926 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node12929 = (inp[2]) ? node12949 : node12930;
												assign node12930 = (inp[13]) ? node12940 : node12931;
													assign node12931 = (inp[7]) ? node12937 : node12932;
														assign node12932 = (inp[10]) ? 4'b1001 : node12933;
															assign node12933 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node12937 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node12940 = (inp[10]) ? 4'b0101 : node12941;
														assign node12941 = (inp[12]) ? node12945 : node12942;
															assign node12942 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node12945 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node12949 = (inp[7]) ? node12969 : node12950;
													assign node12950 = (inp[13]) ? node12958 : node12951;
														assign node12951 = (inp[12]) ? node12955 : node12952;
															assign node12952 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node12955 = (inp[14]) ? 4'b1000 : 4'b0100;
														assign node12958 = (inp[14]) ? node12964 : node12959;
															assign node12959 = (inp[12]) ? 4'b0100 : node12960;
																assign node12960 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node12964 = (inp[12]) ? node12966 : 4'b0100;
																assign node12966 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node12969 = (inp[13]) ? node12977 : node12970;
														assign node12970 = (inp[14]) ? node12972 : 4'b0000;
															assign node12972 = (inp[12]) ? 4'b0000 : node12973;
																assign node12973 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node12977 = (inp[10]) ? node12981 : node12978;
															assign node12978 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node12981 = (inp[12]) ? 4'b0100 : 4'b1100;
									assign node12984 = (inp[10]) ? node13054 : node12985;
										assign node12985 = (inp[4]) ? node13019 : node12986;
											assign node12986 = (inp[3]) ? node13006 : node12987;
												assign node12987 = (inp[13]) ? node12997 : node12988;
													assign node12988 = (inp[12]) ? node12992 : node12989;
														assign node12989 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node12992 = (inp[2]) ? 4'b1100 : node12993;
															assign node12993 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node12997 = (inp[2]) ? node12999 : 4'b0000;
														assign node12999 = (inp[12]) ? node13003 : node13000;
															assign node13000 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node13003 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node13006 = (inp[2]) ? node13012 : node13007;
													assign node13007 = (inp[7]) ? node13009 : 4'b0000;
														assign node13009 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node13012 = (inp[12]) ? node13014 : 4'b0000;
														assign node13014 = (inp[7]) ? node13016 : 4'b0000;
															assign node13016 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node13019 = (inp[13]) ? node13041 : node13020;
												assign node13020 = (inp[7]) ? node13030 : node13021;
													assign node13021 = (inp[3]) ? node13025 : node13022;
														assign node13022 = (inp[2]) ? 4'b1000 : 4'b0100;
														assign node13025 = (inp[2]) ? 4'b0100 : node13026;
															assign node13026 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13030 = (inp[2]) ? node13036 : node13031;
														assign node13031 = (inp[3]) ? node13033 : 4'b0000;
															assign node13033 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13036 = (inp[12]) ? node13038 : 4'b0000;
															assign node13038 = (inp[3]) ? 4'b0000 : 4'b1100;
												assign node13041 = (inp[3]) ? node13047 : node13042;
													assign node13042 = (inp[2]) ? node13044 : 4'b0100;
														assign node13044 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13047 = (inp[12]) ? node13049 : 4'b0100;
														assign node13049 = (inp[2]) ? 4'b0100 : node13050;
															assign node13050 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node13054 = (inp[13]) ? node13084 : node13055;
											assign node13055 = (inp[2]) ? node13071 : node13056;
												assign node13056 = (inp[3]) ? node13064 : node13057;
													assign node13057 = (inp[7]) ? node13061 : node13058;
														assign node13058 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node13061 = (inp[14]) ? 4'b0100 : 4'b1000;
													assign node13064 = (inp[4]) ? node13068 : node13065;
														assign node13065 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node13068 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node13071 = (inp[3]) ? node13077 : node13072;
													assign node13072 = (inp[4]) ? 4'b0000 : node13073;
														assign node13073 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node13077 = (inp[4]) ? node13081 : node13078;
														assign node13078 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node13081 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node13084 = (inp[4]) ? node13092 : node13085;
												assign node13085 = (inp[3]) ? 4'b1000 : node13086;
													assign node13086 = (inp[7]) ? node13088 : 4'b1000;
														assign node13088 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node13092 = (inp[2]) ? node13094 : 4'b1100;
													assign node13094 = (inp[3]) ? 4'b1100 : 4'b1000;
							assign node13097 = (inp[2]) ? 4'b1100 : node13098;
								assign node13098 = (inp[1]) ? node13228 : node13099;
									assign node13099 = (inp[13]) ? node13167 : node13100;
										assign node13100 = (inp[12]) ? node13140 : node13101;
											assign node13101 = (inp[10]) ? node13119 : node13102;
												assign node13102 = (inp[3]) ? node13108 : node13103;
													assign node13103 = (inp[11]) ? 4'b1100 : node13104;
														assign node13104 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node13108 = (inp[4]) ? node13114 : node13109;
														assign node13109 = (inp[14]) ? node13111 : 4'b1001;
															assign node13111 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13114 = (inp[7]) ? 4'b1001 : node13115;
															assign node13115 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node13119 = (inp[3]) ? node13129 : node13120;
													assign node13120 = (inp[7]) ? node13126 : node13121;
														assign node13121 = (inp[14]) ? node13123 : 4'b0001;
															assign node13123 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node13126 = (inp[4]) ? 4'b0001 : 4'b1100;
													assign node13129 = (inp[14]) ? node13135 : node13130;
														assign node13130 = (inp[7]) ? node13132 : 4'b0101;
															assign node13132 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node13135 = (inp[11]) ? 4'b0101 : node13136;
															assign node13136 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node13140 = (inp[3]) ? node13150 : node13141;
												assign node13141 = (inp[4]) ? node13143 : 4'b1100;
													assign node13143 = (inp[7]) ? 4'b1100 : node13144;
														assign node13144 = (inp[11]) ? 4'b1001 : node13145;
															assign node13145 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node13150 = (inp[11]) ? node13162 : node13151;
													assign node13151 = (inp[14]) ? node13157 : node13152;
														assign node13152 = (inp[4]) ? node13154 : 4'b1001;
															assign node13154 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node13157 = (inp[4]) ? node13159 : 4'b1000;
															assign node13159 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node13162 = (inp[4]) ? node13164 : 4'b1001;
														assign node13164 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node13167 = (inp[3]) ? node13199 : node13168;
											assign node13168 = (inp[7]) ? node13184 : node13169;
												assign node13169 = (inp[14]) ? node13175 : node13170;
													assign node13170 = (inp[10]) ? node13172 : 4'b0001;
														assign node13172 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13175 = (inp[11]) ? node13181 : node13176;
														assign node13176 = (inp[12]) ? 4'b0000 : node13177;
															assign node13177 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13181 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node13184 = (inp[4]) ? node13186 : 4'b1100;
													assign node13186 = (inp[11]) ? node13194 : node13187;
														assign node13187 = (inp[14]) ? node13189 : 4'b1001;
															assign node13189 = (inp[10]) ? node13191 : 4'b0000;
																assign node13191 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13194 = (inp[10]) ? node13196 : 4'b0001;
															assign node13196 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node13199 = (inp[7]) ? node13213 : node13200;
												assign node13200 = (inp[14]) ? node13206 : node13201;
													assign node13201 = (inp[10]) ? node13203 : 4'b0101;
														assign node13203 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node13206 = (inp[11]) ? 4'b0101 : node13207;
														assign node13207 = (inp[12]) ? 4'b0100 : node13208;
															assign node13208 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node13213 = (inp[4]) ? node13223 : node13214;
													assign node13214 = (inp[10]) ? node13216 : 4'b0001;
														assign node13216 = (inp[12]) ? node13220 : node13217;
															assign node13217 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node13220 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node13223 = (inp[11]) ? 4'b0101 : node13224;
														assign node13224 = (inp[12]) ? 4'b0101 : 4'b0100;
									assign node13228 = (inp[3]) ? node13294 : node13229;
										assign node13229 = (inp[7]) ? node13265 : node13230;
											assign node13230 = (inp[13]) ? node13246 : node13231;
												assign node13231 = (inp[10]) ? node13241 : node13232;
													assign node13232 = (inp[12]) ? node13238 : node13233;
														assign node13233 = (inp[11]) ? 4'b0000 : node13234;
															assign node13234 = (inp[14]) ? 4'b1100 : 4'b0000;
														assign node13238 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node13241 = (inp[11]) ? 4'b0000 : node13242;
														assign node13242 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node13246 = (inp[11]) ? node13260 : node13247;
													assign node13247 = (inp[14]) ? node13255 : node13248;
														assign node13248 = (inp[4]) ? node13250 : 4'b1000;
															assign node13250 = (inp[12]) ? node13252 : 4'b1000;
																assign node13252 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13255 = (inp[10]) ? node13257 : 4'b0001;
															assign node13257 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13260 = (inp[10]) ? 4'b1000 : node13261;
														assign node13261 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node13265 = (inp[4]) ? node13267 : 4'b1100;
												assign node13267 = (inp[13]) ? node13281 : node13268;
													assign node13268 = (inp[12]) ? node13276 : node13269;
														assign node13269 = (inp[14]) ? node13271 : 4'b0000;
															assign node13271 = (inp[10]) ? 4'b0001 : node13272;
																assign node13272 = (inp[11]) ? 4'b0000 : 4'b1100;
														assign node13276 = (inp[10]) ? node13278 : 4'b1100;
															assign node13278 = (inp[14]) ? 4'b1100 : 4'b0000;
													assign node13281 = (inp[10]) ? node13289 : node13282;
														assign node13282 = (inp[14]) ? node13286 : node13283;
															assign node13283 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13286 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node13289 = (inp[11]) ? 4'b1000 : node13290;
															assign node13290 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node13294 = (inp[4]) ? node13346 : node13295;
											assign node13295 = (inp[7]) ? node13323 : node13296;
												assign node13296 = (inp[11]) ? node13312 : node13297;
													assign node13297 = (inp[14]) ? node13305 : node13298;
														assign node13298 = (inp[13]) ? node13300 : 4'b1000;
															assign node13300 = (inp[10]) ? 4'b1100 : node13301;
																assign node13301 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node13305 = (inp[13]) ? node13309 : node13306;
															assign node13306 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node13309 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node13312 = (inp[13]) ? node13318 : node13313;
														assign node13313 = (inp[10]) ? 4'b0100 : node13314;
															assign node13314 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node13318 = (inp[12]) ? node13320 : 4'b1100;
															assign node13320 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node13323 = (inp[11]) ? node13335 : node13324;
													assign node13324 = (inp[14]) ? node13328 : node13325;
														assign node13325 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node13328 = (inp[12]) ? 4'b0001 : node13329;
															assign node13329 = (inp[13]) ? node13331 : 4'b1001;
																assign node13331 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node13335 = (inp[13]) ? node13341 : node13336;
														assign node13336 = (inp[12]) ? node13338 : 4'b0000;
															assign node13338 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node13341 = (inp[12]) ? node13343 : 4'b1000;
															assign node13343 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node13346 = (inp[11]) ? node13372 : node13347;
												assign node13347 = (inp[14]) ? node13359 : node13348;
													assign node13348 = (inp[13]) ? node13354 : node13349;
														assign node13349 = (inp[10]) ? 4'b0100 : node13350;
															assign node13350 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node13354 = (inp[10]) ? 4'b1100 : node13355;
															assign node13355 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node13359 = (inp[12]) ? node13369 : node13360;
														assign node13360 = (inp[10]) ? node13366 : node13361;
															assign node13361 = (inp[7]) ? 4'b1001 : node13362;
																assign node13362 = (inp[13]) ? 4'b0101 : 4'b1101;
															assign node13366 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node13369 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node13372 = (inp[13]) ? node13378 : node13373;
													assign node13373 = (inp[12]) ? node13375 : 4'b0100;
														assign node13375 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node13378 = (inp[10]) ? 4'b1100 : node13379;
														assign node13379 = (inp[12]) ? 4'b0100 : 4'b1100;
						assign node13384 = (inp[3]) ? node14044 : node13385;
							assign node13385 = (inp[4]) ? node13721 : node13386;
								assign node13386 = (inp[7]) ? node13562 : node13387;
									assign node13387 = (inp[1]) ? node13471 : node13388;
										assign node13388 = (inp[2]) ? node13426 : node13389;
											assign node13389 = (inp[0]) ? node13407 : node13390;
												assign node13390 = (inp[13]) ? node13396 : node13391;
													assign node13391 = (inp[12]) ? node13393 : 4'b0000;
														assign node13393 = (inp[11]) ? 4'b0000 : 4'b1100;
													assign node13396 = (inp[12]) ? node13402 : node13397;
														assign node13397 = (inp[11]) ? node13399 : 4'b0100;
															assign node13399 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node13402 = (inp[11]) ? 4'b0100 : node13403;
															assign node13403 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node13407 = (inp[11]) ? node13415 : node13408;
													assign node13408 = (inp[10]) ? 4'b0001 : node13409;
														assign node13409 = (inp[13]) ? 4'b1001 : node13410;
															assign node13410 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node13415 = (inp[13]) ? node13421 : node13416;
														assign node13416 = (inp[12]) ? 4'b1101 : node13417;
															assign node13417 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13421 = (inp[12]) ? node13423 : 4'b1000;
															assign node13423 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node13426 = (inp[13]) ? node13444 : node13427;
												assign node13427 = (inp[12]) ? node13435 : node13428;
													assign node13428 = (inp[11]) ? 4'b0001 : node13429;
														assign node13429 = (inp[10]) ? node13431 : 4'b1100;
															assign node13431 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node13435 = (inp[0]) ? 4'b1100 : node13436;
														assign node13436 = (inp[10]) ? node13440 : node13437;
															assign node13437 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node13440 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node13444 = (inp[11]) ? node13464 : node13445;
													assign node13445 = (inp[10]) ? node13455 : node13446;
														assign node13446 = (inp[12]) ? 4'b0000 : node13447;
															assign node13447 = (inp[14]) ? node13451 : node13448;
																assign node13448 = (inp[0]) ? 4'b0001 : 4'b1000;
																assign node13451 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node13455 = (inp[0]) ? node13461 : node13456;
															assign node13456 = (inp[14]) ? node13458 : 4'b0100;
																assign node13458 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node13461 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13464 = (inp[12]) ? node13466 : 4'b1001;
														assign node13466 = (inp[10]) ? node13468 : 4'b0001;
															assign node13468 = (inp[0]) ? 4'b0001 : 4'b0101;
										assign node13471 = (inp[11]) ? node13529 : node13472;
											assign node13472 = (inp[13]) ? node13498 : node13473;
												assign node13473 = (inp[0]) ? node13485 : node13474;
													assign node13474 = (inp[10]) ? node13480 : node13475;
														assign node13475 = (inp[14]) ? 4'b0000 : node13476;
															assign node13476 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node13480 = (inp[12]) ? node13482 : 4'b1000;
															assign node13482 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node13485 = (inp[12]) ? node13493 : node13486;
														assign node13486 = (inp[2]) ? node13488 : 4'b0001;
															assign node13488 = (inp[10]) ? node13490 : 4'b1100;
																assign node13490 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node13493 = (inp[10]) ? node13495 : 4'b1100;
															assign node13495 = (inp[14]) ? 4'b1100 : 4'b0000;
												assign node13498 = (inp[12]) ? node13516 : node13499;
													assign node13499 = (inp[2]) ? node13507 : node13500;
														assign node13500 = (inp[14]) ? 4'b0001 : node13501;
															assign node13501 = (inp[10]) ? node13503 : 4'b1100;
																assign node13503 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node13507 = (inp[10]) ? node13513 : node13508;
															assign node13508 = (inp[0]) ? 4'b1000 : node13509;
																assign node13509 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node13513 = (inp[0]) ? 4'b1000 : 4'b1100;
													assign node13516 = (inp[10]) ? node13522 : node13517;
														assign node13517 = (inp[0]) ? node13519 : 4'b1001;
															assign node13519 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node13522 = (inp[2]) ? node13524 : 4'b0001;
															assign node13524 = (inp[0]) ? 4'b1000 : node13525;
																assign node13525 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node13529 = (inp[0]) ? node13547 : node13530;
												assign node13530 = (inp[13]) ? node13538 : node13531;
													assign node13531 = (inp[2]) ? node13533 : 4'b1000;
														assign node13533 = (inp[12]) ? 4'b0000 : node13534;
															assign node13534 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node13538 = (inp[2]) ? node13542 : node13539;
														assign node13539 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node13542 = (inp[10]) ? 4'b1100 : node13543;
															assign node13543 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node13547 = (inp[10]) ? node13557 : node13548;
													assign node13548 = (inp[2]) ? node13550 : 4'b0000;
														assign node13550 = (inp[13]) ? node13554 : node13551;
															assign node13551 = (inp[14]) ? 4'b0000 : 4'b1100;
															assign node13554 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13557 = (inp[13]) ? 4'b1000 : node13558;
														assign node13558 = (inp[2]) ? 4'b0000 : 4'b1000;
									assign node13562 = (inp[13]) ? node13646 : node13563;
										assign node13563 = (inp[0]) ? node13617 : node13564;
											assign node13564 = (inp[10]) ? node13594 : node13565;
												assign node13565 = (inp[11]) ? node13581 : node13566;
													assign node13566 = (inp[2]) ? node13576 : node13567;
														assign node13567 = (inp[1]) ? node13573 : node13568;
															assign node13568 = (inp[12]) ? node13570 : 4'b0100;
																assign node13570 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node13573 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node13576 = (inp[1]) ? node13578 : 4'b1101;
															assign node13578 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node13581 = (inp[2]) ? node13589 : node13582;
														assign node13582 = (inp[1]) ? node13586 : node13583;
															assign node13583 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node13586 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node13589 = (inp[12]) ? node13591 : 4'b0100;
															assign node13591 = (inp[1]) ? 4'b0100 : 4'b1100;
												assign node13594 = (inp[2]) ? node13606 : node13595;
													assign node13595 = (inp[1]) ? node13601 : node13596;
														assign node13596 = (inp[11]) ? 4'b0000 : node13597;
															assign node13597 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node13601 = (inp[11]) ? 4'b1000 : node13602;
															assign node13602 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13606 = (inp[11]) ? node13612 : node13607;
														assign node13607 = (inp[12]) ? 4'b0101 : node13608;
															assign node13608 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node13612 = (inp[1]) ? 4'b0000 : node13613;
															assign node13613 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node13617 = (inp[2]) ? 4'b1100 : node13618;
												assign node13618 = (inp[12]) ? node13634 : node13619;
													assign node13619 = (inp[10]) ? node13627 : node13620;
														assign node13620 = (inp[1]) ? node13624 : node13621;
															assign node13621 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node13624 = (inp[11]) ? 4'b0100 : 4'b1101;
														assign node13627 = (inp[14]) ? node13629 : 4'b0100;
															assign node13629 = (inp[11]) ? 4'b0100 : node13630;
																assign node13630 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node13634 = (inp[1]) ? node13640 : node13635;
														assign node13635 = (inp[11]) ? 4'b1101 : node13636;
															assign node13636 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13640 = (inp[14]) ? 4'b1101 : node13641;
															assign node13641 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node13646 = (inp[0]) ? node13694 : node13647;
											assign node13647 = (inp[2]) ? node13669 : node13648;
												assign node13648 = (inp[10]) ? node13658 : node13649;
													assign node13649 = (inp[1]) ? node13651 : 4'b0000;
														assign node13651 = (inp[14]) ? node13653 : 4'b1000;
															assign node13653 = (inp[11]) ? 4'b1000 : node13654;
																assign node13654 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13658 = (inp[1]) ? node13664 : node13659;
														assign node13659 = (inp[12]) ? node13661 : 4'b0100;
															assign node13661 = (inp[11]) ? 4'b0100 : 4'b1000;
														assign node13664 = (inp[14]) ? node13666 : 4'b1100;
															assign node13666 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node13669 = (inp[1]) ? node13681 : node13670;
													assign node13670 = (inp[11]) ? node13676 : node13671;
														assign node13671 = (inp[14]) ? node13673 : 4'b0000;
															assign node13673 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13676 = (inp[10]) ? 4'b0001 : node13677;
															assign node13677 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13681 = (inp[11]) ? node13689 : node13682;
														assign node13682 = (inp[14]) ? node13686 : node13683;
															assign node13683 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node13686 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node13689 = (inp[10]) ? 4'b1000 : node13690;
															assign node13690 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node13694 = (inp[2]) ? 4'b1100 : node13695;
												assign node13695 = (inp[11]) ? node13711 : node13696;
													assign node13696 = (inp[10]) ? node13706 : node13697;
														assign node13697 = (inp[12]) ? node13703 : node13698;
															assign node13698 = (inp[1]) ? 4'b0001 : node13699;
																assign node13699 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node13703 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node13706 = (inp[1]) ? node13708 : 4'b0001;
															assign node13708 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node13711 = (inp[10]) ? node13715 : node13712;
														assign node13712 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node13715 = (inp[1]) ? 4'b1000 : node13716;
															assign node13716 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node13721 = (inp[1]) ? node13901 : node13722;
									assign node13722 = (inp[2]) ? node13820 : node13723;
										assign node13723 = (inp[11]) ? node13769 : node13724;
											assign node13724 = (inp[10]) ? node13742 : node13725;
												assign node13725 = (inp[0]) ? node13737 : node13726;
													assign node13726 = (inp[14]) ? node13732 : node13727;
														assign node13727 = (inp[12]) ? node13729 : 4'b0001;
															assign node13729 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node13732 = (inp[12]) ? 4'b0100 : node13733;
															assign node13733 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node13737 = (inp[13]) ? node13739 : 4'b1001;
														assign node13739 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node13742 = (inp[13]) ? node13754 : node13743;
													assign node13743 = (inp[7]) ? node13749 : node13744;
														assign node13744 = (inp[14]) ? node13746 : 4'b0101;
															assign node13746 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node13749 = (inp[0]) ? 4'b0001 : node13750;
															assign node13750 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node13754 = (inp[14]) ? node13762 : node13755;
														assign node13755 = (inp[0]) ? 4'b0000 : node13756;
															assign node13756 = (inp[7]) ? 4'b1001 : node13757;
																assign node13757 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13762 = (inp[12]) ? node13766 : node13763;
															assign node13763 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node13766 = (inp[0]) ? 4'b0101 : 4'b0001;
											assign node13769 = (inp[7]) ? node13793 : node13770;
												assign node13770 = (inp[13]) ? node13782 : node13771;
													assign node13771 = (inp[0]) ? node13775 : node13772;
														assign node13772 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node13775 = (inp[10]) ? node13779 : node13776;
															assign node13776 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node13779 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node13782 = (inp[0]) ? node13788 : node13783;
														assign node13783 = (inp[10]) ? 4'b1001 : node13784;
															assign node13784 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13788 = (inp[10]) ? 4'b0001 : node13789;
															assign node13789 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node13793 = (inp[13]) ? node13809 : node13794;
													assign node13794 = (inp[0]) ? node13800 : node13795;
														assign node13795 = (inp[12]) ? 4'b0001 : node13796;
															assign node13796 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13800 = (inp[14]) ? 4'b0000 : node13801;
															assign node13801 = (inp[12]) ? node13805 : node13802;
																assign node13802 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node13805 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node13809 = (inp[0]) ? node13817 : node13810;
														assign node13810 = (inp[12]) ? node13814 : node13811;
															assign node13811 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node13814 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13817 = (inp[10]) ? 4'b0001 : 4'b1000;
										assign node13820 = (inp[0]) ? node13868 : node13821;
											assign node13821 = (inp[12]) ? node13839 : node13822;
												assign node13822 = (inp[10]) ? node13830 : node13823;
													assign node13823 = (inp[7]) ? node13827 : node13824;
														assign node13824 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node13827 = (inp[13]) ? 4'b0000 : 4'b0101;
													assign node13830 = (inp[7]) ? node13836 : node13831;
														assign node13831 = (inp[11]) ? 4'b0001 : node13832;
															assign node13832 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node13836 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node13839 = (inp[11]) ? node13857 : node13840;
													assign node13840 = (inp[13]) ? 4'b1000 : node13841;
														assign node13841 = (inp[14]) ? node13849 : node13842;
															assign node13842 = (inp[7]) ? node13846 : node13843;
																assign node13843 = (inp[10]) ? 4'b1000 : 4'b1100;
																assign node13846 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node13849 = (inp[10]) ? node13853 : node13850;
																assign node13850 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node13853 = (inp[7]) ? 4'b0101 : 4'b1000;
													assign node13857 = (inp[13]) ? node13863 : node13858;
														assign node13858 = (inp[7]) ? node13860 : 4'b0000;
															assign node13860 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node13863 = (inp[10]) ? 4'b1001 : node13864;
															assign node13864 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node13868 = (inp[13]) ? node13886 : node13869;
												assign node13869 = (inp[7]) ? node13881 : node13870;
													assign node13870 = (inp[10]) ? node13876 : node13871;
														assign node13871 = (inp[11]) ? 4'b1001 : node13872;
															assign node13872 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node13876 = (inp[12]) ? 4'b1001 : node13877;
															assign node13877 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node13881 = (inp[10]) ? node13883 : 4'b1100;
														assign node13883 = (inp[12]) ? 4'b1100 : 4'b0001;
												assign node13886 = (inp[10]) ? node13892 : node13887;
													assign node13887 = (inp[14]) ? node13889 : 4'b0001;
														assign node13889 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node13892 = (inp[12]) ? node13898 : node13893;
														assign node13893 = (inp[11]) ? 4'b1001 : node13894;
															assign node13894 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node13898 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node13901 = (inp[11]) ? node14001 : node13902;
										assign node13902 = (inp[2]) ? node13948 : node13903;
											assign node13903 = (inp[10]) ? node13927 : node13904;
												assign node13904 = (inp[13]) ? node13920 : node13905;
													assign node13905 = (inp[14]) ? node13911 : node13906;
														assign node13906 = (inp[0]) ? node13908 : 4'b1000;
															assign node13908 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node13911 = (inp[12]) ? node13917 : node13912;
															assign node13912 = (inp[7]) ? node13914 : 4'b0101;
																assign node13914 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node13917 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node13920 = (inp[0]) ? node13922 : 4'b1001;
														assign node13922 = (inp[12]) ? 4'b1001 : node13923;
															assign node13923 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node13927 = (inp[13]) ? node13939 : node13928;
													assign node13928 = (inp[7]) ? node13932 : node13929;
														assign node13929 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node13932 = (inp[14]) ? 4'b1001 : node13933;
															assign node13933 = (inp[0]) ? 4'b1001 : node13934;
																assign node13934 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node13939 = (inp[14]) ? node13943 : node13940;
														assign node13940 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node13943 = (inp[0]) ? node13945 : 4'b0000;
															assign node13945 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node13948 = (inp[14]) ? node13974 : node13949;
												assign node13949 = (inp[12]) ? node13959 : node13950;
													assign node13950 = (inp[13]) ? 4'b1000 : node13951;
														assign node13951 = (inp[0]) ? 4'b0000 : node13952;
															assign node13952 = (inp[7]) ? node13954 : 4'b1000;
																assign node13954 = (inp[10]) ? 4'b1000 : 4'b0101;
													assign node13959 = (inp[0]) ? node13967 : node13960;
														assign node13960 = (inp[10]) ? 4'b0000 : node13961;
															assign node13961 = (inp[7]) ? node13963 : 4'b0000;
																assign node13963 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node13967 = (inp[13]) ? node13971 : node13968;
															assign node13968 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node13971 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node13974 = (inp[13]) ? node13986 : node13975;
													assign node13975 = (inp[7]) ? node13983 : node13976;
														assign node13976 = (inp[0]) ? node13980 : node13977;
															assign node13977 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13980 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13983 = (inp[0]) ? 4'b1100 : 4'b0100;
													assign node13986 = (inp[0]) ? node13996 : node13987;
														assign node13987 = (inp[7]) ? node13993 : node13988;
															assign node13988 = (inp[10]) ? 4'b0001 : node13989;
																assign node13989 = (inp[12]) ? 4'b0100 : 4'b0001;
															assign node13993 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13996 = (inp[10]) ? node13998 : 4'b0001;
															assign node13998 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node14001 = (inp[10]) ? node14031 : node14002;
											assign node14002 = (inp[2]) ? node14010 : node14003;
												assign node14003 = (inp[7]) ? 4'b0000 : node14004;
													assign node14004 = (inp[13]) ? node14006 : 4'b0100;
														assign node14006 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node14010 = (inp[13]) ? node14024 : node14011;
													assign node14011 = (inp[7]) ? node14017 : node14012;
														assign node14012 = (inp[12]) ? 4'b1000 : node14013;
															assign node14013 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node14017 = (inp[0]) ? node14021 : node14018;
															assign node14018 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node14021 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node14024 = (inp[12]) ? node14026 : 4'b1000;
														assign node14026 = (inp[7]) ? node14028 : 4'b0000;
															assign node14028 = (inp[0]) ? 4'b0000 : 4'b1000;
											assign node14031 = (inp[13]) ? 4'b1000 : node14032;
												assign node14032 = (inp[0]) ? node14038 : node14033;
													assign node14033 = (inp[2]) ? 4'b1000 : node14034;
														assign node14034 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node14038 = (inp[2]) ? 4'b0000 : node14039;
														assign node14039 = (inp[7]) ? 4'b1000 : 4'b0000;
							assign node14044 = (inp[4]) ? node14448 : node14045;
								assign node14045 = (inp[11]) ? node14265 : node14046;
									assign node14046 = (inp[2]) ? node14150 : node14047;
										assign node14047 = (inp[13]) ? node14099 : node14048;
											assign node14048 = (inp[10]) ? node14062 : node14049;
												assign node14049 = (inp[0]) ? node14051 : 4'b0000;
													assign node14051 = (inp[1]) ? node14057 : node14052;
														assign node14052 = (inp[12]) ? node14054 : 4'b0000;
															assign node14054 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node14057 = (inp[12]) ? 4'b0000 : node14058;
															assign node14058 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node14062 = (inp[0]) ? node14084 : node14063;
													assign node14063 = (inp[12]) ? node14075 : node14064;
														assign node14064 = (inp[1]) ? node14070 : node14065;
															assign node14065 = (inp[7]) ? 4'b0000 : node14066;
																assign node14066 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14070 = (inp[7]) ? node14072 : 4'b0001;
																assign node14072 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node14075 = (inp[14]) ? node14081 : node14076;
															assign node14076 = (inp[1]) ? 4'b1000 : node14077;
																assign node14077 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node14081 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node14084 = (inp[7]) ? node14092 : node14085;
														assign node14085 = (inp[14]) ? node14087 : 4'b0000;
															assign node14087 = (inp[1]) ? node14089 : 4'b0000;
																assign node14089 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14092 = (inp[14]) ? 4'b0000 : node14093;
															assign node14093 = (inp[12]) ? node14095 : 4'b1000;
																assign node14095 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node14099 = (inp[10]) ? node14131 : node14100;
												assign node14100 = (inp[0]) ? node14114 : node14101;
													assign node14101 = (inp[1]) ? node14109 : node14102;
														assign node14102 = (inp[7]) ? 4'b0001 : node14103;
															assign node14103 = (inp[12]) ? 4'b0001 : node14104;
																assign node14104 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node14109 = (inp[14]) ? 4'b0000 : node14110;
															assign node14110 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node14114 = (inp[1]) ? node14126 : node14115;
														assign node14115 = (inp[14]) ? node14121 : node14116;
															assign node14116 = (inp[7]) ? 4'b1000 : node14117;
																assign node14117 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node14121 = (inp[12]) ? 4'b1000 : node14122;
																assign node14122 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node14126 = (inp[12]) ? 4'b0000 : node14127;
															assign node14127 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node14131 = (inp[0]) ? node14143 : node14132;
													assign node14132 = (inp[1]) ? node14138 : node14133;
														assign node14133 = (inp[14]) ? node14135 : 4'b0001;
															assign node14135 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14138 = (inp[14]) ? 4'b1001 : node14139;
															assign node14139 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node14143 = (inp[1]) ? node14145 : 4'b1001;
														assign node14145 = (inp[7]) ? 4'b0001 : node14146;
															assign node14146 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node14150 = (inp[13]) ? node14212 : node14151;
											assign node14151 = (inp[10]) ? node14183 : node14152;
												assign node14152 = (inp[12]) ? node14174 : node14153;
													assign node14153 = (inp[7]) ? node14163 : node14154;
														assign node14154 = (inp[0]) ? node14158 : node14155;
															assign node14155 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node14158 = (inp[1]) ? 4'b0001 : node14159;
																assign node14159 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node14163 = (inp[14]) ? node14171 : node14164;
															assign node14164 = (inp[1]) ? node14168 : node14165;
																assign node14165 = (inp[0]) ? 4'b1001 : 4'b0001;
																assign node14168 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node14171 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node14174 = (inp[14]) ? node14180 : node14175;
														assign node14175 = (inp[1]) ? node14177 : 4'b1001;
															assign node14177 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14180 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node14183 = (inp[0]) ? node14193 : node14184;
													assign node14184 = (inp[7]) ? node14188 : node14185;
														assign node14185 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node14188 = (inp[1]) ? 4'b0001 : node14189;
															assign node14189 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14193 = (inp[7]) ? node14199 : node14194;
														assign node14194 = (inp[12]) ? 4'b0001 : node14195;
															assign node14195 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node14199 = (inp[12]) ? node14205 : node14200;
															assign node14200 = (inp[1]) ? node14202 : 4'b0000;
																assign node14202 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node14205 = (inp[14]) ? node14209 : node14206;
																assign node14206 = (inp[1]) ? 4'b0000 : 4'b1001;
																assign node14209 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node14212 = (inp[0]) ? node14240 : node14213;
												assign node14213 = (inp[10]) ? node14225 : node14214;
													assign node14214 = (inp[14]) ? node14220 : node14215;
														assign node14215 = (inp[7]) ? node14217 : 4'b0000;
															assign node14217 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node14220 = (inp[7]) ? node14222 : 4'b0000;
															assign node14222 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node14225 = (inp[7]) ? node14233 : node14226;
														assign node14226 = (inp[12]) ? node14228 : 4'b0000;
															assign node14228 = (inp[14]) ? node14230 : 4'b1001;
																assign node14230 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node14233 = (inp[12]) ? 4'b0000 : node14234;
															assign node14234 = (inp[1]) ? 4'b0001 : node14235;
																assign node14235 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node14240 = (inp[7]) ? node14254 : node14241;
													assign node14241 = (inp[10]) ? node14245 : node14242;
														assign node14242 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14245 = (inp[12]) ? node14249 : node14246;
															assign node14246 = (inp[1]) ? 4'b1000 : 4'b0001;
															assign node14249 = (inp[14]) ? 4'b0001 : node14250;
																assign node14250 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node14254 = (inp[10]) ? node14260 : node14255;
														assign node14255 = (inp[1]) ? node14257 : 4'b0000;
															assign node14257 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node14260 = (inp[1]) ? node14262 : 4'b0001;
															assign node14262 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node14265 = (inp[1]) ? node14365 : node14266;
										assign node14266 = (inp[7]) ? node14312 : node14267;
											assign node14267 = (inp[0]) ? node14293 : node14268;
												assign node14268 = (inp[10]) ? node14282 : node14269;
													assign node14269 = (inp[12]) ? node14275 : node14270;
														assign node14270 = (inp[13]) ? node14272 : 4'b1000;
															assign node14272 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node14275 = (inp[2]) ? node14279 : node14276;
															assign node14276 = (inp[13]) ? 4'b0001 : 4'b1000;
															assign node14279 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node14282 = (inp[13]) ? node14288 : node14283;
														assign node14283 = (inp[12]) ? node14285 : 4'b0001;
															assign node14285 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node14288 = (inp[2]) ? node14290 : 4'b1001;
															assign node14290 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node14293 = (inp[13]) ? node14303 : node14294;
													assign node14294 = (inp[2]) ? node14296 : 4'b0000;
														assign node14296 = (inp[12]) ? node14300 : node14297;
															assign node14297 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node14300 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node14303 = (inp[2]) ? node14307 : node14304;
														assign node14304 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node14307 = (inp[10]) ? 4'b0001 : node14308;
															assign node14308 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node14312 = (inp[2]) ? node14340 : node14313;
												assign node14313 = (inp[13]) ? node14327 : node14314;
													assign node14314 = (inp[10]) ? node14320 : node14315;
														assign node14315 = (inp[0]) ? 4'b1001 : node14316;
															assign node14316 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node14320 = (inp[14]) ? node14324 : node14321;
															assign node14321 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node14324 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node14327 = (inp[12]) ? node14333 : node14328;
														assign node14328 = (inp[10]) ? node14330 : 4'b0000;
															assign node14330 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node14333 = (inp[0]) ? node14337 : node14334;
															assign node14334 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node14337 = (inp[10]) ? 4'b1001 : 4'b0000;
												assign node14340 = (inp[0]) ? node14354 : node14341;
													assign node14341 = (inp[10]) ? node14347 : node14342;
														assign node14342 = (inp[12]) ? node14344 : 4'b0001;
															assign node14344 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node14347 = (inp[13]) ? node14351 : node14348;
															assign node14348 = (inp[14]) ? 4'b0000 : 4'b1000;
															assign node14351 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14354 = (inp[13]) ? node14360 : node14355;
														assign node14355 = (inp[10]) ? node14357 : 4'b1001;
															assign node14357 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14360 = (inp[10]) ? 4'b1000 : node14361;
															assign node14361 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node14365 = (inp[13]) ? node14421 : node14366;
											assign node14366 = (inp[2]) ? node14404 : node14367;
												assign node14367 = (inp[10]) ? node14377 : node14368;
													assign node14368 = (inp[12]) ? node14374 : node14369;
														assign node14369 = (inp[7]) ? 4'b1000 : node14370;
															assign node14370 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node14374 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node14377 = (inp[12]) ? node14391 : node14378;
														assign node14378 = (inp[14]) ? node14386 : node14379;
															assign node14379 = (inp[0]) ? node14383 : node14380;
																assign node14380 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node14383 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node14386 = (inp[7]) ? node14388 : 4'b0000;
																assign node14388 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node14391 = (inp[14]) ? node14397 : node14392;
															assign node14392 = (inp[7]) ? 4'b0000 : node14393;
																assign node14393 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node14397 = (inp[7]) ? node14401 : node14398;
																assign node14398 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node14401 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node14404 = (inp[0]) ? node14406 : 4'b0000;
													assign node14406 = (inp[12]) ? node14412 : node14407;
														assign node14407 = (inp[10]) ? node14409 : 4'b0000;
															assign node14409 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node14412 = (inp[14]) ? node14414 : 4'b1000;
															assign node14414 = (inp[7]) ? node14418 : node14415;
																assign node14415 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node14418 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node14421 = (inp[10]) ? 4'b1000 : node14422;
												assign node14422 = (inp[0]) ? node14440 : node14423;
													assign node14423 = (inp[14]) ? node14433 : node14424;
														assign node14424 = (inp[2]) ? node14428 : node14425;
															assign node14425 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node14428 = (inp[7]) ? 4'b1000 : node14429;
																assign node14429 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14433 = (inp[2]) ? node14435 : 4'b1000;
															assign node14435 = (inp[12]) ? node14437 : 4'b1000;
																assign node14437 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node14440 = (inp[7]) ? node14442 : 4'b0000;
														assign node14442 = (inp[2]) ? 4'b0000 : node14443;
															assign node14443 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node14448 = (inp[13]) ? node14632 : node14449;
									assign node14449 = (inp[1]) ? node14557 : node14450;
										assign node14450 = (inp[10]) ? node14498 : node14451;
											assign node14451 = (inp[2]) ? node14477 : node14452;
												assign node14452 = (inp[0]) ? node14464 : node14453;
													assign node14453 = (inp[12]) ? node14459 : node14454;
														assign node14454 = (inp[7]) ? 4'b1000 : node14455;
															assign node14455 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node14459 = (inp[11]) ? node14461 : 4'b1000;
															assign node14461 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node14464 = (inp[7]) ? node14468 : node14465;
														assign node14465 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node14468 = (inp[11]) ? node14474 : node14469;
															assign node14469 = (inp[14]) ? node14471 : 4'b0000;
																assign node14471 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node14474 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node14477 = (inp[11]) ? node14491 : node14478;
													assign node14478 = (inp[7]) ? node14482 : node14479;
														assign node14479 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14482 = (inp[14]) ? node14488 : node14483;
															assign node14483 = (inp[12]) ? 4'b1001 : node14484;
																assign node14484 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node14488 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node14491 = (inp[7]) ? node14495 : node14492;
														assign node14492 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node14495 = (inp[0]) ? 4'b1000 : 4'b0000;
											assign node14498 = (inp[0]) ? node14530 : node14499;
												assign node14499 = (inp[2]) ? node14509 : node14500;
													assign node14500 = (inp[7]) ? 4'b0001 : node14501;
														assign node14501 = (inp[12]) ? node14505 : node14502;
															assign node14502 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node14505 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node14509 = (inp[14]) ? node14523 : node14510;
														assign node14510 = (inp[12]) ? node14516 : node14511;
															assign node14511 = (inp[7]) ? 4'b1000 : node14512;
																assign node14512 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node14516 = (inp[11]) ? node14520 : node14517;
																assign node14517 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node14520 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node14523 = (inp[7]) ? node14525 : 4'b0000;
															assign node14525 = (inp[12]) ? node14527 : 4'b0001;
																assign node14527 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node14530 = (inp[12]) ? node14542 : node14531;
													assign node14531 = (inp[7]) ? node14539 : node14532;
														assign node14532 = (inp[11]) ? 4'b0000 : node14533;
															assign node14533 = (inp[14]) ? node14535 : 4'b0000;
																assign node14535 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node14539 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node14542 = (inp[2]) ? node14548 : node14543;
														assign node14543 = (inp[11]) ? 4'b0000 : node14544;
															assign node14544 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node14548 = (inp[14]) ? node14550 : 4'b0001;
															assign node14550 = (inp[11]) ? node14554 : node14551;
																assign node14551 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node14554 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node14557 = (inp[11]) ? node14605 : node14558;
											assign node14558 = (inp[14]) ? node14584 : node14559;
												assign node14559 = (inp[2]) ? node14571 : node14560;
													assign node14560 = (inp[0]) ? node14566 : node14561;
														assign node14561 = (inp[7]) ? 4'b0001 : node14562;
															assign node14562 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node14566 = (inp[12]) ? node14568 : 4'b0000;
															assign node14568 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node14571 = (inp[0]) ? node14579 : node14572;
														assign node14572 = (inp[12]) ? 4'b0001 : node14573;
															assign node14573 = (inp[10]) ? 4'b0000 : node14574;
																assign node14574 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node14579 = (inp[12]) ? node14581 : 4'b0001;
															assign node14581 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node14584 = (inp[7]) ? node14596 : node14585;
													assign node14585 = (inp[0]) ? node14589 : node14586;
														assign node14586 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14589 = (inp[12]) ? node14591 : 4'b0001;
															assign node14591 = (inp[2]) ? node14593 : 4'b0001;
																assign node14593 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node14596 = (inp[0]) ? node14600 : node14597;
														assign node14597 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node14600 = (inp[12]) ? 4'b0000 : node14601;
															assign node14601 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node14605 = (inp[10]) ? 4'b0000 : node14606;
												assign node14606 = (inp[2]) ? node14620 : node14607;
													assign node14607 = (inp[7]) ? node14613 : node14608;
														assign node14608 = (inp[12]) ? node14610 : 4'b0000;
															assign node14610 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node14613 = (inp[0]) ? node14617 : node14614;
															assign node14614 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14617 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node14620 = (inp[7]) ? node14626 : node14621;
														assign node14621 = (inp[14]) ? node14623 : 4'b1000;
															assign node14623 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node14626 = (inp[12]) ? 4'b0000 : node14627;
															assign node14627 = (inp[0]) ? 4'b1000 : 4'b0000;
									assign node14632 = (inp[10]) ? node14714 : node14633;
										assign node14633 = (inp[11]) ? node14683 : node14634;
											assign node14634 = (inp[12]) ? node14656 : node14635;
												assign node14635 = (inp[0]) ? node14647 : node14636;
													assign node14636 = (inp[1]) ? node14640 : node14637;
														assign node14637 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node14640 = (inp[14]) ? node14642 : 4'b0001;
															assign node14642 = (inp[2]) ? 4'b0001 : node14643;
																assign node14643 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node14647 = (inp[2]) ? 4'b0000 : node14648;
														assign node14648 = (inp[14]) ? 4'b0001 : node14649;
															assign node14649 = (inp[1]) ? 4'b0000 : node14650;
																assign node14650 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node14656 = (inp[7]) ? node14672 : node14657;
													assign node14657 = (inp[1]) ? node14667 : node14658;
														assign node14658 = (inp[0]) ? node14662 : node14659;
															assign node14659 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node14662 = (inp[2]) ? 4'b0000 : node14663;
																assign node14663 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node14667 = (inp[0]) ? 4'b0001 : node14668;
															assign node14668 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node14672 = (inp[14]) ? 4'b0000 : node14673;
														assign node14673 = (inp[1]) ? 4'b0000 : node14674;
															assign node14674 = (inp[2]) ? node14678 : node14675;
																assign node14675 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node14678 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node14683 = (inp[1]) ? 4'b0000 : node14684;
												assign node14684 = (inp[14]) ? node14704 : node14685;
													assign node14685 = (inp[7]) ? node14695 : node14686;
														assign node14686 = (inp[2]) ? node14690 : node14687;
															assign node14687 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node14690 = (inp[0]) ? 4'b0001 : node14691;
																assign node14691 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node14695 = (inp[2]) ? 4'b0000 : node14696;
															assign node14696 = (inp[12]) ? node14700 : node14697;
																assign node14697 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node14700 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node14704 = (inp[2]) ? node14706 : 4'b0000;
														assign node14706 = (inp[12]) ? node14710 : node14707;
															assign node14707 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node14710 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node14714 = (inp[1]) ? 4'b0000 : node14715;
											assign node14715 = (inp[11]) ? 4'b0000 : node14716;
												assign node14716 = (inp[14]) ? node14728 : node14717;
													assign node14717 = (inp[7]) ? node14719 : 4'b0000;
														assign node14719 = (inp[12]) ? node14721 : 4'b0000;
															assign node14721 = (inp[0]) ? node14725 : node14722;
																assign node14722 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node14725 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node14728 = (inp[7]) ? node14738 : node14729;
														assign node14729 = (inp[2]) ? node14733 : node14730;
															assign node14730 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node14733 = (inp[0]) ? 4'b0001 : node14734;
																assign node14734 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node14738 = (inp[12]) ? 4'b0000 : node14739;
															assign node14739 = (inp[2]) ? node14743 : node14740;
																assign node14740 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node14743 = (inp[0]) ? 4'b0001 : 4'b0000;
				assign node14749 = (inp[0]) ? node16703 : node14750;
					assign node14750 = (inp[6]) ? node15330 : node14751;
						assign node14751 = (inp[5]) ? node14873 : node14752;
							assign node14752 = (inp[3]) ? node14754 : 4'b1010;
								assign node14754 = (inp[2]) ? 4'b1010 : node14755;
									assign node14755 = (inp[4]) ? node14809 : node14756;
										assign node14756 = (inp[7]) ? 4'b1010 : node14757;
											assign node14757 = (inp[13]) ? node14785 : node14758;
												assign node14758 = (inp[12]) ? node14778 : node14759;
													assign node14759 = (inp[10]) ? node14767 : node14760;
														assign node14760 = (inp[1]) ? node14762 : 4'b1010;
															assign node14762 = (inp[11]) ? 4'b0000 : node14763;
																assign node14763 = (inp[14]) ? 4'b1010 : 4'b0000;
														assign node14767 = (inp[1]) ? node14773 : node14768;
															assign node14768 = (inp[11]) ? 4'b0001 : node14769;
																assign node14769 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14773 = (inp[11]) ? 4'b0000 : node14774;
																assign node14774 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node14778 = (inp[14]) ? 4'b1010 : node14779;
														assign node14779 = (inp[10]) ? node14781 : 4'b1010;
															assign node14781 = (inp[1]) ? 4'b0000 : 4'b1010;
												assign node14785 = (inp[1]) ? node14797 : node14786;
													assign node14786 = (inp[10]) ? node14792 : node14787;
														assign node14787 = (inp[14]) ? node14789 : 4'b0001;
															assign node14789 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node14792 = (inp[12]) ? 4'b0001 : node14793;
															assign node14793 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14797 = (inp[11]) ? node14803 : node14798;
														assign node14798 = (inp[14]) ? node14800 : 4'b1000;
															assign node14800 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node14803 = (inp[10]) ? 4'b1000 : node14804;
															assign node14804 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node14809 = (inp[1]) ? node14843 : node14810;
											assign node14810 = (inp[13]) ? node14830 : node14811;
												assign node14811 = (inp[7]) ? node14821 : node14812;
													assign node14812 = (inp[12]) ? node14816 : node14813;
														assign node14813 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node14816 = (inp[14]) ? node14818 : 4'b1001;
															assign node14818 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node14821 = (inp[10]) ? node14823 : 4'b1010;
														assign node14823 = (inp[12]) ? 4'b1010 : node14824;
															assign node14824 = (inp[11]) ? 4'b0001 : node14825;
																assign node14825 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node14830 = (inp[14]) ? node14836 : node14831;
													assign node14831 = (inp[12]) ? 4'b0001 : node14832;
														assign node14832 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14836 = (inp[11]) ? node14840 : node14837;
														assign node14837 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14840 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node14843 = (inp[14]) ? node14855 : node14844;
												assign node14844 = (inp[13]) ? node14850 : node14845;
													assign node14845 = (inp[10]) ? 4'b0000 : node14846;
														assign node14846 = (inp[7]) ? 4'b1010 : 4'b0000;
													assign node14850 = (inp[10]) ? 4'b1000 : node14851;
														assign node14851 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node14855 = (inp[11]) ? node14867 : node14856;
													assign node14856 = (inp[13]) ? node14862 : node14857;
														assign node14857 = (inp[10]) ? 4'b0001 : node14858;
															assign node14858 = (inp[7]) ? 4'b1010 : 4'b1001;
														assign node14862 = (inp[12]) ? 4'b0001 : node14863;
															assign node14863 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14867 = (inp[13]) ? node14869 : 4'b0000;
														assign node14869 = (inp[12]) ? 4'b0000 : 4'b1000;
							assign node14873 = (inp[2]) ? node15201 : node14874;
								assign node14874 = (inp[1]) ? node15038 : node14875;
									assign node14875 = (inp[14]) ? node14949 : node14876;
										assign node14876 = (inp[13]) ? node14908 : node14877;
											assign node14877 = (inp[10]) ? node14887 : node14878;
												assign node14878 = (inp[3]) ? node14882 : node14879;
													assign node14879 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node14882 = (inp[7]) ? 4'b1101 : node14883;
														assign node14883 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node14887 = (inp[12]) ? node14901 : node14888;
													assign node14888 = (inp[11]) ? node14894 : node14889;
														assign node14889 = (inp[3]) ? node14891 : 4'b0101;
															assign node14891 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node14894 = (inp[7]) ? node14896 : 4'b0001;
															assign node14896 = (inp[3]) ? 4'b0101 : node14897;
																assign node14897 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node14901 = (inp[3]) ? node14903 : 4'b1001;
														assign node14903 = (inp[4]) ? node14905 : 4'b1101;
															assign node14905 = (inp[11]) ? 4'b1001 : 4'b1101;
											assign node14908 = (inp[10]) ? node14920 : node14909;
												assign node14909 = (inp[3]) ? node14915 : node14910;
													assign node14910 = (inp[4]) ? 4'b0101 : node14911;
														assign node14911 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node14915 = (inp[7]) ? node14917 : 4'b0001;
														assign node14917 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node14920 = (inp[12]) ? node14932 : node14921;
													assign node14921 = (inp[11]) ? 4'b1001 : node14922;
														assign node14922 = (inp[3]) ? node14928 : node14923;
															assign node14923 = (inp[4]) ? 4'b1101 : node14924;
																assign node14924 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node14928 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node14932 = (inp[11]) ? node14940 : node14933;
														assign node14933 = (inp[4]) ? 4'b0001 : node14934;
															assign node14934 = (inp[7]) ? node14936 : 4'b0001;
																assign node14936 = (inp[3]) ? 4'b0101 : 4'b0001;
														assign node14940 = (inp[3]) ? node14946 : node14941;
															assign node14941 = (inp[7]) ? node14943 : 4'b0101;
																assign node14943 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node14946 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node14949 = (inp[11]) ? node14989 : node14950;
											assign node14950 = (inp[13]) ? node14974 : node14951;
												assign node14951 = (inp[10]) ? node14963 : node14952;
													assign node14952 = (inp[3]) ? node14958 : node14953;
														assign node14953 = (inp[4]) ? node14955 : 4'b1000;
															assign node14955 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node14958 = (inp[7]) ? 4'b1100 : node14959;
															assign node14959 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node14963 = (inp[12]) ? node14967 : node14964;
														assign node14964 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node14967 = (inp[3]) ? node14971 : node14968;
															assign node14968 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node14971 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node14974 = (inp[10]) ? node14982 : node14975;
													assign node14975 = (inp[3]) ? node14977 : 4'b0100;
														assign node14977 = (inp[4]) ? 4'b0000 : node14978;
															assign node14978 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node14982 = (inp[12]) ? 4'b0100 : node14983;
														assign node14983 = (inp[4]) ? node14985 : 4'b1100;
															assign node14985 = (inp[3]) ? 4'b1000 : 4'b1100;
											assign node14989 = (inp[13]) ? node15015 : node14990;
												assign node14990 = (inp[12]) ? node15004 : node14991;
													assign node14991 = (inp[10]) ? node14995 : node14992;
														assign node14992 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node14995 = (inp[4]) ? node15001 : node14996;
															assign node14996 = (inp[3]) ? node14998 : 4'b0001;
																assign node14998 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node15001 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node15004 = (inp[4]) ? node15008 : node15005;
														assign node15005 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node15008 = (inp[7]) ? node15012 : node15009;
															assign node15009 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node15012 = (inp[3]) ? 4'b1101 : 4'b1001;
												assign node15015 = (inp[10]) ? node15023 : node15016;
													assign node15016 = (inp[3]) ? 4'b0001 : node15017;
														assign node15017 = (inp[7]) ? node15019 : 4'b0101;
															assign node15019 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node15023 = (inp[12]) ? node15031 : node15024;
														assign node15024 = (inp[3]) ? 4'b1001 : node15025;
															assign node15025 = (inp[7]) ? node15027 : 4'b1101;
																assign node15027 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node15031 = (inp[4]) ? 4'b0101 : node15032;
															assign node15032 = (inp[3]) ? 4'b0101 : node15033;
																assign node15033 = (inp[7]) ? 4'b0001 : 4'b0101;
									assign node15038 = (inp[11]) ? node15136 : node15039;
										assign node15039 = (inp[14]) ? node15081 : node15040;
											assign node15040 = (inp[13]) ? node15058 : node15041;
												assign node15041 = (inp[10]) ? node15049 : node15042;
													assign node15042 = (inp[12]) ? node15044 : 4'b0100;
														assign node15044 = (inp[7]) ? 4'b1100 : node15045;
															assign node15045 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node15049 = (inp[3]) ? node15053 : node15050;
														assign node15050 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15053 = (inp[7]) ? node15055 : 4'b0000;
															assign node15055 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node15058 = (inp[12]) ? node15070 : node15059;
													assign node15059 = (inp[3]) ? node15065 : node15060;
														assign node15060 = (inp[4]) ? 4'b1100 : node15061;
															assign node15061 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node15065 = (inp[7]) ? node15067 : 4'b1000;
															assign node15067 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node15070 = (inp[10]) ? node15078 : node15071;
														assign node15071 = (inp[4]) ? node15075 : node15072;
															assign node15072 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node15075 = (inp[3]) ? 4'b0000 : 4'b0100;
														assign node15078 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node15081 = (inp[13]) ? node15115 : node15082;
												assign node15082 = (inp[12]) ? node15104 : node15083;
													assign node15083 = (inp[10]) ? node15093 : node15084;
														assign node15084 = (inp[3]) ? node15090 : node15085;
															assign node15085 = (inp[4]) ? node15087 : 4'b1001;
																assign node15087 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node15090 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node15093 = (inp[3]) ? node15099 : node15094;
															assign node15094 = (inp[4]) ? 4'b0101 : node15095;
																assign node15095 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node15099 = (inp[7]) ? node15101 : 4'b0001;
																assign node15101 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node15104 = (inp[3]) ? node15110 : node15105;
														assign node15105 = (inp[4]) ? node15107 : 4'b1001;
															assign node15107 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node15110 = (inp[4]) ? node15112 : 4'b1101;
															assign node15112 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node15115 = (inp[12]) ? node15125 : node15116;
													assign node15116 = (inp[10]) ? node15118 : 4'b0001;
														assign node15118 = (inp[7]) ? node15122 : node15119;
															assign node15119 = (inp[3]) ? 4'b1001 : 4'b1101;
															assign node15122 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node15125 = (inp[3]) ? node15131 : node15126;
														assign node15126 = (inp[4]) ? 4'b0101 : node15127;
															assign node15127 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node15131 = (inp[4]) ? 4'b0001 : node15132;
															assign node15132 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node15136 = (inp[13]) ? node15166 : node15137;
											assign node15137 = (inp[12]) ? node15149 : node15138;
												assign node15138 = (inp[3]) ? node15144 : node15139;
													assign node15139 = (inp[4]) ? 4'b0100 : node15140;
														assign node15140 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node15144 = (inp[4]) ? 4'b0000 : node15145;
														assign node15145 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node15149 = (inp[10]) ? node15157 : node15150;
													assign node15150 = (inp[4]) ? node15152 : 4'b1100;
														assign node15152 = (inp[7]) ? 4'b1000 : node15153;
															assign node15153 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node15157 = (inp[7]) ? node15159 : 4'b0100;
														assign node15159 = (inp[4]) ? node15163 : node15160;
															assign node15160 = (inp[3]) ? 4'b0100 : 4'b0000;
															assign node15163 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node15166 = (inp[10]) ? node15190 : node15167;
												assign node15167 = (inp[12]) ? node15179 : node15168;
													assign node15168 = (inp[3]) ? node15174 : node15169;
														assign node15169 = (inp[7]) ? node15171 : 4'b1100;
															assign node15171 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node15174 = (inp[7]) ? node15176 : 4'b1000;
															assign node15176 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node15179 = (inp[3]) ? node15185 : node15180;
														assign node15180 = (inp[4]) ? 4'b0100 : node15181;
															assign node15181 = (inp[14]) ? 4'b0000 : 4'b0100;
														assign node15185 = (inp[14]) ? node15187 : 4'b0000;
															assign node15187 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node15190 = (inp[3]) ? node15196 : node15191;
													assign node15191 = (inp[4]) ? 4'b1100 : node15192;
														assign node15192 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node15196 = (inp[7]) ? node15198 : 4'b1000;
														assign node15198 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node15201 = (inp[3]) ? node15203 : 4'b1010;
									assign node15203 = (inp[4]) ? node15253 : node15204;
										assign node15204 = (inp[7]) ? 4'b1010 : node15205;
											assign node15205 = (inp[13]) ? node15227 : node15206;
												assign node15206 = (inp[12]) ? node15220 : node15207;
													assign node15207 = (inp[10]) ? node15211 : node15208;
														assign node15208 = (inp[1]) ? 4'b0000 : 4'b1010;
														assign node15211 = (inp[14]) ? node15213 : 4'b0000;
															assign node15213 = (inp[1]) ? node15217 : node15214;
																assign node15214 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node15217 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node15220 = (inp[14]) ? 4'b1010 : node15221;
														assign node15221 = (inp[10]) ? node15223 : 4'b1010;
															assign node15223 = (inp[1]) ? 4'b0000 : 4'b1010;
												assign node15227 = (inp[12]) ? node15239 : node15228;
													assign node15228 = (inp[10]) ? node15234 : node15229;
														assign node15229 = (inp[1]) ? 4'b1000 : node15230;
															assign node15230 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15234 = (inp[1]) ? 4'b1001 : node15235;
															assign node15235 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node15239 = (inp[1]) ? node15245 : node15240;
														assign node15240 = (inp[11]) ? 4'b0001 : node15241;
															assign node15241 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node15245 = (inp[10]) ? 4'b1000 : node15246;
															assign node15246 = (inp[14]) ? node15248 : 4'b0000;
																assign node15248 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node15253 = (inp[1]) ? node15291 : node15254;
											assign node15254 = (inp[13]) ? node15280 : node15255;
												assign node15255 = (inp[7]) ? node15271 : node15256;
													assign node15256 = (inp[11]) ? node15266 : node15257;
														assign node15257 = (inp[14]) ? node15263 : node15258;
															assign node15258 = (inp[12]) ? 4'b1001 : node15259;
																assign node15259 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node15263 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node15266 = (inp[12]) ? 4'b1001 : node15267;
															assign node15267 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node15271 = (inp[10]) ? node15273 : 4'b1010;
														assign node15273 = (inp[12]) ? 4'b1010 : node15274;
															assign node15274 = (inp[11]) ? 4'b0001 : node15275;
																assign node15275 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node15280 = (inp[11]) ? node15286 : node15281;
													assign node15281 = (inp[14]) ? 4'b0000 : node15282;
														assign node15282 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15286 = (inp[10]) ? node15288 : 4'b0001;
														assign node15288 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node15291 = (inp[11]) ? node15317 : node15292;
												assign node15292 = (inp[14]) ? node15306 : node15293;
													assign node15293 = (inp[13]) ? node15301 : node15294;
														assign node15294 = (inp[12]) ? node15296 : 4'b0000;
															assign node15296 = (inp[10]) ? 4'b0000 : node15297;
																assign node15297 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node15301 = (inp[12]) ? node15303 : 4'b1000;
															assign node15303 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node15306 = (inp[12]) ? node15314 : node15307;
														assign node15307 = (inp[10]) ? node15311 : node15308;
															assign node15308 = (inp[7]) ? 4'b1010 : 4'b1001;
															assign node15311 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node15314 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node15317 = (inp[13]) ? node15325 : node15318;
													assign node15318 = (inp[10]) ? 4'b0000 : node15319;
														assign node15319 = (inp[12]) ? node15321 : 4'b0000;
															assign node15321 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node15325 = (inp[10]) ? 4'b1000 : node15326;
														assign node15326 = (inp[12]) ? 4'b0000 : 4'b1000;
						assign node15330 = (inp[5]) ? node16014 : node15331;
							assign node15331 = (inp[11]) ? node15721 : node15332;
								assign node15332 = (inp[3]) ? node15534 : node15333;
									assign node15333 = (inp[7]) ? node15445 : node15334;
										assign node15334 = (inp[2]) ? node15390 : node15335;
											assign node15335 = (inp[4]) ? node15373 : node15336;
												assign node15336 = (inp[13]) ? node15354 : node15337;
													assign node15337 = (inp[10]) ? node15347 : node15338;
														assign node15338 = (inp[14]) ? node15344 : node15339;
															assign node15339 = (inp[1]) ? node15341 : 4'b1001;
																assign node15341 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node15344 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node15347 = (inp[14]) ? node15349 : 4'b0100;
															assign node15349 = (inp[12]) ? 4'b1001 : node15350;
																assign node15350 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node15354 = (inp[10]) ? node15364 : node15355;
														assign node15355 = (inp[12]) ? node15361 : node15356;
															assign node15356 = (inp[1]) ? 4'b1100 : node15357;
																assign node15357 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node15361 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node15364 = (inp[12]) ? node15368 : node15365;
															assign node15365 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node15368 = (inp[14]) ? node15370 : 4'b1100;
																assign node15370 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node15373 = (inp[10]) ? node15385 : node15374;
													assign node15374 = (inp[12]) ? node15378 : node15375;
														assign node15375 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node15378 = (inp[13]) ? 4'b1001 : node15379;
															assign node15379 = (inp[14]) ? 4'b1100 : node15380;
																assign node15380 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node15385 = (inp[1]) ? node15387 : 4'b0001;
														assign node15387 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node15390 = (inp[13]) ? node15424 : node15391;
												assign node15391 = (inp[4]) ? node15405 : node15392;
													assign node15392 = (inp[12]) ? node15398 : node15393;
														assign node15393 = (inp[14]) ? node15395 : 4'b1001;
															assign node15395 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node15398 = (inp[10]) ? 4'b1001 : node15399;
															assign node15399 = (inp[1]) ? node15401 : 4'b1001;
																assign node15401 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node15405 = (inp[12]) ? node15415 : node15406;
														assign node15406 = (inp[10]) ? node15412 : node15407;
															assign node15407 = (inp[14]) ? 4'b1101 : node15408;
																assign node15408 = (inp[1]) ? 4'b0100 : 4'b1101;
															assign node15412 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node15415 = (inp[14]) ? node15421 : node15416;
															assign node15416 = (inp[1]) ? node15418 : 4'b1101;
																assign node15418 = (inp[10]) ? 4'b0100 : 4'b1100;
															assign node15421 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node15424 = (inp[12]) ? node15438 : node15425;
													assign node15425 = (inp[10]) ? node15431 : node15426;
														assign node15426 = (inp[1]) ? 4'b1100 : node15427;
															assign node15427 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node15431 = (inp[1]) ? node15435 : node15432;
															assign node15432 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node15435 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node15438 = (inp[1]) ? node15442 : node15439;
														assign node15439 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node15442 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node15445 = (inp[4]) ? node15491 : node15446;
											assign node15446 = (inp[13]) ? node15472 : node15447;
												assign node15447 = (inp[12]) ? node15463 : node15448;
													assign node15448 = (inp[10]) ? node15456 : node15449;
														assign node15449 = (inp[14]) ? node15453 : node15450;
															assign node15450 = (inp[1]) ? 4'b0000 : 4'b1001;
															assign node15453 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node15456 = (inp[1]) ? node15460 : node15457;
															assign node15457 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node15460 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node15463 = (inp[14]) ? node15469 : node15464;
														assign node15464 = (inp[1]) ? node15466 : 4'b1001;
															assign node15466 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node15469 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node15472 = (inp[1]) ? node15484 : node15473;
													assign node15473 = (inp[14]) ? node15479 : node15474;
														assign node15474 = (inp[10]) ? node15476 : 4'b0001;
															assign node15476 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15479 = (inp[12]) ? 4'b0000 : node15480;
															assign node15480 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node15484 = (inp[14]) ? node15486 : 4'b1000;
														assign node15486 = (inp[2]) ? node15488 : 4'b0001;
															assign node15488 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node15491 = (inp[13]) ? node15513 : node15492;
												assign node15492 = (inp[1]) ? node15506 : node15493;
													assign node15493 = (inp[14]) ? node15499 : node15494;
														assign node15494 = (inp[12]) ? 4'b1001 : node15495;
															assign node15495 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node15499 = (inp[2]) ? node15501 : 4'b1000;
															assign node15501 = (inp[10]) ? node15503 : 4'b1000;
																assign node15503 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node15506 = (inp[14]) ? node15508 : 4'b0100;
														assign node15508 = (inp[10]) ? node15510 : 4'b1001;
															assign node15510 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node15513 = (inp[10]) ? node15523 : node15514;
													assign node15514 = (inp[12]) ? node15520 : node15515;
														assign node15515 = (inp[1]) ? 4'b0001 : node15516;
															assign node15516 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node15520 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node15523 = (inp[2]) ? node15529 : node15524;
														assign node15524 = (inp[12]) ? 4'b0001 : node15525;
															assign node15525 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node15529 = (inp[1]) ? 4'b1100 : node15530;
															assign node15530 = (inp[12]) ? 4'b0101 : 4'b1101;
									assign node15534 = (inp[10]) ? node15620 : node15535;
										assign node15535 = (inp[2]) ? node15567 : node15536;
											assign node15536 = (inp[12]) ? node15556 : node15537;
												assign node15537 = (inp[1]) ? node15545 : node15538;
													assign node15538 = (inp[4]) ? 4'b1101 : node15539;
														assign node15539 = (inp[14]) ? 4'b1001 : node15540;
															assign node15540 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node15545 = (inp[4]) ? node15551 : node15546;
														assign node15546 = (inp[13]) ? 4'b0101 : node15547;
															assign node15547 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node15551 = (inp[7]) ? node15553 : 4'b0001;
															assign node15553 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node15556 = (inp[4]) ? node15562 : node15557;
													assign node15557 = (inp[7]) ? 4'b1001 : node15558;
														assign node15558 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node15562 = (inp[13]) ? node15564 : 4'b1101;
														assign node15564 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node15567 = (inp[13]) ? node15595 : node15568;
												assign node15568 = (inp[4]) ? node15578 : node15569;
													assign node15569 = (inp[1]) ? node15573 : node15570;
														assign node15570 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node15573 = (inp[14]) ? 4'b1101 : node15574;
															assign node15574 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node15578 = (inp[7]) ? node15586 : node15579;
														assign node15579 = (inp[12]) ? node15581 : 4'b0001;
															assign node15581 = (inp[1]) ? 4'b1001 : node15582;
																assign node15582 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15586 = (inp[12]) ? node15590 : node15587;
															assign node15587 = (inp[1]) ? 4'b0000 : 4'b1101;
															assign node15590 = (inp[1]) ? node15592 : 4'b1100;
																assign node15592 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node15595 = (inp[4]) ? node15609 : node15596;
													assign node15596 = (inp[7]) ? node15602 : node15597;
														assign node15597 = (inp[1]) ? 4'b0001 : node15598;
															assign node15598 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15602 = (inp[14]) ? node15606 : node15603;
															assign node15603 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node15606 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node15609 = (inp[7]) ? node15615 : node15610;
														assign node15610 = (inp[12]) ? 4'b1001 : node15611;
															assign node15611 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node15615 = (inp[1]) ? 4'b0001 : node15616;
															assign node15616 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node15620 = (inp[4]) ? node15678 : node15621;
											assign node15621 = (inp[2]) ? node15639 : node15622;
												assign node15622 = (inp[7]) ? node15628 : node15623;
													assign node15623 = (inp[12]) ? 4'b0101 : node15624;
														assign node15624 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node15628 = (inp[13]) ? node15634 : node15629;
														assign node15629 = (inp[12]) ? 4'b0001 : node15630;
															assign node15630 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node15634 = (inp[12]) ? 4'b0101 : node15635;
															assign node15635 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node15639 = (inp[7]) ? node15661 : node15640;
													assign node15640 = (inp[13]) ? node15650 : node15641;
														assign node15641 = (inp[12]) ? node15643 : 4'b0000;
															assign node15643 = (inp[14]) ? node15647 : node15644;
																assign node15644 = (inp[1]) ? 4'b0000 : 4'b1101;
																assign node15647 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node15650 = (inp[12]) ? node15656 : node15651;
															assign node15651 = (inp[14]) ? node15653 : 4'b1000;
																assign node15653 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node15656 = (inp[1]) ? 4'b1000 : node15657;
																assign node15657 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node15661 = (inp[13]) ? node15671 : node15662;
														assign node15662 = (inp[1]) ? node15668 : node15663;
															assign node15663 = (inp[14]) ? 4'b0100 : node15664;
																assign node15664 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node15668 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node15671 = (inp[1]) ? node15675 : node15672;
															assign node15672 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node15675 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node15678 = (inp[1]) ? node15692 : node15679;
												assign node15679 = (inp[13]) ? node15687 : node15680;
													assign node15680 = (inp[7]) ? node15682 : 4'b0001;
														assign node15682 = (inp[12]) ? 4'b1101 : node15683;
															assign node15683 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node15687 = (inp[2]) ? 4'b0001 : node15688;
														assign node15688 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node15692 = (inp[12]) ? node15708 : node15693;
													assign node15693 = (inp[13]) ? node15703 : node15694;
														assign node15694 = (inp[2]) ? node15700 : node15695;
															assign node15695 = (inp[7]) ? 4'b1101 : node15696;
																assign node15696 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node15700 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node15703 = (inp[14]) ? node15705 : 4'b1001;
															assign node15705 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node15708 = (inp[13]) ? node15716 : node15709;
														assign node15709 = (inp[7]) ? node15711 : 4'b0001;
															assign node15711 = (inp[14]) ? 4'b1101 : node15712;
																assign node15712 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node15716 = (inp[14]) ? node15718 : 4'b0001;
															assign node15718 = (inp[2]) ? 4'b0001 : 4'b0000;
								assign node15721 = (inp[1]) ? node15873 : node15722;
									assign node15722 = (inp[3]) ? node15788 : node15723;
										assign node15723 = (inp[13]) ? node15753 : node15724;
											assign node15724 = (inp[12]) ? node15744 : node15725;
												assign node15725 = (inp[10]) ? node15737 : node15726;
													assign node15726 = (inp[2]) ? node15732 : node15727;
														assign node15727 = (inp[7]) ? 4'b1001 : node15728;
															assign node15728 = (inp[4]) ? 4'b0000 : 4'b1001;
														assign node15732 = (inp[7]) ? 4'b1001 : node15733;
															assign node15733 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node15737 = (inp[7]) ? node15741 : node15738;
														assign node15738 = (inp[4]) ? 4'b1000 : 4'b0101;
														assign node15741 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node15744 = (inp[7]) ? 4'b1001 : node15745;
													assign node15745 = (inp[4]) ? node15747 : 4'b1001;
														assign node15747 = (inp[10]) ? node15749 : 4'b1101;
															assign node15749 = (inp[2]) ? 4'b1101 : 4'b0000;
											assign node15753 = (inp[2]) ? node15779 : node15754;
												assign node15754 = (inp[4]) ? node15764 : node15755;
													assign node15755 = (inp[7]) ? node15759 : node15756;
														assign node15756 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node15759 = (inp[12]) ? 4'b0001 : node15760;
															assign node15760 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node15764 = (inp[7]) ? node15774 : node15765;
														assign node15765 = (inp[14]) ? node15767 : 4'b1000;
															assign node15767 = (inp[12]) ? node15771 : node15768;
																assign node15768 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node15771 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node15774 = (inp[10]) ? node15776 : 4'b0101;
															assign node15776 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node15779 = (inp[10]) ? node15785 : node15780;
													assign node15780 = (inp[7]) ? node15782 : 4'b0101;
														assign node15782 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node15785 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node15788 = (inp[4]) ? node15816 : node15789;
											assign node15789 = (inp[2]) ? node15811 : node15790;
												assign node15790 = (inp[7]) ? node15802 : node15791;
													assign node15791 = (inp[13]) ? node15795 : node15792;
														assign node15792 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node15795 = (inp[10]) ? node15799 : node15796;
															assign node15796 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node15799 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node15802 = (inp[12]) ? 4'b1000 : node15803;
														assign node15803 = (inp[10]) ? node15807 : node15804;
															assign node15804 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node15807 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node15811 = (inp[13]) ? node15813 : 4'b1101;
													assign node15813 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node15816 = (inp[13]) ? node15852 : node15817;
												assign node15817 = (inp[7]) ? node15837 : node15818;
													assign node15818 = (inp[14]) ? node15830 : node15819;
														assign node15819 = (inp[2]) ? node15825 : node15820;
															assign node15820 = (inp[12]) ? 4'b0000 : node15821;
																assign node15821 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15825 = (inp[12]) ? node15827 : 4'b0000;
																assign node15827 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node15830 = (inp[12]) ? node15834 : node15831;
															assign node15831 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15834 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node15837 = (inp[2]) ? node15847 : node15838;
														assign node15838 = (inp[14]) ? node15844 : node15839;
															assign node15839 = (inp[12]) ? 4'b1100 : node15840;
																assign node15840 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node15844 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node15847 = (inp[10]) ? node15849 : 4'b1101;
															assign node15849 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node15852 = (inp[2]) ? node15862 : node15853;
													assign node15853 = (inp[10]) ? 4'b0001 : node15854;
														assign node15854 = (inp[7]) ? node15858 : node15855;
															assign node15855 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node15858 = (inp[12]) ? 4'b1100 : 4'b0000;
													assign node15862 = (inp[12]) ? node15866 : node15863;
														assign node15863 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node15866 = (inp[7]) ? node15870 : node15867;
															assign node15867 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node15870 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node15873 = (inp[13]) ? node15965 : node15874;
										assign node15874 = (inp[12]) ? node15926 : node15875;
											assign node15875 = (inp[10]) ? node15903 : node15876;
												assign node15876 = (inp[3]) ? node15886 : node15877;
													assign node15877 = (inp[7]) ? node15883 : node15878;
														assign node15878 = (inp[2]) ? 4'b0100 : node15879;
															assign node15879 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node15883 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node15886 = (inp[7]) ? node15892 : node15887;
														assign node15887 = (inp[4]) ? 4'b0000 : node15888;
															assign node15888 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node15892 = (inp[14]) ? node15898 : node15893;
															assign node15893 = (inp[2]) ? node15895 : 4'b0100;
																assign node15895 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node15898 = (inp[4]) ? 4'b0000 : node15899;
																assign node15899 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node15903 = (inp[3]) ? node15913 : node15904;
													assign node15904 = (inp[4]) ? node15908 : node15905;
														assign node15905 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15908 = (inp[2]) ? 4'b0100 : node15909;
															assign node15909 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node15913 = (inp[7]) ? node15921 : node15914;
														assign node15914 = (inp[4]) ? node15918 : node15915;
															assign node15915 = (inp[2]) ? 4'b0000 : 4'b1100;
															assign node15918 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node15921 = (inp[2]) ? 4'b0100 : node15922;
															assign node15922 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node15926 = (inp[10]) ? node15944 : node15927;
												assign node15927 = (inp[3]) ? node15937 : node15928;
													assign node15928 = (inp[4]) ? node15930 : 4'b1000;
														assign node15930 = (inp[2]) ? node15934 : node15931;
															assign node15931 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node15934 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node15937 = (inp[7]) ? 4'b1100 : node15938;
														assign node15938 = (inp[4]) ? 4'b0000 : node15939;
															assign node15939 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node15944 = (inp[7]) ? node15956 : node15945;
													assign node15945 = (inp[4]) ? node15951 : node15946;
														assign node15946 = (inp[3]) ? node15948 : 4'b0100;
															assign node15948 = (inp[2]) ? 4'b0000 : 4'b1100;
														assign node15951 = (inp[3]) ? 4'b1000 : node15952;
															assign node15952 = (inp[2]) ? 4'b0100 : 4'b1000;
													assign node15956 = (inp[4]) ? node15960 : node15957;
														assign node15957 = (inp[3]) ? 4'b0100 : 4'b0000;
														assign node15960 = (inp[3]) ? node15962 : 4'b0100;
															assign node15962 = (inp[2]) ? 4'b0000 : 4'b1100;
										assign node15965 = (inp[10]) ? node15999 : node15966;
											assign node15966 = (inp[4]) ? node15986 : node15967;
												assign node15967 = (inp[12]) ? node15983 : node15968;
													assign node15968 = (inp[2]) ? node15972 : node15969;
														assign node15969 = (inp[3]) ? 4'b0100 : 4'b1100;
														assign node15972 = (inp[14]) ? node15978 : node15973;
															assign node15973 = (inp[3]) ? node15975 : 4'b1000;
																assign node15975 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node15978 = (inp[3]) ? 4'b1100 : node15979;
																assign node15979 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node15983 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node15986 = (inp[2]) ? node15994 : node15987;
													assign node15987 = (inp[3]) ? node15989 : 4'b0000;
														assign node15989 = (inp[12]) ? node15991 : 4'b0000;
															assign node15991 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node15994 = (inp[3]) ? 4'b0000 : node15995;
														assign node15995 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node15999 = (inp[4]) ? node16009 : node16000;
												assign node16000 = (inp[7]) ? node16006 : node16001;
													assign node16001 = (inp[3]) ? node16003 : 4'b1100;
														assign node16003 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node16006 = (inp[3]) ? 4'b1100 : 4'b1000;
												assign node16009 = (inp[3]) ? 4'b1000 : node16010;
													assign node16010 = (inp[2]) ? 4'b1100 : 4'b1000;
							assign node16014 = (inp[3]) ? node16396 : node16015;
								assign node16015 = (inp[11]) ? node16243 : node16016;
									assign node16016 = (inp[4]) ? node16114 : node16017;
										assign node16017 = (inp[2]) ? node16077 : node16018;
											assign node16018 = (inp[13]) ? node16054 : node16019;
												assign node16019 = (inp[7]) ? node16037 : node16020;
													assign node16020 = (inp[1]) ? node16032 : node16021;
														assign node16021 = (inp[14]) ? node16027 : node16022;
															assign node16022 = (inp[12]) ? 4'b1000 : node16023;
																assign node16023 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node16027 = (inp[10]) ? node16029 : 4'b1001;
																assign node16029 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node16032 = (inp[14]) ? 4'b0100 : node16033;
															assign node16033 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node16037 = (inp[14]) ? node16045 : node16038;
														assign node16038 = (inp[1]) ? node16042 : node16039;
															assign node16039 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node16042 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node16045 = (inp[1]) ? node16051 : node16046;
															assign node16046 = (inp[12]) ? node16048 : 4'b1001;
																assign node16048 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node16051 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node16054 = (inp[7]) ? node16064 : node16055;
													assign node16055 = (inp[12]) ? node16059 : node16056;
														assign node16056 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node16059 = (inp[1]) ? 4'b0000 : node16060;
															assign node16060 = (inp[10]) ? 4'b1000 : 4'b0100;
													assign node16064 = (inp[10]) ? node16070 : node16065;
														assign node16065 = (inp[1]) ? 4'b1101 : node16066;
															assign node16066 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node16070 = (inp[12]) ? node16074 : node16071;
															assign node16071 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node16074 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node16077 = (inp[10]) ? node16089 : node16078;
												assign node16078 = (inp[12]) ? 4'b1001 : node16079;
													assign node16079 = (inp[1]) ? node16083 : node16080;
														assign node16080 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node16083 = (inp[14]) ? 4'b0101 : node16084;
															assign node16084 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node16089 = (inp[1]) ? node16103 : node16090;
													assign node16090 = (inp[14]) ? node16096 : node16091;
														assign node16091 = (inp[7]) ? node16093 : 4'b0000;
															assign node16093 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node16096 = (inp[12]) ? 4'b0101 : node16097;
															assign node16097 = (inp[7]) ? 4'b0101 : node16098;
																assign node16098 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node16103 = (inp[12]) ? node16109 : node16104;
														assign node16104 = (inp[7]) ? 4'b1001 : node16105;
															assign node16105 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node16109 = (inp[13]) ? 4'b0000 : node16110;
															assign node16110 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node16114 = (inp[7]) ? node16178 : node16115;
											assign node16115 = (inp[10]) ? node16149 : node16116;
												assign node16116 = (inp[2]) ? node16130 : node16117;
													assign node16117 = (inp[1]) ? node16125 : node16118;
														assign node16118 = (inp[12]) ? node16122 : node16119;
															assign node16119 = (inp[13]) ? 4'b1001 : 4'b0100;
															assign node16122 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node16125 = (inp[12]) ? 4'b0100 : node16126;
															assign node16126 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node16130 = (inp[13]) ? node16140 : node16131;
														assign node16131 = (inp[1]) ? node16137 : node16132;
															assign node16132 = (inp[14]) ? 4'b1001 : node16133;
																assign node16133 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node16137 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node16140 = (inp[1]) ? node16146 : node16141;
															assign node16141 = (inp[12]) ? node16143 : 4'b0000;
																assign node16143 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node16146 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node16149 = (inp[2]) ? node16163 : node16150;
													assign node16150 = (inp[13]) ? node16160 : node16151;
														assign node16151 = (inp[1]) ? node16155 : node16152;
															assign node16152 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node16155 = (inp[14]) ? 4'b1001 : node16156;
																assign node16156 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16160 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16163 = (inp[13]) ? node16171 : node16164;
														assign node16164 = (inp[12]) ? node16168 : node16165;
															assign node16165 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node16168 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node16171 = (inp[1]) ? node16175 : node16172;
															assign node16172 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node16175 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node16178 = (inp[1]) ? node16208 : node16179;
												assign node16179 = (inp[13]) ? node16191 : node16180;
													assign node16180 = (inp[2]) ? node16184 : node16181;
														assign node16181 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node16184 = (inp[10]) ? node16186 : 4'b1101;
															assign node16186 = (inp[14]) ? node16188 : 4'b1000;
																assign node16188 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16191 = (inp[14]) ? node16197 : node16192;
														assign node16192 = (inp[10]) ? 4'b1001 : node16193;
															assign node16193 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16197 = (inp[2]) ? node16203 : node16198;
															assign node16198 = (inp[12]) ? node16200 : 4'b1000;
																assign node16200 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node16203 = (inp[12]) ? node16205 : 4'b0000;
																assign node16205 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node16208 = (inp[13]) ? node16230 : node16209;
													assign node16209 = (inp[14]) ? node16219 : node16210;
														assign node16210 = (inp[2]) ? node16214 : node16211;
															assign node16211 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node16214 = (inp[12]) ? node16216 : 4'b0001;
																assign node16216 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node16219 = (inp[10]) ? node16225 : node16220;
															assign node16220 = (inp[12]) ? 4'b0000 : node16221;
																assign node16221 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node16225 = (inp[2]) ? node16227 : 4'b1100;
																assign node16227 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node16230 = (inp[2]) ? node16240 : node16231;
														assign node16231 = (inp[14]) ? node16235 : node16232;
															assign node16232 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node16235 = (inp[12]) ? node16237 : 4'b0001;
																assign node16237 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node16240 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node16243 = (inp[1]) ? node16327 : node16244;
										assign node16244 = (inp[13]) ? node16290 : node16245;
											assign node16245 = (inp[7]) ? node16271 : node16246;
												assign node16246 = (inp[4]) ? node16260 : node16247;
													assign node16247 = (inp[2]) ? node16253 : node16248;
														assign node16248 = (inp[10]) ? 4'b1101 : node16249;
															assign node16249 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node16253 = (inp[10]) ? node16257 : node16254;
															assign node16254 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node16257 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node16260 = (inp[2]) ? node16266 : node16261;
														assign node16261 = (inp[10]) ? node16263 : 4'b0100;
															assign node16263 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16266 = (inp[12]) ? 4'b1001 : node16267;
															assign node16267 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node16271 = (inp[4]) ? node16281 : node16272;
													assign node16272 = (inp[2]) ? node16276 : node16273;
														assign node16273 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16276 = (inp[12]) ? node16278 : 4'b1000;
															assign node16278 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node16281 = (inp[2]) ? node16285 : node16282;
														assign node16282 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node16285 = (inp[10]) ? 4'b1001 : node16286;
															assign node16286 = (inp[12]) ? 4'b1100 : 4'b0001;
											assign node16290 = (inp[4]) ? node16310 : node16291;
												assign node16291 = (inp[10]) ? node16305 : node16292;
													assign node16292 = (inp[7]) ? node16298 : node16293;
														assign node16293 = (inp[2]) ? node16295 : 4'b0000;
															assign node16295 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node16298 = (inp[2]) ? node16302 : node16299;
															assign node16299 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node16302 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node16305 = (inp[2]) ? node16307 : 4'b0000;
														assign node16307 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node16310 = (inp[10]) ? node16320 : node16311;
													assign node16311 = (inp[7]) ? node16315 : node16312;
														assign node16312 = (inp[2]) ? 4'b0000 : 4'b1001;
														assign node16315 = (inp[12]) ? node16317 : 4'b1001;
															assign node16317 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node16320 = (inp[2]) ? 4'b0000 : node16321;
														assign node16321 = (inp[12]) ? node16323 : 4'b0000;
															assign node16323 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node16327 = (inp[13]) ? node16363 : node16328;
											assign node16328 = (inp[7]) ? node16346 : node16329;
												assign node16329 = (inp[4]) ? node16335 : node16330;
													assign node16330 = (inp[10]) ? node16332 : 4'b0100;
														assign node16332 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node16335 = (inp[10]) ? node16343 : node16336;
														assign node16336 = (inp[2]) ? node16340 : node16337;
															assign node16337 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node16340 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16343 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node16346 = (inp[10]) ? node16358 : node16347;
													assign node16347 = (inp[12]) ? node16353 : node16348;
														assign node16348 = (inp[2]) ? node16350 : 4'b1000;
															assign node16350 = (inp[4]) ? 4'b1000 : 4'b0000;
														assign node16353 = (inp[4]) ? node16355 : 4'b0000;
															assign node16355 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node16358 = (inp[4]) ? 4'b0000 : node16359;
														assign node16359 = (inp[2]) ? 4'b1000 : 4'b0100;
											assign node16363 = (inp[10]) ? node16389 : node16364;
												assign node16364 = (inp[7]) ? node16376 : node16365;
													assign node16365 = (inp[14]) ? node16371 : node16366;
														assign node16366 = (inp[2]) ? 4'b1000 : node16367;
															assign node16367 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node16371 = (inp[4]) ? 4'b0000 : node16372;
															assign node16372 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node16376 = (inp[4]) ? node16382 : node16377;
														assign node16377 = (inp[12]) ? node16379 : 4'b0100;
															assign node16379 = (inp[14]) ? 4'b1100 : 4'b0100;
														assign node16382 = (inp[2]) ? node16386 : node16383;
															assign node16383 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node16386 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node16389 = (inp[7]) ? node16391 : 4'b1000;
													assign node16391 = (inp[2]) ? node16393 : 4'b1000;
														assign node16393 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node16396 = (inp[4]) ? node16554 : node16397;
									assign node16397 = (inp[1]) ? node16481 : node16398;
										assign node16398 = (inp[11]) ? node16442 : node16399;
											assign node16399 = (inp[2]) ? node16421 : node16400;
												assign node16400 = (inp[7]) ? node16410 : node16401;
													assign node16401 = (inp[13]) ? node16403 : 4'b0000;
														assign node16403 = (inp[14]) ? node16407 : node16404;
															assign node16404 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node16407 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node16410 = (inp[10]) ? node16416 : node16411;
														assign node16411 = (inp[13]) ? 4'b0000 : node16412;
															assign node16412 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16416 = (inp[13]) ? 4'b1001 : node16417;
															assign node16417 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node16421 = (inp[12]) ? node16433 : node16422;
													assign node16422 = (inp[13]) ? node16430 : node16423;
														assign node16423 = (inp[14]) ? 4'b0000 : node16424;
															assign node16424 = (inp[7]) ? node16426 : 4'b0001;
																assign node16426 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node16430 = (inp[10]) ? 4'b1000 : 4'b0001;
													assign node16433 = (inp[10]) ? node16439 : node16434;
														assign node16434 = (inp[13]) ? node16436 : 4'b1000;
															assign node16436 = (inp[14]) ? 4'b0000 : 4'b1001;
														assign node16439 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node16442 = (inp[10]) ? node16464 : node16443;
												assign node16443 = (inp[7]) ? node16451 : node16444;
													assign node16444 = (inp[13]) ? node16446 : 4'b0001;
														assign node16446 = (inp[2]) ? node16448 : 4'b0001;
															assign node16448 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node16451 = (inp[12]) ? node16459 : node16452;
														assign node16452 = (inp[2]) ? node16456 : node16453;
															assign node16453 = (inp[13]) ? 4'b0001 : 4'b1000;
															assign node16456 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node16459 = (inp[2]) ? 4'b0000 : node16460;
															assign node16460 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node16464 = (inp[7]) ? node16474 : node16465;
													assign node16465 = (inp[13]) ? node16471 : node16466;
														assign node16466 = (inp[2]) ? node16468 : 4'b1000;
															assign node16468 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node16471 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node16474 = (inp[2]) ? node16476 : 4'b0001;
														assign node16476 = (inp[13]) ? 4'b1001 : node16477;
															assign node16477 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node16481 = (inp[11]) ? node16527 : node16482;
											assign node16482 = (inp[10]) ? node16516 : node16483;
												assign node16483 = (inp[13]) ? node16503 : node16484;
													assign node16484 = (inp[2]) ? node16494 : node16485;
														assign node16485 = (inp[12]) ? node16489 : node16486;
															assign node16486 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16489 = (inp[14]) ? node16491 : 4'b1001;
																assign node16491 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node16494 = (inp[12]) ? node16500 : node16495;
															assign node16495 = (inp[14]) ? node16497 : 4'b1000;
																assign node16497 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node16500 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node16503 = (inp[12]) ? node16511 : node16504;
														assign node16504 = (inp[2]) ? node16506 : 4'b1001;
															assign node16506 = (inp[14]) ? node16508 : 4'b1001;
																assign node16508 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node16511 = (inp[7]) ? node16513 : 4'b0001;
															assign node16513 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node16516 = (inp[2]) ? node16522 : node16517;
													assign node16517 = (inp[12]) ? node16519 : 4'b0000;
														assign node16519 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node16522 = (inp[13]) ? 4'b0000 : node16523;
														assign node16523 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node16527 = (inp[10]) ? node16545 : node16528;
												assign node16528 = (inp[13]) ? node16536 : node16529;
													assign node16529 = (inp[2]) ? node16533 : node16530;
														assign node16530 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16533 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node16536 = (inp[7]) ? 4'b0000 : node16537;
														assign node16537 = (inp[14]) ? 4'b1000 : node16538;
															assign node16538 = (inp[2]) ? node16540 : 4'b0000;
																assign node16540 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node16545 = (inp[13]) ? 4'b1000 : node16546;
													assign node16546 = (inp[2]) ? node16550 : node16547;
														assign node16547 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node16550 = (inp[7]) ? 4'b0000 : 4'b1000;
									assign node16554 = (inp[13]) ? node16648 : node16555;
										assign node16555 = (inp[10]) ? node16613 : node16556;
											assign node16556 = (inp[1]) ? node16580 : node16557;
												assign node16557 = (inp[11]) ? node16567 : node16558;
													assign node16558 = (inp[12]) ? node16562 : node16559;
														assign node16559 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node16562 = (inp[7]) ? node16564 : 4'b0001;
															assign node16564 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node16567 = (inp[7]) ? node16573 : node16568;
														assign node16568 = (inp[2]) ? 4'b1000 : node16569;
															assign node16569 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16573 = (inp[2]) ? node16577 : node16574;
															assign node16574 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node16577 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node16580 = (inp[11]) ? node16602 : node16581;
													assign node16581 = (inp[7]) ? node16591 : node16582;
														assign node16582 = (inp[14]) ? node16586 : node16583;
															assign node16583 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node16586 = (inp[12]) ? 4'b1000 : node16587;
																assign node16587 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node16591 = (inp[12]) ? node16597 : node16592;
															assign node16592 = (inp[14]) ? node16594 : 4'b1001;
																assign node16594 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node16597 = (inp[2]) ? 4'b0001 : node16598;
																assign node16598 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node16602 = (inp[12]) ? node16608 : node16603;
														assign node16603 = (inp[2]) ? node16605 : 4'b0000;
															assign node16605 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node16608 = (inp[2]) ? node16610 : 4'b1000;
															assign node16610 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node16613 = (inp[11]) ? node16641 : node16614;
												assign node16614 = (inp[2]) ? node16622 : node16615;
													assign node16615 = (inp[7]) ? 4'b0001 : node16616;
														assign node16616 = (inp[1]) ? 4'b0000 : node16617;
															assign node16617 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node16622 = (inp[7]) ? node16632 : node16623;
														assign node16623 = (inp[12]) ? node16629 : node16624;
															assign node16624 = (inp[14]) ? 4'b0001 : node16625;
																assign node16625 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node16629 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node16632 = (inp[12]) ? node16636 : node16633;
															assign node16633 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node16636 = (inp[14]) ? 4'b0000 : node16637;
																assign node16637 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node16641 = (inp[1]) ? 4'b0000 : node16642;
													assign node16642 = (inp[7]) ? 4'b0000 : node16643;
														assign node16643 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node16648 = (inp[12]) ? node16662 : node16649;
											assign node16649 = (inp[1]) ? 4'b0000 : node16650;
												assign node16650 = (inp[11]) ? 4'b0000 : node16651;
													assign node16651 = (inp[7]) ? 4'b0000 : node16652;
														assign node16652 = (inp[10]) ? node16656 : node16653;
															assign node16653 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node16656 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node16662 = (inp[10]) ? node16694 : node16663;
												assign node16663 = (inp[14]) ? node16683 : node16664;
													assign node16664 = (inp[7]) ? node16676 : node16665;
														assign node16665 = (inp[11]) ? node16671 : node16666;
															assign node16666 = (inp[1]) ? 4'b0001 : node16667;
																assign node16667 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node16671 = (inp[1]) ? 4'b0000 : node16672;
																assign node16672 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node16676 = (inp[1]) ? node16680 : node16677;
															assign node16677 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node16680 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node16683 = (inp[1]) ? 4'b0000 : node16684;
														assign node16684 = (inp[7]) ? node16686 : 4'b0000;
															assign node16686 = (inp[11]) ? node16690 : node16687;
																assign node16687 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node16690 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node16694 = (inp[14]) ? node16696 : 4'b0000;
													assign node16696 = (inp[11]) ? 4'b0000 : node16697;
														assign node16697 = (inp[2]) ? node16699 : 4'b0001;
															assign node16699 = (inp[7]) ? 4'b0000 : 4'b0001;
					assign node16703 = (inp[6]) ? node16705 : 4'b1000;
						assign node16705 = (inp[2]) ? node17209 : node16706;
							assign node16706 = (inp[5]) ? node16830 : node16707;
								assign node16707 = (inp[3]) ? node16709 : 4'b1000;
									assign node16709 = (inp[4]) ? node16757 : node16710;
										assign node16710 = (inp[7]) ? 4'b1000 : node16711;
											assign node16711 = (inp[1]) ? node16729 : node16712;
												assign node16712 = (inp[13]) ? node16716 : node16713;
													assign node16713 = (inp[10]) ? 4'b0001 : 4'b1000;
													assign node16716 = (inp[12]) ? node16724 : node16717;
														assign node16717 = (inp[10]) ? node16719 : 4'b0000;
															assign node16719 = (inp[11]) ? 4'b1001 : node16720;
																assign node16720 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node16724 = (inp[14]) ? node16726 : 4'b0001;
															assign node16726 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node16729 = (inp[14]) ? node16741 : node16730;
													assign node16730 = (inp[13]) ? node16736 : node16731;
														assign node16731 = (inp[12]) ? node16733 : 4'b0000;
															assign node16733 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node16736 = (inp[10]) ? 4'b1000 : node16737;
															assign node16737 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16741 = (inp[11]) ? node16747 : node16742;
														assign node16742 = (inp[13]) ? 4'b0001 : node16743;
															assign node16743 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node16747 = (inp[12]) ? node16751 : node16748;
															assign node16748 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node16751 = (inp[13]) ? 4'b0000 : node16752;
																assign node16752 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node16757 = (inp[1]) ? node16795 : node16758;
											assign node16758 = (inp[13]) ? node16778 : node16759;
												assign node16759 = (inp[7]) ? node16773 : node16760;
													assign node16760 = (inp[10]) ? node16766 : node16761;
														assign node16761 = (inp[14]) ? node16763 : 4'b1001;
															assign node16763 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node16766 = (inp[12]) ? node16768 : 4'b0001;
															assign node16768 = (inp[14]) ? node16770 : 4'b1001;
																assign node16770 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16773 = (inp[12]) ? 4'b1000 : node16774;
														assign node16774 = (inp[10]) ? 4'b0001 : 4'b1000;
												assign node16778 = (inp[14]) ? node16784 : node16779;
													assign node16779 = (inp[12]) ? 4'b0001 : node16780;
														assign node16780 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node16784 = (inp[11]) ? node16790 : node16785;
														assign node16785 = (inp[10]) ? node16787 : 4'b0000;
															assign node16787 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node16790 = (inp[12]) ? 4'b0001 : node16791;
															assign node16791 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node16795 = (inp[11]) ? node16819 : node16796;
												assign node16796 = (inp[14]) ? node16806 : node16797;
													assign node16797 = (inp[10]) ? node16803 : node16798;
														assign node16798 = (inp[13]) ? 4'b0000 : node16799;
															assign node16799 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16803 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node16806 = (inp[13]) ? node16814 : node16807;
														assign node16807 = (inp[12]) ? node16811 : node16808;
															assign node16808 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node16811 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node16814 = (inp[10]) ? node16816 : 4'b0001;
															assign node16816 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node16819 = (inp[13]) ? node16825 : node16820;
													assign node16820 = (inp[12]) ? node16822 : 4'b0000;
														assign node16822 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node16825 = (inp[12]) ? node16827 : 4'b1000;
														assign node16827 = (inp[10]) ? 4'b1000 : 4'b0000;
								assign node16830 = (inp[3]) ? node17034 : node16831;
									assign node16831 = (inp[1]) ? node16929 : node16832;
										assign node16832 = (inp[13]) ? node16876 : node16833;
											assign node16833 = (inp[10]) ? node16847 : node16834;
												assign node16834 = (inp[14]) ? node16840 : node16835;
													assign node16835 = (inp[7]) ? 4'b1001 : node16836;
														assign node16836 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node16840 = (inp[11]) ? 4'b1001 : node16841;
														assign node16841 = (inp[12]) ? node16843 : 4'b1000;
															assign node16843 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node16847 = (inp[12]) ? node16865 : node16848;
													assign node16848 = (inp[11]) ? node16856 : node16849;
														assign node16849 = (inp[14]) ? 4'b0000 : node16850;
															assign node16850 = (inp[7]) ? node16852 : 4'b0001;
																assign node16852 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node16856 = (inp[14]) ? 4'b0101 : node16857;
															assign node16857 = (inp[7]) ? node16861 : node16858;
																assign node16858 = (inp[4]) ? 4'b1000 : 4'b0101;
																assign node16861 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16865 = (inp[14]) ? node16867 : 4'b1001;
														assign node16867 = (inp[7]) ? node16873 : node16868;
															assign node16868 = (inp[4]) ? node16870 : 4'b1001;
																assign node16870 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node16873 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node16876 = (inp[4]) ? node16900 : node16877;
												assign node16877 = (inp[7]) ? node16885 : node16878;
													assign node16878 = (inp[11]) ? node16880 : 4'b1101;
														assign node16880 = (inp[10]) ? node16882 : 4'b0101;
															assign node16882 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node16885 = (inp[14]) ? node16891 : node16886;
														assign node16886 = (inp[12]) ? 4'b0001 : node16887;
															assign node16887 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node16891 = (inp[11]) ? node16897 : node16892;
															assign node16892 = (inp[10]) ? node16894 : 4'b0000;
																assign node16894 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node16897 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node16900 = (inp[11]) ? node16908 : node16901;
													assign node16901 = (inp[10]) ? 4'b0001 : node16902;
														assign node16902 = (inp[7]) ? node16904 : 4'b1001;
															assign node16904 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node16908 = (inp[7]) ? node16922 : node16909;
														assign node16909 = (inp[14]) ? node16915 : node16910;
															assign node16910 = (inp[12]) ? node16912 : 4'b1000;
																assign node16912 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node16915 = (inp[10]) ? node16919 : node16916;
																assign node16916 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node16919 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16922 = (inp[10]) ? node16926 : node16923;
															assign node16923 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node16926 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node16929 = (inp[11]) ? node16989 : node16930;
											assign node16930 = (inp[14]) ? node16962 : node16931;
												assign node16931 = (inp[4]) ? node16951 : node16932;
													assign node16932 = (inp[7]) ? node16942 : node16933;
														assign node16933 = (inp[13]) ? node16937 : node16934;
															assign node16934 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node16937 = (inp[10]) ? 4'b1100 : node16938;
																assign node16938 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node16942 = (inp[12]) ? node16946 : node16943;
															assign node16943 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node16946 = (inp[10]) ? 4'b1000 : node16947;
																assign node16947 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node16951 = (inp[10]) ? 4'b1001 : node16952;
														assign node16952 = (inp[12]) ? node16956 : node16953;
															assign node16953 = (inp[7]) ? 4'b0100 : 4'b0001;
															assign node16956 = (inp[13]) ? 4'b0100 : node16957;
																assign node16957 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node16962 = (inp[13]) ? node16974 : node16963;
													assign node16963 = (inp[12]) ? 4'b1001 : node16964;
														assign node16964 = (inp[10]) ? node16970 : node16965;
															assign node16965 = (inp[4]) ? node16967 : 4'b1001;
																assign node16967 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node16970 = (inp[4]) ? 4'b1001 : 4'b0001;
													assign node16974 = (inp[7]) ? node16984 : node16975;
														assign node16975 = (inp[4]) ? node16979 : node16976;
															assign node16976 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node16979 = (inp[12]) ? 4'b1001 : node16980;
																assign node16980 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node16984 = (inp[10]) ? 4'b0001 : node16985;
															assign node16985 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node16989 = (inp[12]) ? node17013 : node16990;
												assign node16990 = (inp[13]) ? node17006 : node16991;
													assign node16991 = (inp[10]) ? node16999 : node16992;
														assign node16992 = (inp[4]) ? node16996 : node16993;
															assign node16993 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node16996 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node16999 = (inp[14]) ? 4'b1000 : node17000;
															assign node17000 = (inp[7]) ? node17002 : 4'b0100;
																assign node17002 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node17006 = (inp[4]) ? node17010 : node17007;
														assign node17007 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node17010 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node17013 = (inp[10]) ? node17027 : node17014;
													assign node17014 = (inp[13]) ? node17022 : node17015;
														assign node17015 = (inp[14]) ? node17017 : 4'b0000;
															assign node17017 = (inp[4]) ? node17019 : 4'b1000;
																assign node17019 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17022 = (inp[4]) ? 4'b0000 : node17023;
															assign node17023 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node17027 = (inp[13]) ? 4'b1000 : node17028;
														assign node17028 = (inp[7]) ? node17030 : 4'b1000;
															assign node17030 = (inp[4]) ? 4'b0100 : 4'b0000;
									assign node17034 = (inp[4]) ? node17130 : node17035;
										assign node17035 = (inp[11]) ? node17085 : node17036;
											assign node17036 = (inp[13]) ? node17064 : node17037;
												assign node17037 = (inp[7]) ? node17057 : node17038;
													assign node17038 = (inp[12]) ? node17048 : node17039;
														assign node17039 = (inp[1]) ? node17045 : node17040;
															assign node17040 = (inp[14]) ? 4'b1001 : node17041;
																assign node17041 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node17045 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17048 = (inp[10]) ? node17050 : 4'b1001;
															assign node17050 = (inp[14]) ? node17054 : node17051;
																assign node17051 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node17054 = (inp[1]) ? 4'b1000 : 4'b0001;
													assign node17057 = (inp[10]) ? 4'b0001 : node17058;
														assign node17058 = (inp[14]) ? node17060 : 4'b1001;
															assign node17060 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node17064 = (inp[14]) ? node17072 : node17065;
													assign node17065 = (inp[12]) ? 4'b0000 : node17066;
														assign node17066 = (inp[1]) ? node17068 : 4'b0000;
															assign node17068 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node17072 = (inp[12]) ? node17080 : node17073;
														assign node17073 = (inp[1]) ? 4'b0001 : node17074;
															assign node17074 = (inp[7]) ? node17076 : 4'b0000;
																assign node17076 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node17080 = (inp[1]) ? node17082 : 4'b0001;
															assign node17082 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node17085 = (inp[1]) ? node17117 : node17086;
												assign node17086 = (inp[13]) ? node17100 : node17087;
													assign node17087 = (inp[7]) ? node17093 : node17088;
														assign node17088 = (inp[10]) ? 4'b1001 : node17089;
															assign node17089 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node17093 = (inp[14]) ? 4'b1000 : node17094;
															assign node17094 = (inp[10]) ? node17096 : 4'b0000;
																assign node17096 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17100 = (inp[14]) ? node17108 : node17101;
														assign node17101 = (inp[7]) ? node17105 : node17102;
															assign node17102 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node17105 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node17108 = (inp[7]) ? node17112 : node17109;
															assign node17109 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node17112 = (inp[10]) ? 4'b0000 : node17113;
																assign node17113 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node17117 = (inp[13]) ? node17125 : node17118;
													assign node17118 = (inp[10]) ? 4'b0000 : node17119;
														assign node17119 = (inp[7]) ? 4'b0000 : node17120;
															assign node17120 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17125 = (inp[7]) ? node17127 : 4'b1000;
														assign node17127 = (inp[14]) ? 4'b0000 : 4'b1000;
										assign node17130 = (inp[13]) ? node17178 : node17131;
											assign node17131 = (inp[1]) ? node17157 : node17132;
												assign node17132 = (inp[7]) ? node17144 : node17133;
													assign node17133 = (inp[11]) ? node17137 : node17134;
														assign node17134 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node17137 = (inp[10]) ? node17141 : node17138;
															assign node17138 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node17141 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node17144 = (inp[11]) ? 4'b0001 : node17145;
														assign node17145 = (inp[10]) ? node17151 : node17146;
															assign node17146 = (inp[12]) ? 4'b1000 : node17147;
																assign node17147 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17151 = (inp[14]) ? 4'b1001 : node17152;
																assign node17152 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node17157 = (inp[11]) ? node17171 : node17158;
													assign node17158 = (inp[10]) ? node17166 : node17159;
														assign node17159 = (inp[14]) ? node17161 : 4'b1000;
															assign node17161 = (inp[7]) ? node17163 : 4'b0000;
																assign node17163 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node17166 = (inp[7]) ? 4'b0000 : node17167;
															assign node17167 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node17171 = (inp[7]) ? 4'b0000 : node17172;
														assign node17172 = (inp[10]) ? 4'b0000 : node17173;
															assign node17173 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node17178 = (inp[11]) ? 4'b0000 : node17179;
												assign node17179 = (inp[10]) ? node17195 : node17180;
													assign node17180 = (inp[1]) ? node17186 : node17181;
														assign node17181 = (inp[7]) ? node17183 : 4'b0000;
															assign node17183 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node17186 = (inp[14]) ? node17190 : node17187;
															assign node17187 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node17190 = (inp[7]) ? node17192 : 4'b0001;
																assign node17192 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node17195 = (inp[1]) ? 4'b0000 : node17196;
														assign node17196 = (inp[12]) ? node17202 : node17197;
															assign node17197 = (inp[7]) ? 4'b0001 : node17198;
																assign node17198 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node17202 = (inp[7]) ? 4'b0000 : node17203;
																assign node17203 = (inp[14]) ? 4'b0000 : 4'b0001;
							assign node17209 = (inp[3]) ? node17211 : 4'b1000;
								assign node17211 = (inp[5]) ? node17213 : 4'b1000;
									assign node17213 = (inp[4]) ? node17263 : node17214;
										assign node17214 = (inp[7]) ? 4'b1000 : node17215;
											assign node17215 = (inp[1]) ? node17233 : node17216;
												assign node17216 = (inp[13]) ? node17224 : node17217;
													assign node17217 = (inp[10]) ? node17219 : 4'b1000;
														assign node17219 = (inp[12]) ? 4'b1000 : node17220;
															assign node17220 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17224 = (inp[11]) ? node17228 : node17225;
														assign node17225 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17228 = (inp[10]) ? node17230 : 4'b0001;
															assign node17230 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node17233 = (inp[12]) ? node17245 : node17234;
													assign node17234 = (inp[13]) ? node17240 : node17235;
														assign node17235 = (inp[11]) ? 4'b0000 : node17236;
															assign node17236 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node17240 = (inp[14]) ? node17242 : 4'b1000;
															assign node17242 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node17245 = (inp[11]) ? node17249 : node17246;
														assign node17246 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node17249 = (inp[14]) ? node17257 : node17250;
															assign node17250 = (inp[13]) ? node17254 : node17251;
																assign node17251 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node17254 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node17257 = (inp[10]) ? node17259 : 4'b0000;
																assign node17259 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node17263 = (inp[13]) ? node17307 : node17264;
											assign node17264 = (inp[10]) ? node17284 : node17265;
												assign node17265 = (inp[7]) ? node17279 : node17266;
													assign node17266 = (inp[12]) ? node17274 : node17267;
														assign node17267 = (inp[11]) ? 4'b0000 : node17268;
															assign node17268 = (inp[1]) ? 4'b0001 : node17269;
																assign node17269 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node17274 = (inp[14]) ? node17276 : 4'b1001;
															assign node17276 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node17279 = (inp[12]) ? 4'b1000 : node17280;
														assign node17280 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node17284 = (inp[11]) ? node17298 : node17285;
													assign node17285 = (inp[7]) ? node17293 : node17286;
														assign node17286 = (inp[12]) ? 4'b0001 : node17287;
															assign node17287 = (inp[14]) ? node17289 : 4'b0001;
																assign node17289 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node17293 = (inp[12]) ? 4'b1000 : node17294;
															assign node17294 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node17298 = (inp[1]) ? 4'b0000 : node17299;
														assign node17299 = (inp[12]) ? node17303 : node17300;
															assign node17300 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node17303 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node17307 = (inp[11]) ? node17335 : node17308;
												assign node17308 = (inp[10]) ? node17324 : node17309;
													assign node17309 = (inp[7]) ? node17315 : node17310;
														assign node17310 = (inp[14]) ? node17312 : 4'b0000;
															assign node17312 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node17315 = (inp[14]) ? node17321 : node17316;
															assign node17316 = (inp[1]) ? node17318 : 4'b0001;
																assign node17318 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node17321 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node17324 = (inp[1]) ? 4'b0000 : node17325;
														assign node17325 = (inp[12]) ? node17331 : node17326;
															assign node17326 = (inp[7]) ? 4'b0000 : node17327;
																assign node17327 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17331 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node17335 = (inp[1]) ? 4'b0000 : node17336;
													assign node17336 = (inp[10]) ? 4'b0000 : node17337;
														assign node17337 = (inp[7]) ? node17339 : 4'b0000;
															assign node17339 = (inp[12]) ? 4'b0001 : 4'b0000;
			assign node17344 = (inp[15]) ? node20358 : node17345;
				assign node17345 = (inp[6]) ? node18069 : node17346;
					assign node17346 = (inp[0]) ? 4'b0100 : node17347;
						assign node17347 = (inp[2]) ? node17799 : node17348;
							assign node17348 = (inp[3]) ? node17592 : node17349;
								assign node17349 = (inp[5]) ? node17441 : node17350;
									assign node17350 = (inp[7]) ? node17412 : node17351;
										assign node17351 = (inp[4]) ? node17373 : node17352;
											assign node17352 = (inp[13]) ? node17354 : 4'b0110;
												assign node17354 = (inp[12]) ? node17368 : node17355;
													assign node17355 = (inp[10]) ? node17359 : node17356;
														assign node17356 = (inp[1]) ? 4'b0000 : 4'b0110;
														assign node17359 = (inp[11]) ? node17365 : node17360;
															assign node17360 = (inp[14]) ? node17362 : 4'b0000;
																assign node17362 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node17365 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node17368 = (inp[1]) ? node17370 : 4'b0110;
														assign node17370 = (inp[10]) ? 4'b0000 : 4'b0110;
											assign node17373 = (inp[1]) ? node17397 : node17374;
												assign node17374 = (inp[11]) ? node17386 : node17375;
													assign node17375 = (inp[14]) ? node17381 : node17376;
														assign node17376 = (inp[13]) ? 4'b1001 : node17377;
															assign node17377 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node17381 = (inp[13]) ? 4'b1000 : node17382;
															assign node17382 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17386 = (inp[13]) ? node17392 : node17387;
														assign node17387 = (inp[12]) ? 4'b0001 : node17388;
															assign node17388 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node17392 = (inp[12]) ? 4'b1001 : node17393;
															assign node17393 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node17397 = (inp[14]) ? node17405 : node17398;
													assign node17398 = (inp[13]) ? 4'b0000 : node17399;
														assign node17399 = (inp[12]) ? node17401 : 4'b1000;
															assign node17401 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node17405 = (inp[11]) ? 4'b1000 : node17406;
														assign node17406 = (inp[13]) ? 4'b1001 : node17407;
															assign node17407 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node17412 = (inp[4]) ? node17414 : 4'b0110;
											assign node17414 = (inp[13]) ? node17416 : 4'b0110;
												assign node17416 = (inp[12]) ? node17432 : node17417;
													assign node17417 = (inp[10]) ? node17423 : node17418;
														assign node17418 = (inp[1]) ? node17420 : 4'b0110;
															assign node17420 = (inp[11]) ? 4'b0000 : 4'b0110;
														assign node17423 = (inp[11]) ? node17429 : node17424;
															assign node17424 = (inp[14]) ? node17426 : 4'b0000;
																assign node17426 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node17429 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node17432 = (inp[10]) ? node17434 : 4'b0110;
														assign node17434 = (inp[1]) ? node17436 : 4'b0110;
															assign node17436 = (inp[11]) ? 4'b0000 : node17437;
																assign node17437 = (inp[14]) ? 4'b0110 : 4'b0000;
									assign node17441 = (inp[1]) ? node17501 : node17442;
										assign node17442 = (inp[13]) ? node17466 : node17443;
											assign node17443 = (inp[12]) ? node17457 : node17444;
												assign node17444 = (inp[10]) ? node17450 : node17445;
													assign node17445 = (inp[14]) ? node17447 : 4'b0101;
														assign node17447 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node17450 = (inp[14]) ? node17452 : 4'b1101;
														assign node17452 = (inp[4]) ? node17454 : 4'b1101;
															assign node17454 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node17457 = (inp[4]) ? node17463 : node17458;
													assign node17458 = (inp[11]) ? 4'b0101 : node17459;
														assign node17459 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node17463 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node17466 = (inp[10]) ? node17482 : node17467;
												assign node17467 = (inp[14]) ? node17473 : node17468;
													assign node17468 = (inp[7]) ? 4'b1101 : node17469;
														assign node17469 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node17473 = (inp[11]) ? node17479 : node17474;
														assign node17474 = (inp[7]) ? 4'b1100 : node17475;
															assign node17475 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node17479 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node17482 = (inp[12]) ? node17494 : node17483;
													assign node17483 = (inp[4]) ? node17489 : node17484;
														assign node17484 = (inp[7]) ? 4'b0101 : node17485;
															assign node17485 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17489 = (inp[11]) ? 4'b0001 : node17490;
															assign node17490 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17494 = (inp[14]) ? node17496 : 4'b1101;
														assign node17496 = (inp[11]) ? node17498 : 4'b1100;
															assign node17498 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node17501 = (inp[4]) ? node17541 : node17502;
											assign node17502 = (inp[13]) ? node17520 : node17503;
												assign node17503 = (inp[10]) ? node17515 : node17504;
													assign node17504 = (inp[12]) ? node17510 : node17505;
														assign node17505 = (inp[14]) ? node17507 : 4'b1100;
															assign node17507 = (inp[11]) ? 4'b1100 : 4'b0101;
														assign node17510 = (inp[14]) ? node17512 : 4'b0100;
															assign node17512 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node17515 = (inp[14]) ? node17517 : 4'b1100;
														assign node17517 = (inp[7]) ? 4'b1100 : 4'b0101;
												assign node17520 = (inp[7]) ? node17528 : node17521;
													assign node17521 = (inp[12]) ? node17523 : 4'b0000;
														assign node17523 = (inp[10]) ? node17525 : 4'b1100;
															assign node17525 = (inp[11]) ? 4'b0000 : 4'b1101;
													assign node17528 = (inp[10]) ? 4'b0100 : node17529;
														assign node17529 = (inp[12]) ? node17535 : node17530;
															assign node17530 = (inp[14]) ? node17532 : 4'b0100;
																assign node17532 = (inp[11]) ? 4'b0100 : 4'b1101;
															assign node17535 = (inp[11]) ? 4'b1100 : node17536;
																assign node17536 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node17541 = (inp[7]) ? node17563 : node17542;
												assign node17542 = (inp[11]) ? node17552 : node17543;
													assign node17543 = (inp[14]) ? node17547 : node17544;
														assign node17544 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node17547 = (inp[12]) ? node17549 : 4'b1001;
															assign node17549 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node17552 = (inp[13]) ? node17558 : node17553;
														assign node17553 = (inp[12]) ? node17555 : 4'b1000;
															assign node17555 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17558 = (inp[12]) ? node17560 : 4'b0000;
															assign node17560 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node17563 = (inp[13]) ? node17577 : node17564;
													assign node17564 = (inp[12]) ? node17570 : node17565;
														assign node17565 = (inp[11]) ? 4'b1100 : node17566;
															assign node17566 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node17570 = (inp[10]) ? node17572 : 4'b0100;
															assign node17572 = (inp[14]) ? node17574 : 4'b1100;
																assign node17574 = (inp[11]) ? 4'b1100 : 4'b0101;
													assign node17577 = (inp[10]) ? node17585 : node17578;
														assign node17578 = (inp[12]) ? 4'b1100 : node17579;
															assign node17579 = (inp[14]) ? node17581 : 4'b0000;
																assign node17581 = (inp[11]) ? 4'b0000 : 4'b1101;
														assign node17585 = (inp[14]) ? node17587 : 4'b0000;
															assign node17587 = (inp[11]) ? 4'b0000 : node17588;
																assign node17588 = (inp[12]) ? 4'b1101 : 4'b0001;
								assign node17592 = (inp[1]) ? node17688 : node17593;
									assign node17593 = (inp[13]) ? node17635 : node17594;
										assign node17594 = (inp[7]) ? node17622 : node17595;
											assign node17595 = (inp[4]) ? node17609 : node17596;
												assign node17596 = (inp[10]) ? node17602 : node17597;
													assign node17597 = (inp[14]) ? node17599 : 4'b0001;
														assign node17599 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node17602 = (inp[12]) ? 4'b0001 : node17603;
														assign node17603 = (inp[11]) ? 4'b1001 : node17604;
															assign node17604 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node17609 = (inp[10]) ? node17615 : node17610;
													assign node17610 = (inp[14]) ? node17612 : 4'b0101;
														assign node17612 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node17615 = (inp[12]) ? 4'b0101 : node17616;
														assign node17616 = (inp[14]) ? node17618 : 4'b1101;
															assign node17618 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node17622 = (inp[14]) ? node17628 : node17623;
												assign node17623 = (inp[12]) ? 4'b0001 : node17624;
													assign node17624 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node17628 = (inp[11]) ? node17630 : 4'b0000;
													assign node17630 = (inp[12]) ? 4'b0001 : node17631;
														assign node17631 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node17635 = (inp[7]) ? node17665 : node17636;
											assign node17636 = (inp[4]) ? node17648 : node17637;
												assign node17637 = (inp[12]) ? node17643 : node17638;
													assign node17638 = (inp[10]) ? 4'b0101 : node17639;
														assign node17639 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node17643 = (inp[14]) ? node17645 : 4'b1001;
														assign node17645 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node17648 = (inp[14]) ? node17654 : node17649;
													assign node17649 = (inp[12]) ? 4'b1101 : node17650;
														assign node17650 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node17654 = (inp[11]) ? node17660 : node17655;
														assign node17655 = (inp[12]) ? 4'b1100 : node17656;
															assign node17656 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node17660 = (inp[10]) ? node17662 : 4'b1101;
															assign node17662 = (inp[12]) ? 4'b1101 : 4'b0101;
											assign node17665 = (inp[11]) ? node17681 : node17666;
												assign node17666 = (inp[14]) ? node17674 : node17667;
													assign node17667 = (inp[12]) ? 4'b1001 : node17668;
														assign node17668 = (inp[10]) ? node17670 : 4'b1001;
															assign node17670 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node17674 = (inp[12]) ? 4'b1000 : node17675;
														assign node17675 = (inp[10]) ? node17677 : 4'b1000;
															assign node17677 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node17681 = (inp[10]) ? node17683 : 4'b1001;
													assign node17683 = (inp[12]) ? 4'b1001 : node17684;
														assign node17684 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node17688 = (inp[4]) ? node17734 : node17689;
										assign node17689 = (inp[11]) ? node17717 : node17690;
											assign node17690 = (inp[14]) ? node17704 : node17691;
												assign node17691 = (inp[13]) ? node17697 : node17692;
													assign node17692 = (inp[10]) ? 4'b1000 : node17693;
														assign node17693 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17697 = (inp[10]) ? node17701 : node17698;
														assign node17698 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node17701 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node17704 = (inp[13]) ? node17710 : node17705;
													assign node17705 = (inp[12]) ? 4'b0001 : node17706;
														assign node17706 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node17710 = (inp[10]) ? node17712 : 4'b1001;
														assign node17712 = (inp[12]) ? 4'b1001 : node17713;
															assign node17713 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node17717 = (inp[13]) ? node17723 : node17718;
												assign node17718 = (inp[10]) ? 4'b1000 : node17719;
													assign node17719 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node17723 = (inp[7]) ? node17729 : node17724;
													assign node17724 = (inp[12]) ? node17726 : 4'b0100;
														assign node17726 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node17729 = (inp[12]) ? node17731 : 4'b0000;
														assign node17731 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node17734 = (inp[7]) ? node17768 : node17735;
											assign node17735 = (inp[11]) ? node17757 : node17736;
												assign node17736 = (inp[14]) ? node17746 : node17737;
													assign node17737 = (inp[13]) ? node17741 : node17738;
														assign node17738 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node17741 = (inp[12]) ? node17743 : 4'b0100;
															assign node17743 = (inp[5]) ? 4'b0100 : 4'b1100;
													assign node17746 = (inp[13]) ? node17752 : node17747;
														assign node17747 = (inp[10]) ? node17749 : 4'b0101;
															assign node17749 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node17752 = (inp[10]) ? node17754 : 4'b1101;
															assign node17754 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node17757 = (inp[13]) ? node17763 : node17758;
													assign node17758 = (inp[12]) ? node17760 : 4'b1100;
														assign node17760 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node17763 = (inp[12]) ? node17765 : 4'b0100;
														assign node17765 = (inp[10]) ? 4'b0100 : 4'b1100;
											assign node17768 = (inp[13]) ? node17782 : node17769;
												assign node17769 = (inp[10]) ? node17777 : node17770;
													assign node17770 = (inp[12]) ? 4'b0000 : node17771;
														assign node17771 = (inp[14]) ? node17773 : 4'b1000;
															assign node17773 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node17777 = (inp[14]) ? node17779 : 4'b1000;
														assign node17779 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node17782 = (inp[12]) ? node17788 : node17783;
													assign node17783 = (inp[14]) ? node17785 : 4'b0100;
														assign node17785 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node17788 = (inp[10]) ? node17794 : node17789;
														assign node17789 = (inp[11]) ? 4'b1000 : node17790;
															assign node17790 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node17794 = (inp[14]) ? node17796 : 4'b0100;
															assign node17796 = (inp[11]) ? 4'b0100 : 4'b1001;
							assign node17799 = (inp[5]) ? node17801 : 4'b0110;
								assign node17801 = (inp[3]) ? node17897 : node17802;
									assign node17802 = (inp[4]) ? node17826 : node17803;
										assign node17803 = (inp[7]) ? 4'b0110 : node17804;
											assign node17804 = (inp[13]) ? node17806 : 4'b0110;
												assign node17806 = (inp[12]) ? node17820 : node17807;
													assign node17807 = (inp[10]) ? node17815 : node17808;
														assign node17808 = (inp[1]) ? node17810 : 4'b0110;
															assign node17810 = (inp[14]) ? node17812 : 4'b0000;
																assign node17812 = (inp[11]) ? 4'b0000 : 4'b0110;
														assign node17815 = (inp[1]) ? node17817 : 4'b0001;
															assign node17817 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node17820 = (inp[1]) ? node17822 : 4'b0110;
														assign node17822 = (inp[10]) ? 4'b0000 : 4'b0110;
										assign node17826 = (inp[7]) ? node17876 : node17827;
											assign node17827 = (inp[1]) ? node17853 : node17828;
												assign node17828 = (inp[11]) ? node17842 : node17829;
													assign node17829 = (inp[14]) ? node17833 : node17830;
														assign node17830 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node17833 = (inp[12]) ? 4'b0000 : node17834;
															assign node17834 = (inp[13]) ? node17838 : node17835;
																assign node17835 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node17838 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node17842 = (inp[13]) ? node17848 : node17843;
														assign node17843 = (inp[12]) ? 4'b0001 : node17844;
															assign node17844 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node17848 = (inp[10]) ? node17850 : 4'b1001;
															assign node17850 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node17853 = (inp[14]) ? node17865 : node17854;
													assign node17854 = (inp[13]) ? node17860 : node17855;
														assign node17855 = (inp[12]) ? node17857 : 4'b1000;
															assign node17857 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17860 = (inp[12]) ? node17862 : 4'b0000;
															assign node17862 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node17865 = (inp[11]) ? node17873 : node17866;
														assign node17866 = (inp[10]) ? node17868 : 4'b0001;
															assign node17868 = (inp[13]) ? node17870 : 4'b1001;
																assign node17870 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node17873 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node17876 = (inp[13]) ? node17878 : 4'b0110;
												assign node17878 = (inp[12]) ? node17892 : node17879;
													assign node17879 = (inp[10]) ? node17883 : node17880;
														assign node17880 = (inp[1]) ? 4'b0000 : 4'b0110;
														assign node17883 = (inp[14]) ? node17885 : 4'b0000;
															assign node17885 = (inp[1]) ? node17889 : node17886;
																assign node17886 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node17889 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node17892 = (inp[11]) ? node17894 : 4'b0110;
														assign node17894 = (inp[1]) ? 4'b0000 : 4'b0110;
									assign node17897 = (inp[4]) ? node17975 : node17898;
										assign node17898 = (inp[1]) ? node17938 : node17899;
											assign node17899 = (inp[14]) ? node17913 : node17900;
												assign node17900 = (inp[13]) ? node17906 : node17901;
													assign node17901 = (inp[10]) ? node17903 : 4'b0001;
														assign node17903 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node17906 = (inp[12]) ? 4'b1001 : node17907;
														assign node17907 = (inp[10]) ? node17909 : 4'b1001;
															assign node17909 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node17913 = (inp[11]) ? node17927 : node17914;
													assign node17914 = (inp[13]) ? node17920 : node17915;
														assign node17915 = (inp[12]) ? 4'b0000 : node17916;
															assign node17916 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17920 = (inp[10]) ? node17922 : 4'b1000;
															assign node17922 = (inp[12]) ? 4'b1000 : node17923;
																assign node17923 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node17927 = (inp[13]) ? node17933 : node17928;
														assign node17928 = (inp[10]) ? node17930 : 4'b0001;
															assign node17930 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node17933 = (inp[10]) ? node17935 : 4'b1001;
															assign node17935 = (inp[12]) ? 4'b1001 : 4'b0101;
											assign node17938 = (inp[11]) ? node17958 : node17939;
												assign node17939 = (inp[14]) ? node17947 : node17940;
													assign node17940 = (inp[10]) ? 4'b1000 : node17941;
														assign node17941 = (inp[12]) ? node17943 : 4'b0000;
															assign node17943 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node17947 = (inp[13]) ? node17953 : node17948;
														assign node17948 = (inp[12]) ? 4'b0001 : node17949;
															assign node17949 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node17953 = (inp[12]) ? 4'b1001 : node17954;
															assign node17954 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node17958 = (inp[13]) ? node17964 : node17959;
													assign node17959 = (inp[12]) ? node17961 : 4'b1000;
														assign node17961 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node17964 = (inp[7]) ? node17970 : node17965;
														assign node17965 = (inp[12]) ? node17967 : 4'b0100;
															assign node17967 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node17970 = (inp[10]) ? 4'b0000 : node17971;
															assign node17971 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node17975 = (inp[7]) ? node18027 : node17976;
											assign node17976 = (inp[1]) ? node17998 : node17977;
												assign node17977 = (inp[13]) ? node17989 : node17978;
													assign node17978 = (inp[10]) ? node17980 : 4'b0101;
														assign node17980 = (inp[12]) ? node17984 : node17981;
															assign node17981 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node17984 = (inp[14]) ? node17986 : 4'b0101;
																assign node17986 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node17989 = (inp[11]) ? node17993 : node17990;
														assign node17990 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node17993 = (inp[12]) ? 4'b1101 : node17994;
															assign node17994 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node17998 = (inp[11]) ? node18018 : node17999;
													assign node17999 = (inp[14]) ? node18009 : node18000;
														assign node18000 = (inp[13]) ? node18004 : node18001;
															assign node18001 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18004 = (inp[12]) ? node18006 : 4'b0100;
																assign node18006 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node18009 = (inp[10]) ? node18011 : 4'b1101;
															assign node18011 = (inp[12]) ? node18015 : node18012;
																assign node18012 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node18015 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node18018 = (inp[13]) ? node18022 : node18019;
														assign node18019 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node18022 = (inp[10]) ? 4'b0100 : node18023;
															assign node18023 = (inp[14]) ? 4'b0100 : 4'b1100;
											assign node18027 = (inp[1]) ? node18049 : node18028;
												assign node18028 = (inp[11]) ? node18038 : node18029;
													assign node18029 = (inp[14]) ? node18031 : 4'b1001;
														assign node18031 = (inp[13]) ? node18033 : 4'b0000;
															assign node18033 = (inp[10]) ? node18035 : 4'b1000;
																assign node18035 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node18038 = (inp[13]) ? node18044 : node18039;
														assign node18039 = (inp[12]) ? 4'b0001 : node18040;
															assign node18040 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18044 = (inp[10]) ? node18046 : 4'b1001;
															assign node18046 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node18049 = (inp[13]) ? node18059 : node18050;
													assign node18050 = (inp[12]) ? node18056 : node18051;
														assign node18051 = (inp[14]) ? node18053 : 4'b1000;
															assign node18053 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node18056 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18059 = (inp[12]) ? node18063 : node18060;
														assign node18060 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node18063 = (inp[14]) ? 4'b1001 : node18064;
															assign node18064 = (inp[10]) ? 4'b0100 : 4'b1000;
					assign node18069 = (inp[5]) ? node19025 : node18070;
						assign node18070 = (inp[0]) ? node18760 : node18071;
							assign node18071 = (inp[11]) ? node18475 : node18072;
								assign node18072 = (inp[3]) ? node18276 : node18073;
									assign node18073 = (inp[4]) ? node18181 : node18074;
										assign node18074 = (inp[7]) ? node18136 : node18075;
											assign node18075 = (inp[13]) ? node18101 : node18076;
												assign node18076 = (inp[10]) ? node18086 : node18077;
													assign node18077 = (inp[1]) ? node18081 : node18078;
														assign node18078 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node18081 = (inp[14]) ? 4'b0101 : node18082;
															assign node18082 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node18086 = (inp[12]) ? node18094 : node18087;
														assign node18087 = (inp[1]) ? node18091 : node18088;
															assign node18088 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node18091 = (inp[2]) ? 4'b1100 : 4'b0001;
														assign node18094 = (inp[14]) ? node18098 : node18095;
															assign node18095 = (inp[1]) ? 4'b1100 : 4'b0101;
															assign node18098 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node18101 = (inp[2]) ? node18111 : node18102;
													assign node18102 = (inp[10]) ? node18108 : node18103;
														assign node18103 = (inp[1]) ? node18105 : 4'b0001;
															assign node18105 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18108 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node18111 = (inp[12]) ? node18123 : node18112;
														assign node18112 = (inp[10]) ? node18118 : node18113;
															assign node18113 = (inp[14]) ? node18115 : 4'b0000;
																assign node18115 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node18118 = (inp[14]) ? 4'b0001 : node18119;
																assign node18119 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node18123 = (inp[10]) ? node18131 : node18124;
															assign node18124 = (inp[14]) ? node18128 : node18125;
																assign node18125 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node18128 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node18131 = (inp[1]) ? 4'b0000 : node18132;
																assign node18132 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node18136 = (inp[13]) ? node18160 : node18137;
												assign node18137 = (inp[10]) ? node18147 : node18138;
													assign node18138 = (inp[12]) ? 4'b0100 : node18139;
														assign node18139 = (inp[14]) ? node18143 : node18140;
															assign node18140 = (inp[1]) ? 4'b1100 : 4'b0101;
															assign node18143 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node18147 = (inp[12]) ? node18155 : node18148;
														assign node18148 = (inp[14]) ? node18152 : node18149;
															assign node18149 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node18152 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node18155 = (inp[14]) ? node18157 : 4'b1100;
															assign node18157 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node18160 = (inp[12]) ? node18172 : node18161;
													assign node18161 = (inp[2]) ? node18163 : 4'b0100;
														assign node18163 = (inp[10]) ? node18169 : node18164;
															assign node18164 = (inp[14]) ? node18166 : 4'b1101;
																assign node18166 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node18169 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node18172 = (inp[1]) ? node18176 : node18173;
														assign node18173 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node18176 = (inp[14]) ? 4'b1101 : node18177;
															assign node18177 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node18181 = (inp[2]) ? node18219 : node18182;
											assign node18182 = (inp[7]) ? node18206 : node18183;
												assign node18183 = (inp[13]) ? node18195 : node18184;
													assign node18184 = (inp[10]) ? node18190 : node18185;
														assign node18185 = (inp[12]) ? 4'b0001 : node18186;
															assign node18186 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node18190 = (inp[12]) ? 4'b1001 : node18191;
															assign node18191 = (inp[1]) ? 4'b0101 : 4'b1001;
													assign node18195 = (inp[10]) ? node18201 : node18196;
														assign node18196 = (inp[12]) ? 4'b0101 : node18197;
															assign node18197 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node18201 = (inp[12]) ? 4'b1101 : node18202;
															assign node18202 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node18206 = (inp[10]) ? node18212 : node18207;
													assign node18207 = (inp[1]) ? node18209 : 4'b0001;
														assign node18209 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node18212 = (inp[1]) ? node18214 : 4'b1001;
														assign node18214 = (inp[12]) ? 4'b1001 : node18215;
															assign node18215 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node18219 = (inp[7]) ? node18239 : node18220;
												assign node18220 = (inp[14]) ? node18226 : node18221;
													assign node18221 = (inp[1]) ? node18223 : 4'b0001;
														assign node18223 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node18226 = (inp[1]) ? node18230 : node18227;
														assign node18227 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18230 = (inp[12]) ? 4'b1001 : node18231;
															assign node18231 = (inp[10]) ? node18235 : node18232;
																assign node18232 = (inp[13]) ? 4'b1001 : 4'b0001;
																assign node18235 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node18239 = (inp[13]) ? node18257 : node18240;
													assign node18240 = (inp[10]) ? node18250 : node18241;
														assign node18241 = (inp[1]) ? node18245 : node18242;
															assign node18242 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node18245 = (inp[14]) ? 4'b0101 : node18246;
																assign node18246 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node18250 = (inp[14]) ? node18254 : node18251;
															assign node18251 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node18254 = (inp[12]) ? 4'b0101 : 4'b1100;
													assign node18257 = (inp[12]) ? node18265 : node18258;
														assign node18258 = (inp[1]) ? 4'b0000 : node18259;
															assign node18259 = (inp[10]) ? 4'b0000 : node18260;
																assign node18260 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node18265 = (inp[10]) ? node18271 : node18266;
															assign node18266 = (inp[1]) ? 4'b1101 : node18267;
																assign node18267 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node18271 = (inp[1]) ? node18273 : 4'b1101;
																assign node18273 = (inp[14]) ? 4'b1101 : 4'b0000;
									assign node18276 = (inp[2]) ? node18386 : node18277;
										assign node18277 = (inp[4]) ? node18313 : node18278;
											assign node18278 = (inp[13]) ? node18292 : node18279;
												assign node18279 = (inp[10]) ? node18285 : node18280;
													assign node18280 = (inp[12]) ? 4'b0101 : node18281;
														assign node18281 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node18285 = (inp[12]) ? 4'b1101 : node18286;
														assign node18286 = (inp[1]) ? node18288 : 4'b1101;
															assign node18288 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node18292 = (inp[7]) ? node18308 : node18293;
													assign node18293 = (inp[14]) ? node18303 : node18294;
														assign node18294 = (inp[10]) ? node18300 : node18295;
															assign node18295 = (inp[12]) ? 4'b0001 : node18296;
																assign node18296 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node18300 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node18303 = (inp[12]) ? node18305 : 4'b1001;
															assign node18305 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18308 = (inp[10]) ? 4'b1101 : node18309;
														assign node18309 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node18313 = (inp[13]) ? node18347 : node18314;
												assign node18314 = (inp[12]) ? node18328 : node18315;
													assign node18315 = (inp[1]) ? node18323 : node18316;
														assign node18316 = (inp[14]) ? 4'b0001 : node18317;
															assign node18317 = (inp[7]) ? node18319 : 4'b1000;
																assign node18319 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node18323 = (inp[10]) ? node18325 : 4'b1001;
															assign node18325 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18328 = (inp[7]) ? node18338 : node18329;
														assign node18329 = (inp[14]) ? node18335 : node18330;
															assign node18330 = (inp[1]) ? node18332 : 4'b0000;
																assign node18332 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node18335 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18338 = (inp[10]) ? node18340 : 4'b0001;
															assign node18340 = (inp[14]) ? node18344 : node18341;
																assign node18341 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node18344 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node18347 = (inp[7]) ? node18371 : node18348;
													assign node18348 = (inp[1]) ? node18360 : node18349;
														assign node18349 = (inp[14]) ? node18355 : node18350;
															assign node18350 = (inp[12]) ? 4'b1000 : node18351;
																assign node18351 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node18355 = (inp[10]) ? node18357 : 4'b1001;
																assign node18357 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node18360 = (inp[14]) ? node18366 : node18361;
															assign node18361 = (inp[12]) ? node18363 : 4'b0101;
																assign node18363 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node18366 = (inp[12]) ? node18368 : 4'b0100;
																assign node18368 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node18371 = (inp[1]) ? node18375 : node18372;
														assign node18372 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node18375 = (inp[14]) ? node18381 : node18376;
															assign node18376 = (inp[12]) ? 4'b1001 : node18377;
																assign node18377 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node18381 = (inp[10]) ? node18383 : 4'b0000;
																assign node18383 = (inp[12]) ? 4'b1000 : 4'b0100;
										assign node18386 = (inp[4]) ? node18440 : node18387;
											assign node18387 = (inp[13]) ? node18415 : node18388;
												assign node18388 = (inp[12]) ? node18406 : node18389;
													assign node18389 = (inp[14]) ? node18397 : node18390;
														assign node18390 = (inp[1]) ? node18392 : 4'b1001;
															assign node18392 = (inp[7]) ? 4'b1000 : node18393;
																assign node18393 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node18397 = (inp[1]) ? node18401 : node18398;
															assign node18398 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node18401 = (inp[7]) ? node18403 : 4'b0001;
																assign node18403 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18406 = (inp[14]) ? node18412 : node18407;
														assign node18407 = (inp[1]) ? node18409 : 4'b0001;
															assign node18409 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18412 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node18415 = (inp[14]) ? node18433 : node18416;
													assign node18416 = (inp[1]) ? node18422 : node18417;
														assign node18417 = (inp[7]) ? node18419 : 4'b1001;
															assign node18419 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node18422 = (inp[7]) ? node18428 : node18423;
															assign node18423 = (inp[10]) ? node18425 : 4'b0001;
																assign node18425 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node18428 = (inp[12]) ? 4'b0000 : node18429;
																assign node18429 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node18433 = (inp[1]) ? 4'b1001 : node18434;
														assign node18434 = (inp[7]) ? 4'b1000 : node18435;
															assign node18435 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node18440 = (inp[7]) ? node18462 : node18441;
												assign node18441 = (inp[13]) ? node18453 : node18442;
													assign node18442 = (inp[14]) ? node18444 : 4'b1001;
														assign node18444 = (inp[10]) ? node18450 : node18445;
															assign node18445 = (inp[12]) ? 4'b0001 : node18446;
																assign node18446 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node18450 = (inp[1]) ? 4'b0101 : 4'b1001;
													assign node18453 = (inp[1]) ? node18457 : node18454;
														assign node18454 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node18457 = (inp[10]) ? 4'b0101 : node18458;
															assign node18458 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node18462 = (inp[10]) ? node18468 : node18463;
													assign node18463 = (inp[12]) ? 4'b0001 : node18464;
														assign node18464 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node18468 = (inp[12]) ? 4'b1001 : node18469;
														assign node18469 = (inp[1]) ? node18471 : 4'b1001;
															assign node18471 = (inp[13]) ? 4'b0101 : 4'b0001;
								assign node18475 = (inp[1]) ? node18643 : node18476;
									assign node18476 = (inp[3]) ? node18552 : node18477;
										assign node18477 = (inp[2]) ? node18521 : node18478;
											assign node18478 = (inp[4]) ? node18498 : node18479;
												assign node18479 = (inp[7]) ? node18491 : node18480;
													assign node18480 = (inp[13]) ? node18486 : node18481;
														assign node18481 = (inp[12]) ? 4'b0101 : node18482;
															assign node18482 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node18486 = (inp[12]) ? 4'b0000 : node18487;
															assign node18487 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node18491 = (inp[13]) ? 4'b1101 : node18492;
														assign node18492 = (inp[12]) ? 4'b0101 : node18493;
															assign node18493 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node18498 = (inp[13]) ? node18512 : node18499;
													assign node18499 = (inp[7]) ? node18505 : node18500;
														assign node18500 = (inp[10]) ? 4'b0100 : node18501;
															assign node18501 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18505 = (inp[10]) ? node18509 : node18506;
															assign node18506 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node18509 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node18512 = (inp[10]) ? node18518 : node18513;
														assign node18513 = (inp[7]) ? 4'b1000 : node18514;
															assign node18514 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node18518 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node18521 = (inp[7]) ? node18543 : node18522;
												assign node18522 = (inp[4]) ? node18532 : node18523;
													assign node18523 = (inp[13]) ? node18527 : node18524;
														assign node18524 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node18527 = (inp[12]) ? 4'b1101 : node18528;
															assign node18528 = (inp[10]) ? 4'b0001 : 4'b1101;
													assign node18532 = (inp[13]) ? node18538 : node18533;
														assign node18533 = (inp[10]) ? node18535 : 4'b0001;
															assign node18535 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18538 = (inp[12]) ? 4'b1001 : node18539;
															assign node18539 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node18543 = (inp[13]) ? node18549 : node18544;
													assign node18544 = (inp[12]) ? 4'b0101 : node18545;
														assign node18545 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node18549 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node18552 = (inp[2]) ? node18598 : node18553;
											assign node18553 = (inp[4]) ? node18583 : node18554;
												assign node18554 = (inp[13]) ? node18570 : node18555;
													assign node18555 = (inp[14]) ? node18563 : node18556;
														assign node18556 = (inp[10]) ? node18560 : node18557;
															assign node18557 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18560 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node18563 = (inp[10]) ? node18567 : node18564;
															assign node18564 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18567 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node18570 = (inp[7]) ? node18578 : node18571;
														assign node18571 = (inp[14]) ? node18573 : 4'b0000;
															assign node18573 = (inp[12]) ? node18575 : 4'b1000;
																assign node18575 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18578 = (inp[12]) ? node18580 : 4'b0000;
															assign node18580 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node18583 = (inp[13]) ? node18593 : node18584;
													assign node18584 = (inp[10]) ? 4'b0001 : node18585;
														assign node18585 = (inp[7]) ? node18589 : node18586;
															assign node18586 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node18589 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node18593 = (inp[7]) ? 4'b1001 : node18594;
														assign node18594 = (inp[10]) ? 4'b1101 : 4'b1001;
											assign node18598 = (inp[4]) ? node18620 : node18599;
												assign node18599 = (inp[13]) ? node18609 : node18600;
													assign node18600 = (inp[10]) ? node18602 : 4'b0001;
														assign node18602 = (inp[7]) ? node18606 : node18603;
															assign node18603 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node18606 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node18609 = (inp[7]) ? node18615 : node18610;
														assign node18610 = (inp[12]) ? 4'b0000 : node18611;
															assign node18611 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node18615 = (inp[12]) ? 4'b1001 : node18616;
															assign node18616 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node18620 = (inp[13]) ? node18628 : node18621;
													assign node18621 = (inp[12]) ? node18625 : node18622;
														assign node18622 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node18625 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18628 = (inp[7]) ? node18638 : node18629;
														assign node18629 = (inp[14]) ? node18631 : 4'b0100;
															assign node18631 = (inp[12]) ? node18635 : node18632;
																assign node18632 = (inp[10]) ? 4'b0100 : 4'b1100;
																assign node18635 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node18638 = (inp[10]) ? node18640 : 4'b1000;
															assign node18640 = (inp[12]) ? 4'b1000 : 4'b0100;
									assign node18643 = (inp[10]) ? node18715 : node18644;
										assign node18644 = (inp[4]) ? node18674 : node18645;
											assign node18645 = (inp[2]) ? node18655 : node18646;
												assign node18646 = (inp[13]) ? node18652 : node18647;
													assign node18647 = (inp[12]) ? node18649 : 4'b1100;
														assign node18649 = (inp[3]) ? 4'b1100 : 4'b0100;
													assign node18652 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node18655 = (inp[3]) ? node18665 : node18656;
													assign node18656 = (inp[12]) ? node18662 : node18657;
														assign node18657 = (inp[13]) ? node18659 : 4'b1100;
															assign node18659 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node18662 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node18665 = (inp[7]) ? node18669 : node18666;
														assign node18666 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18669 = (inp[12]) ? node18671 : 4'b0000;
															assign node18671 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node18674 = (inp[3]) ? node18694 : node18675;
												assign node18675 = (inp[2]) ? node18681 : node18676;
													assign node18676 = (inp[7]) ? 4'b1000 : node18677;
														assign node18677 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node18681 = (inp[7]) ? node18687 : node18682;
														assign node18682 = (inp[12]) ? node18684 : 4'b0000;
															assign node18684 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node18687 = (inp[13]) ? node18691 : node18688;
															assign node18688 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18691 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node18694 = (inp[7]) ? node18706 : node18695;
													assign node18695 = (inp[13]) ? node18701 : node18696;
														assign node18696 = (inp[12]) ? 4'b1000 : node18697;
															assign node18697 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node18701 = (inp[12]) ? node18703 : 4'b1100;
															assign node18703 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node18706 = (inp[2]) ? 4'b1000 : node18707;
														assign node18707 = (inp[12]) ? node18711 : node18708;
															assign node18708 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node18711 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node18715 = (inp[13]) ? node18747 : node18716;
											assign node18716 = (inp[7]) ? node18734 : node18717;
												assign node18717 = (inp[4]) ? node18723 : node18718;
													assign node18718 = (inp[3]) ? 4'b0000 : node18719;
														assign node18719 = (inp[2]) ? 4'b1100 : 4'b0000;
													assign node18723 = (inp[12]) ? node18729 : node18724;
														assign node18724 = (inp[3]) ? node18726 : 4'b1000;
															assign node18726 = (inp[2]) ? 4'b0100 : 4'b1000;
														assign node18729 = (inp[2]) ? 4'b0100 : node18730;
															assign node18730 = (inp[14]) ? 4'b0100 : 4'b1000;
												assign node18734 = (inp[3]) ? node18740 : node18735;
													assign node18735 = (inp[2]) ? 4'b1100 : node18736;
														assign node18736 = (inp[4]) ? 4'b0000 : 4'b1100;
													assign node18740 = (inp[2]) ? node18744 : node18741;
														assign node18741 = (inp[4]) ? 4'b1000 : 4'b0100;
														assign node18744 = (inp[4]) ? 4'b0000 : 4'b1000;
											assign node18747 = (inp[4]) ? node18755 : node18748;
												assign node18748 = (inp[2]) ? node18750 : 4'b0000;
													assign node18750 = (inp[3]) ? 4'b0000 : node18751;
														assign node18751 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node18755 = (inp[3]) ? 4'b0100 : node18756;
													assign node18756 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node18760 = (inp[2]) ? 4'b0100 : node18761;
								assign node18761 = (inp[3]) ? node18865 : node18762;
									assign node18762 = (inp[4]) ? node18788 : node18763;
										assign node18763 = (inp[13]) ? node18765 : 4'b0100;
											assign node18765 = (inp[7]) ? 4'b0100 : node18766;
												assign node18766 = (inp[12]) ? node18780 : node18767;
													assign node18767 = (inp[10]) ? node18773 : node18768;
														assign node18768 = (inp[14]) ? node18770 : 4'b0000;
															assign node18770 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node18773 = (inp[1]) ? node18775 : 4'b0001;
															assign node18775 = (inp[11]) ? 4'b0000 : node18776;
																assign node18776 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18780 = (inp[10]) ? node18782 : 4'b0100;
														assign node18782 = (inp[1]) ? node18784 : 4'b0100;
															assign node18784 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node18788 = (inp[7]) ? node18844 : node18789;
											assign node18789 = (inp[1]) ? node18813 : node18790;
												assign node18790 = (inp[13]) ? node18804 : node18791;
													assign node18791 = (inp[12]) ? 4'b0001 : node18792;
														assign node18792 = (inp[10]) ? node18798 : node18793;
															assign node18793 = (inp[11]) ? 4'b0001 : node18794;
																assign node18794 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18798 = (inp[11]) ? 4'b1001 : node18799;
																assign node18799 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18804 = (inp[10]) ? node18810 : node18805;
														assign node18805 = (inp[12]) ? 4'b1001 : node18806;
															assign node18806 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18810 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node18813 = (inp[11]) ? node18825 : node18814;
													assign node18814 = (inp[14]) ? node18822 : node18815;
														assign node18815 = (inp[13]) ? node18817 : 4'b1000;
															assign node18817 = (inp[10]) ? 4'b0000 : node18818;
																assign node18818 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node18822 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node18825 = (inp[14]) ? node18833 : node18826;
														assign node18826 = (inp[12]) ? node18828 : 4'b0000;
															assign node18828 = (inp[10]) ? 4'b0000 : node18829;
																assign node18829 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node18833 = (inp[13]) ? node18839 : node18834;
															assign node18834 = (inp[10]) ? 4'b1000 : node18835;
																assign node18835 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node18839 = (inp[10]) ? 4'b0000 : node18840;
																assign node18840 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node18844 = (inp[13]) ? node18846 : 4'b0100;
												assign node18846 = (inp[1]) ? node18852 : node18847;
													assign node18847 = (inp[12]) ? 4'b0100 : node18848;
														assign node18848 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node18852 = (inp[12]) ? node18858 : node18853;
														assign node18853 = (inp[11]) ? 4'b0000 : node18854;
															assign node18854 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18858 = (inp[14]) ? node18860 : 4'b0000;
															assign node18860 = (inp[10]) ? node18862 : 4'b0100;
																assign node18862 = (inp[11]) ? 4'b0000 : 4'b0100;
									assign node18865 = (inp[1]) ? node18953 : node18866;
										assign node18866 = (inp[11]) ? node18916 : node18867;
											assign node18867 = (inp[14]) ? node18891 : node18868;
												assign node18868 = (inp[4]) ? node18880 : node18869;
													assign node18869 = (inp[13]) ? node18875 : node18870;
														assign node18870 = (inp[12]) ? 4'b0001 : node18871;
															assign node18871 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18875 = (inp[10]) ? node18877 : 4'b1001;
															assign node18877 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node18880 = (inp[7]) ? node18886 : node18881;
														assign node18881 = (inp[12]) ? 4'b1101 : node18882;
															assign node18882 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node18886 = (inp[13]) ? 4'b1001 : node18887;
															assign node18887 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node18891 = (inp[13]) ? node18901 : node18892;
													assign node18892 = (inp[12]) ? node18896 : node18893;
														assign node18893 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18896 = (inp[7]) ? 4'b0000 : node18897;
															assign node18897 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node18901 = (inp[12]) ? node18911 : node18902;
														assign node18902 = (inp[10]) ? node18906 : node18903;
															assign node18903 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node18906 = (inp[7]) ? node18908 : 4'b0100;
																assign node18908 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node18911 = (inp[7]) ? 4'b1000 : node18912;
															assign node18912 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node18916 = (inp[7]) ? node18940 : node18917;
												assign node18917 = (inp[4]) ? node18927 : node18918;
													assign node18918 = (inp[13]) ? node18924 : node18919;
														assign node18919 = (inp[10]) ? node18921 : 4'b0001;
															assign node18921 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18924 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node18927 = (inp[13]) ? node18935 : node18928;
														assign node18928 = (inp[14]) ? 4'b0101 : node18929;
															assign node18929 = (inp[10]) ? node18931 : 4'b0101;
																assign node18931 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node18935 = (inp[12]) ? 4'b1101 : node18936;
															assign node18936 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node18940 = (inp[13]) ? node18946 : node18941;
													assign node18941 = (inp[12]) ? 4'b0001 : node18942;
														assign node18942 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18946 = (inp[12]) ? 4'b1001 : node18947;
														assign node18947 = (inp[10]) ? node18949 : 4'b1001;
															assign node18949 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node18953 = (inp[11]) ? node18989 : node18954;
											assign node18954 = (inp[14]) ? node18974 : node18955;
												assign node18955 = (inp[7]) ? node18961 : node18956;
													assign node18956 = (inp[13]) ? 4'b0100 : node18957;
														assign node18957 = (inp[4]) ? 4'b0100 : 4'b1000;
													assign node18961 = (inp[13]) ? node18965 : node18962;
														assign node18962 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18965 = (inp[4]) ? node18969 : node18966;
															assign node18966 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node18969 = (inp[10]) ? 4'b0100 : node18970;
																assign node18970 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node18974 = (inp[13]) ? node18980 : node18975;
													assign node18975 = (inp[12]) ? 4'b0001 : node18976;
														assign node18976 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node18980 = (inp[4]) ? node18982 : 4'b1001;
														assign node18982 = (inp[12]) ? node18986 : node18983;
															assign node18983 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node18986 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node18989 = (inp[4]) ? node19007 : node18990;
												assign node18990 = (inp[13]) ? node18996 : node18991;
													assign node18991 = (inp[12]) ? node18993 : 4'b1000;
														assign node18993 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18996 = (inp[7]) ? node19002 : node18997;
														assign node18997 = (inp[12]) ? node18999 : 4'b0100;
															assign node18999 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node19002 = (inp[10]) ? 4'b0000 : node19003;
															assign node19003 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node19007 = (inp[13]) ? node19019 : node19008;
													assign node19008 = (inp[7]) ? node19014 : node19009;
														assign node19009 = (inp[10]) ? 4'b1100 : node19010;
															assign node19010 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19014 = (inp[12]) ? node19016 : 4'b1000;
															assign node19016 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node19019 = (inp[10]) ? 4'b0100 : node19020;
														assign node19020 = (inp[12]) ? 4'b1100 : 4'b0100;
						assign node19025 = (inp[3]) ? node19643 : node19026;
							assign node19026 = (inp[4]) ? node19320 : node19027;
								assign node19027 = (inp[13]) ? node19149 : node19028;
									assign node19028 = (inp[0]) ? node19110 : node19029;
										assign node19029 = (inp[10]) ? node19063 : node19030;
											assign node19030 = (inp[11]) ? node19046 : node19031;
												assign node19031 = (inp[2]) ? node19041 : node19032;
													assign node19032 = (inp[1]) ? node19038 : node19033;
														assign node19033 = (inp[14]) ? 4'b0101 : node19034;
															assign node19034 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19038 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node19041 = (inp[12]) ? 4'b0101 : node19042;
														assign node19042 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node19046 = (inp[1]) ? node19054 : node19047;
													assign node19047 = (inp[12]) ? node19051 : node19048;
														assign node19048 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19051 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node19054 = (inp[7]) ? node19060 : node19055;
														assign node19055 = (inp[12]) ? node19057 : 4'b0000;
															assign node19057 = (inp[14]) ? 4'b1100 : 4'b0000;
														assign node19060 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node19063 = (inp[7]) ? node19087 : node19064;
												assign node19064 = (inp[2]) ? node19074 : node19065;
													assign node19065 = (inp[1]) ? node19069 : node19066;
														assign node19066 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node19069 = (inp[11]) ? 4'b0000 : node19070;
															assign node19070 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19074 = (inp[1]) ? node19080 : node19075;
														assign node19075 = (inp[14]) ? 4'b0001 : node19076;
															assign node19076 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node19080 = (inp[11]) ? 4'b1000 : node19081;
															assign node19081 = (inp[12]) ? node19083 : 4'b1001;
																assign node19083 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node19087 = (inp[11]) ? node19101 : node19088;
													assign node19088 = (inp[2]) ? node19096 : node19089;
														assign node19089 = (inp[12]) ? node19091 : 4'b0000;
															assign node19091 = (inp[1]) ? node19093 : 4'b1101;
																assign node19093 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node19096 = (inp[14]) ? node19098 : 4'b1101;
															assign node19098 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node19101 = (inp[2]) ? node19105 : node19102;
														assign node19102 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node19105 = (inp[12]) ? node19107 : 4'b0100;
															assign node19107 = (inp[1]) ? 4'b0100 : 4'b1100;
										assign node19110 = (inp[2]) ? 4'b0100 : node19111;
											assign node19111 = (inp[1]) ? node19129 : node19112;
												assign node19112 = (inp[14]) ? node19118 : node19113;
													assign node19113 = (inp[12]) ? 4'b0101 : node19114;
														assign node19114 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node19118 = (inp[11]) ? node19124 : node19119;
														assign node19119 = (inp[12]) ? 4'b0100 : node19120;
															assign node19120 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node19124 = (inp[10]) ? node19126 : 4'b0101;
															assign node19126 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node19129 = (inp[10]) ? node19137 : node19130;
													assign node19130 = (inp[12]) ? node19132 : 4'b1100;
														assign node19132 = (inp[14]) ? node19134 : 4'b0100;
															assign node19134 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19137 = (inp[7]) ? node19143 : node19138;
														assign node19138 = (inp[11]) ? 4'b0000 : node19139;
															assign node19139 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node19143 = (inp[11]) ? 4'b1100 : node19144;
															assign node19144 = (inp[14]) ? 4'b0101 : 4'b1100;
									assign node19149 = (inp[1]) ? node19231 : node19150;
										assign node19150 = (inp[0]) ? node19196 : node19151;
											assign node19151 = (inp[2]) ? node19165 : node19152;
												assign node19152 = (inp[10]) ? node19156 : node19153;
													assign node19153 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node19156 = (inp[7]) ? node19162 : node19157;
														assign node19157 = (inp[12]) ? node19159 : 4'b1100;
															assign node19159 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node19162 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node19165 = (inp[10]) ? node19187 : node19166;
													assign node19166 = (inp[7]) ? node19176 : node19167;
														assign node19167 = (inp[12]) ? node19171 : node19168;
															assign node19168 = (inp[14]) ? 4'b1001 : 4'b0001;
															assign node19171 = (inp[11]) ? 4'b1001 : node19172;
																assign node19172 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node19176 = (inp[12]) ? node19184 : node19177;
															assign node19177 = (inp[14]) ? node19181 : node19178;
																assign node19178 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node19181 = (inp[11]) ? 4'b0001 : 4'b0101;
															assign node19184 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19187 = (inp[14]) ? node19191 : node19188;
														assign node19188 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19191 = (inp[12]) ? node19193 : 4'b1001;
															assign node19193 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node19196 = (inp[2]) ? node19220 : node19197;
												assign node19197 = (inp[7]) ? node19211 : node19198;
													assign node19198 = (inp[11]) ? node19202 : node19199;
														assign node19199 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19202 = (inp[14]) ? 4'b0000 : node19203;
															assign node19203 = (inp[10]) ? node19207 : node19204;
																assign node19204 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node19207 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19211 = (inp[10]) ? node19213 : 4'b1101;
														assign node19213 = (inp[12]) ? node19217 : node19214;
															assign node19214 = (inp[11]) ? 4'b0000 : 4'b0100;
															assign node19217 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node19220 = (inp[10]) ? node19222 : 4'b0100;
													assign node19222 = (inp[7]) ? 4'b0100 : node19223;
														assign node19223 = (inp[12]) ? 4'b0100 : node19224;
															assign node19224 = (inp[11]) ? 4'b0001 : node19225;
																assign node19225 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node19231 = (inp[11]) ? node19291 : node19232;
											assign node19232 = (inp[12]) ? node19270 : node19233;
												assign node19233 = (inp[10]) ? node19253 : node19234;
													assign node19234 = (inp[14]) ? node19246 : node19235;
														assign node19235 = (inp[2]) ? node19241 : node19236;
															assign node19236 = (inp[0]) ? 4'b1001 : node19237;
																assign node19237 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node19241 = (inp[0]) ? node19243 : 4'b0001;
																assign node19243 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node19246 = (inp[0]) ? 4'b0100 : node19247;
															assign node19247 = (inp[2]) ? 4'b0000 : node19248;
																assign node19248 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node19253 = (inp[2]) ? node19259 : node19254;
														assign node19254 = (inp[0]) ? 4'b0001 : node19255;
															assign node19255 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node19259 = (inp[14]) ? node19267 : node19260;
															assign node19260 = (inp[0]) ? node19264 : node19261;
																assign node19261 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node19264 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node19267 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node19270 = (inp[0]) ? node19282 : node19271;
													assign node19271 = (inp[2]) ? node19277 : node19272;
														assign node19272 = (inp[7]) ? 4'b1000 : node19273;
															assign node19273 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node19277 = (inp[10]) ? 4'b1001 : node19278;
															assign node19278 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19282 = (inp[2]) ? node19288 : node19283;
														assign node19283 = (inp[10]) ? node19285 : 4'b0001;
															assign node19285 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node19288 = (inp[14]) ? 4'b0100 : 4'b0000;
											assign node19291 = (inp[7]) ? node19307 : node19292;
												assign node19292 = (inp[0]) ? node19300 : node19293;
													assign node19293 = (inp[10]) ? node19297 : node19294;
														assign node19294 = (inp[2]) ? 4'b1000 : 4'b0100;
														assign node19297 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node19300 = (inp[10]) ? 4'b0000 : node19301;
														assign node19301 = (inp[2]) ? node19303 : 4'b1000;
															assign node19303 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node19307 = (inp[0]) ? node19311 : node19308;
													assign node19308 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node19311 = (inp[10]) ? node19317 : node19312;
														assign node19312 = (inp[2]) ? 4'b0100 : node19313;
															assign node19313 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node19317 = (inp[2]) ? 4'b0100 : 4'b0000;
								assign node19320 = (inp[2]) ? node19492 : node19321;
									assign node19321 = (inp[11]) ? node19423 : node19322;
										assign node19322 = (inp[10]) ? node19370 : node19323;
											assign node19323 = (inp[0]) ? node19347 : node19324;
												assign node19324 = (inp[13]) ? node19338 : node19325;
													assign node19325 = (inp[7]) ? node19331 : node19326;
														assign node19326 = (inp[1]) ? 4'b0000 : node19327;
															assign node19327 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19331 = (inp[12]) ? node19333 : 4'b1100;
															assign node19333 = (inp[1]) ? node19335 : 4'b0100;
																assign node19335 = (inp[14]) ? 4'b1100 : 4'b0000;
													assign node19338 = (inp[1]) ? 4'b0001 : node19339;
														assign node19339 = (inp[7]) ? node19343 : node19340;
															assign node19340 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node19343 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node19347 = (inp[12]) ? node19361 : node19348;
													assign node19348 = (inp[1]) ? node19354 : node19349;
														assign node19349 = (inp[13]) ? node19351 : 4'b0001;
															assign node19351 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node19354 = (inp[13]) ? node19356 : 4'b1001;
															assign node19356 = (inp[7]) ? 4'b1001 : node19357;
																assign node19357 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19361 = (inp[7]) ? 4'b0001 : node19362;
														assign node19362 = (inp[1]) ? node19364 : 4'b0101;
															assign node19364 = (inp[14]) ? node19366 : 4'b0001;
																assign node19366 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node19370 = (inp[12]) ? node19406 : node19371;
												assign node19371 = (inp[0]) ? node19397 : node19372;
													assign node19372 = (inp[7]) ? node19386 : node19373;
														assign node19373 = (inp[13]) ? node19381 : node19374;
															assign node19374 = (inp[1]) ? node19378 : node19375;
																assign node19375 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node19378 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node19381 = (inp[1]) ? node19383 : 4'b0000;
																assign node19383 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node19386 = (inp[13]) ? node19394 : node19387;
															assign node19387 = (inp[14]) ? node19391 : node19388;
																assign node19388 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node19391 = (inp[1]) ? 4'b0001 : 4'b1000;
															assign node19394 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node19397 = (inp[1]) ? node19399 : 4'b1001;
														assign node19399 = (inp[13]) ? node19403 : node19400;
															assign node19400 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node19403 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node19406 = (inp[1]) ? node19416 : node19407;
													assign node19407 = (inp[7]) ? node19413 : node19408;
														assign node19408 = (inp[13]) ? node19410 : 4'b1001;
															assign node19410 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node19413 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node19416 = (inp[14]) ? node19418 : 4'b1001;
														assign node19418 = (inp[7]) ? 4'b1001 : node19419;
															assign node19419 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node19423 = (inp[10]) ? node19457 : node19424;
											assign node19424 = (inp[1]) ? node19444 : node19425;
												assign node19425 = (inp[13]) ? node19433 : node19426;
													assign node19426 = (inp[7]) ? node19430 : node19427;
														assign node19427 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node19430 = (inp[0]) ? 4'b1000 : 4'b1100;
													assign node19433 = (inp[7]) ? node19441 : node19434;
														assign node19434 = (inp[0]) ? node19438 : node19435;
															assign node19435 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19438 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node19441 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node19444 = (inp[12]) ? node19446 : 4'b1000;
													assign node19446 = (inp[7]) ? node19452 : node19447;
														assign node19447 = (inp[0]) ? node19449 : 4'b1000;
															assign node19449 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node19452 = (inp[0]) ? 4'b1000 : node19453;
															assign node19453 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node19457 = (inp[1]) ? node19481 : node19458;
												assign node19458 = (inp[7]) ? node19466 : node19459;
													assign node19459 = (inp[13]) ? node19463 : node19460;
														assign node19460 = (inp[12]) ? 4'b1001 : 4'b0100;
														assign node19463 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node19466 = (inp[13]) ? node19474 : node19467;
														assign node19467 = (inp[12]) ? node19471 : node19468;
															assign node19468 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node19471 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node19474 = (inp[0]) ? node19478 : node19475;
															assign node19475 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19478 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node19481 = (inp[7]) ? node19487 : node19482;
													assign node19482 = (inp[0]) ? node19484 : 4'b0000;
														assign node19484 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node19487 = (inp[0]) ? 4'b0000 : node19488;
														assign node19488 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node19492 = (inp[7]) ? node19588 : node19493;
										assign node19493 = (inp[1]) ? node19543 : node19494;
											assign node19494 = (inp[11]) ? node19520 : node19495;
												assign node19495 = (inp[0]) ? node19511 : node19496;
													assign node19496 = (inp[13]) ? node19504 : node19497;
														assign node19497 = (inp[10]) ? node19501 : node19498;
															assign node19498 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node19501 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19504 = (inp[10]) ? node19508 : node19505;
															assign node19505 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19508 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19511 = (inp[14]) ? node19513 : 4'b1001;
														assign node19513 = (inp[13]) ? 4'b1000 : node19514;
															assign node19514 = (inp[10]) ? node19516 : 4'b0000;
																assign node19516 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node19520 = (inp[0]) ? node19532 : node19521;
													assign node19521 = (inp[13]) ? node19527 : node19522;
														assign node19522 = (inp[10]) ? 4'b1000 : node19523;
															assign node19523 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node19527 = (inp[10]) ? node19529 : 4'b1000;
															assign node19529 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node19532 = (inp[13]) ? node19538 : node19533;
														assign node19533 = (inp[10]) ? node19535 : 4'b0001;
															assign node19535 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19538 = (inp[12]) ? 4'b1001 : node19539;
															assign node19539 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node19543 = (inp[11]) ? node19571 : node19544;
												assign node19544 = (inp[12]) ? node19556 : node19545;
													assign node19545 = (inp[0]) ? node19551 : node19546;
														assign node19546 = (inp[13]) ? node19548 : 4'b0000;
															assign node19548 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node19551 = (inp[14]) ? 4'b0001 : node19552;
															assign node19552 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node19556 = (inp[0]) ? node19566 : node19557;
														assign node19557 = (inp[13]) ? node19561 : node19558;
															assign node19558 = (inp[14]) ? 4'b1000 : 4'b1101;
															assign node19561 = (inp[14]) ? node19563 : 4'b1000;
																assign node19563 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node19566 = (inp[14]) ? 4'b0001 : node19567;
															assign node19567 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node19571 = (inp[0]) ? node19577 : node19572;
													assign node19572 = (inp[10]) ? 4'b0000 : node19573;
														assign node19573 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node19577 = (inp[13]) ? node19583 : node19578;
														assign node19578 = (inp[12]) ? node19580 : 4'b1000;
															assign node19580 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19583 = (inp[10]) ? 4'b0000 : node19584;
															assign node19584 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node19588 = (inp[0]) ? node19624 : node19589;
											assign node19589 = (inp[13]) ? node19613 : node19590;
												assign node19590 = (inp[10]) ? node19604 : node19591;
													assign node19591 = (inp[1]) ? node19599 : node19592;
														assign node19592 = (inp[12]) ? node19596 : node19593;
															assign node19593 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node19596 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19599 = (inp[14]) ? 4'b1000 : node19600;
															assign node19600 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node19604 = (inp[1]) ? node19606 : 4'b0101;
														assign node19606 = (inp[11]) ? 4'b0000 : node19607;
															assign node19607 = (inp[14]) ? node19609 : 4'b0101;
																assign node19609 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node19613 = (inp[1]) ? node19619 : node19614;
													assign node19614 = (inp[11]) ? 4'b1000 : node19615;
														assign node19615 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node19619 = (inp[11]) ? 4'b0000 : node19620;
														assign node19620 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node19624 = (inp[13]) ? node19626 : 4'b0100;
												assign node19626 = (inp[10]) ? node19632 : node19627;
													assign node19627 = (inp[1]) ? node19629 : 4'b0100;
														assign node19629 = (inp[14]) ? 4'b0100 : 4'b0000;
													assign node19632 = (inp[12]) ? node19636 : node19633;
														assign node19633 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node19636 = (inp[1]) ? node19638 : 4'b0100;
															assign node19638 = (inp[11]) ? 4'b0000 : node19639;
																assign node19639 = (inp[14]) ? 4'b0100 : 4'b0000;
							assign node19643 = (inp[4]) ? node20035 : node19644;
								assign node19644 = (inp[11]) ? node19890 : node19645;
									assign node19645 = (inp[2]) ? node19773 : node19646;
										assign node19646 = (inp[1]) ? node19716 : node19647;
											assign node19647 = (inp[0]) ? node19681 : node19648;
												assign node19648 = (inp[10]) ? node19662 : node19649;
													assign node19649 = (inp[7]) ? node19655 : node19650;
														assign node19650 = (inp[12]) ? node19652 : 4'b1001;
															assign node19652 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node19655 = (inp[13]) ? node19659 : node19656;
															assign node19656 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node19659 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19662 = (inp[12]) ? node19670 : node19663;
														assign node19663 = (inp[13]) ? 4'b0000 : node19664;
															assign node19664 = (inp[7]) ? 4'b1000 : node19665;
																assign node19665 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19670 = (inp[14]) ? node19676 : node19671;
															assign node19671 = (inp[7]) ? node19673 : 4'b1000;
																assign node19673 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node19676 = (inp[13]) ? node19678 : 4'b1000;
																assign node19678 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node19681 = (inp[12]) ? node19697 : node19682;
													assign node19682 = (inp[10]) ? node19694 : node19683;
														assign node19683 = (inp[14]) ? node19689 : node19684;
															assign node19684 = (inp[13]) ? node19686 : 4'b1000;
																assign node19686 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node19689 = (inp[13]) ? node19691 : 4'b0001;
																assign node19691 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node19694 = (inp[13]) ? 4'b0001 : 4'b1000;
													assign node19697 = (inp[7]) ? node19707 : node19698;
														assign node19698 = (inp[10]) ? node19702 : node19699;
															assign node19699 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node19702 = (inp[13]) ? node19704 : 4'b0000;
																assign node19704 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19707 = (inp[10]) ? node19711 : node19708;
															assign node19708 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node19711 = (inp[14]) ? 4'b1001 : node19712;
																assign node19712 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node19716 = (inp[10]) ? node19740 : node19717;
												assign node19717 = (inp[14]) ? node19731 : node19718;
													assign node19718 = (inp[7]) ? node19724 : node19719;
														assign node19719 = (inp[0]) ? 4'b1000 : node19720;
															assign node19720 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node19724 = (inp[12]) ? node19726 : 4'b1001;
															assign node19726 = (inp[0]) ? 4'b1001 : node19727;
																assign node19727 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node19731 = (inp[13]) ? node19733 : 4'b1000;
														assign node19733 = (inp[0]) ? node19737 : node19734;
															assign node19734 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node19737 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node19740 = (inp[12]) ? node19754 : node19741;
													assign node19741 = (inp[14]) ? node19749 : node19742;
														assign node19742 = (inp[7]) ? node19746 : node19743;
															assign node19743 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node19746 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node19749 = (inp[0]) ? node19751 : 4'b0001;
															assign node19751 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node19754 = (inp[13]) ? node19766 : node19755;
														assign node19755 = (inp[14]) ? node19761 : node19756;
															assign node19756 = (inp[7]) ? 4'b0001 : node19757;
																assign node19757 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node19761 = (inp[7]) ? 4'b1000 : node19762;
																assign node19762 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node19766 = (inp[0]) ? node19768 : 4'b0001;
															assign node19768 = (inp[14]) ? 4'b1001 : node19769;
																assign node19769 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node19773 = (inp[13]) ? node19825 : node19774;
											assign node19774 = (inp[14]) ? node19798 : node19775;
												assign node19775 = (inp[1]) ? node19785 : node19776;
													assign node19776 = (inp[0]) ? 4'b0001 : node19777;
														assign node19777 = (inp[12]) ? node19781 : node19778;
															assign node19778 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node19781 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node19785 = (inp[0]) ? node19791 : node19786;
														assign node19786 = (inp[7]) ? node19788 : 4'b0001;
															assign node19788 = (inp[10]) ? 4'b1001 : 4'b0000;
														assign node19791 = (inp[10]) ? node19795 : node19792;
															assign node19792 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19795 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node19798 = (inp[1]) ? node19814 : node19799;
													assign node19799 = (inp[0]) ? node19809 : node19800;
														assign node19800 = (inp[10]) ? node19804 : node19801;
															assign node19801 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19804 = (inp[12]) ? node19806 : 4'b0001;
																assign node19806 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node19809 = (inp[12]) ? 4'b0000 : node19810;
															assign node19810 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node19814 = (inp[0]) ? node19818 : node19815;
														assign node19815 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node19818 = (inp[12]) ? 4'b0001 : node19819;
															assign node19819 = (inp[10]) ? node19821 : 4'b0001;
																assign node19821 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node19825 = (inp[0]) ? node19857 : node19826;
												assign node19826 = (inp[10]) ? node19844 : node19827;
													assign node19827 = (inp[7]) ? node19833 : node19828;
														assign node19828 = (inp[1]) ? 4'b1000 : node19829;
															assign node19829 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node19833 = (inp[12]) ? node19841 : node19834;
															assign node19834 = (inp[14]) ? node19838 : node19835;
																assign node19835 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node19838 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node19841 = (inp[1]) ? 4'b1001 : 4'b0000;
													assign node19844 = (inp[7]) ? node19852 : node19845;
														assign node19845 = (inp[12]) ? 4'b0001 : node19846;
															assign node19846 = (inp[14]) ? node19848 : 4'b1001;
																assign node19848 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node19852 = (inp[14]) ? node19854 : 4'b1000;
															assign node19854 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node19857 = (inp[12]) ? node19877 : node19858;
													assign node19858 = (inp[14]) ? node19870 : node19859;
														assign node19859 = (inp[10]) ? node19865 : node19860;
															assign node19860 = (inp[1]) ? 4'b1001 : node19861;
																assign node19861 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node19865 = (inp[7]) ? 4'b0001 : node19866;
																assign node19866 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node19870 = (inp[1]) ? node19874 : node19871;
															assign node19871 = (inp[7]) ? 4'b0000 : 4'b1001;
															assign node19874 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node19877 = (inp[7]) ? node19881 : node19878;
														assign node19878 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19881 = (inp[14]) ? node19887 : node19882;
															assign node19882 = (inp[1]) ? node19884 : 4'b1001;
																assign node19884 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node19887 = (inp[1]) ? 4'b1001 : 4'b1000;
									assign node19890 = (inp[1]) ? node19976 : node19891;
										assign node19891 = (inp[13]) ? node19927 : node19892;
											assign node19892 = (inp[0]) ? node19916 : node19893;
												assign node19893 = (inp[10]) ? node19905 : node19894;
													assign node19894 = (inp[7]) ? node19900 : node19895;
														assign node19895 = (inp[2]) ? node19897 : 4'b0000;
															assign node19897 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node19900 = (inp[12]) ? 4'b1001 : node19901;
															assign node19901 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node19905 = (inp[12]) ? node19911 : node19906;
														assign node19906 = (inp[14]) ? node19908 : 4'b1001;
															assign node19908 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node19911 = (inp[2]) ? 4'b0000 : node19912;
															assign node19912 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node19916 = (inp[2]) ? 4'b0001 : node19917;
													assign node19917 = (inp[12]) ? node19921 : node19918;
														assign node19918 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node19921 = (inp[7]) ? 4'b0001 : node19922;
															assign node19922 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node19927 = (inp[12]) ? node19949 : node19928;
												assign node19928 = (inp[2]) ? node19940 : node19929;
													assign node19929 = (inp[10]) ? node19933 : node19930;
														assign node19930 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node19933 = (inp[0]) ? node19937 : node19934;
															assign node19934 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node19937 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node19940 = (inp[7]) ? node19944 : node19941;
														assign node19941 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node19944 = (inp[10]) ? node19946 : 4'b1001;
															assign node19946 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node19949 = (inp[0]) ? node19963 : node19950;
													assign node19950 = (inp[10]) ? node19956 : node19951;
														assign node19951 = (inp[2]) ? node19953 : 4'b0000;
															assign node19953 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node19956 = (inp[7]) ? node19960 : node19957;
															assign node19957 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node19960 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node19963 = (inp[7]) ? node19971 : node19964;
														assign node19964 = (inp[14]) ? 4'b0000 : node19965;
															assign node19965 = (inp[2]) ? node19967 : 4'b0000;
																assign node19967 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19971 = (inp[10]) ? 4'b0001 : node19972;
															assign node19972 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node19976 = (inp[2]) ? node19996 : node19977;
											assign node19977 = (inp[12]) ? node19979 : 4'b0000;
												assign node19979 = (inp[0]) ? node19987 : node19980;
													assign node19980 = (inp[13]) ? 4'b0000 : node19981;
														assign node19981 = (inp[10]) ? node19983 : 4'b0000;
															assign node19983 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node19987 = (inp[10]) ? 4'b0000 : node19988;
														assign node19988 = (inp[14]) ? node19990 : 4'b1000;
															assign node19990 = (inp[7]) ? 4'b0000 : node19991;
																assign node19991 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node19996 = (inp[10]) ? node20022 : node19997;
												assign node19997 = (inp[7]) ? node20009 : node19998;
													assign node19998 = (inp[14]) ? 4'b1000 : node19999;
														assign node19999 = (inp[0]) ? node20003 : node20000;
															assign node20000 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node20003 = (inp[12]) ? node20005 : 4'b1000;
																assign node20005 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node20009 = (inp[0]) ? node20015 : node20010;
														assign node20010 = (inp[12]) ? 4'b0000 : node20011;
															assign node20011 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node20015 = (inp[14]) ? 4'b0000 : node20016;
															assign node20016 = (inp[12]) ? node20018 : 4'b1000;
																assign node20018 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node20022 = (inp[13]) ? 4'b0000 : node20023;
													assign node20023 = (inp[12]) ? node20029 : node20024;
														assign node20024 = (inp[0]) ? node20026 : 4'b0000;
															assign node20026 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node20029 = (inp[14]) ? 4'b1000 : node20030;
															assign node20030 = (inp[0]) ? 4'b0000 : 4'b1000;
								assign node20035 = (inp[13]) ? node20237 : node20036;
									assign node20036 = (inp[10]) ? node20152 : node20037;
										assign node20037 = (inp[11]) ? node20105 : node20038;
											assign node20038 = (inp[12]) ? node20070 : node20039;
												assign node20039 = (inp[1]) ? node20051 : node20040;
													assign node20040 = (inp[14]) ? node20048 : node20041;
														assign node20041 = (inp[0]) ? node20043 : 4'b0000;
															assign node20043 = (inp[7]) ? node20045 : 4'b1000;
																assign node20045 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node20048 = (inp[0]) ? 4'b0001 : 4'b1001;
													assign node20051 = (inp[7]) ? node20063 : node20052;
														assign node20052 = (inp[0]) ? node20058 : node20053;
															assign node20053 = (inp[2]) ? node20055 : 4'b1001;
																assign node20055 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node20058 = (inp[14]) ? node20060 : 4'b0000;
																assign node20060 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node20063 = (inp[0]) ? node20065 : 4'b1000;
															assign node20065 = (inp[14]) ? node20067 : 4'b1001;
																assign node20067 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node20070 = (inp[14]) ? node20092 : node20071;
													assign node20071 = (inp[1]) ? node20085 : node20072;
														assign node20072 = (inp[7]) ? node20080 : node20073;
															assign node20073 = (inp[0]) ? node20077 : node20074;
																assign node20074 = (inp[2]) ? 4'b1000 : 4'b0000;
																assign node20077 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node20080 = (inp[2]) ? 4'b1001 : node20081;
																assign node20081 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20085 = (inp[0]) ? node20089 : node20086;
															assign node20086 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node20089 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node20092 = (inp[1]) ? node20098 : node20093;
														assign node20093 = (inp[0]) ? 4'b0001 : node20094;
															assign node20094 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node20098 = (inp[7]) ? node20100 : 4'b0001;
															assign node20100 = (inp[0]) ? 4'b0000 : node20101;
																assign node20101 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node20105 = (inp[1]) ? node20129 : node20106;
												assign node20106 = (inp[2]) ? node20116 : node20107;
													assign node20107 = (inp[7]) ? node20111 : node20108;
														assign node20108 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20111 = (inp[12]) ? 4'b1000 : node20112;
															assign node20112 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node20116 = (inp[12]) ? node20124 : node20117;
														assign node20117 = (inp[0]) ? node20121 : node20118;
															assign node20118 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node20121 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node20124 = (inp[7]) ? node20126 : 4'b1000;
															assign node20126 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node20129 = (inp[0]) ? node20141 : node20130;
													assign node20130 = (inp[7]) ? node20136 : node20131;
														assign node20131 = (inp[12]) ? node20133 : 4'b0000;
															assign node20133 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node20136 = (inp[12]) ? node20138 : 4'b1000;
															assign node20138 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node20141 = (inp[7]) ? node20147 : node20142;
														assign node20142 = (inp[2]) ? 4'b0000 : node20143;
															assign node20143 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node20147 = (inp[12]) ? node20149 : 4'b0000;
															assign node20149 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node20152 = (inp[11]) ? node20216 : node20153;
											assign node20153 = (inp[1]) ? node20179 : node20154;
												assign node20154 = (inp[14]) ? node20164 : node20155;
													assign node20155 = (inp[2]) ? node20159 : node20156;
														assign node20156 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20159 = (inp[0]) ? node20161 : 4'b0000;
															assign node20161 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20164 = (inp[7]) ? node20168 : node20165;
														assign node20165 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node20168 = (inp[2]) ? node20174 : node20169;
															assign node20169 = (inp[12]) ? 4'b1000 : node20170;
																assign node20170 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node20174 = (inp[12]) ? node20176 : 4'b1001;
																assign node20176 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node20179 = (inp[0]) ? node20197 : node20180;
													assign node20180 = (inp[2]) ? node20192 : node20181;
														assign node20181 = (inp[7]) ? node20187 : node20182;
															assign node20182 = (inp[12]) ? 4'b0001 : node20183;
																assign node20183 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20187 = (inp[14]) ? node20189 : 4'b0000;
																assign node20189 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node20192 = (inp[7]) ? 4'b0001 : node20193;
															assign node20193 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node20197 = (inp[12]) ? node20207 : node20198;
														assign node20198 = (inp[7]) ? node20204 : node20199;
															assign node20199 = (inp[14]) ? node20201 : 4'b1000;
																assign node20201 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node20204 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20207 = (inp[2]) ? node20209 : 4'b0000;
															assign node20209 = (inp[7]) ? node20213 : node20210;
																assign node20210 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node20213 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node20216 = (inp[1]) ? 4'b0000 : node20217;
												assign node20217 = (inp[0]) ? node20225 : node20218;
													assign node20218 = (inp[14]) ? 4'b0000 : node20219;
														assign node20219 = (inp[2]) ? node20221 : 4'b0000;
															assign node20221 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node20225 = (inp[7]) ? node20231 : node20226;
														assign node20226 = (inp[2]) ? node20228 : 4'b0001;
															assign node20228 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node20231 = (inp[12]) ? 4'b0001 : node20232;
															assign node20232 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node20237 = (inp[11]) ? node20331 : node20238;
										assign node20238 = (inp[10]) ? node20292 : node20239;
											assign node20239 = (inp[0]) ? node20269 : node20240;
												assign node20240 = (inp[1]) ? node20256 : node20241;
													assign node20241 = (inp[7]) ? node20251 : node20242;
														assign node20242 = (inp[12]) ? 4'b0001 : node20243;
															assign node20243 = (inp[2]) ? node20247 : node20244;
																assign node20244 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node20247 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20251 = (inp[14]) ? node20253 : 4'b0000;
															assign node20253 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node20256 = (inp[12]) ? node20262 : node20257;
														assign node20257 = (inp[14]) ? node20259 : 4'b0000;
															assign node20259 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node20262 = (inp[2]) ? node20264 : 4'b0000;
															assign node20264 = (inp[14]) ? 4'b0000 : node20265;
																assign node20265 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node20269 = (inp[1]) ? node20281 : node20270;
													assign node20270 = (inp[7]) ? node20276 : node20271;
														assign node20271 = (inp[2]) ? node20273 : 4'b0000;
															assign node20273 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20276 = (inp[14]) ? node20278 : 4'b0001;
															assign node20278 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node20281 = (inp[7]) ? node20289 : node20282;
														assign node20282 = (inp[12]) ? node20284 : 4'b0001;
															assign node20284 = (inp[2]) ? node20286 : 4'b0001;
																assign node20286 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20289 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node20292 = (inp[1]) ? 4'b0000 : node20293;
												assign node20293 = (inp[12]) ? node20313 : node20294;
													assign node20294 = (inp[2]) ? node20306 : node20295;
														assign node20295 = (inp[7]) ? node20301 : node20296;
															assign node20296 = (inp[0]) ? node20298 : 4'b0001;
																assign node20298 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node20301 = (inp[0]) ? node20303 : 4'b0000;
																assign node20303 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20306 = (inp[7]) ? node20308 : 4'b0000;
															assign node20308 = (inp[0]) ? 4'b0000 : node20309;
																assign node20309 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node20313 = (inp[2]) ? node20323 : node20314;
														assign node20314 = (inp[7]) ? node20320 : node20315;
															assign node20315 = (inp[14]) ? 4'b0000 : node20316;
																assign node20316 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20320 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20323 = (inp[14]) ? node20325 : 4'b0001;
															assign node20325 = (inp[7]) ? node20327 : 4'b0001;
																assign node20327 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node20331 = (inp[1]) ? 4'b0000 : node20332;
											assign node20332 = (inp[10]) ? 4'b0000 : node20333;
												assign node20333 = (inp[0]) ? node20345 : node20334;
													assign node20334 = (inp[2]) ? node20340 : node20335;
														assign node20335 = (inp[12]) ? node20337 : 4'b0000;
															assign node20337 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node20340 = (inp[7]) ? 4'b0001 : node20341;
															assign node20341 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node20345 = (inp[12]) ? node20351 : node20346;
														assign node20346 = (inp[7]) ? 4'b0000 : node20347;
															assign node20347 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node20351 = (inp[7]) ? node20353 : 4'b0000;
															assign node20353 = (inp[14]) ? 4'b0000 : 4'b0001;
				assign node20358 = (inp[0]) ? node22220 : node20359;
					assign node20359 = (inp[6]) ? node20901 : node20360;
						assign node20360 = (inp[2]) ? node20804 : node20361;
							assign node20361 = (inp[5]) ? node20447 : node20362;
								assign node20362 = (inp[3]) ? node20364 : 4'b0010;
									assign node20364 = (inp[7]) ? node20428 : node20365;
										assign node20365 = (inp[4]) ? node20389 : node20366;
											assign node20366 = (inp[13]) ? node20368 : 4'b0010;
												assign node20368 = (inp[10]) ? node20374 : node20369;
													assign node20369 = (inp[1]) ? node20371 : 4'b0010;
														assign node20371 = (inp[14]) ? 4'b0010 : 4'b0000;
													assign node20374 = (inp[12]) ? node20386 : node20375;
														assign node20375 = (inp[1]) ? node20381 : node20376;
															assign node20376 = (inp[14]) ? node20378 : 4'b0001;
																assign node20378 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20381 = (inp[14]) ? node20383 : 4'b0000;
																assign node20383 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node20386 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node20389 = (inp[1]) ? node20413 : node20390;
												assign node20390 = (inp[13]) ? node20404 : node20391;
													assign node20391 = (inp[14]) ? node20397 : node20392;
														assign node20392 = (inp[10]) ? node20394 : 4'b0001;
															assign node20394 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20397 = (inp[11]) ? 4'b0001 : node20398;
															assign node20398 = (inp[12]) ? 4'b0000 : node20399;
																assign node20399 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node20404 = (inp[11]) ? 4'b1001 : node20405;
														assign node20405 = (inp[14]) ? 4'b1000 : node20406;
															assign node20406 = (inp[10]) ? node20408 : 4'b1001;
																assign node20408 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node20413 = (inp[13]) ? node20419 : node20414;
													assign node20414 = (inp[10]) ? 4'b1000 : node20415;
														assign node20415 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20419 = (inp[12]) ? node20425 : node20420;
														assign node20420 = (inp[11]) ? 4'b0000 : node20421;
															assign node20421 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20425 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node20428 = (inp[13]) ? node20430 : 4'b0010;
											assign node20430 = (inp[4]) ? node20432 : 4'b0010;
												assign node20432 = (inp[12]) ? 4'b0010 : node20433;
													assign node20433 = (inp[10]) ? node20437 : node20434;
														assign node20434 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node20437 = (inp[14]) ? node20439 : 4'b0000;
															assign node20439 = (inp[1]) ? node20443 : node20440;
																assign node20440 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node20443 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node20447 = (inp[1]) ? node20621 : node20448;
									assign node20448 = (inp[13]) ? node20536 : node20449;
										assign node20449 = (inp[11]) ? node20499 : node20450;
											assign node20450 = (inp[14]) ? node20476 : node20451;
												assign node20451 = (inp[10]) ? node20461 : node20452;
													assign node20452 = (inp[7]) ? node20458 : node20453;
														assign node20453 = (inp[12]) ? node20455 : 4'b0001;
															assign node20455 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node20458 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node20461 = (inp[12]) ? node20469 : node20462;
														assign node20462 = (inp[3]) ? node20464 : 4'b1001;
															assign node20464 = (inp[4]) ? node20466 : 4'b1101;
																assign node20466 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node20469 = (inp[4]) ? node20473 : node20470;
															assign node20470 = (inp[3]) ? 4'b0101 : 4'b0001;
															assign node20473 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node20476 = (inp[10]) ? node20488 : node20477;
													assign node20477 = (inp[3]) ? node20483 : node20478;
														assign node20478 = (inp[7]) ? 4'b0000 : node20479;
															assign node20479 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node20483 = (inp[4]) ? node20485 : 4'b0100;
															assign node20485 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node20488 = (inp[12]) ? node20496 : node20489;
														assign node20489 = (inp[4]) ? node20491 : 4'b1100;
															assign node20491 = (inp[3]) ? 4'b1000 : node20492;
																assign node20492 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node20496 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node20499 = (inp[3]) ? node20517 : node20500;
												assign node20500 = (inp[10]) ? node20506 : node20501;
													assign node20501 = (inp[4]) ? node20503 : 4'b0001;
														assign node20503 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node20506 = (inp[12]) ? node20512 : node20507;
														assign node20507 = (inp[4]) ? node20509 : 4'b1001;
															assign node20509 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node20512 = (inp[7]) ? 4'b0001 : node20513;
															assign node20513 = (inp[14]) ? 4'b0001 : 4'b0101;
												assign node20517 = (inp[4]) ? node20523 : node20518;
													assign node20518 = (inp[10]) ? node20520 : 4'b0101;
														assign node20520 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node20523 = (inp[7]) ? node20529 : node20524;
														assign node20524 = (inp[12]) ? 4'b0001 : node20525;
															assign node20525 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node20529 = (inp[14]) ? 4'b0101 : node20530;
															assign node20530 = (inp[10]) ? node20532 : 4'b0101;
																assign node20532 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node20536 = (inp[14]) ? node20564 : node20537;
											assign node20537 = (inp[10]) ? node20549 : node20538;
												assign node20538 = (inp[3]) ? node20544 : node20539;
													assign node20539 = (inp[4]) ? node20541 : 4'b1001;
														assign node20541 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node20544 = (inp[7]) ? 4'b1101 : node20545;
														assign node20545 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node20549 = (inp[12]) ? node20559 : node20550;
													assign node20550 = (inp[3]) ? node20554 : node20551;
														assign node20551 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node20554 = (inp[4]) ? 4'b0001 : node20555;
															assign node20555 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node20559 = (inp[3]) ? node20561 : 4'b1001;
														assign node20561 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node20564 = (inp[11]) ? node20596 : node20565;
												assign node20565 = (inp[10]) ? node20577 : node20566;
													assign node20566 = (inp[3]) ? node20572 : node20567;
														assign node20567 = (inp[4]) ? node20569 : 4'b1000;
															assign node20569 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node20572 = (inp[4]) ? node20574 : 4'b1100;
															assign node20574 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node20577 = (inp[12]) ? node20587 : node20578;
														assign node20578 = (inp[4]) ? 4'b0000 : node20579;
															assign node20579 = (inp[3]) ? node20583 : node20580;
																assign node20580 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node20583 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node20587 = (inp[4]) ? node20591 : node20588;
															assign node20588 = (inp[3]) ? 4'b1100 : 4'b1000;
															assign node20591 = (inp[3]) ? 4'b1000 : node20592;
																assign node20592 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node20596 = (inp[10]) ? node20608 : node20597;
													assign node20597 = (inp[3]) ? node20603 : node20598;
														assign node20598 = (inp[4]) ? node20600 : 4'b1001;
															assign node20600 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node20603 = (inp[4]) ? node20605 : 4'b1101;
															assign node20605 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node20608 = (inp[12]) ? node20612 : node20609;
														assign node20609 = (inp[3]) ? 4'b0001 : 4'b0101;
														assign node20612 = (inp[4]) ? node20614 : 4'b1001;
															assign node20614 = (inp[7]) ? node20618 : node20615;
																assign node20615 = (inp[3]) ? 4'b1001 : 4'b1101;
																assign node20618 = (inp[3]) ? 4'b1101 : 4'b1001;
									assign node20621 = (inp[11]) ? node20731 : node20622;
										assign node20622 = (inp[14]) ? node20674 : node20623;
											assign node20623 = (inp[13]) ? node20649 : node20624;
												assign node20624 = (inp[3]) ? node20638 : node20625;
													assign node20625 = (inp[12]) ? node20631 : node20626;
														assign node20626 = (inp[4]) ? node20628 : 4'b1000;
															assign node20628 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node20631 = (inp[10]) ? node20633 : 4'b0000;
															assign node20633 = (inp[4]) ? node20635 : 4'b1000;
																assign node20635 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node20638 = (inp[10]) ? 4'b1100 : node20639;
														assign node20639 = (inp[12]) ? node20645 : node20640;
															assign node20640 = (inp[7]) ? 4'b1100 : node20641;
																assign node20641 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node20645 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node20649 = (inp[10]) ? node20663 : node20650;
													assign node20650 = (inp[12]) ? node20654 : node20651;
														assign node20651 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node20654 = (inp[7]) ? node20660 : node20655;
															assign node20655 = (inp[3]) ? 4'b1000 : node20656;
																assign node20656 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node20660 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node20663 = (inp[3]) ? node20669 : node20664;
														assign node20664 = (inp[4]) ? 4'b0100 : node20665;
															assign node20665 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20669 = (inp[7]) ? node20671 : 4'b0000;
															assign node20671 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node20674 = (inp[13]) ? node20708 : node20675;
												assign node20675 = (inp[10]) ? node20689 : node20676;
													assign node20676 = (inp[3]) ? node20684 : node20677;
														assign node20677 = (inp[12]) ? node20679 : 4'b0001;
															assign node20679 = (inp[4]) ? node20681 : 4'b0001;
																assign node20681 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node20684 = (inp[7]) ? 4'b0101 : node20685;
															assign node20685 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node20689 = (inp[12]) ? node20701 : node20690;
														assign node20690 = (inp[3]) ? node20696 : node20691;
															assign node20691 = (inp[7]) ? 4'b1001 : node20692;
																assign node20692 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node20696 = (inp[4]) ? node20698 : 4'b1101;
																assign node20698 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node20701 = (inp[7]) ? node20705 : node20702;
															assign node20702 = (inp[3]) ? 4'b0001 : 4'b0101;
															assign node20705 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node20708 = (inp[10]) ? node20720 : node20709;
													assign node20709 = (inp[3]) ? node20715 : node20710;
														assign node20710 = (inp[7]) ? 4'b1001 : node20711;
															assign node20711 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node20715 = (inp[7]) ? 4'b1101 : node20716;
															assign node20716 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node20720 = (inp[12]) ? node20728 : node20721;
														assign node20721 = (inp[3]) ? node20725 : node20722;
															assign node20722 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node20725 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node20728 = (inp[3]) ? 4'b1101 : 4'b1001;
										assign node20731 = (inp[13]) ? node20765 : node20732;
											assign node20732 = (inp[10]) ? node20754 : node20733;
												assign node20733 = (inp[12]) ? node20743 : node20734;
													assign node20734 = (inp[3]) ? node20736 : 4'b1000;
														assign node20736 = (inp[14]) ? node20738 : 4'b1000;
															assign node20738 = (inp[7]) ? 4'b1100 : node20739;
																assign node20739 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node20743 = (inp[3]) ? node20749 : node20744;
														assign node20744 = (inp[7]) ? 4'b0000 : node20745;
															assign node20745 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node20749 = (inp[4]) ? node20751 : 4'b0100;
															assign node20751 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node20754 = (inp[3]) ? node20760 : node20755;
													assign node20755 = (inp[4]) ? node20757 : 4'b1000;
														assign node20757 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node20760 = (inp[4]) ? node20762 : 4'b1100;
														assign node20762 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node20765 = (inp[12]) ? node20777 : node20766;
												assign node20766 = (inp[3]) ? node20772 : node20767;
													assign node20767 = (inp[4]) ? 4'b0100 : node20768;
														assign node20768 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node20772 = (inp[4]) ? 4'b0000 : node20773;
														assign node20773 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node20777 = (inp[10]) ? node20795 : node20778;
													assign node20778 = (inp[4]) ? node20782 : node20779;
														assign node20779 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node20782 = (inp[14]) ? node20788 : node20783;
															assign node20783 = (inp[3]) ? node20785 : 4'b1100;
																assign node20785 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node20788 = (inp[7]) ? node20792 : node20789;
																assign node20789 = (inp[3]) ? 4'b1000 : 4'b1100;
																assign node20792 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node20795 = (inp[4]) ? 4'b0100 : node20796;
														assign node20796 = (inp[7]) ? node20800 : node20797;
															assign node20797 = (inp[3]) ? 4'b0000 : 4'b0100;
															assign node20800 = (inp[3]) ? 4'b0100 : 4'b0000;
							assign node20804 = (inp[3]) ? node20806 : 4'b0010;
								assign node20806 = (inp[5]) ? node20808 : 4'b0010;
									assign node20808 = (inp[4]) ? node20832 : node20809;
										assign node20809 = (inp[13]) ? node20811 : 4'b0010;
											assign node20811 = (inp[7]) ? 4'b0010 : node20812;
												assign node20812 = (inp[12]) ? node20822 : node20813;
													assign node20813 = (inp[10]) ? node20819 : node20814;
														assign node20814 = (inp[1]) ? node20816 : 4'b0010;
															assign node20816 = (inp[14]) ? 4'b0010 : 4'b0000;
														assign node20819 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node20822 = (inp[1]) ? node20824 : 4'b0010;
														assign node20824 = (inp[10]) ? node20826 : 4'b0010;
															assign node20826 = (inp[11]) ? 4'b0000 : node20827;
																assign node20827 = (inp[14]) ? 4'b0010 : 4'b0000;
										assign node20832 = (inp[7]) ? node20880 : node20833;
											assign node20833 = (inp[1]) ? node20861 : node20834;
												assign node20834 = (inp[11]) ? node20850 : node20835;
													assign node20835 = (inp[14]) ? node20839 : node20836;
														assign node20836 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node20839 = (inp[13]) ? node20845 : node20840;
															assign node20840 = (inp[12]) ? 4'b0000 : node20841;
																assign node20841 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node20845 = (inp[12]) ? 4'b1000 : node20846;
																assign node20846 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node20850 = (inp[13]) ? node20856 : node20851;
														assign node20851 = (inp[10]) ? node20853 : 4'b0001;
															assign node20853 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20856 = (inp[12]) ? 4'b1001 : node20857;
															assign node20857 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node20861 = (inp[14]) ? node20871 : node20862;
													assign node20862 = (inp[10]) ? node20868 : node20863;
														assign node20863 = (inp[12]) ? node20865 : 4'b1000;
															assign node20865 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node20868 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node20871 = (inp[11]) ? node20875 : node20872;
														assign node20872 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20875 = (inp[13]) ? node20877 : 4'b1000;
															assign node20877 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node20880 = (inp[13]) ? node20882 : 4'b0010;
												assign node20882 = (inp[12]) ? node20894 : node20883;
													assign node20883 = (inp[10]) ? node20889 : node20884;
														assign node20884 = (inp[14]) ? 4'b0010 : node20885;
															assign node20885 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node20889 = (inp[1]) ? node20891 : 4'b0001;
															assign node20891 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node20894 = (inp[11]) ? node20896 : 4'b0010;
														assign node20896 = (inp[10]) ? node20898 : 4'b0010;
															assign node20898 = (inp[1]) ? 4'b0000 : 4'b0010;
						assign node20901 = (inp[5]) ? node21513 : node20902;
							assign node20902 = (inp[1]) ? node21196 : node20903;
								assign node20903 = (inp[3]) ? node21035 : node20904;
									assign node20904 = (inp[13]) ? node20952 : node20905;
										assign node20905 = (inp[14]) ? node20923 : node20906;
											assign node20906 = (inp[12]) ? node20918 : node20907;
												assign node20907 = (inp[10]) ? node20913 : node20908;
													assign node20908 = (inp[4]) ? node20910 : 4'b0001;
														assign node20910 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node20913 = (inp[7]) ? 4'b1001 : node20914;
														assign node20914 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node20918 = (inp[7]) ? 4'b0001 : node20919;
													assign node20919 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node20923 = (inp[11]) ? node20937 : node20924;
												assign node20924 = (inp[7]) ? node20932 : node20925;
													assign node20925 = (inp[4]) ? node20927 : 4'b0000;
														assign node20927 = (inp[12]) ? 4'b0100 : node20928;
															assign node20928 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node20932 = (inp[12]) ? 4'b0000 : node20933;
														assign node20933 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node20937 = (inp[7]) ? node20947 : node20938;
													assign node20938 = (inp[4]) ? node20942 : node20939;
														assign node20939 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node20942 = (inp[12]) ? 4'b0101 : node20943;
															assign node20943 = (inp[10]) ? 4'b0000 : 4'b0101;
													assign node20947 = (inp[10]) ? node20949 : 4'b0001;
														assign node20949 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node20952 = (inp[12]) ? node20998 : node20953;
											assign node20953 = (inp[10]) ? node20979 : node20954;
												assign node20954 = (inp[14]) ? node20966 : node20955;
													assign node20955 = (inp[2]) ? node20961 : node20956;
														assign node20956 = (inp[4]) ? node20958 : 4'b1001;
															assign node20958 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node20961 = (inp[4]) ? node20963 : 4'b1001;
															assign node20963 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node20966 = (inp[11]) ? node20974 : node20967;
														assign node20967 = (inp[7]) ? 4'b1000 : node20968;
															assign node20968 = (inp[2]) ? 4'b1100 : node20969;
																assign node20969 = (inp[4]) ? 4'b0001 : 4'b1000;
														assign node20974 = (inp[4]) ? node20976 : 4'b1001;
															assign node20976 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node20979 = (inp[7]) ? node20987 : node20980;
													assign node20980 = (inp[11]) ? 4'b0101 : node20981;
														assign node20981 = (inp[2]) ? 4'b0100 : node20982;
															assign node20982 = (inp[4]) ? 4'b1001 : 4'b0100;
													assign node20987 = (inp[4]) ? node20993 : node20988;
														assign node20988 = (inp[11]) ? 4'b0001 : node20989;
															assign node20989 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20993 = (inp[11]) ? 4'b0000 : node20994;
															assign node20994 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node20998 = (inp[14]) ? node21010 : node20999;
												assign node20999 = (inp[4]) ? node21001 : 4'b1001;
													assign node21001 = (inp[7]) ? 4'b1001 : node21002;
														assign node21002 = (inp[2]) ? 4'b1101 : node21003;
															assign node21003 = (inp[11]) ? node21005 : 4'b1001;
																assign node21005 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node21010 = (inp[11]) ? node21024 : node21011;
													assign node21011 = (inp[2]) ? node21019 : node21012;
														assign node21012 = (inp[4]) ? node21014 : 4'b1000;
															assign node21014 = (inp[7]) ? 4'b1000 : node21015;
																assign node21015 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node21019 = (inp[10]) ? 4'b1000 : node21020;
															assign node21020 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node21024 = (inp[7]) ? 4'b1001 : node21025;
														assign node21025 = (inp[2]) ? node21031 : node21026;
															assign node21026 = (inp[4]) ? node21028 : 4'b1001;
																assign node21028 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node21031 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node21035 = (inp[10]) ? node21105 : node21036;
										assign node21036 = (inp[11]) ? node21068 : node21037;
											assign node21037 = (inp[2]) ? node21049 : node21038;
												assign node21038 = (inp[4]) ? node21044 : node21039;
													assign node21039 = (inp[13]) ? node21041 : 4'b0001;
														assign node21041 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node21044 = (inp[7]) ? 4'b0101 : node21045;
														assign node21045 = (inp[14]) ? 4'b0101 : 4'b0000;
												assign node21049 = (inp[14]) ? node21057 : node21050;
													assign node21050 = (inp[13]) ? node21052 : 4'b0101;
														assign node21052 = (inp[7]) ? 4'b1101 : node21053;
															assign node21053 = (inp[4]) ? 4'b0001 : 4'b1101;
													assign node21057 = (inp[7]) ? node21065 : node21058;
														assign node21058 = (inp[4]) ? node21062 : node21059;
															assign node21059 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node21062 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node21065 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node21068 = (inp[2]) ? node21092 : node21069;
												assign node21069 = (inp[12]) ? node21081 : node21070;
													assign node21070 = (inp[4]) ? node21076 : node21071;
														assign node21071 = (inp[7]) ? 4'b1000 : node21072;
															assign node21072 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node21076 = (inp[13]) ? node21078 : 4'b1100;
															assign node21078 = (inp[7]) ? 4'b1100 : 4'b0001;
													assign node21081 = (inp[4]) ? node21087 : node21082;
														assign node21082 = (inp[13]) ? node21084 : 4'b0000;
															assign node21084 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21087 = (inp[7]) ? 4'b0100 : node21088;
															assign node21088 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node21092 = (inp[13]) ? node21098 : node21093;
													assign node21093 = (inp[7]) ? 4'b0101 : node21094;
														assign node21094 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node21098 = (inp[7]) ? 4'b1101 : node21099;
														assign node21099 = (inp[4]) ? node21101 : 4'b1101;
															assign node21101 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node21105 = (inp[11]) ? node21155 : node21106;
											assign node21106 = (inp[2]) ? node21120 : node21107;
												assign node21107 = (inp[4]) ? node21113 : node21108;
													assign node21108 = (inp[7]) ? 4'b1001 : node21109;
														assign node21109 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node21113 = (inp[7]) ? 4'b1101 : node21114;
														assign node21114 = (inp[13]) ? node21116 : 4'b1101;
															assign node21116 = (inp[12]) ? 4'b0001 : 4'b1000;
												assign node21120 = (inp[14]) ? node21138 : node21121;
													assign node21121 = (inp[4]) ? node21131 : node21122;
														assign node21122 = (inp[7]) ? node21124 : 4'b1101;
															assign node21124 = (inp[13]) ? node21128 : node21125;
																assign node21125 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node21128 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node21131 = (inp[7]) ? node21133 : 4'b1001;
															assign node21133 = (inp[12]) ? 4'b1101 : node21134;
																assign node21134 = (inp[13]) ? 4'b0001 : 4'b1101;
													assign node21138 = (inp[4]) ? node21148 : node21139;
														assign node21139 = (inp[13]) ? node21143 : node21140;
															assign node21140 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node21143 = (inp[12]) ? 4'b1100 : node21144;
																assign node21144 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node21148 = (inp[7]) ? 4'b1100 : node21149;
															assign node21149 = (inp[13]) ? 4'b1001 : node21150;
																assign node21150 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node21155 = (inp[2]) ? node21179 : node21156;
												assign node21156 = (inp[12]) ? node21168 : node21157;
													assign node21157 = (inp[4]) ? node21163 : node21158;
														assign node21158 = (inp[7]) ? node21160 : 4'b0100;
															assign node21160 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node21163 = (inp[13]) ? node21165 : 4'b0000;
															assign node21165 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node21168 = (inp[4]) ? node21174 : node21169;
														assign node21169 = (inp[13]) ? node21171 : 4'b1000;
															assign node21171 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node21174 = (inp[13]) ? node21176 : 4'b1100;
															assign node21176 = (inp[7]) ? 4'b1100 : 4'b1001;
												assign node21179 = (inp[4]) ? node21189 : node21180;
													assign node21180 = (inp[13]) ? node21184 : node21181;
														assign node21181 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node21184 = (inp[12]) ? 4'b1101 : node21185;
															assign node21185 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node21189 = (inp[12]) ? node21191 : 4'b0000;
														assign node21191 = (inp[7]) ? node21193 : 4'b1000;
															assign node21193 = (inp[13]) ? 4'b1101 : 4'b0101;
								assign node21196 = (inp[11]) ? node21416 : node21197;
									assign node21197 = (inp[14]) ? node21311 : node21198;
										assign node21198 = (inp[3]) ? node21250 : node21199;
											assign node21199 = (inp[4]) ? node21213 : node21200;
												assign node21200 = (inp[13]) ? node21206 : node21201;
													assign node21201 = (inp[10]) ? 4'b1000 : node21202;
														assign node21202 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node21206 = (inp[12]) ? node21210 : node21207;
														assign node21207 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21210 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node21213 = (inp[2]) ? node21237 : node21214;
													assign node21214 = (inp[12]) ? node21228 : node21215;
														assign node21215 = (inp[10]) ? node21223 : node21216;
															assign node21216 = (inp[7]) ? node21220 : node21217;
																assign node21217 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node21220 = (inp[13]) ? 4'b0100 : 4'b1000;
															assign node21223 = (inp[7]) ? node21225 : 4'b0001;
																assign node21225 = (inp[13]) ? 4'b0001 : 4'b1000;
														assign node21228 = (inp[7]) ? node21232 : node21229;
															assign node21229 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node21232 = (inp[10]) ? node21234 : 4'b1000;
																assign node21234 = (inp[13]) ? 4'b0100 : 4'b1000;
													assign node21237 = (inp[13]) ? node21243 : node21238;
														assign node21238 = (inp[10]) ? 4'b1100 : node21239;
															assign node21239 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node21243 = (inp[10]) ? 4'b0100 : node21244;
															assign node21244 = (inp[12]) ? node21246 : 4'b0100;
																assign node21246 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node21250 = (inp[2]) ? node21284 : node21251;
												assign node21251 = (inp[4]) ? node21271 : node21252;
													assign node21252 = (inp[13]) ? node21262 : node21253;
														assign node21253 = (inp[7]) ? 4'b0001 : node21254;
															assign node21254 = (inp[12]) ? node21258 : node21255;
																assign node21255 = (inp[10]) ? 4'b0101 : 4'b1001;
																assign node21258 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node21262 = (inp[7]) ? node21264 : 4'b0101;
															assign node21264 = (inp[12]) ? node21268 : node21265;
																assign node21265 = (inp[10]) ? 4'b0101 : 4'b1001;
																assign node21268 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node21271 = (inp[7]) ? node21277 : node21272;
														assign node21272 = (inp[13]) ? 4'b0001 : node21273;
															assign node21273 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node21277 = (inp[12]) ? node21281 : node21278;
															assign node21278 = (inp[10]) ? 4'b0001 : 4'b1101;
															assign node21281 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node21284 = (inp[4]) ? node21296 : node21285;
													assign node21285 = (inp[12]) ? node21291 : node21286;
														assign node21286 = (inp[13]) ? node21288 : 4'b1100;
															assign node21288 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node21291 = (inp[13]) ? 4'b1100 : node21292;
															assign node21292 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node21296 = (inp[7]) ? node21308 : node21297;
														assign node21297 = (inp[13]) ? node21305 : node21298;
															assign node21298 = (inp[12]) ? node21302 : node21299;
																assign node21299 = (inp[10]) ? 4'b0001 : 4'b1000;
																assign node21302 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node21305 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21308 = (inp[12]) ? 4'b0000 : 4'b1100;
										assign node21311 = (inp[13]) ? node21351 : node21312;
											assign node21312 = (inp[3]) ? node21330 : node21313;
												assign node21313 = (inp[10]) ? node21319 : node21314;
													assign node21314 = (inp[7]) ? 4'b0001 : node21315;
														assign node21315 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node21319 = (inp[12]) ? node21325 : node21320;
														assign node21320 = (inp[4]) ? node21322 : 4'b1001;
															assign node21322 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node21325 = (inp[7]) ? 4'b0001 : node21326;
															assign node21326 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node21330 = (inp[2]) ? node21346 : node21331;
													assign node21331 = (inp[4]) ? node21337 : node21332;
														assign node21332 = (inp[10]) ? 4'b0101 : node21333;
															assign node21333 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21337 = (inp[12]) ? node21343 : node21338;
															assign node21338 = (inp[10]) ? node21340 : 4'b1101;
																assign node21340 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node21343 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node21346 = (inp[7]) ? 4'b0101 : node21347;
														assign node21347 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node21351 = (inp[12]) ? node21387 : node21352;
												assign node21352 = (inp[10]) ? node21364 : node21353;
													assign node21353 = (inp[3]) ? node21359 : node21354;
														assign node21354 = (inp[4]) ? node21356 : 4'b1001;
															assign node21356 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node21359 = (inp[7]) ? 4'b1101 : node21360;
															assign node21360 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node21364 = (inp[4]) ? node21378 : node21365;
														assign node21365 = (inp[2]) ? node21371 : node21366;
															assign node21366 = (inp[7]) ? node21368 : 4'b0101;
																assign node21368 = (inp[3]) ? 4'b0101 : 4'b0001;
															assign node21371 = (inp[3]) ? node21375 : node21372;
																assign node21372 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node21375 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node21378 = (inp[7]) ? node21382 : node21379;
															assign node21379 = (inp[3]) ? 4'b0001 : 4'b0101;
															assign node21382 = (inp[2]) ? 4'b0001 : node21383;
																assign node21383 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node21387 = (inp[2]) ? node21405 : node21388;
													assign node21388 = (inp[10]) ? node21398 : node21389;
														assign node21389 = (inp[3]) ? node21393 : node21390;
															assign node21390 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node21393 = (inp[7]) ? node21395 : 4'b0000;
																assign node21395 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node21398 = (inp[4]) ? 4'b1000 : node21399;
															assign node21399 = (inp[3]) ? node21401 : 4'b1001;
																assign node21401 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node21405 = (inp[3]) ? node21411 : node21406;
														assign node21406 = (inp[4]) ? node21408 : 4'b1001;
															assign node21408 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node21411 = (inp[4]) ? node21413 : 4'b1101;
															assign node21413 = (inp[7]) ? 4'b1101 : 4'b1001;
									assign node21416 = (inp[10]) ? node21476 : node21417;
										assign node21417 = (inp[3]) ? node21449 : node21418;
											assign node21418 = (inp[7]) ? node21434 : node21419;
												assign node21419 = (inp[4]) ? node21427 : node21420;
													assign node21420 = (inp[13]) ? node21424 : node21421;
														assign node21421 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21424 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node21427 = (inp[13]) ? node21431 : node21428;
														assign node21428 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node21431 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node21434 = (inp[4]) ? node21442 : node21435;
													assign node21435 = (inp[13]) ? node21439 : node21436;
														assign node21436 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21439 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node21442 = (inp[12]) ? node21446 : node21443;
														assign node21443 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node21446 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node21449 = (inp[2]) ? node21457 : node21450;
												assign node21450 = (inp[4]) ? 4'b1100 : node21451;
													assign node21451 = (inp[13]) ? node21453 : 4'b1000;
														assign node21453 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node21457 = (inp[7]) ? node21463 : node21458;
													assign node21458 = (inp[4]) ? 4'b1000 : node21459;
														assign node21459 = (inp[13]) ? 4'b0000 : 4'b1100;
													assign node21463 = (inp[4]) ? node21471 : node21464;
														assign node21464 = (inp[13]) ? node21468 : node21465;
															assign node21465 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node21468 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node21471 = (inp[12]) ? node21473 : 4'b0000;
															assign node21473 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node21476 = (inp[13]) ? node21498 : node21477;
											assign node21477 = (inp[3]) ? node21485 : node21478;
												assign node21478 = (inp[4]) ? node21480 : 4'b1000;
													assign node21480 = (inp[7]) ? 4'b1000 : node21481;
														assign node21481 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node21485 = (inp[2]) ? node21493 : node21486;
													assign node21486 = (inp[4]) ? node21490 : node21487;
														assign node21487 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21490 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node21493 = (inp[7]) ? 4'b1100 : node21494;
														assign node21494 = (inp[4]) ? 4'b0000 : 4'b1100;
											assign node21498 = (inp[4]) ? node21508 : node21499;
												assign node21499 = (inp[3]) ? node21503 : node21500;
													assign node21500 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node21503 = (inp[7]) ? 4'b0100 : node21504;
														assign node21504 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node21508 = (inp[3]) ? 4'b0000 : node21509;
													assign node21509 = (inp[2]) ? 4'b0100 : 4'b0000;
							assign node21513 = (inp[3]) ? node21867 : node21514;
								assign node21514 = (inp[11]) ? node21726 : node21515;
									assign node21515 = (inp[2]) ? node21623 : node21516;
										assign node21516 = (inp[4]) ? node21578 : node21517;
											assign node21517 = (inp[13]) ? node21547 : node21518;
												assign node21518 = (inp[7]) ? node21534 : node21519;
													assign node21519 = (inp[10]) ? node21525 : node21520;
														assign node21520 = (inp[1]) ? 4'b1000 : node21521;
															assign node21521 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21525 = (inp[1]) ? node21531 : node21526;
															assign node21526 = (inp[14]) ? node21528 : 4'b0100;
																assign node21528 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node21531 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node21534 = (inp[10]) ? node21540 : node21535;
														assign node21535 = (inp[1]) ? 4'b1001 : node21536;
															assign node21536 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21540 = (inp[12]) ? node21544 : node21541;
															assign node21541 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21544 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node21547 = (inp[10]) ? node21561 : node21548;
													assign node21548 = (inp[1]) ? node21554 : node21549;
														assign node21549 = (inp[14]) ? 4'b1101 : node21550;
															assign node21550 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node21554 = (inp[14]) ? node21556 : 4'b0101;
															assign node21556 = (inp[12]) ? 4'b0100 : node21557;
																assign node21557 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node21561 = (inp[7]) ? node21569 : node21562;
														assign node21562 = (inp[1]) ? node21566 : node21563;
															assign node21563 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21566 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node21569 = (inp[12]) ? node21575 : node21570;
															assign node21570 = (inp[1]) ? 4'b0000 : node21571;
																assign node21571 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21575 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node21578 = (inp[13]) ? node21600 : node21579;
												assign node21579 = (inp[12]) ? node21589 : node21580;
													assign node21580 = (inp[1]) ? node21584 : node21581;
														assign node21581 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node21584 = (inp[10]) ? node21586 : 4'b0100;
															assign node21586 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node21589 = (inp[1]) ? node21593 : node21590;
														assign node21590 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21593 = (inp[7]) ? 4'b1000 : node21594;
															assign node21594 = (inp[10]) ? node21596 : 4'b1000;
																assign node21596 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node21600 = (inp[1]) ? node21618 : node21601;
													assign node21601 = (inp[14]) ? node21611 : node21602;
														assign node21602 = (inp[12]) ? node21604 : 4'b0001;
															assign node21604 = (inp[10]) ? node21608 : node21605;
																assign node21605 = (inp[7]) ? 4'b0100 : 4'b1001;
																assign node21608 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node21611 = (inp[7]) ? node21613 : 4'b1000;
															assign node21613 = (inp[12]) ? node21615 : 4'b0000;
																assign node21615 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node21618 = (inp[14]) ? 4'b1001 : node21619;
														assign node21619 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node21623 = (inp[4]) ? node21661 : node21624;
											assign node21624 = (inp[10]) ? node21642 : node21625;
												assign node21625 = (inp[13]) ? node21631 : node21626;
													assign node21626 = (inp[1]) ? node21628 : 4'b0001;
														assign node21628 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node21631 = (inp[7]) ? node21637 : node21632;
														assign node21632 = (inp[12]) ? 4'b0101 : node21633;
															assign node21633 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node21637 = (inp[1]) ? node21639 : 4'b0001;
															assign node21639 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node21642 = (inp[12]) ? node21656 : node21643;
													assign node21643 = (inp[1]) ? node21649 : node21644;
														assign node21644 = (inp[7]) ? 4'b1001 : node21645;
															assign node21645 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node21649 = (inp[13]) ? node21653 : node21650;
															assign node21650 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node21653 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node21656 = (inp[13]) ? node21658 : 4'b1001;
														assign node21658 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node21661 = (inp[10]) ? node21691 : node21662;
												assign node21662 = (inp[13]) ? node21674 : node21663;
													assign node21663 = (inp[7]) ? node21669 : node21664;
														assign node21664 = (inp[1]) ? node21666 : 4'b0001;
															assign node21666 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node21669 = (inp[1]) ? node21671 : 4'b0101;
															assign node21671 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21674 = (inp[1]) ? node21680 : node21675;
														assign node21675 = (inp[14]) ? 4'b1001 : node21676;
															assign node21676 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node21680 = (inp[14]) ? node21688 : node21681;
															assign node21681 = (inp[12]) ? node21685 : node21682;
																assign node21682 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node21685 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node21688 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node21691 = (inp[13]) ? node21703 : node21692;
													assign node21692 = (inp[14]) ? node21696 : node21693;
														assign node21693 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node21696 = (inp[1]) ? node21700 : node21697;
															assign node21697 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node21700 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node21703 = (inp[7]) ? node21719 : node21704;
														assign node21704 = (inp[14]) ? node21712 : node21705;
															assign node21705 = (inp[12]) ? node21709 : node21706;
																assign node21706 = (inp[1]) ? 4'b0000 : 4'b1000;
																assign node21709 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node21712 = (inp[12]) ? node21716 : node21713;
																assign node21713 = (inp[1]) ? 4'b0000 : 4'b1000;
																assign node21716 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node21719 = (inp[1]) ? 4'b1000 : node21720;
															assign node21720 = (inp[12]) ? 4'b0001 : node21721;
																assign node21721 = (inp[14]) ? 4'b1001 : 4'b1000;
									assign node21726 = (inp[1]) ? node21804 : node21727;
										assign node21727 = (inp[4]) ? node21769 : node21728;
											assign node21728 = (inp[2]) ? node21744 : node21729;
												assign node21729 = (inp[13]) ? node21737 : node21730;
													assign node21730 = (inp[10]) ? node21734 : node21731;
														assign node21731 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21734 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node21737 = (inp[10]) ? node21741 : node21738;
														assign node21738 = (inp[7]) ? 4'b1001 : 4'b0101;
														assign node21741 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node21744 = (inp[13]) ? node21754 : node21745;
													assign node21745 = (inp[12]) ? node21751 : node21746;
														assign node21746 = (inp[10]) ? node21748 : 4'b1000;
															assign node21748 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21751 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node21754 = (inp[7]) ? node21762 : node21755;
														assign node21755 = (inp[12]) ? node21759 : node21756;
															assign node21756 = (inp[10]) ? 4'b0100 : 4'b1100;
															assign node21759 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node21762 = (inp[10]) ? node21766 : node21763;
															assign node21763 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21766 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node21769 = (inp[13]) ? node21785 : node21770;
												assign node21770 = (inp[2]) ? node21778 : node21771;
													assign node21771 = (inp[7]) ? 4'b1000 : node21772;
														assign node21772 = (inp[12]) ? node21774 : 4'b0001;
															assign node21774 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node21778 = (inp[10]) ? 4'b0001 : node21779;
														assign node21779 = (inp[7]) ? node21781 : 4'b0001;
															assign node21781 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node21785 = (inp[10]) ? node21793 : node21786;
													assign node21786 = (inp[2]) ? node21788 : 4'b0001;
														assign node21788 = (inp[12]) ? 4'b1001 : node21789;
															assign node21789 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node21793 = (inp[7]) ? node21799 : node21794;
														assign node21794 = (inp[2]) ? 4'b1000 : node21795;
															assign node21795 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21799 = (inp[2]) ? 4'b1001 : node21800;
															assign node21800 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node21804 = (inp[13]) ? node21840 : node21805;
											assign node21805 = (inp[2]) ? node21825 : node21806;
												assign node21806 = (inp[4]) ? node21816 : node21807;
													assign node21807 = (inp[7]) ? 4'b1000 : node21808;
														assign node21808 = (inp[12]) ? node21812 : node21809;
															assign node21809 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node21812 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node21816 = (inp[12]) ? node21818 : 4'b0100;
														assign node21818 = (inp[7]) ? node21822 : node21819;
															assign node21819 = (inp[14]) ? 4'b0100 : 4'b1000;
															assign node21822 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node21825 = (inp[4]) ? node21831 : node21826;
													assign node21826 = (inp[10]) ? node21828 : 4'b1000;
														assign node21828 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node21831 = (inp[12]) ? node21835 : node21832;
														assign node21832 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node21835 = (inp[10]) ? 4'b1000 : node21836;
															assign node21836 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node21840 = (inp[10]) ? node21862 : node21841;
												assign node21841 = (inp[4]) ? node21851 : node21842;
													assign node21842 = (inp[2]) ? node21848 : node21843;
														assign node21843 = (inp[7]) ? node21845 : 4'b0000;
															assign node21845 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node21848 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node21851 = (inp[12]) ? node21859 : node21852;
														assign node21852 = (inp[2]) ? node21856 : node21853;
															assign node21853 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node21856 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node21859 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node21862 = (inp[7]) ? node21864 : 4'b0000;
													assign node21864 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node21867 = (inp[11]) ? node22093 : node21868;
									assign node21868 = (inp[4]) ? node21976 : node21869;
										assign node21869 = (inp[12]) ? node21933 : node21870;
											assign node21870 = (inp[13]) ? node21902 : node21871;
												assign node21871 = (inp[1]) ? node21885 : node21872;
													assign node21872 = (inp[2]) ? node21880 : node21873;
														assign node21873 = (inp[14]) ? node21877 : node21874;
															assign node21874 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node21877 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node21880 = (inp[14]) ? 4'b1000 : node21881;
															assign node21881 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node21885 = (inp[14]) ? node21895 : node21886;
														assign node21886 = (inp[2]) ? node21892 : node21887;
															assign node21887 = (inp[7]) ? 4'b0001 : node21888;
																assign node21888 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node21892 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node21895 = (inp[2]) ? 4'b0001 : node21896;
															assign node21896 = (inp[7]) ? node21898 : 4'b1000;
																assign node21898 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21902 = (inp[1]) ? node21918 : node21903;
													assign node21903 = (inp[10]) ? node21911 : node21904;
														assign node21904 = (inp[14]) ? node21908 : node21905;
															assign node21905 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node21908 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node21911 = (inp[14]) ? 4'b0001 : node21912;
															assign node21912 = (inp[7]) ? node21914 : 4'b0000;
																assign node21914 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node21918 = (inp[10]) ? node21928 : node21919;
														assign node21919 = (inp[2]) ? node21923 : node21920;
															assign node21920 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node21923 = (inp[7]) ? 4'b0001 : node21924;
																assign node21924 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node21928 = (inp[7]) ? node21930 : 4'b1000;
															assign node21930 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node21933 = (inp[2]) ? node21955 : node21934;
												assign node21934 = (inp[7]) ? node21948 : node21935;
													assign node21935 = (inp[1]) ? node21943 : node21936;
														assign node21936 = (inp[14]) ? node21940 : node21937;
															assign node21937 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node21940 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node21943 = (inp[13]) ? 4'b0000 : node21944;
															assign node21944 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node21948 = (inp[13]) ? node21950 : 4'b0001;
														assign node21950 = (inp[10]) ? 4'b0001 : node21951;
															assign node21951 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node21955 = (inp[13]) ? node21971 : node21956;
													assign node21956 = (inp[10]) ? node21964 : node21957;
														assign node21957 = (inp[1]) ? node21959 : 4'b0000;
															assign node21959 = (inp[14]) ? 4'b1000 : node21960;
																assign node21960 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node21964 = (inp[1]) ? node21968 : node21965;
															assign node21965 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node21968 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node21971 = (inp[10]) ? node21973 : 4'b0001;
														assign node21973 = (inp[1]) ? 4'b1000 : 4'b1001;
										assign node21976 = (inp[13]) ? node22040 : node21977;
											assign node21977 = (inp[10]) ? node22005 : node21978;
												assign node21978 = (inp[12]) ? node21996 : node21979;
													assign node21979 = (inp[2]) ? node21991 : node21980;
														assign node21980 = (inp[14]) ? node21986 : node21981;
															assign node21981 = (inp[7]) ? 4'b0001 : node21982;
																assign node21982 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node21986 = (inp[7]) ? 4'b0000 : node21987;
																assign node21987 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node21991 = (inp[1]) ? node21993 : 4'b1000;
															assign node21993 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node21996 = (inp[1]) ? node21998 : 4'b1000;
														assign node21998 = (inp[7]) ? node22000 : 4'b0001;
															assign node22000 = (inp[14]) ? 4'b1001 : node22001;
																assign node22001 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node22005 = (inp[7]) ? node22023 : node22006;
													assign node22006 = (inp[14]) ? node22016 : node22007;
														assign node22007 = (inp[12]) ? node22009 : 4'b0001;
															assign node22009 = (inp[1]) ? node22013 : node22010;
																assign node22010 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node22013 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22016 = (inp[1]) ? 4'b0000 : node22017;
															assign node22017 = (inp[2]) ? 4'b0000 : node22018;
																assign node22018 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node22023 = (inp[1]) ? node22035 : node22024;
														assign node22024 = (inp[2]) ? node22032 : node22025;
															assign node22025 = (inp[12]) ? node22029 : node22026;
																assign node22026 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node22029 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22032 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22035 = (inp[2]) ? 4'b0001 : node22036;
															assign node22036 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node22040 = (inp[10]) ? node22074 : node22041;
												assign node22041 = (inp[1]) ? node22061 : node22042;
													assign node22042 = (inp[2]) ? node22052 : node22043;
														assign node22043 = (inp[7]) ? node22047 : node22044;
															assign node22044 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22047 = (inp[14]) ? node22049 : 4'b0000;
																assign node22049 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node22052 = (inp[12]) ? node22058 : node22053;
															assign node22053 = (inp[7]) ? 4'b0000 : node22054;
																assign node22054 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22058 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node22061 = (inp[2]) ? node22067 : node22062;
														assign node22062 = (inp[7]) ? node22064 : 4'b0001;
															assign node22064 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22067 = (inp[7]) ? node22069 : 4'b0000;
															assign node22069 = (inp[12]) ? node22071 : 4'b0001;
																assign node22071 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node22074 = (inp[1]) ? 4'b0000 : node22075;
													assign node22075 = (inp[14]) ? node22083 : node22076;
														assign node22076 = (inp[2]) ? node22078 : 4'b0001;
															assign node22078 = (inp[12]) ? 4'b0000 : node22079;
																assign node22079 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node22083 = (inp[2]) ? node22087 : node22084;
															assign node22084 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node22087 = (inp[7]) ? node22089 : 4'b0000;
																assign node22089 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node22093 = (inp[1]) ? node22165 : node22094;
										assign node22094 = (inp[13]) ? node22136 : node22095;
											assign node22095 = (inp[12]) ? node22117 : node22096;
												assign node22096 = (inp[2]) ? node22106 : node22097;
													assign node22097 = (inp[10]) ? node22101 : node22098;
														assign node22098 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node22101 = (inp[7]) ? node22103 : 4'b0000;
															assign node22103 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node22106 = (inp[10]) ? node22112 : node22107;
														assign node22107 = (inp[4]) ? node22109 : 4'b1000;
															assign node22109 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node22112 = (inp[7]) ? 4'b0001 : node22113;
															assign node22113 = (inp[4]) ? 4'b1000 : 4'b0001;
												assign node22117 = (inp[4]) ? node22127 : node22118;
													assign node22118 = (inp[10]) ? node22120 : 4'b1000;
														assign node22120 = (inp[2]) ? node22124 : node22121;
															assign node22121 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node22124 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22127 = (inp[7]) ? node22131 : node22128;
														assign node22128 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node22131 = (inp[10]) ? node22133 : 4'b0001;
															assign node22133 = (inp[2]) ? 4'b1000 : 4'b0001;
											assign node22136 = (inp[4]) ? node22152 : node22137;
												assign node22137 = (inp[7]) ? node22143 : node22138;
													assign node22138 = (inp[2]) ? node22140 : 4'b1001;
														assign node22140 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node22143 = (inp[2]) ? node22149 : node22144;
														assign node22144 = (inp[10]) ? node22146 : 4'b0000;
															assign node22146 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node22149 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node22152 = (inp[10]) ? 4'b0000 : node22153;
													assign node22153 = (inp[12]) ? node22159 : node22154;
														assign node22154 = (inp[7]) ? 4'b0000 : node22155;
															assign node22155 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22159 = (inp[2]) ? node22161 : 4'b0000;
															assign node22161 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node22165 = (inp[4]) ? node22201 : node22166;
											assign node22166 = (inp[10]) ? node22194 : node22167;
												assign node22167 = (inp[13]) ? node22177 : node22168;
													assign node22168 = (inp[2]) ? node22172 : node22169;
														assign node22169 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22172 = (inp[7]) ? 4'b0000 : node22173;
															assign node22173 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node22177 = (inp[14]) ? node22185 : node22178;
														assign node22178 = (inp[12]) ? node22180 : 4'b1000;
															assign node22180 = (inp[7]) ? 4'b1000 : node22181;
																assign node22181 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node22185 = (inp[2]) ? node22189 : node22186;
															assign node22186 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node22189 = (inp[12]) ? node22191 : 4'b1000;
																assign node22191 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node22194 = (inp[2]) ? node22196 : 4'b0000;
													assign node22196 = (inp[13]) ? 4'b0000 : node22197;
														assign node22197 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node22201 = (inp[10]) ? 4'b0000 : node22202;
												assign node22202 = (inp[13]) ? 4'b0000 : node22203;
													assign node22203 = (inp[14]) ? node22211 : node22204;
														assign node22204 = (inp[7]) ? 4'b0000 : node22205;
															assign node22205 = (inp[2]) ? 4'b0000 : node22206;
																assign node22206 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22211 = (inp[12]) ? node22213 : 4'b0000;
															assign node22213 = (inp[7]) ? node22215 : 4'b0000;
																assign node22215 = (inp[2]) ? 4'b1000 : 4'b0000;
					assign node22220 = (inp[6]) ? node22222 : 4'b0000;
						assign node22222 = (inp[2]) ? node22684 : node22223;
							assign node22223 = (inp[5]) ? node22299 : node22224;
								assign node22224 = (inp[3]) ? node22226 : 4'b0000;
									assign node22226 = (inp[7]) ? node22284 : node22227;
										assign node22227 = (inp[4]) ? node22239 : node22228;
											assign node22228 = (inp[13]) ? node22230 : 4'b0000;
												assign node22230 = (inp[10]) ? node22232 : 4'b0000;
													assign node22232 = (inp[12]) ? 4'b0000 : node22233;
														assign node22233 = (inp[1]) ? node22235 : 4'b0001;
															assign node22235 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node22239 = (inp[1]) ? node22261 : node22240;
												assign node22240 = (inp[14]) ? node22250 : node22241;
													assign node22241 = (inp[13]) ? node22245 : node22242;
														assign node22242 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22245 = (inp[12]) ? 4'b1001 : node22246;
															assign node22246 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node22250 = (inp[11]) ? node22256 : node22251;
														assign node22251 = (inp[13]) ? node22253 : 4'b0000;
															assign node22253 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node22256 = (inp[13]) ? node22258 : 4'b0001;
															assign node22258 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node22261 = (inp[14]) ? node22271 : node22262;
													assign node22262 = (inp[13]) ? node22266 : node22263;
														assign node22263 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22266 = (inp[12]) ? node22268 : 4'b0000;
															assign node22268 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node22271 = (inp[11]) ? node22279 : node22272;
														assign node22272 = (inp[13]) ? node22274 : 4'b0001;
															assign node22274 = (inp[10]) ? node22276 : 4'b1001;
																assign node22276 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node22279 = (inp[13]) ? node22281 : 4'b1000;
															assign node22281 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node22284 = (inp[13]) ? node22286 : 4'b0000;
											assign node22286 = (inp[1]) ? 4'b0000 : node22287;
												assign node22287 = (inp[4]) ? node22289 : 4'b0000;
													assign node22289 = (inp[12]) ? 4'b0000 : node22290;
														assign node22290 = (inp[11]) ? 4'b0001 : node22291;
															assign node22291 = (inp[10]) ? node22293 : 4'b0000;
																assign node22293 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node22299 = (inp[1]) ? node22505 : node22300;
									assign node22300 = (inp[3]) ? node22400 : node22301;
										assign node22301 = (inp[14]) ? node22341 : node22302;
											assign node22302 = (inp[13]) ? node22320 : node22303;
												assign node22303 = (inp[12]) ? node22315 : node22304;
													assign node22304 = (inp[10]) ? node22310 : node22305;
														assign node22305 = (inp[7]) ? 4'b0001 : node22306;
															assign node22306 = (inp[11]) ? 4'b0101 : 4'b0001;
														assign node22310 = (inp[4]) ? node22312 : 4'b1001;
															assign node22312 = (inp[11]) ? 4'b0000 : 4'b1001;
													assign node22315 = (inp[4]) ? node22317 : 4'b0001;
														assign node22317 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node22320 = (inp[12]) ? node22328 : node22321;
													assign node22321 = (inp[10]) ? node22323 : 4'b1001;
														assign node22323 = (inp[7]) ? node22325 : 4'b0101;
															assign node22325 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node22328 = (inp[7]) ? 4'b1001 : node22329;
														assign node22329 = (inp[10]) ? node22335 : node22330;
															assign node22330 = (inp[4]) ? node22332 : 4'b1001;
																assign node22332 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22335 = (inp[4]) ? node22337 : 4'b1001;
																assign node22337 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node22341 = (inp[11]) ? node22367 : node22342;
												assign node22342 = (inp[13]) ? node22356 : node22343;
													assign node22343 = (inp[7]) ? node22351 : node22344;
														assign node22344 = (inp[4]) ? node22346 : 4'b0000;
															assign node22346 = (inp[10]) ? node22348 : 4'b0100;
																assign node22348 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node22351 = (inp[12]) ? 4'b0000 : node22352;
															assign node22352 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node22356 = (inp[7]) ? node22362 : node22357;
														assign node22357 = (inp[4]) ? node22359 : 4'b1000;
															assign node22359 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node22362 = (inp[12]) ? 4'b1000 : node22363;
															assign node22363 = (inp[10]) ? 4'b0100 : 4'b1000;
												assign node22367 = (inp[13]) ? node22383 : node22368;
													assign node22368 = (inp[7]) ? node22378 : node22369;
														assign node22369 = (inp[4]) ? node22373 : node22370;
															assign node22370 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node22373 = (inp[12]) ? 4'b0101 : node22374;
																assign node22374 = (inp[10]) ? 4'b0000 : 4'b0101;
														assign node22378 = (inp[10]) ? node22380 : 4'b0001;
															assign node22380 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node22383 = (inp[4]) ? node22389 : node22384;
														assign node22384 = (inp[10]) ? node22386 : 4'b1001;
															assign node22386 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node22389 = (inp[7]) ? node22395 : node22390;
															assign node22390 = (inp[10]) ? 4'b0000 : node22391;
																assign node22391 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22395 = (inp[10]) ? node22397 : 4'b1001;
																assign node22397 = (inp[12]) ? 4'b1001 : 4'b0000;
										assign node22400 = (inp[4]) ? node22444 : node22401;
											assign node22401 = (inp[10]) ? node22425 : node22402;
												assign node22402 = (inp[11]) ? node22414 : node22403;
													assign node22403 = (inp[13]) ? node22405 : 4'b0001;
														assign node22405 = (inp[7]) ? node22409 : node22406;
															assign node22406 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node22409 = (inp[14]) ? 4'b0001 : node22410;
																assign node22410 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node22414 = (inp[13]) ? node22418 : node22415;
														assign node22415 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22418 = (inp[7]) ? node22422 : node22419;
															assign node22419 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node22422 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node22425 = (inp[7]) ? node22431 : node22426;
													assign node22426 = (inp[11]) ? node22428 : 4'b0000;
														assign node22428 = (inp[13]) ? 4'b1000 : 4'b0001;
													assign node22431 = (inp[11]) ? node22439 : node22432;
														assign node22432 = (inp[14]) ? node22436 : node22433;
															assign node22433 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node22436 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22439 = (inp[13]) ? 4'b1001 : node22440;
															assign node22440 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node22444 = (inp[13]) ? node22474 : node22445;
												assign node22445 = (inp[10]) ? node22463 : node22446;
													assign node22446 = (inp[7]) ? node22458 : node22447;
														assign node22447 = (inp[12]) ? node22453 : node22448;
															assign node22448 = (inp[11]) ? 4'b0000 : node22449;
																assign node22449 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node22453 = (inp[11]) ? 4'b1001 : node22454;
																assign node22454 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22458 = (inp[12]) ? node22460 : 4'b1000;
															assign node22460 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node22463 = (inp[11]) ? 4'b0000 : node22464;
														assign node22464 = (inp[14]) ? node22468 : node22465;
															assign node22465 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node22468 = (inp[7]) ? node22470 : 4'b0001;
																assign node22470 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node22474 = (inp[10]) ? node22494 : node22475;
													assign node22475 = (inp[11]) ? node22481 : node22476;
														assign node22476 = (inp[12]) ? node22478 : 4'b0000;
															assign node22478 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node22481 = (inp[14]) ? node22487 : node22482;
															assign node22482 = (inp[12]) ? 4'b0001 : node22483;
																assign node22483 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node22487 = (inp[7]) ? node22491 : node22488;
																assign node22488 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node22491 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node22494 = (inp[11]) ? 4'b0000 : node22495;
														assign node22495 = (inp[12]) ? node22497 : 4'b0000;
															assign node22497 = (inp[14]) ? node22501 : node22498;
																assign node22498 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node22501 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node22505 = (inp[11]) ? node22613 : node22506;
										assign node22506 = (inp[4]) ? node22566 : node22507;
											assign node22507 = (inp[10]) ? node22537 : node22508;
												assign node22508 = (inp[7]) ? node22522 : node22509;
													assign node22509 = (inp[14]) ? node22519 : node22510;
														assign node22510 = (inp[3]) ? node22516 : node22511;
															assign node22511 = (inp[12]) ? node22513 : 4'b1000;
																assign node22513 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node22516 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22519 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node22522 = (inp[13]) ? node22532 : node22523;
														assign node22523 = (inp[14]) ? node22527 : node22524;
															assign node22524 = (inp[3]) ? 4'b0001 : 4'b0000;
															assign node22527 = (inp[3]) ? node22529 : 4'b0001;
																assign node22529 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22532 = (inp[3]) ? node22534 : 4'b1001;
															assign node22534 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node22537 = (inp[12]) ? node22547 : node22538;
													assign node22538 = (inp[13]) ? node22544 : node22539;
														assign node22539 = (inp[3]) ? node22541 : 4'b1000;
															assign node22541 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node22544 = (inp[3]) ? 4'b0000 : 4'b0100;
													assign node22547 = (inp[7]) ? node22555 : node22548;
														assign node22548 = (inp[13]) ? 4'b1000 : node22549;
															assign node22549 = (inp[3]) ? node22551 : 4'b1000;
																assign node22551 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22555 = (inp[3]) ? node22561 : node22556;
															assign node22556 = (inp[14]) ? 4'b1001 : node22557;
																assign node22557 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node22561 = (inp[13]) ? node22563 : 4'b1001;
																assign node22563 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node22566 = (inp[3]) ? node22592 : node22567;
												assign node22567 = (inp[14]) ? node22585 : node22568;
													assign node22568 = (inp[13]) ? node22578 : node22569;
														assign node22569 = (inp[7]) ? 4'b1000 : node22570;
															assign node22570 = (inp[10]) ? node22574 : node22571;
																assign node22571 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node22574 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node22578 = (inp[7]) ? node22580 : 4'b0001;
															assign node22580 = (inp[10]) ? node22582 : 4'b0100;
																assign node22582 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node22585 = (inp[12]) ? node22587 : 4'b0001;
														assign node22587 = (inp[13]) ? node22589 : 4'b0101;
															assign node22589 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node22592 = (inp[13]) ? node22604 : node22593;
													assign node22593 = (inp[7]) ? node22599 : node22594;
														assign node22594 = (inp[10]) ? node22596 : 4'b0001;
															assign node22596 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node22599 = (inp[14]) ? node22601 : 4'b0000;
															assign node22601 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node22604 = (inp[7]) ? node22606 : 4'b0000;
														assign node22606 = (inp[12]) ? 4'b0000 : node22607;
															assign node22607 = (inp[10]) ? 4'b0000 : node22608;
																assign node22608 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node22613 = (inp[13]) ? node22659 : node22614;
											assign node22614 = (inp[4]) ? node22632 : node22615;
												assign node22615 = (inp[12]) ? node22625 : node22616;
													assign node22616 = (inp[3]) ? node22618 : 4'b1000;
														assign node22618 = (inp[10]) ? node22622 : node22619;
															assign node22619 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node22622 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node22625 = (inp[3]) ? node22629 : node22626;
														assign node22626 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22629 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node22632 = (inp[10]) ? node22654 : node22633;
													assign node22633 = (inp[3]) ? node22641 : node22634;
														assign node22634 = (inp[7]) ? node22638 : node22635;
															assign node22635 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node22638 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22641 = (inp[14]) ? node22649 : node22642;
															assign node22642 = (inp[7]) ? node22646 : node22643;
																assign node22643 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node22646 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22649 = (inp[12]) ? 4'b1000 : node22650;
																assign node22650 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node22654 = (inp[7]) ? node22656 : 4'b0000;
														assign node22656 = (inp[3]) ? 4'b0000 : 4'b1000;
											assign node22659 = (inp[3]) ? node22675 : node22660;
												assign node22660 = (inp[10]) ? node22670 : node22661;
													assign node22661 = (inp[12]) ? 4'b1000 : node22662;
														assign node22662 = (inp[4]) ? node22666 : node22663;
															assign node22663 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node22666 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node22670 = (inp[7]) ? 4'b0000 : node22671;
														assign node22671 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node22675 = (inp[7]) ? node22677 : 4'b0000;
													assign node22677 = (inp[4]) ? 4'b0000 : node22678;
														assign node22678 = (inp[12]) ? 4'b0000 : node22679;
															assign node22679 = (inp[10]) ? 4'b0000 : 4'b1000;
							assign node22684 = (inp[5]) ? node22686 : 4'b0000;
								assign node22686 = (inp[3]) ? node22688 : 4'b0000;
									assign node22688 = (inp[7]) ? node22740 : node22689;
										assign node22689 = (inp[4]) ? node22705 : node22690;
											assign node22690 = (inp[13]) ? node22692 : 4'b0000;
												assign node22692 = (inp[10]) ? node22694 : 4'b0000;
													assign node22694 = (inp[12]) ? 4'b0000 : node22695;
														assign node22695 = (inp[1]) ? node22701 : node22696;
															assign node22696 = (inp[11]) ? 4'b0001 : node22697;
																assign node22697 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22701 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node22705 = (inp[11]) ? node22731 : node22706;
												assign node22706 = (inp[12]) ? node22720 : node22707;
													assign node22707 = (inp[13]) ? node22715 : node22708;
														assign node22708 = (inp[10]) ? node22712 : node22709;
															assign node22709 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node22712 = (inp[14]) ? 4'b1000 : 4'b0001;
														assign node22715 = (inp[1]) ? 4'b0000 : node22716;
															assign node22716 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node22720 = (inp[1]) ? node22726 : node22721;
														assign node22721 = (inp[13]) ? 4'b0001 : node22722;
															assign node22722 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22726 = (inp[14]) ? node22728 : 4'b0000;
															assign node22728 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node22731 = (inp[1]) ? 4'b0000 : node22732;
													assign node22732 = (inp[10]) ? 4'b0000 : node22733;
														assign node22733 = (inp[13]) ? node22735 : 4'b0001;
															assign node22735 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node22740 = (inp[12]) ? 4'b0000 : node22741;
											assign node22741 = (inp[10]) ? node22743 : 4'b0000;
												assign node22743 = (inp[11]) ? 4'b0000 : node22744;
													assign node22744 = (inp[4]) ? node22746 : 4'b0000;
														assign node22746 = (inp[1]) ? 4'b0000 : node22747;
															assign node22747 = (inp[13]) ? 4'b0001 : 4'b0000;

endmodule