module dtc_split66_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node841;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node938;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node978;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1034;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1068;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;

	assign outp = (inp[6]) ? node232 : node1;
		assign node1 = (inp[7]) ? node51 : node2;
			assign node2 = (inp[0]) ? node4 : 3'b000;
				assign node4 = (inp[9]) ? 3'b000 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[10]) ? 3'b000 : node7;
							assign node7 = (inp[8]) ? node9 : 3'b000;
								assign node9 = (inp[3]) ? node27 : node10;
									assign node10 = (inp[5]) ? node18 : node11;
										assign node11 = (inp[4]) ? 3'b000 : node12;
											assign node12 = (inp[11]) ? 3'b000 : node13;
												assign node13 = (inp[2]) ? 3'b000 : 3'b100;
										assign node18 = (inp[4]) ? 3'b100 : node19;
											assign node19 = (inp[11]) ? node23 : node20;
												assign node20 = (inp[2]) ? 3'b000 : 3'b100;
												assign node23 = (inp[2]) ? 3'b100 : 3'b000;
									assign node27 = (inp[4]) ? node43 : node28;
										assign node28 = (inp[5]) ? node36 : node29;
											assign node29 = (inp[11]) ? node33 : node30;
												assign node30 = (inp[2]) ? 3'b000 : 3'b100;
												assign node33 = (inp[2]) ? 3'b100 : 3'b000;
											assign node36 = (inp[11]) ? node40 : node37;
												assign node37 = (inp[2]) ? 3'b000 : 3'b100;
												assign node40 = (inp[2]) ? 3'b100 : 3'b000;
										assign node43 = (inp[11]) ? node45 : 3'b100;
											assign node45 = (inp[2]) ? 3'b100 : 3'b000;
			assign node51 = (inp[9]) ? node197 : node52;
				assign node52 = (inp[0]) ? node130 : node53;
					assign node53 = (inp[10]) ? node97 : node54;
						assign node54 = (inp[1]) ? node58 : node55;
							assign node55 = (inp[11]) ? 3'b001 : 3'b101;
							assign node58 = (inp[8]) ? node74 : node59;
								assign node59 = (inp[3]) ? node67 : node60;
									assign node60 = (inp[11]) ? 3'b010 : node61;
										assign node61 = (inp[2]) ? node63 : 3'b110;
											assign node63 = (inp[4]) ? 3'b010 : 3'b110;
									assign node67 = (inp[2]) ? node71 : node68;
										assign node68 = (inp[11]) ? 3'b010 : 3'b110;
										assign node71 = (inp[11]) ? 3'b110 : 3'b010;
								assign node74 = (inp[11]) ? node86 : node75;
									assign node75 = (inp[4]) ? 3'b001 : node76;
										assign node76 = (inp[2]) ? node82 : node77;
											assign node77 = (inp[5]) ? 3'b001 : node78;
												assign node78 = (inp[3]) ? 3'b001 : 3'b101;
											assign node82 = (inp[3]) ? 3'b110 : 3'b001;
									assign node86 = (inp[4]) ? 3'b110 : node87;
										assign node87 = (inp[5]) ? node93 : node88;
											assign node88 = (inp[3]) ? 3'b110 : node89;
												assign node89 = (inp[2]) ? 3'b110 : 3'b001;
											assign node93 = (inp[2]) ? 3'b010 : 3'b110;
						assign node97 = (inp[1]) ? node99 : 3'b110;
							assign node99 = (inp[8]) ? node103 : node100;
								assign node100 = (inp[11]) ? 3'b000 : 3'b100;
								assign node103 = (inp[11]) ? node117 : node104;
									assign node104 = (inp[2]) ? node110 : node105;
										assign node105 = (inp[5]) ? 3'b010 : node106;
											assign node106 = (inp[3]) ? 3'b010 : 3'b110;
										assign node110 = (inp[3]) ? node112 : 3'b010;
											assign node112 = (inp[4]) ? 3'b100 : node113;
												assign node113 = (inp[5]) ? 3'b100 : 3'b010;
									assign node117 = (inp[4]) ? 3'b100 : node118;
										assign node118 = (inp[5]) ? node124 : node119;
											assign node119 = (inp[2]) ? 3'b110 : node120;
												assign node120 = (inp[3]) ? 3'b110 : 3'b010;
											assign node124 = (inp[2]) ? node126 : 3'b100;
												assign node126 = (inp[3]) ? 3'b000 : 3'b010;
					assign node130 = (inp[10]) ? node184 : node131;
						assign node131 = (inp[1]) ? node159 : node132;
							assign node132 = (inp[8]) ? node148 : node133;
								assign node133 = (inp[11]) ? node141 : node134;
									assign node134 = (inp[2]) ? node136 : 3'b010;
										assign node136 = (inp[4]) ? 3'b100 : node137;
											assign node137 = (inp[3]) ? 3'b100 : 3'b010;
									assign node141 = (inp[2]) ? node143 : 3'b100;
										assign node143 = (inp[4]) ? 3'b010 : node144;
											assign node144 = (inp[3]) ? 3'b010 : 3'b100;
								assign node148 = (inp[2]) ? node152 : node149;
									assign node149 = (inp[11]) ? 3'b010 : 3'b110;
									assign node152 = (inp[11]) ? node154 : 3'b010;
										assign node154 = (inp[3]) ? 3'b100 : node155;
											assign node155 = (inp[4]) ? 3'b100 : 3'b010;
							assign node159 = (inp[8]) ? node167 : node160;
								assign node160 = (inp[2]) ? 3'b000 : node161;
									assign node161 = (inp[3]) ? 3'b000 : node162;
										assign node162 = (inp[11]) ? 3'b000 : 3'b100;
								assign node167 = (inp[5]) ? node177 : node168;
									assign node168 = (inp[11]) ? node172 : node169;
										assign node169 = (inp[2]) ? 3'b100 : 3'b010;
										assign node172 = (inp[2]) ? 3'b000 : node173;
											assign node173 = (inp[3]) ? 3'b000 : 3'b100;
									assign node177 = (inp[4]) ? node179 : 3'b100;
										assign node179 = (inp[11]) ? node181 : 3'b100;
											assign node181 = (inp[3]) ? 3'b000 : 3'b100;
						assign node184 = (inp[11]) ? 3'b000 : node185;
							assign node185 = (inp[1]) ? 3'b000 : node186;
								assign node186 = (inp[8]) ? node188 : 3'b000;
									assign node188 = (inp[2]) ? node190 : 3'b100;
										assign node190 = (inp[4]) ? 3'b000 : node191;
											assign node191 = (inp[3]) ? 3'b000 : 3'b100;
				assign node197 = (inp[0]) ? 3'b000 : node198;
					assign node198 = (inp[10]) ? 3'b000 : node199;
						assign node199 = (inp[1]) ? node207 : node200;
							assign node200 = (inp[2]) ? node204 : node201;
								assign node201 = (inp[11]) ? 3'b110 : 3'b010;
								assign node204 = (inp[11]) ? 3'b000 : 3'b100;
							assign node207 = (inp[8]) ? node209 : 3'b000;
								assign node209 = (inp[3]) ? node219 : node210;
									assign node210 = (inp[4]) ? 3'b000 : node211;
										assign node211 = (inp[2]) ? node215 : node212;
											assign node212 = (inp[11]) ? 3'b000 : 3'b100;
											assign node215 = (inp[11]) ? 3'b100 : 3'b000;
									assign node219 = (inp[11]) ? node225 : node220;
										assign node220 = (inp[4]) ? node222 : 3'b000;
											assign node222 = (inp[2]) ? 3'b100 : 3'b000;
										assign node225 = (inp[4]) ? node227 : 3'b100;
											assign node227 = (inp[2]) ? 3'b000 : 3'b100;
		assign node232 = (inp[9]) ? node756 : node233;
			assign node233 = (inp[0]) ? node461 : node234;
				assign node234 = (inp[7]) ? node388 : node235;
					assign node235 = (inp[10]) ? node311 : node236;
						assign node236 = (inp[1]) ? node266 : node237;
							assign node237 = (inp[11]) ? node253 : node238;
								assign node238 = (inp[8]) ? node244 : node239;
									assign node239 = (inp[3]) ? 3'b011 : node240;
										assign node240 = (inp[2]) ? 3'b011 : 3'b111;
									assign node244 = (inp[2]) ? 3'b111 : node245;
										assign node245 = (inp[3]) ? node247 : 3'b011;
											assign node247 = (inp[4]) ? 3'b111 : node248;
												assign node248 = (inp[5]) ? 3'b111 : 3'b011;
								assign node253 = (inp[8]) ? node259 : node254;
									assign node254 = (inp[3]) ? 3'b101 : node255;
										assign node255 = (inp[2]) ? 3'b101 : 3'b001;
									assign node259 = (inp[2]) ? 3'b011 : node260;
										assign node260 = (inp[3]) ? node262 : 3'b111;
											assign node262 = (inp[4]) ? 3'b011 : 3'b111;
							assign node266 = (inp[8]) ? node288 : node267;
								assign node267 = (inp[11]) ? node277 : node268;
									assign node268 = (inp[2]) ? node274 : node269;
										assign node269 = (inp[3]) ? 3'b101 : node270;
											assign node270 = (inp[4]) ? 3'b101 : 3'b110;
										assign node274 = (inp[3]) ? 3'b001 : 3'b101;
									assign node277 = (inp[5]) ? 3'b001 : node278;
										assign node278 = (inp[2]) ? node284 : node279;
											assign node279 = (inp[3]) ? 3'b001 : node280;
												assign node280 = (inp[4]) ? 3'b001 : 3'b101;
											assign node284 = (inp[4]) ? 3'b110 : 3'b001;
								assign node288 = (inp[11]) ? node300 : node289;
									assign node289 = (inp[2]) ? node295 : node290;
										assign node290 = (inp[4]) ? 3'b011 : node291;
											assign node291 = (inp[3]) ? 3'b011 : 3'b101;
										assign node295 = (inp[3]) ? node297 : 3'b011;
											assign node297 = (inp[5]) ? 3'b011 : 3'b101;
									assign node300 = (inp[3]) ? node306 : node301;
										assign node301 = (inp[5]) ? 3'b101 : node302;
											assign node302 = (inp[2]) ? 3'b101 : 3'b011;
										assign node306 = (inp[5]) ? node308 : 3'b101;
											assign node308 = (inp[2]) ? 3'b001 : 3'b101;
						assign node311 = (inp[1]) ? node345 : node312;
							assign node312 = (inp[8]) ? node334 : node313;
								assign node313 = (inp[11]) ? node323 : node314;
									assign node314 = (inp[2]) ? 3'b001 : node315;
										assign node315 = (inp[3]) ? 3'b001 : node316;
											assign node316 = (inp[5]) ? node318 : 3'b101;
												assign node318 = (inp[4]) ? 3'b101 : 3'b001;
									assign node323 = (inp[3]) ? node331 : node324;
										assign node324 = (inp[2]) ? node326 : 3'b001;
											assign node326 = (inp[5]) ? 3'b010 : node327;
												assign node327 = (inp[4]) ? 3'b101 : 3'b111;
										assign node331 = (inp[2]) ? 3'b111 : 3'b110;
								assign node334 = (inp[11]) ? node338 : node335;
									assign node335 = (inp[2]) ? 3'b101 : 3'b011;
									assign node338 = (inp[2]) ? 3'b001 : node339;
										assign node339 = (inp[4]) ? node341 : 3'b101;
											assign node341 = (inp[3]) ? 3'b001 : 3'b101;
							assign node345 = (inp[8]) ? node363 : node346;
								assign node346 = (inp[11]) ? node358 : node347;
									assign node347 = (inp[2]) ? node353 : node348;
										assign node348 = (inp[4]) ? 3'b110 : node349;
											assign node349 = (inp[3]) ? 3'b110 : 3'b001;
										assign node353 = (inp[3]) ? node355 : 3'b110;
											assign node355 = (inp[4]) ? 3'b010 : 3'b110;
									assign node358 = (inp[2]) ? node360 : 3'b010;
										assign node360 = (inp[3]) ? 3'b100 : 3'b010;
								assign node363 = (inp[11]) ? node377 : node364;
									assign node364 = (inp[2]) ? node370 : node365;
										assign node365 = (inp[4]) ? 3'b001 : node366;
											assign node366 = (inp[5]) ? 3'b001 : 3'b101;
										assign node370 = (inp[4]) ? node372 : 3'b001;
											assign node372 = (inp[5]) ? 3'b110 : node373;
												assign node373 = (inp[3]) ? 3'b101 : 3'b001;
									assign node377 = (inp[4]) ? node381 : node378;
										assign node378 = (inp[2]) ? 3'b110 : 3'b010;
										assign node381 = (inp[3]) ? node383 : 3'b001;
											assign node383 = (inp[5]) ? node385 : 3'b001;
												assign node385 = (inp[2]) ? 3'b010 : 3'b110;
					assign node388 = (inp[10]) ? node408 : node389;
						assign node389 = (inp[8]) ? 3'b111 : node390;
							assign node390 = (inp[1]) ? node392 : 3'b111;
								assign node392 = (inp[11]) ? node398 : node393;
									assign node393 = (inp[3]) ? 3'b111 : node394;
										assign node394 = (inp[2]) ? 3'b111 : 3'b011;
									assign node398 = (inp[5]) ? node400 : 3'b011;
										assign node400 = (inp[3]) ? node404 : node401;
											assign node401 = (inp[2]) ? 3'b011 : 3'b111;
											assign node404 = (inp[2]) ? 3'b101 : 3'b011;
						assign node408 = (inp[1]) ? node438 : node409;
							assign node409 = (inp[11]) ? node415 : node410;
								assign node410 = (inp[8]) ? 3'b111 : node411;
									assign node411 = (inp[2]) ? 3'b011 : 3'b111;
								assign node415 = (inp[5]) ? node425 : node416;
									assign node416 = (inp[2]) ? node420 : node417;
										assign node417 = (inp[8]) ? 3'b111 : 3'b011;
										assign node420 = (inp[4]) ? node422 : 3'b011;
											assign node422 = (inp[8]) ? 3'b011 : 3'b111;
									assign node425 = (inp[8]) ? node435 : node426;
										assign node426 = (inp[4]) ? node430 : node427;
											assign node427 = (inp[3]) ? 3'b001 : 3'b011;
											assign node430 = (inp[2]) ? 3'b101 : node431;
												assign node431 = (inp[3]) ? 3'b101 : 3'b011;
										assign node435 = (inp[2]) ? 3'b011 : 3'b111;
							assign node438 = (inp[11]) ? node450 : node439;
								assign node439 = (inp[8]) ? node445 : node440;
									assign node440 = (inp[2]) ? 3'b101 : node441;
										assign node441 = (inp[3]) ? 3'b101 : 3'b011;
									assign node445 = (inp[3]) ? 3'b011 : node446;
										assign node446 = (inp[2]) ? 3'b011 : 3'b111;
								assign node450 = (inp[8]) ? node456 : node451;
									assign node451 = (inp[3]) ? 3'b001 : node452;
										assign node452 = (inp[2]) ? 3'b001 : 3'b101;
									assign node456 = (inp[3]) ? 3'b101 : node457;
										assign node457 = (inp[2]) ? 3'b101 : 3'b001;
				assign node461 = (inp[7]) ? node587 : node462;
					assign node462 = (inp[10]) ? node534 : node463;
						assign node463 = (inp[8]) ? node501 : node464;
							assign node464 = (inp[11]) ? node482 : node465;
								assign node465 = (inp[1]) ? node473 : node466;
									assign node466 = (inp[2]) ? node468 : 3'b001;
										assign node468 = (inp[3]) ? 3'b110 : node469;
											assign node469 = (inp[4]) ? 3'b110 : 3'b001;
									assign node473 = (inp[2]) ? 3'b010 : node474;
										assign node474 = (inp[4]) ? node476 : 3'b110;
											assign node476 = (inp[3]) ? 3'b010 : node477;
												assign node477 = (inp[5]) ? 3'b110 : 3'b010;
								assign node482 = (inp[1]) ? node490 : node483;
									assign node483 = (inp[2]) ? node485 : 3'b110;
										assign node485 = (inp[3]) ? 3'b010 : node486;
											assign node486 = (inp[4]) ? 3'b010 : 3'b110;
									assign node490 = (inp[2]) ? node496 : node491;
										assign node491 = (inp[3]) ? node493 : 3'b010;
											assign node493 = (inp[5]) ? 3'b100 : 3'b010;
										assign node496 = (inp[5]) ? 3'b100 : node497;
											assign node497 = (inp[4]) ? 3'b010 : 3'b100;
							assign node501 = (inp[1]) ? node521 : node502;
								assign node502 = (inp[3]) ? node514 : node503;
									assign node503 = (inp[11]) ? node509 : node504;
										assign node504 = (inp[2]) ? node506 : 3'b101;
											assign node506 = (inp[4]) ? 3'b001 : 3'b101;
										assign node509 = (inp[2]) ? node511 : 3'b001;
											assign node511 = (inp[4]) ? 3'b101 : 3'b001;
									assign node514 = (inp[11]) ? node518 : node515;
										assign node515 = (inp[2]) ? 3'b001 : 3'b101;
										assign node518 = (inp[2]) ? 3'b110 : 3'b001;
								assign node521 = (inp[11]) ? node529 : node522;
									assign node522 = (inp[2]) ? 3'b110 : node523;
										assign node523 = (inp[5]) ? node525 : 3'b001;
											assign node525 = (inp[4]) ? 3'b110 : 3'b001;
									assign node529 = (inp[4]) ? node531 : 3'b110;
										assign node531 = (inp[2]) ? 3'b010 : 3'b110;
						assign node534 = (inp[1]) ? node560 : node535;
							assign node535 = (inp[11]) ? node547 : node536;
								assign node536 = (inp[8]) ? node542 : node537;
									assign node537 = (inp[3]) ? node539 : 3'b010;
										assign node539 = (inp[2]) ? 3'b100 : 3'b010;
									assign node542 = (inp[2]) ? node544 : 3'b110;
										assign node544 = (inp[3]) ? 3'b010 : 3'b110;
								assign node547 = (inp[8]) ? node553 : node548;
									assign node548 = (inp[5]) ? node550 : 3'b000;
										assign node550 = (inp[4]) ? 3'b100 : 3'b000;
									assign node553 = (inp[2]) ? 3'b100 : node554;
										assign node554 = (inp[3]) ? 3'b010 : node555;
											assign node555 = (inp[4]) ? 3'b010 : 3'b110;
							assign node560 = (inp[4]) ? node572 : node561;
								assign node561 = (inp[8]) ? node563 : 3'b100;
									assign node563 = (inp[11]) ? node569 : node564;
										assign node564 = (inp[2]) ? node566 : 3'b010;
											assign node566 = (inp[3]) ? 3'b100 : 3'b110;
										assign node569 = (inp[2]) ? 3'b000 : 3'b100;
								assign node572 = (inp[8]) ? node580 : node573;
									assign node573 = (inp[3]) ? 3'b000 : node574;
										assign node574 = (inp[2]) ? 3'b000 : node575;
											assign node575 = (inp[11]) ? 3'b000 : 3'b100;
									assign node580 = (inp[2]) ? node584 : node581;
										assign node581 = (inp[11]) ? 3'b100 : 3'b010;
										assign node584 = (inp[11]) ? 3'b000 : 3'b100;
					assign node587 = (inp[10]) ? node685 : node588;
						assign node588 = (inp[1]) ? node630 : node589;
							assign node589 = (inp[8]) ? node617 : node590;
								assign node590 = (inp[2]) ? node606 : node591;
									assign node591 = (inp[11]) ? node599 : node592;
										assign node592 = (inp[3]) ? 3'b011 : node593;
											assign node593 = (inp[5]) ? node595 : 3'b101;
												assign node595 = (inp[4]) ? 3'b011 : 3'b001;
										assign node599 = (inp[4]) ? 3'b101 : node600;
											assign node600 = (inp[3]) ? 3'b101 : node601;
												assign node601 = (inp[5]) ? 3'b111 : 3'b011;
									assign node606 = (inp[11]) ? node612 : node607;
										assign node607 = (inp[3]) ? 3'b101 : node608;
											assign node608 = (inp[4]) ? 3'b101 : 3'b111;
										assign node612 = (inp[5]) ? 3'b001 : node613;
											assign node613 = (inp[4]) ? 3'b001 : 3'b101;
								assign node617 = (inp[4]) ? node623 : node618;
									assign node618 = (inp[2]) ? 3'b011 : node619;
										assign node619 = (inp[11]) ? 3'b011 : 3'b111;
									assign node623 = (inp[11]) ? node627 : node624;
										assign node624 = (inp[2]) ? 3'b011 : 3'b111;
										assign node627 = (inp[2]) ? 3'b101 : 3'b011;
							assign node630 = (inp[4]) ? node644 : node631;
								assign node631 = (inp[2]) ? node637 : node632;
									assign node632 = (inp[8]) ? 3'b101 : node633;
										assign node633 = (inp[11]) ? 3'b001 : 3'b101;
									assign node637 = (inp[11]) ? node641 : node638;
										assign node638 = (inp[8]) ? 3'b101 : 3'b001;
										assign node641 = (inp[8]) ? 3'b001 : 3'b111;
								assign node644 = (inp[3]) ? node666 : node645;
									assign node645 = (inp[5]) ? node657 : node646;
										assign node646 = (inp[11]) ? node652 : node647;
											assign node647 = (inp[2]) ? node649 : 3'b011;
												assign node649 = (inp[8]) ? 3'b101 : 3'b001;
											assign node652 = (inp[2]) ? 3'b111 : node653;
												assign node653 = (inp[8]) ? 3'b101 : 3'b001;
										assign node657 = (inp[8]) ? node663 : node658;
											assign node658 = (inp[2]) ? 3'b001 : node659;
												assign node659 = (inp[11]) ? 3'b001 : 3'b101;
											assign node663 = (inp[2]) ? 3'b001 : 3'b011;
									assign node666 = (inp[5]) ? node680 : node667;
										assign node667 = (inp[8]) ? node675 : node668;
											assign node668 = (inp[2]) ? node672 : node669;
												assign node669 = (inp[11]) ? 3'b001 : 3'b101;
												assign node672 = (inp[11]) ? 3'b111 : 3'b001;
											assign node675 = (inp[2]) ? node677 : 3'b011;
												assign node677 = (inp[11]) ? 3'b001 : 3'b101;
										assign node680 = (inp[2]) ? node682 : 3'b101;
											assign node682 = (inp[11]) ? 3'b001 : 3'b101;
						assign node685 = (inp[1]) ? node731 : node686;
							assign node686 = (inp[2]) ? node714 : node687;
								assign node687 = (inp[3]) ? node697 : node688;
									assign node688 = (inp[5]) ? 3'b101 : node689;
										assign node689 = (inp[8]) ? node693 : node690;
											assign node690 = (inp[11]) ? 3'b101 : 3'b001;
											assign node693 = (inp[11]) ? 3'b001 : 3'b101;
									assign node697 = (inp[5]) ? node707 : node698;
										assign node698 = (inp[4]) ? node700 : 3'b001;
											assign node700 = (inp[8]) ? node704 : node701;
												assign node701 = (inp[11]) ? 3'b101 : 3'b001;
												assign node704 = (inp[11]) ? 3'b001 : 3'b101;
										assign node707 = (inp[11]) ? node711 : node708;
											assign node708 = (inp[8]) ? 3'b101 : 3'b001;
											assign node711 = (inp[8]) ? 3'b001 : 3'b110;
								assign node714 = (inp[4]) ? node722 : node715;
									assign node715 = (inp[11]) ? node719 : node716;
										assign node716 = (inp[8]) ? 3'b101 : 3'b001;
										assign node719 = (inp[8]) ? 3'b010 : 3'b101;
									assign node722 = (inp[8]) ? node726 : node723;
										assign node723 = (inp[11]) ? 3'b010 : 3'b110;
										assign node726 = (inp[11]) ? 3'b110 : node727;
											assign node727 = (inp[3]) ? 3'b001 : 3'b101;
							assign node731 = (inp[8]) ? node739 : node732;
								assign node732 = (inp[2]) ? node736 : node733;
									assign node733 = (inp[11]) ? 3'b010 : 3'b110;
									assign node736 = (inp[11]) ? 3'b100 : 3'b010;
								assign node739 = (inp[11]) ? node751 : node740;
									assign node740 = (inp[2]) ? node746 : node741;
										assign node741 = (inp[4]) ? 3'b001 : node742;
											assign node742 = (inp[3]) ? 3'b001 : 3'b000;
										assign node746 = (inp[3]) ? node748 : 3'b111;
											assign node748 = (inp[4]) ? 3'b110 : 3'b111;
									assign node751 = (inp[2]) ? 3'b010 : node752;
										assign node752 = (inp[4]) ? 3'b110 : 3'b111;
			assign node756 = (inp[0]) ? node1014 : node757;
				assign node757 = (inp[7]) ? node873 : node758;
					assign node758 = (inp[10]) ? node826 : node759;
						assign node759 = (inp[11]) ? node803 : node760;
							assign node760 = (inp[8]) ? node774 : node761;
								assign node761 = (inp[1]) ? node767 : node762;
									assign node762 = (inp[2]) ? 3'b010 : node763;
										assign node763 = (inp[3]) ? 3'b010 : 3'b110;
									assign node767 = (inp[3]) ? 3'b100 : node768;
										assign node768 = (inp[2]) ? 3'b100 : node769;
											assign node769 = (inp[4]) ? 3'b100 : 3'b010;
								assign node774 = (inp[4]) ? node784 : node775;
									assign node775 = (inp[1]) ? node779 : node776;
										assign node776 = (inp[2]) ? 3'b110 : 3'b001;
										assign node779 = (inp[2]) ? 3'b010 : node780;
											assign node780 = (inp[3]) ? 3'b010 : 3'b110;
									assign node784 = (inp[1]) ? node798 : node785;
										assign node785 = (inp[3]) ? node793 : node786;
											assign node786 = (inp[2]) ? node790 : node787;
												assign node787 = (inp[5]) ? 3'b010 : 3'b110;
												assign node790 = (inp[5]) ? 3'b110 : 3'b010;
											assign node793 = (inp[2]) ? node795 : 3'b110;
												assign node795 = (inp[5]) ? 3'b110 : 3'b010;
										assign node798 = (inp[2]) ? 3'b010 : node799;
											assign node799 = (inp[3]) ? 3'b010 : 3'b110;
							assign node803 = (inp[8]) ? node819 : node804;
								assign node804 = (inp[1]) ? node810 : node805;
									assign node805 = (inp[2]) ? 3'b100 : node806;
										assign node806 = (inp[3]) ? 3'b100 : 3'b000;
									assign node810 = (inp[2]) ? 3'b000 : node811;
										assign node811 = (inp[3]) ? 3'b000 : node812;
											assign node812 = (inp[5]) ? node814 : 3'b100;
												assign node814 = (inp[4]) ? 3'b000 : 3'b100;
								assign node819 = (inp[1]) ? 3'b100 : node820;
									assign node820 = (inp[2]) ? 3'b010 : node821;
										assign node821 = (inp[4]) ? 3'b110 : 3'b101;
						assign node826 = (inp[1]) ? node864 : node827;
							assign node827 = (inp[11]) ? node837 : node828;
								assign node828 = (inp[8]) ? node832 : node829;
									assign node829 = (inp[2]) ? 3'b000 : 3'b100;
									assign node832 = (inp[2]) ? node834 : 3'b010;
										assign node834 = (inp[3]) ? 3'b100 : 3'b110;
								assign node837 = (inp[4]) ? node857 : node838;
									assign node838 = (inp[3]) ? node844 : node839;
										assign node839 = (inp[5]) ? node841 : 3'b100;
											assign node841 = (inp[2]) ? 3'b000 : 3'b100;
										assign node844 = (inp[5]) ? node852 : node845;
											assign node845 = (inp[2]) ? node849 : node846;
												assign node846 = (inp[8]) ? 3'b100 : 3'b000;
												assign node849 = (inp[8]) ? 3'b000 : 3'b100;
											assign node852 = (inp[8]) ? 3'b100 : node853;
												assign node853 = (inp[2]) ? 3'b100 : 3'b000;
									assign node857 = (inp[2]) ? node861 : node858;
										assign node858 = (inp[8]) ? 3'b100 : 3'b000;
										assign node861 = (inp[8]) ? 3'b000 : 3'b100;
							assign node864 = (inp[4]) ? node866 : 3'b000;
								assign node866 = (inp[8]) ? node868 : 3'b000;
									assign node868 = (inp[3]) ? 3'b000 : node869;
										assign node869 = (inp[11]) ? 3'b000 : 3'b100;
					assign node873 = (inp[10]) ? node953 : node874;
						assign node874 = (inp[1]) ? node910 : node875;
							assign node875 = (inp[8]) ? node895 : node876;
								assign node876 = (inp[2]) ? node886 : node877;
									assign node877 = (inp[5]) ? node879 : 3'b101;
										assign node879 = (inp[4]) ? 3'b001 : node880;
											assign node880 = (inp[11]) ? node882 : 3'b101;
												assign node882 = (inp[3]) ? 3'b001 : 3'b101;
									assign node886 = (inp[11]) ? 3'b110 : node887;
										assign node887 = (inp[5]) ? 3'b001 : node888;
											assign node888 = (inp[3]) ? node890 : 3'b101;
												assign node890 = (inp[4]) ? 3'b101 : 3'b001;
								assign node895 = (inp[11]) ? node903 : node896;
									assign node896 = (inp[2]) ? node898 : 3'b011;
										assign node898 = (inp[4]) ? 3'b101 : node899;
											assign node899 = (inp[3]) ? 3'b101 : 3'b011;
									assign node903 = (inp[2]) ? 3'b001 : node904;
										assign node904 = (inp[3]) ? 3'b101 : node905;
											assign node905 = (inp[4]) ? 3'b101 : 3'b001;
							assign node910 = (inp[11]) ? node932 : node911;
								assign node911 = (inp[8]) ? node925 : node912;
									assign node912 = (inp[2]) ? 3'b110 : node913;
										assign node913 = (inp[3]) ? node919 : node914;
											assign node914 = (inp[5]) ? node916 : 3'b001;
												assign node916 = (inp[4]) ? 3'b001 : 3'b110;
											assign node919 = (inp[5]) ? 3'b110 : node920;
												assign node920 = (inp[4]) ? 3'b110 : 3'b001;
									assign node925 = (inp[2]) ? 3'b001 : node926;
										assign node926 = (inp[5]) ? 3'b101 : node927;
											assign node927 = (inp[3]) ? 3'b001 : 3'b101;
								assign node932 = (inp[4]) ? node942 : node933;
									assign node933 = (inp[5]) ? 3'b110 : node934;
										assign node934 = (inp[8]) ? node938 : node935;
											assign node935 = (inp[2]) ? 3'b001 : 3'b110;
											assign node938 = (inp[2]) ? 3'b110 : 3'b010;
									assign node942 = (inp[8]) ? node948 : node943;
										assign node943 = (inp[2]) ? 3'b010 : node944;
											assign node944 = (inp[3]) ? 3'b010 : 3'b110;
										assign node948 = (inp[3]) ? 3'b110 : node949;
											assign node949 = (inp[2]) ? 3'b110 : 3'b010;
						assign node953 = (inp[1]) ? node973 : node954;
							assign node954 = (inp[11]) ? node966 : node955;
								assign node955 = (inp[2]) ? node959 : node956;
									assign node956 = (inp[8]) ? 3'b001 : 3'b110;
									assign node959 = (inp[8]) ? node961 : 3'b010;
										assign node961 = (inp[4]) ? 3'b110 : node962;
											assign node962 = (inp[3]) ? 3'b110 : 3'b111;
								assign node966 = (inp[2]) ? node970 : node967;
									assign node967 = (inp[8]) ? 3'b110 : 3'b010;
									assign node970 = (inp[8]) ? 3'b010 : 3'b100;
							assign node973 = (inp[8]) ? node989 : node974;
								assign node974 = (inp[11]) ? node982 : node975;
									assign node975 = (inp[2]) ? 3'b100 : node976;
										assign node976 = (inp[3]) ? node978 : 3'b010;
											assign node978 = (inp[4]) ? 3'b100 : 3'b000;
									assign node982 = (inp[2]) ? 3'b000 : node983;
										assign node983 = (inp[3]) ? node985 : 3'b100;
											assign node985 = (inp[4]) ? 3'b000 : 3'b100;
								assign node989 = (inp[4]) ? node1005 : node990;
									assign node990 = (inp[3]) ? 3'b010 : node991;
										assign node991 = (inp[5]) ? node999 : node992;
											assign node992 = (inp[11]) ? node996 : node993;
												assign node993 = (inp[2]) ? 3'b010 : 3'b100;
												assign node996 = (inp[2]) ? 3'b100 : 3'b010;
											assign node999 = (inp[2]) ? node1001 : 3'b100;
												assign node1001 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1005 = (inp[2]) ? node1011 : node1006;
										assign node1006 = (inp[5]) ? node1008 : 3'b010;
											assign node1008 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1011 = (inp[5]) ? 3'b010 : 3'b100;
				assign node1014 = (inp[7]) ? node1040 : node1015;
					assign node1015 = (inp[10]) ? 3'b000 : node1016;
						assign node1016 = (inp[8]) ? node1018 : 3'b000;
							assign node1018 = (inp[1]) ? 3'b000 : node1019;
								assign node1019 = (inp[4]) ? node1031 : node1020;
									assign node1020 = (inp[11]) ? node1026 : node1021;
										assign node1021 = (inp[3]) ? 3'b100 : node1022;
											assign node1022 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1026 = (inp[3]) ? 3'b010 : node1027;
											assign node1027 = (inp[2]) ? 3'b010 : 3'b100;
									assign node1031 = (inp[11]) ? 3'b000 : node1032;
										assign node1032 = (inp[3]) ? node1034 : 3'b100;
											assign node1034 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1040 = (inp[10]) ? node1116 : node1041;
						assign node1041 = (inp[1]) ? node1071 : node1042;
							assign node1042 = (inp[8]) ? node1058 : node1043;
								assign node1043 = (inp[4]) ? node1045 : 3'b010;
									assign node1045 = (inp[2]) ? node1051 : node1046;
										assign node1046 = (inp[5]) ? node1048 : 3'b010;
											assign node1048 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1051 = (inp[3]) ? node1053 : 3'b100;
											assign node1053 = (inp[5]) ? node1055 : 3'b000;
												assign node1055 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1058 = (inp[4]) ? node1064 : node1059;
									assign node1059 = (inp[2]) ? node1061 : 3'b110;
										assign node1061 = (inp[11]) ? 3'b100 : 3'b110;
									assign node1064 = (inp[2]) ? node1068 : node1065;
										assign node1065 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1068 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1071 = (inp[11]) ? node1085 : node1072;
								assign node1072 = (inp[8]) ? node1076 : node1073;
									assign node1073 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1076 = (inp[2]) ? node1080 : node1077;
										assign node1077 = (inp[3]) ? 3'b010 : 3'b000;
										assign node1080 = (inp[3]) ? node1082 : 3'b110;
											assign node1082 = (inp[4]) ? 3'b100 : 3'b110;
								assign node1085 = (inp[5]) ? node1103 : node1086;
									assign node1086 = (inp[4]) ? node1098 : node1087;
										assign node1087 = (inp[3]) ? node1093 : node1088;
											assign node1088 = (inp[8]) ? 3'b000 : node1089;
												assign node1089 = (inp[2]) ? 3'b100 : 3'b000;
											assign node1093 = (inp[8]) ? 3'b100 : node1094;
												assign node1094 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1098 = (inp[2]) ? node1100 : 3'b100;
											assign node1100 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1103 = (inp[3]) ? node1105 : 3'b000;
										assign node1105 = (inp[4]) ? node1111 : node1106;
											assign node1106 = (inp[2]) ? 3'b000 : node1107;
												assign node1107 = (inp[8]) ? 3'b100 : 3'b000;
											assign node1111 = (inp[8]) ? 3'b000 : node1112;
												assign node1112 = (inp[2]) ? 3'b100 : 3'b000;
						assign node1116 = (inp[1]) ? 3'b000 : node1117;
							assign node1117 = (inp[8]) ? node1119 : 3'b000;
								assign node1119 = (inp[11]) ? node1127 : node1120;
									assign node1120 = (inp[3]) ? 3'b100 : node1121;
										assign node1121 = (inp[2]) ? 3'b100 : node1122;
											assign node1122 = (inp[4]) ? 3'b010 : 3'b000;
									assign node1127 = (inp[2]) ? 3'b000 : node1128;
										assign node1128 = (inp[3]) ? 3'b000 : 3'b100;

endmodule