module dtc_split33_bm95 (
	input  wire [11-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node159;

	assign outp = (inp[5]) ? node2 : 3'b000;
		assign node2 = (inp[8]) ? node56 : node3;
			assign node3 = (inp[6]) ? node27 : node4;
				assign node4 = (inp[0]) ? 3'b001 : node5;
					assign node5 = (inp[9]) ? node7 : 3'b011;
						assign node7 = (inp[3]) ? node15 : node8;
							assign node8 = (inp[4]) ? node10 : 3'b101;
								assign node10 = (inp[1]) ? node12 : 3'b011;
									assign node12 = (inp[7]) ? 3'b101 : 3'b001;
							assign node15 = (inp[1]) ? node17 : 3'b011;
								assign node17 = (inp[7]) ? node19 : 3'b001;
									assign node19 = (inp[2]) ? node23 : node20;
										assign node20 = (inp[10]) ? 3'b001 : 3'b101;
										assign node23 = (inp[10]) ? 3'b101 : 3'b001;
				assign node27 = (inp[0]) ? node29 : 3'b111;
					assign node29 = (inp[9]) ? node31 : 3'b110;
						assign node31 = (inp[7]) ? node43 : node32;
							assign node32 = (inp[1]) ? 3'b110 : node33;
								assign node33 = (inp[3]) ? node37 : node34;
									assign node34 = (inp[2]) ? 3'b110 : 3'b001;
									assign node37 = (inp[4]) ? 3'b110 : node38;
										assign node38 = (inp[10]) ? 3'b000 : 3'b110;
							assign node43 = (inp[3]) ? node49 : node44;
								assign node44 = (inp[2]) ? node46 : 3'b001;
									assign node46 = (inp[10]) ? 3'b001 : 3'b110;
								assign node49 = (inp[2]) ? node51 : 3'b110;
									assign node51 = (inp[10]) ? node53 : 3'b001;
										assign node53 = (inp[1]) ? 3'b001 : 3'b110;
			assign node56 = (inp[0]) ? node144 : node57;
				assign node57 = (inp[9]) ? node91 : node58;
					assign node58 = (inp[6]) ? node60 : 3'b010;
						assign node60 = (inp[1]) ? node78 : node61;
							assign node61 = (inp[10]) ? node73 : node62;
								assign node62 = (inp[2]) ? node68 : node63;
									assign node63 = (inp[7]) ? 3'b011 : node64;
										assign node64 = (inp[3]) ? 3'b101 : 3'b111;
									assign node68 = (inp[7]) ? 3'b101 : node69;
										assign node69 = (inp[4]) ? 3'b001 : 3'b011;
								assign node73 = (inp[7]) ? 3'b001 : node74;
									assign node74 = (inp[2]) ? 3'b111 : 3'b001;
							assign node78 = (inp[10]) ? node84 : node79;
								assign node79 = (inp[2]) ? 3'b011 : node80;
									assign node80 = (inp[3]) ? 3'b001 : 3'b101;
								assign node84 = (inp[7]) ? 3'b110 : node85;
									assign node85 = (inp[3]) ? 3'b010 : node86;
										assign node86 = (inp[2]) ? 3'b010 : 3'b110;
					assign node91 = (inp[7]) ? node123 : node92;
						assign node92 = (inp[1]) ? node112 : node93;
							assign node93 = (inp[6]) ? node105 : node94;
								assign node94 = (inp[3]) ? node100 : node95;
									assign node95 = (inp[2]) ? 3'b100 : node96;
										assign node96 = (inp[10]) ? 3'b000 : 3'b100;
									assign node100 = (inp[4]) ? node102 : 3'b000;
										assign node102 = (inp[10]) ? 3'b100 : 3'b000;
								assign node105 = (inp[4]) ? 3'b010 : node106;
									assign node106 = (inp[10]) ? 3'b000 : node107;
										assign node107 = (inp[2]) ? 3'b000 : 3'b100;
							assign node112 = (inp[6]) ? node114 : 3'b000;
								assign node114 = (inp[10]) ? node118 : node115;
									assign node115 = (inp[2]) ? 3'b000 : 3'b010;
									assign node118 = (inp[3]) ? 3'b000 : node119;
										assign node119 = (inp[2]) ? 3'b000 : 3'b100;
						assign node123 = (inp[1]) ? node131 : node124;
							assign node124 = (inp[10]) ? 3'b010 : node125;
								assign node125 = (inp[2]) ? 3'b100 : node126;
									assign node126 = (inp[6]) ? 3'b001 : 3'b010;
							assign node131 = (inp[10]) ? node139 : node132;
								assign node132 = (inp[3]) ? node136 : node133;
									assign node133 = (inp[6]) ? 3'b110 : 3'b100;
									assign node136 = (inp[6]) ? 3'b010 : 3'b000;
								assign node139 = (inp[6]) ? 3'b100 : node140;
									assign node140 = (inp[4]) ? 3'b000 : 3'b100;
				assign node144 = (inp[6]) ? node146 : 3'b000;
					assign node146 = (inp[9]) ? 3'b000 : node147;
						assign node147 = (inp[10]) ? node153 : node148;
							assign node148 = (inp[1]) ? 3'b000 : node149;
								assign node149 = (inp[3]) ? 3'b010 : 3'b110;
							assign node153 = (inp[1]) ? node157 : node154;
								assign node154 = (inp[2]) ? 3'b100 : 3'b000;
								assign node157 = (inp[3]) ? node159 : 3'b000;
									assign node159 = (inp[4]) ? 3'b100 : 3'b000;

endmodule