module dtc_split875_bm65 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node25;
	wire [4-1:0] node26;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node38;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node49;
	wire [4-1:0] node51;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node60;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node67;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node79;
	wire [4-1:0] node80;
	wire [4-1:0] node83;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node113;
	wire [4-1:0] node115;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node127;
	wire [4-1:0] node130;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node167;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node191;
	wire [4-1:0] node193;
	wire [4-1:0] node195;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node204;
	wire [4-1:0] node207;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node239;
	wire [4-1:0] node241;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node259;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node328;
	wire [4-1:0] node331;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node335;
	wire [4-1:0] node338;
	wire [4-1:0] node339;
	wire [4-1:0] node343;
	wire [4-1:0] node345;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node356;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node377;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node387;
	wire [4-1:0] node389;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node413;
	wire [4-1:0] node415;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node447;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node461;
	wire [4-1:0] node462;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node471;
	wire [4-1:0] node474;
	wire [4-1:0] node477;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node487;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node493;
	wire [4-1:0] node494;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node507;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node523;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node532;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node551;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node564;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node573;
	wire [4-1:0] node575;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node582;
	wire [4-1:0] node585;
	wire [4-1:0] node587;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node651;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node658;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node664;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node687;
	wire [4-1:0] node689;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node695;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node701;
	wire [4-1:0] node704;
	wire [4-1:0] node705;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node713;
	wire [4-1:0] node715;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node736;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node746;
	wire [4-1:0] node747;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node757;
	wire [4-1:0] node759;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node783;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node797;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node825;
	wire [4-1:0] node827;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node848;
	wire [4-1:0] node849;
	wire [4-1:0] node851;
	wire [4-1:0] node853;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node865;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node876;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node910;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node932;
	wire [4-1:0] node934;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node952;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node983;
	wire [4-1:0] node984;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node992;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1004;
	wire [4-1:0] node1007;
	wire [4-1:0] node1009;
	wire [4-1:0] node1012;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1018;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1052;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1059;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1131;
	wire [4-1:0] node1133;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1150;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1176;
	wire [4-1:0] node1178;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1187;
	wire [4-1:0] node1189;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1194;
	wire [4-1:0] node1196;
	wire [4-1:0] node1198;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1212;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1252;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1262;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1284;
	wire [4-1:0] node1286;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1296;
	wire [4-1:0] node1298;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1312;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1318;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1334;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1344;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1365;
	wire [4-1:0] node1366;
	wire [4-1:0] node1370;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1374;
	wire [4-1:0] node1378;
	wire [4-1:0] node1380;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1387;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1398;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1418;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1431;
	wire [4-1:0] node1435;
	wire [4-1:0] node1437;
	wire [4-1:0] node1439;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1455;
	wire [4-1:0] node1457;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1469;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1488;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1500;
	wire [4-1:0] node1501;
	wire [4-1:0] node1505;
	wire [4-1:0] node1507;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1513;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1520;
	wire [4-1:0] node1523;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1530;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1544;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1555;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1561;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1574;
	wire [4-1:0] node1576;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1582;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1592;
	wire [4-1:0] node1594;
	wire [4-1:0] node1597;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1606;
	wire [4-1:0] node1608;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1622;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1632;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1638;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1657;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1666;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1674;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1679;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1693;
	wire [4-1:0] node1696;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1715;
	wire [4-1:0] node1718;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1727;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1735;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1745;
	wire [4-1:0] node1748;
	wire [4-1:0] node1751;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1757;
	wire [4-1:0] node1760;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1765;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1772;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1782;
	wire [4-1:0] node1785;
	wire [4-1:0] node1786;
	wire [4-1:0] node1787;
	wire [4-1:0] node1791;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1809;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1814;
	wire [4-1:0] node1817;
	wire [4-1:0] node1819;
	wire [4-1:0] node1822;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1833;
	wire [4-1:0] node1836;
	wire [4-1:0] node1837;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1854;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1889;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1896;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1901;
	wire [4-1:0] node1902;
	wire [4-1:0] node1904;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1911;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1922;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1929;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1938;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1946;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1957;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1963;
	wire [4-1:0] node1966;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1973;
	wire [4-1:0] node1976;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1982;
	wire [4-1:0] node1985;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1992;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2013;
	wire [4-1:0] node2016;
	wire [4-1:0] node2017;
	wire [4-1:0] node2019;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2035;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2047;
	wire [4-1:0] node2049;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2062;
	wire [4-1:0] node2063;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2069;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2076;
	wire [4-1:0] node2079;
	wire [4-1:0] node2080;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2098;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2104;
	wire [4-1:0] node2106;
	wire [4-1:0] node2108;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2123;
	wire [4-1:0] node2125;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2141;
	wire [4-1:0] node2144;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2177;
	wire [4-1:0] node2180;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2187;
	wire [4-1:0] node2190;
	wire [4-1:0] node2191;
	wire [4-1:0] node2192;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2208;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2213;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2230;
	wire [4-1:0] node2232;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2244;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2279;
	wire [4-1:0] node2281;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2288;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2296;
	wire [4-1:0] node2297;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2305;
	wire [4-1:0] node2306;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2310;
	wire [4-1:0] node2313;
	wire [4-1:0] node2314;
	wire [4-1:0] node2316;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2325;
	wire [4-1:0] node2328;
	wire [4-1:0] node2329;
	wire [4-1:0] node2330;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2341;
	wire [4-1:0] node2342;
	wire [4-1:0] node2345;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2353;
	wire [4-1:0] node2356;
	wire [4-1:0] node2357;
	wire [4-1:0] node2360;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2366;
	wire [4-1:0] node2369;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2382;
	wire [4-1:0] node2385;
	wire [4-1:0] node2388;
	wire [4-1:0] node2389;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2398;
	wire [4-1:0] node2399;
	wire [4-1:0] node2402;
	wire [4-1:0] node2405;
	wire [4-1:0] node2406;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2416;
	wire [4-1:0] node2417;
	wire [4-1:0] node2419;
	wire [4-1:0] node2422;
	wire [4-1:0] node2425;
	wire [4-1:0] node2427;
	wire [4-1:0] node2428;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2435;
	wire [4-1:0] node2437;
	wire [4-1:0] node2440;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2463;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2482;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2493;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2501;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2518;
	wire [4-1:0] node2520;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2526;
	wire [4-1:0] node2529;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2537;
	wire [4-1:0] node2538;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2543;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2554;
	wire [4-1:0] node2557;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2563;
	wire [4-1:0] node2566;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2573;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2585;
	wire [4-1:0] node2586;
	wire [4-1:0] node2587;
	wire [4-1:0] node2588;
	wire [4-1:0] node2590;
	wire [4-1:0] node2593;
	wire [4-1:0] node2594;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2601;
	wire [4-1:0] node2604;
	wire [4-1:0] node2606;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2618;
	wire [4-1:0] node2620;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2627;
	wire [4-1:0] node2628;
	wire [4-1:0] node2632;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2635;
	wire [4-1:0] node2636;
	wire [4-1:0] node2640;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2652;
	wire [4-1:0] node2654;
	wire [4-1:0] node2657;
	wire [4-1:0] node2658;
	wire [4-1:0] node2659;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2673;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2686;
	wire [4-1:0] node2687;
	wire [4-1:0] node2689;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2695;
	wire [4-1:0] node2698;
	wire [4-1:0] node2700;
	wire [4-1:0] node2703;
	wire [4-1:0] node2704;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2710;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2724;
	wire [4-1:0] node2725;
	wire [4-1:0] node2728;
	wire [4-1:0] node2731;
	wire [4-1:0] node2732;
	wire [4-1:0] node2733;
	wire [4-1:0] node2735;
	wire [4-1:0] node2738;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2746;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2753;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2758;
	wire [4-1:0] node2759;
	wire [4-1:0] node2760;
	wire [4-1:0] node2763;
	wire [4-1:0] node2766;
	wire [4-1:0] node2768;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2783;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2788;
	wire [4-1:0] node2789;
	wire [4-1:0] node2793;
	wire [4-1:0] node2794;
	wire [4-1:0] node2797;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2807;
	wire [4-1:0] node2811;
	wire [4-1:0] node2812;
	wire [4-1:0] node2813;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2819;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2826;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2833;
	wire [4-1:0] node2834;
	wire [4-1:0] node2838;
	wire [4-1:0] node2839;
	wire [4-1:0] node2840;
	wire [4-1:0] node2843;
	wire [4-1:0] node2846;
	wire [4-1:0] node2847;
	wire [4-1:0] node2849;
	wire [4-1:0] node2852;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2862;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2869;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2876;
	wire [4-1:0] node2877;
	wire [4-1:0] node2881;
	wire [4-1:0] node2882;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2888;
	wire [4-1:0] node2890;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2910;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2919;
	wire [4-1:0] node2920;
	wire [4-1:0] node2921;
	wire [4-1:0] node2923;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2930;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2936;
	wire [4-1:0] node2939;
	wire [4-1:0] node2940;
	wire [4-1:0] node2944;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2947;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2960;
	wire [4-1:0] node2963;
	wire [4-1:0] node2964;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2974;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2981;
	wire [4-1:0] node2984;
	wire [4-1:0] node2985;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2993;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2997;
	wire [4-1:0] node2998;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3010;
	wire [4-1:0] node3012;
	wire [4-1:0] node3013;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3021;
	wire [4-1:0] node3024;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3036;
	wire [4-1:0] node3039;
	wire [4-1:0] node3040;
	wire [4-1:0] node3042;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3054;
	wire [4-1:0] node3055;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3060;
	wire [4-1:0] node3063;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3070;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3075;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3082;
	wire [4-1:0] node3085;
	wire [4-1:0] node3086;
	wire [4-1:0] node3087;
	wire [4-1:0] node3089;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3102;
	wire [4-1:0] node3105;
	wire [4-1:0] node3106;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3114;
	wire [4-1:0] node3116;
	wire [4-1:0] node3118;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3130;
	wire [4-1:0] node3133;
	wire [4-1:0] node3136;
	wire [4-1:0] node3137;
	wire [4-1:0] node3140;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3147;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3152;
	wire [4-1:0] node3156;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3171;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3180;
	wire [4-1:0] node3181;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3186;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3197;
	wire [4-1:0] node3198;
	wire [4-1:0] node3202;
	wire [4-1:0] node3204;
	wire [4-1:0] node3207;
	wire [4-1:0] node3209;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3214;
	wire [4-1:0] node3218;
	wire [4-1:0] node3219;
	wire [4-1:0] node3221;
	wire [4-1:0] node3224;
	wire [4-1:0] node3226;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3240;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3246;
	wire [4-1:0] node3250;
	wire [4-1:0] node3251;
	wire [4-1:0] node3255;
	wire [4-1:0] node3256;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3270;
	wire [4-1:0] node3272;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3282;
	wire [4-1:0] node3283;
	wire [4-1:0] node3284;
	wire [4-1:0] node3286;
	wire [4-1:0] node3289;
	wire [4-1:0] node3291;
	wire [4-1:0] node3294;
	wire [4-1:0] node3296;
	wire [4-1:0] node3298;
	wire [4-1:0] node3301;
	wire [4-1:0] node3302;
	wire [4-1:0] node3304;
	wire [4-1:0] node3307;
	wire [4-1:0] node3309;
	wire [4-1:0] node3312;
	wire [4-1:0] node3313;
	wire [4-1:0] node3314;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3328;
	wire [4-1:0] node3330;
	wire [4-1:0] node3333;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3337;
	wire [4-1:0] node3339;
	wire [4-1:0] node3342;
	wire [4-1:0] node3344;
	wire [4-1:0] node3346;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3352;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3357;
	wire [4-1:0] node3361;
	wire [4-1:0] node3363;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3373;
	wire [4-1:0] node3377;
	wire [4-1:0] node3378;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3385;
	wire [4-1:0] node3387;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3395;
	wire [4-1:0] node3397;
	wire [4-1:0] node3400;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3404;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3410;
	wire [4-1:0] node3414;
	wire [4-1:0] node3415;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3422;
	wire [4-1:0] node3424;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3430;
	wire [4-1:0] node3433;
	wire [4-1:0] node3435;
	wire [4-1:0] node3438;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3446;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3455;
	wire [4-1:0] node3457;
	wire [4-1:0] node3458;
	wire [4-1:0] node3459;
	wire [4-1:0] node3463;
	wire [4-1:0] node3465;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3471;
	wire [4-1:0] node3473;
	wire [4-1:0] node3476;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3488;
	wire [4-1:0] node3489;
	wire [4-1:0] node3493;
	wire [4-1:0] node3495;
	wire [4-1:0] node3499;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3505;
	wire [4-1:0] node3506;
	wire [4-1:0] node3507;
	wire [4-1:0] node3508;
	wire [4-1:0] node3509;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3517;
	wire [4-1:0] node3520;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3526;
	wire [4-1:0] node3529;
	wire [4-1:0] node3530;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3546;
	wire [4-1:0] node3549;
	wire [4-1:0] node3551;
	wire [4-1:0] node3554;
	wire [4-1:0] node3555;
	wire [4-1:0] node3556;
	wire [4-1:0] node3560;
	wire [4-1:0] node3562;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3570;
	wire [4-1:0] node3572;
	wire [4-1:0] node3576;
	wire [4-1:0] node3577;
	wire [4-1:0] node3581;
	wire [4-1:0] node3582;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3588;
	wire [4-1:0] node3590;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3596;
	wire [4-1:0] node3599;
	wire [4-1:0] node3601;
	wire [4-1:0] node3604;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3607;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3614;
	wire [4-1:0] node3615;
	wire [4-1:0] node3620;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3623;
	wire [4-1:0] node3627;
	wire [4-1:0] node3629;
	wire [4-1:0] node3632;
	wire [4-1:0] node3633;
	wire [4-1:0] node3638;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3641;
	wire [4-1:0] node3642;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3650;
	wire [4-1:0] node3653;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3658;
	wire [4-1:0] node3661;
	wire [4-1:0] node3664;
	wire [4-1:0] node3665;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3674;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3681;
	wire [4-1:0] node3684;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3694;
	wire [4-1:0] node3695;
	wire [4-1:0] node3697;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3705;
	wire [4-1:0] node3709;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3716;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3725;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3733;
	wire [4-1:0] node3734;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3744;
	wire [4-1:0] node3746;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3761;
	wire [4-1:0] node3762;
	wire [4-1:0] node3765;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3773;
	wire [4-1:0] node3774;
	wire [4-1:0] node3777;
	wire [4-1:0] node3778;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3785;
	wire [4-1:0] node3786;
	wire [4-1:0] node3788;
	wire [4-1:0] node3790;
	wire [4-1:0] node3793;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3805;
	wire [4-1:0] node3807;
	wire [4-1:0] node3810;
	wire [4-1:0] node3812;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3825;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3833;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3840;
	wire [4-1:0] node3844;
	wire [4-1:0] node3846;
	wire [4-1:0] node3849;
	wire [4-1:0] node3850;
	wire [4-1:0] node3852;
	wire [4-1:0] node3855;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3861;
	wire [4-1:0] node3862;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3870;
	wire [4-1:0] node3872;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3883;
	wire [4-1:0] node3884;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3891;
	wire [4-1:0] node3892;
	wire [4-1:0] node3897;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3917;
	wire [4-1:0] node3918;
	wire [4-1:0] node3919;
	wire [4-1:0] node3921;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3928;
	wire [4-1:0] node3931;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3936;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3943;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3948;
	wire [4-1:0] node3951;
	wire [4-1:0] node3954;
	wire [4-1:0] node3955;
	wire [4-1:0] node3958;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3963;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3968;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3975;
	wire [4-1:0] node3978;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3987;
	wire [4-1:0] node3991;
	wire [4-1:0] node3992;
	wire [4-1:0] node3993;
	wire [4-1:0] node3996;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4003;
	wire [4-1:0] node4006;
	wire [4-1:0] node4007;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4013;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4022;
	wire [4-1:0] node4024;
	wire [4-1:0] node4027;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4037;
	wire [4-1:0] node4038;
	wire [4-1:0] node4040;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4066;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4069;
	wire [4-1:0] node4072;
	wire [4-1:0] node4075;
	wire [4-1:0] node4076;
	wire [4-1:0] node4079;
	wire [4-1:0] node4082;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4095;
	wire [4-1:0] node4096;
	wire [4-1:0] node4097;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4109;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4124;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4132;
	wire [4-1:0] node4133;
	wire [4-1:0] node4134;
	wire [4-1:0] node4135;
	wire [4-1:0] node4139;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4145;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4151;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4159;
	wire [4-1:0] node4160;
	wire [4-1:0] node4161;
	wire [4-1:0] node4162;
	wire [4-1:0] node4165;
	wire [4-1:0] node4166;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4176;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4182;
	wire [4-1:0] node4184;
	wire [4-1:0] node4187;
	wire [4-1:0] node4188;
	wire [4-1:0] node4189;
	wire [4-1:0] node4192;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4200;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4205;
	wire [4-1:0] node4208;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4213;
	wire [4-1:0] node4216;
	wire [4-1:0] node4217;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4227;
	wire [4-1:0] node4230;
	wire [4-1:0] node4233;
	wire [4-1:0] node4234;
	wire [4-1:0] node4236;
	wire [4-1:0] node4239;
	wire [4-1:0] node4241;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4249;
	wire [4-1:0] node4253;
	wire [4-1:0] node4254;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4261;
	wire [4-1:0] node4264;
	wire [4-1:0] node4265;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4270;
	wire [4-1:0] node4274;
	wire [4-1:0] node4275;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4282;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4301;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4309;
	wire [4-1:0] node4312;
	wire [4-1:0] node4315;
	wire [4-1:0] node4317;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4332;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4347;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4353;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4361;
	wire [4-1:0] node4363;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4370;
	wire [4-1:0] node4373;
	wire [4-1:0] node4374;
	wire [4-1:0] node4377;
	wire [4-1:0] node4378;
	wire [4-1:0] node4381;
	wire [4-1:0] node4384;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4390;
	wire [4-1:0] node4391;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4397;
	wire [4-1:0] node4401;
	wire [4-1:0] node4402;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4409;
	wire [4-1:0] node4412;
	wire [4-1:0] node4415;
	wire [4-1:0] node4416;
	wire [4-1:0] node4420;
	wire [4-1:0] node4423;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4428;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4436;
	wire [4-1:0] node4439;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4444;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4456;
	wire [4-1:0] node4459;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4466;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4482;
	wire [4-1:0] node4485;
	wire [4-1:0] node4486;
	wire [4-1:0] node4487;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4495;
	wire [4-1:0] node4498;
	wire [4-1:0] node4499;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4513;
	wire [4-1:0] node4516;
	wire [4-1:0] node4518;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4528;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4538;
	wire [4-1:0] node4542;
	wire [4-1:0] node4543;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4550;
	wire [4-1:0] node4552;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4558;
	wire [4-1:0] node4561;
	wire [4-1:0] node4562;
	wire [4-1:0] node4567;
	wire [4-1:0] node4568;
	wire [4-1:0] node4569;
	wire [4-1:0] node4570;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4573;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4576;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4585;
	wire [4-1:0] node4586;
	wire [4-1:0] node4587;
	wire [4-1:0] node4591;
	wire [4-1:0] node4593;
	wire [4-1:0] node4596;
	wire [4-1:0] node4597;
	wire [4-1:0] node4598;
	wire [4-1:0] node4601;
	wire [4-1:0] node4604;
	wire [4-1:0] node4606;
	wire [4-1:0] node4609;
	wire [4-1:0] node4610;
	wire [4-1:0] node4611;
	wire [4-1:0] node4612;
	wire [4-1:0] node4613;
	wire [4-1:0] node4616;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4628;
	wire [4-1:0] node4630;
	wire [4-1:0] node4633;
	wire [4-1:0] node4634;
	wire [4-1:0] node4635;
	wire [4-1:0] node4636;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4651;
	wire [4-1:0] node4653;
	wire [4-1:0] node4656;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4660;
	wire [4-1:0] node4664;
	wire [4-1:0] node4665;
	wire [4-1:0] node4669;
	wire [4-1:0] node4670;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4683;
	wire [4-1:0] node4686;
	wire [4-1:0] node4689;
	wire [4-1:0] node4690;
	wire [4-1:0] node4692;
	wire [4-1:0] node4695;
	wire [4-1:0] node4698;
	wire [4-1:0] node4699;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4705;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4711;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4715;
	wire [4-1:0] node4718;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4725;
	wire [4-1:0] node4727;
	wire [4-1:0] node4728;
	wire [4-1:0] node4731;
	wire [4-1:0] node4734;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4738;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4745;
	wire [4-1:0] node4748;
	wire [4-1:0] node4749;
	wire [4-1:0] node4750;
	wire [4-1:0] node4753;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4760;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4770;
	wire [4-1:0] node4773;
	wire [4-1:0] node4775;
	wire [4-1:0] node4778;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4782;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4789;
	wire [4-1:0] node4792;
	wire [4-1:0] node4794;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4800;
	wire [4-1:0] node4803;
	wire [4-1:0] node4804;
	wire [4-1:0] node4807;
	wire [4-1:0] node4810;
	wire [4-1:0] node4811;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4814;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4820;
	wire [4-1:0] node4823;
	wire [4-1:0] node4826;
	wire [4-1:0] node4829;
	wire [4-1:0] node4830;
	wire [4-1:0] node4832;
	wire [4-1:0] node4834;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4841;
	wire [4-1:0] node4842;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4848;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4854;
	wire [4-1:0] node4856;
	wire [4-1:0] node4859;
	wire [4-1:0] node4861;
	wire [4-1:0] node4863;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4872;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4880;
	wire [4-1:0] node4881;
	wire [4-1:0] node4884;
	wire [4-1:0] node4887;
	wire [4-1:0] node4888;
	wire [4-1:0] node4889;
	wire [4-1:0] node4891;
	wire [4-1:0] node4894;
	wire [4-1:0] node4895;
	wire [4-1:0] node4896;
	wire [4-1:0] node4899;
	wire [4-1:0] node4903;
	wire [4-1:0] node4904;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4911;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4918;
	wire [4-1:0] node4919;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4926;
	wire [4-1:0] node4929;
	wire [4-1:0] node4930;
	wire [4-1:0] node4932;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4943;
	wire [4-1:0] node4945;
	wire [4-1:0] node4949;
	wire [4-1:0] node4950;
	wire [4-1:0] node4951;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4958;
	wire [4-1:0] node4961;
	wire [4-1:0] node4962;
	wire [4-1:0] node4963;
	wire [4-1:0] node4966;
	wire [4-1:0] node4967;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4974;
	wire [4-1:0] node4977;
	wire [4-1:0] node4980;
	wire [4-1:0] node4981;
	wire [4-1:0] node4982;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4989;
	wire [4-1:0] node4990;
	wire [4-1:0] node4993;
	wire [4-1:0] node4996;
	wire [4-1:0] node4997;
	wire [4-1:0] node4998;
	wire [4-1:0] node5000;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5009;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5013;
	wire [4-1:0] node5014;
	wire [4-1:0] node5015;
	wire [4-1:0] node5016;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5028;
	wire [4-1:0] node5029;
	wire [4-1:0] node5033;
	wire [4-1:0] node5035;
	wire [4-1:0] node5038;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5042;
	wire [4-1:0] node5045;
	wire [4-1:0] node5046;
	wire [4-1:0] node5048;
	wire [4-1:0] node5051;
	wire [4-1:0] node5052;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5072;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5075;
	wire [4-1:0] node5077;
	wire [4-1:0] node5081;
	wire [4-1:0] node5082;
	wire [4-1:0] node5086;
	wire [4-1:0] node5087;
	wire [4-1:0] node5088;
	wire [4-1:0] node5089;
	wire [4-1:0] node5094;
	wire [4-1:0] node5096;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5102;
	wire [4-1:0] node5103;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5116;
	wire [4-1:0] node5117;
	wire [4-1:0] node5121;
	wire [4-1:0] node5122;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5130;
	wire [4-1:0] node5131;
	wire [4-1:0] node5135;
	wire [4-1:0] node5137;
	wire [4-1:0] node5140;
	wire [4-1:0] node5141;
	wire [4-1:0] node5144;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5154;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5161;
	wire [4-1:0] node5162;
	wire [4-1:0] node5163;
	wire [4-1:0] node5164;
	wire [4-1:0] node5165;
	wire [4-1:0] node5167;
	wire [4-1:0] node5168;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5176;
	wire [4-1:0] node5180;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5186;
	wire [4-1:0] node5189;
	wire [4-1:0] node5190;
	wire [4-1:0] node5191;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5197;
	wire [4-1:0] node5200;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5208;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5214;
	wire [4-1:0] node5218;
	wire [4-1:0] node5219;
	wire [4-1:0] node5223;
	wire [4-1:0] node5224;
	wire [4-1:0] node5227;
	wire [4-1:0] node5230;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5237;
	wire [4-1:0] node5240;
	wire [4-1:0] node5243;
	wire [4-1:0] node5244;
	wire [4-1:0] node5245;
	wire [4-1:0] node5246;
	wire [4-1:0] node5250;
	wire [4-1:0] node5251;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5258;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5265;
	wire [4-1:0] node5266;
	wire [4-1:0] node5267;
	wire [4-1:0] node5270;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5276;
	wire [4-1:0] node5279;
	wire [4-1:0] node5281;
	wire [4-1:0] node5284;
	wire [4-1:0] node5285;
	wire [4-1:0] node5288;
	wire [4-1:0] node5290;
	wire [4-1:0] node5292;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5300;
	wire [4-1:0] node5303;
	wire [4-1:0] node5306;
	wire [4-1:0] node5307;
	wire [4-1:0] node5310;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5320;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5329;
	wire [4-1:0] node5331;
	wire [4-1:0] node5334;
	wire [4-1:0] node5335;
	wire [4-1:0] node5337;
	wire [4-1:0] node5340;
	wire [4-1:0] node5341;
	wire [4-1:0] node5344;
	wire [4-1:0] node5347;
	wire [4-1:0] node5348;
	wire [4-1:0] node5349;
	wire [4-1:0] node5350;
	wire [4-1:0] node5351;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5360;
	wire [4-1:0] node5363;
	wire [4-1:0] node5364;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5369;
	wire [4-1:0] node5372;
	wire [4-1:0] node5374;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5379;
	wire [4-1:0] node5381;
	wire [4-1:0] node5384;
	wire [4-1:0] node5385;
	wire [4-1:0] node5389;
	wire [4-1:0] node5390;
	wire [4-1:0] node5391;
	wire [4-1:0] node5395;
	wire [4-1:0] node5397;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5403;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5407;
	wire [4-1:0] node5408;
	wire [4-1:0] node5411;
	wire [4-1:0] node5414;
	wire [4-1:0] node5415;
	wire [4-1:0] node5418;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5428;
	wire [4-1:0] node5431;
	wire [4-1:0] node5433;
	wire [4-1:0] node5435;
	wire [4-1:0] node5438;
	wire [4-1:0] node5439;
	wire [4-1:0] node5440;
	wire [4-1:0] node5442;
	wire [4-1:0] node5444;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5449;
	wire [4-1:0] node5453;
	wire [4-1:0] node5454;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5465;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5470;
	wire [4-1:0] node5473;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5484;
	wire [4-1:0] node5485;
	wire [4-1:0] node5489;
	wire [4-1:0] node5491;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5500;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5507;
	wire [4-1:0] node5510;
	wire [4-1:0] node5511;
	wire [4-1:0] node5514;
	wire [4-1:0] node5517;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5523;
	wire [4-1:0] node5526;
	wire [4-1:0] node5528;
	wire [4-1:0] node5531;
	wire [4-1:0] node5532;
	wire [4-1:0] node5533;
	wire [4-1:0] node5537;
	wire [4-1:0] node5539;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5544;
	wire [4-1:0] node5545;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5549;
	wire [4-1:0] node5552;
	wire [4-1:0] node5553;
	wire [4-1:0] node5557;
	wire [4-1:0] node5559;
	wire [4-1:0] node5562;
	wire [4-1:0] node5564;
	wire [4-1:0] node5566;
	wire [4-1:0] node5567;
	wire [4-1:0] node5570;
	wire [4-1:0] node5573;
	wire [4-1:0] node5574;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5580;
	wire [4-1:0] node5583;
	wire [4-1:0] node5584;
	wire [4-1:0] node5585;
	wire [4-1:0] node5588;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5596;
	wire [4-1:0] node5597;
	wire [4-1:0] node5598;
	wire [4-1:0] node5599;
	wire [4-1:0] node5601;
	wire [4-1:0] node5604;
	wire [4-1:0] node5606;
	wire [4-1:0] node5609;
	wire [4-1:0] node5610;
	wire [4-1:0] node5611;
	wire [4-1:0] node5613;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5625;
	wire [4-1:0] node5627;
	wire [4-1:0] node5631;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5634;
	wire [4-1:0] node5635;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5638;
	wire [4-1:0] node5642;
	wire [4-1:0] node5644;
	wire [4-1:0] node5645;
	wire [4-1:0] node5649;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5653;
	wire [4-1:0] node5657;
	wire [4-1:0] node5659;
	wire [4-1:0] node5661;
	wire [4-1:0] node5664;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5667;
	wire [4-1:0] node5668;
	wire [4-1:0] node5671;
	wire [4-1:0] node5675;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5682;
	wire [4-1:0] node5683;
	wire [4-1:0] node5685;
	wire [4-1:0] node5686;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5694;
	wire [4-1:0] node5697;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5700;
	wire [4-1:0] node5702;
	wire [4-1:0] node5705;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5722;
	wire [4-1:0] node5723;
	wire [4-1:0] node5725;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5737;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5744;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5750;
	wire [4-1:0] node5754;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5760;
	wire [4-1:0] node5761;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5768;
	wire [4-1:0] node5771;
	wire [4-1:0] node5773;
	wire [4-1:0] node5776;
	wire [4-1:0] node5777;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5783;
	wire [4-1:0] node5786;
	wire [4-1:0] node5787;
	wire [4-1:0] node5788;
	wire [4-1:0] node5791;
	wire [4-1:0] node5795;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5800;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5808;
	wire [4-1:0] node5809;
	wire [4-1:0] node5812;
	wire [4-1:0] node5815;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5818;
	wire [4-1:0] node5822;
	wire [4-1:0] node5823;
	wire [4-1:0] node5826;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5834;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5840;
	wire [4-1:0] node5842;
	wire [4-1:0] node5844;
	wire [4-1:0] node5845;
	wire [4-1:0] node5849;
	wire [4-1:0] node5850;
	wire [4-1:0] node5851;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5859;
	wire [4-1:0] node5861;
	wire [4-1:0] node5864;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5868;
	wire [4-1:0] node5870;
	wire [4-1:0] node5873;
	wire [4-1:0] node5876;
	wire [4-1:0] node5877;
	wire [4-1:0] node5878;
	wire [4-1:0] node5881;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5887;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5895;
	wire [4-1:0] node5897;
	wire [4-1:0] node5900;
	wire [4-1:0] node5901;
	wire [4-1:0] node5903;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5910;
	wire [4-1:0] node5912;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5918;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5926;
	wire [4-1:0] node5930;
	wire [4-1:0] node5931;
	wire [4-1:0] node5932;
	wire [4-1:0] node5935;
	wire [4-1:0] node5938;
	wire [4-1:0] node5939;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5945;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5959;
	wire [4-1:0] node5961;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5970;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5981;
	wire [4-1:0] node5984;
	wire [4-1:0] node5985;
	wire [4-1:0] node5988;
	wire [4-1:0] node5991;
	wire [4-1:0] node5992;
	wire [4-1:0] node5993;
	wire [4-1:0] node5994;
	wire [4-1:0] node5995;
	wire [4-1:0] node5997;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6003;
	wire [4-1:0] node6008;
	wire [4-1:0] node6009;
	wire [4-1:0] node6011;
	wire [4-1:0] node6013;
	wire [4-1:0] node6016;
	wire [4-1:0] node6017;
	wire [4-1:0] node6019;
	wire [4-1:0] node6022;
	wire [4-1:0] node6023;
	wire [4-1:0] node6028;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6036;
	wire [4-1:0] node6037;
	wire [4-1:0] node6041;
	wire [4-1:0] node6045;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6050;
	wire [4-1:0] node6052;
	wire [4-1:0] node6055;
	wire [4-1:0] node6056;
	wire [4-1:0] node6059;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6064;
	wire [4-1:0] node6065;
	wire [4-1:0] node6068;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6074;
	wire [4-1:0] node6078;
	wire [4-1:0] node6079;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6085;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6091;
	wire [4-1:0] node6094;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6102;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6107;
	wire [4-1:0] node6110;
	wire [4-1:0] node6113;
	wire [4-1:0] node6114;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6121;
	wire [4-1:0] node6123;
	wire [4-1:0] node6126;
	wire [4-1:0] node6127;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6134;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6140;
	wire [4-1:0] node6143;
	wire [4-1:0] node6144;
	wire [4-1:0] node6147;
	wire [4-1:0] node6150;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6157;
	wire [4-1:0] node6158;
	wire [4-1:0] node6160;
	wire [4-1:0] node6163;
	wire [4-1:0] node6165;
	wire [4-1:0] node6168;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6174;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6186;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6194;
	wire [4-1:0] node6195;
	wire [4-1:0] node6196;
	wire [4-1:0] node6201;
	wire [4-1:0] node6202;
	wire [4-1:0] node6203;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6209;
	wire [4-1:0] node6211;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6216;
	wire [4-1:0] node6220;
	wire [4-1:0] node6222;
	wire [4-1:0] node6225;
	wire [4-1:0] node6226;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6231;
	wire [4-1:0] node6234;
	wire [4-1:0] node6236;
	wire [4-1:0] node6239;
	wire [4-1:0] node6241;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6247;
	wire [4-1:0] node6249;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6257;
	wire [4-1:0] node6258;
	wire [4-1:0] node6260;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6267;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6272;
	wire [4-1:0] node6273;
	wire [4-1:0] node6277;
	wire [4-1:0] node6279;
	wire [4-1:0] node6282;
	wire [4-1:0] node6283;
	wire [4-1:0] node6285;
	wire [4-1:0] node6288;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6296;
	wire [4-1:0] node6297;
	wire [4-1:0] node6298;
	wire [4-1:0] node6299;
	wire [4-1:0] node6301;
	wire [4-1:0] node6304;
	wire [4-1:0] node6306;
	wire [4-1:0] node6310;
	wire [4-1:0] node6311;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6317;
	wire [4-1:0] node6320;
	wire [4-1:0] node6321;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6329;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6334;
	wire [4-1:0] node6337;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6343;
	wire [4-1:0] node6346;
	wire [4-1:0] node6347;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6363;
	wire [4-1:0] node6365;
	wire [4-1:0] node6366;
	wire [4-1:0] node6370;
	wire [4-1:0] node6371;
	wire [4-1:0] node6372;
	wire [4-1:0] node6373;
	wire [4-1:0] node6376;
	wire [4-1:0] node6379;
	wire [4-1:0] node6380;
	wire [4-1:0] node6381;
	wire [4-1:0] node6383;
	wire [4-1:0] node6386;
	wire [4-1:0] node6389;
	wire [4-1:0] node6390;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6398;
	wire [4-1:0] node6399;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6402;
	wire [4-1:0] node6406;
	wire [4-1:0] node6407;
	wire [4-1:0] node6411;
	wire [4-1:0] node6412;
	wire [4-1:0] node6414;
	wire [4-1:0] node6417;
	wire [4-1:0] node6420;
	wire [4-1:0] node6421;
	wire [4-1:0] node6422;
	wire [4-1:0] node6425;
	wire [4-1:0] node6428;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6433;
	wire [4-1:0] node6436;
	wire [4-1:0] node6437;
	wire [4-1:0] node6440;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6450;
	wire [4-1:0] node6454;
	wire [4-1:0] node6455;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6463;
	wire [4-1:0] node6464;
	wire [4-1:0] node6465;
	wire [4-1:0] node6468;
	wire [4-1:0] node6471;
	wire [4-1:0] node6473;
	wire [4-1:0] node6476;
	wire [4-1:0] node6477;
	wire [4-1:0] node6478;
	wire [4-1:0] node6479;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6487;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6493;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6500;
	wire [4-1:0] node6504;
	wire [4-1:0] node6505;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6510;
	wire [4-1:0] node6512;
	wire [4-1:0] node6515;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6522;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6527;
	wire [4-1:0] node6529;
	wire [4-1:0] node6532;
	wire [4-1:0] node6533;
	wire [4-1:0] node6534;
	wire [4-1:0] node6537;
	wire [4-1:0] node6540;
	wire [4-1:0] node6541;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6548;
	wire [4-1:0] node6550;
	wire [4-1:0] node6554;
	wire [4-1:0] node6555;
	wire [4-1:0] node6556;
	wire [4-1:0] node6559;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6566;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6571;
	wire [4-1:0] node6574;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6579;
	wire [4-1:0] node6582;
	wire [4-1:0] node6585;
	wire [4-1:0] node6587;
	wire [4-1:0] node6590;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6593;
	wire [4-1:0] node6594;
	wire [4-1:0] node6598;
	wire [4-1:0] node6600;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6609;
	wire [4-1:0] node6612;
	wire [4-1:0] node6613;
	wire [4-1:0] node6616;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6631;
	wire [4-1:0] node6634;
	wire [4-1:0] node6635;
	wire [4-1:0] node6639;
	wire [4-1:0] node6641;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6652;
	wire [4-1:0] node6653;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6662;
	wire [4-1:0] node6664;
	wire [4-1:0] node6668;
	wire [4-1:0] node6669;
	wire [4-1:0] node6671;
	wire [4-1:0] node6675;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6682;
	wire [4-1:0] node6683;
	wire [4-1:0] node6687;
	wire [4-1:0] node6689;
	wire [4-1:0] node6691;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6704;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6720;
	wire [4-1:0] node6721;
	wire [4-1:0] node6723;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6734;
	wire [4-1:0] node6735;
	wire [4-1:0] node6738;
	wire [4-1:0] node6741;
	wire [4-1:0] node6743;
	wire [4-1:0] node6746;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6754;
	wire [4-1:0] node6756;
	wire [4-1:0] node6759;
	wire [4-1:0] node6761;
	wire [4-1:0] node6762;
	wire [4-1:0] node6763;
	wire [4-1:0] node6766;
	wire [4-1:0] node6769;
	wire [4-1:0] node6771;
	wire [4-1:0] node6774;
	wire [4-1:0] node6775;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6782;
	wire [4-1:0] node6785;
	wire [4-1:0] node6786;
	wire [4-1:0] node6790;
	wire [4-1:0] node6791;
	wire [4-1:0] node6792;
	wire [4-1:0] node6793;
	wire [4-1:0] node6796;
	wire [4-1:0] node6799;
	wire [4-1:0] node6801;
	wire [4-1:0] node6804;
	wire [4-1:0] node6806;
	wire [4-1:0] node6808;
	wire [4-1:0] node6813;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6817;
	wire [4-1:0] node6818;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6821;
	wire [4-1:0] node6823;
	wire [4-1:0] node6824;
	wire [4-1:0] node6825;
	wire [4-1:0] node6826;
	wire [4-1:0] node6829;
	wire [4-1:0] node6831;
	wire [4-1:0] node6835;
	wire [4-1:0] node6836;
	wire [4-1:0] node6837;
	wire [4-1:0] node6839;
	wire [4-1:0] node6843;
	wire [4-1:0] node6844;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6853;
	wire [4-1:0] node6855;
	wire [4-1:0] node6858;
	wire [4-1:0] node6859;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6867;
	wire [4-1:0] node6868;
	wire [4-1:0] node6870;
	wire [4-1:0] node6871;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6880;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6888;
	wire [4-1:0] node6890;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6900;
	wire [4-1:0] node6902;
	wire [4-1:0] node6905;
	wire [4-1:0] node6907;
	wire [4-1:0] node6910;
	wire [4-1:0] node6912;
	wire [4-1:0] node6915;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6924;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6933;
	wire [4-1:0] node6937;
	wire [4-1:0] node6939;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6944;
	wire [4-1:0] node6945;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6951;
	wire [4-1:0] node6952;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6962;
	wire [4-1:0] node6963;
	wire [4-1:0] node6967;
	wire [4-1:0] node6968;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6980;
	wire [4-1:0] node6981;
	wire [4-1:0] node6982;
	wire [4-1:0] node6983;
	wire [4-1:0] node6985;
	wire [4-1:0] node6988;
	wire [4-1:0] node6991;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node7002;
	wire [4-1:0] node7003;
	wire [4-1:0] node7005;
	wire [4-1:0] node7006;
	wire [4-1:0] node7010;
	wire [4-1:0] node7012;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7023;
	wire [4-1:0] node7025;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7032;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7040;
	wire [4-1:0] node7041;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7049;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7054;
	wire [4-1:0] node7058;
	wire [4-1:0] node7060;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7065;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7074;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7094;
	wire [4-1:0] node7095;
	wire [4-1:0] node7099;
	wire [4-1:0] node7100;
	wire [4-1:0] node7102;
	wire [4-1:0] node7103;
	wire [4-1:0] node7107;
	wire [4-1:0] node7109;
	wire [4-1:0] node7112;
	wire [4-1:0] node7113;
	wire [4-1:0] node7114;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7120;
	wire [4-1:0] node7124;
	wire [4-1:0] node7125;
	wire [4-1:0] node7126;
	wire [4-1:0] node7130;
	wire [4-1:0] node7132;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7138;
	wire [4-1:0] node7139;
	wire [4-1:0] node7143;
	wire [4-1:0] node7145;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7150;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7162;
	wire [4-1:0] node7163;
	wire [4-1:0] node7164;
	wire [4-1:0] node7166;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7177;
	wire [4-1:0] node7180;
	wire [4-1:0] node7182;
	wire [4-1:0] node7186;
	wire [4-1:0] node7187;
	wire [4-1:0] node7188;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7191;
	wire [4-1:0] node7192;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7198;
	wire [4-1:0] node7199;
	wire [4-1:0] node7200;
	wire [4-1:0] node7204;
	wire [4-1:0] node7206;
	wire [4-1:0] node7209;
	wire [4-1:0] node7210;
	wire [4-1:0] node7212;
	wire [4-1:0] node7215;
	wire [4-1:0] node7216;
	wire [4-1:0] node7217;
	wire [4-1:0] node7221;
	wire [4-1:0] node7222;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7230;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7236;
	wire [4-1:0] node7237;
	wire [4-1:0] node7241;
	wire [4-1:0] node7243;
	wire [4-1:0] node7246;
	wire [4-1:0] node7248;
	wire [4-1:0] node7250;
	wire [4-1:0] node7253;
	wire [4-1:0] node7254;
	wire [4-1:0] node7255;
	wire [4-1:0] node7256;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7263;
	wire [4-1:0] node7266;
	wire [4-1:0] node7267;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7278;
	wire [4-1:0] node7279;
	wire [4-1:0] node7283;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7291;
	wire [4-1:0] node7292;
	wire [4-1:0] node7293;
	wire [4-1:0] node7295;
	wire [4-1:0] node7298;
	wire [4-1:0] node7301;
	wire [4-1:0] node7302;
	wire [4-1:0] node7304;
	wire [4-1:0] node7307;
	wire [4-1:0] node7308;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7315;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7321;
	wire [4-1:0] node7325;
	wire [4-1:0] node7326;
	wire [4-1:0] node7327;
	wire [4-1:0] node7329;
	wire [4-1:0] node7331;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7337;
	wire [4-1:0] node7339;
	wire [4-1:0] node7342;
	wire [4-1:0] node7345;
	wire [4-1:0] node7347;
	wire [4-1:0] node7348;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7360;
	wire [4-1:0] node7362;
	wire [4-1:0] node7365;
	wire [4-1:0] node7366;
	wire [4-1:0] node7370;
	wire [4-1:0] node7371;
	wire [4-1:0] node7373;
	wire [4-1:0] node7376;
	wire [4-1:0] node7377;
	wire [4-1:0] node7379;
	wire [4-1:0] node7382;
	wire [4-1:0] node7384;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7389;
	wire [4-1:0] node7390;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7396;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7402;
	wire [4-1:0] node7404;
	wire [4-1:0] node7407;
	wire [4-1:0] node7409;
	wire [4-1:0] node7410;
	wire [4-1:0] node7412;
	wire [4-1:0] node7416;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7422;
	wire [4-1:0] node7423;
	wire [4-1:0] node7424;
	wire [4-1:0] node7428;
	wire [4-1:0] node7429;
	wire [4-1:0] node7433;
	wire [4-1:0] node7434;
	wire [4-1:0] node7435;
	wire [4-1:0] node7436;
	wire [4-1:0] node7438;
	wire [4-1:0] node7439;
	wire [4-1:0] node7443;
	wire [4-1:0] node7444;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7450;
	wire [4-1:0] node7451;
	wire [4-1:0] node7455;
	wire [4-1:0] node7457;
	wire [4-1:0] node7460;
	wire [4-1:0] node7461;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7468;
	wire [4-1:0] node7469;
	wire [4-1:0] node7473;
	wire [4-1:0] node7474;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7481;
	wire [4-1:0] node7482;
	wire [4-1:0] node7483;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7495;
	wire [4-1:0] node7497;
	wire [4-1:0] node7498;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7505;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7512;
	wire [4-1:0] node7515;
	wire [4-1:0] node7516;
	wire [4-1:0] node7517;
	wire [4-1:0] node7520;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7527;
	wire [4-1:0] node7529;
	wire [4-1:0] node7531;
	wire [4-1:0] node7533;
	wire [4-1:0] node7536;
	wire [4-1:0] node7537;
	wire [4-1:0] node7538;
	wire [4-1:0] node7540;
	wire [4-1:0] node7543;
	wire [4-1:0] node7544;
	wire [4-1:0] node7545;
	wire [4-1:0] node7549;
	wire [4-1:0] node7552;
	wire [4-1:0] node7553;
	wire [4-1:0] node7554;
	wire [4-1:0] node7555;
	wire [4-1:0] node7559;
	wire [4-1:0] node7561;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7567;
	wire [4-1:0] node7570;
	wire [4-1:0] node7572;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7582;
	wire [4-1:0] node7585;
	wire [4-1:0] node7586;
	wire [4-1:0] node7590;
	wire [4-1:0] node7591;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7605;
	wire [4-1:0] node7607;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7615;
	wire [4-1:0] node7617;
	wire [4-1:0] node7620;
	wire [4-1:0] node7622;
	wire [4-1:0] node7624;
	wire [4-1:0] node7626;
	wire [4-1:0] node7629;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7633;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7639;
	wire [4-1:0] node7642;
	wire [4-1:0] node7644;
	wire [4-1:0] node7647;
	wire [4-1:0] node7648;
	wire [4-1:0] node7649;
	wire [4-1:0] node7651;
	wire [4-1:0] node7654;
	wire [4-1:0] node7656;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7664;
	wire [4-1:0] node7665;
	wire [4-1:0] node7666;
	wire [4-1:0] node7667;
	wire [4-1:0] node7668;
	wire [4-1:0] node7669;
	wire [4-1:0] node7671;
	wire [4-1:0] node7674;
	wire [4-1:0] node7675;
	wire [4-1:0] node7679;
	wire [4-1:0] node7681;
	wire [4-1:0] node7684;
	wire [4-1:0] node7685;
	wire [4-1:0] node7687;
	wire [4-1:0] node7689;
	wire [4-1:0] node7693;
	wire [4-1:0] node7694;
	wire [4-1:0] node7695;
	wire [4-1:0] node7696;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7710;
	wire [4-1:0] node7711;
	wire [4-1:0] node7712;
	wire [4-1:0] node7713;
	wire [4-1:0] node7714;
	wire [4-1:0] node7716;
	wire [4-1:0] node7720;
	wire [4-1:0] node7721;
	wire [4-1:0] node7725;
	wire [4-1:0] node7726;
	wire [4-1:0] node7727;
	wire [4-1:0] node7728;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7742;
	wire [4-1:0] node7743;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7750;
	wire [4-1:0] node7752;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7760;
	wire [4-1:0] node7761;
	wire [4-1:0] node7762;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7774;
	wire [4-1:0] node7775;
	wire [4-1:0] node7778;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7783;
	wire [4-1:0] node7787;
	wire [4-1:0] node7788;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7795;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7800;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7810;
	wire [4-1:0] node7811;
	wire [4-1:0] node7815;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7819;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7826;
	wire [4-1:0] node7827;
	wire [4-1:0] node7828;
	wire [4-1:0] node7831;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7841;
	wire [4-1:0] node7842;
	wire [4-1:0] node7843;
	wire [4-1:0] node7844;
	wire [4-1:0] node7848;
	wire [4-1:0] node7850;
	wire [4-1:0] node7853;
	wire [4-1:0] node7854;
	wire [4-1:0] node7858;
	wire [4-1:0] node7859;
	wire [4-1:0] node7860;
	wire [4-1:0] node7861;
	wire [4-1:0] node7862;
	wire [4-1:0] node7863;
	wire [4-1:0] node7866;
	wire [4-1:0] node7867;
	wire [4-1:0] node7871;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7876;
	wire [4-1:0] node7879;
	wire [4-1:0] node7881;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7889;
	wire [4-1:0] node7890;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7899;
	wire [4-1:0] node7902;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7912;
	wire [4-1:0] node7913;
	wire [4-1:0] node7916;
	wire [4-1:0] node7919;
	wire [4-1:0] node7920;
	wire [4-1:0] node7923;
	wire [4-1:0] node7926;
	wire [4-1:0] node7927;
	wire [4-1:0] node7928;
	wire [4-1:0] node7931;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7938;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7945;
	wire [4-1:0] node7948;
	wire [4-1:0] node7951;
	wire [4-1:0] node7952;
	wire [4-1:0] node7953;
	wire [4-1:0] node7956;
	wire [4-1:0] node7959;
	wire [4-1:0] node7961;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7967;
	wire [4-1:0] node7969;
	wire [4-1:0] node7972;
	wire [4-1:0] node7975;
	wire [4-1:0] node7976;
	wire [4-1:0] node7977;
	wire [4-1:0] node7980;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7987;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7992;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7997;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8004;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8009;
	wire [4-1:0] node8012;
	wire [4-1:0] node8015;
	wire [4-1:0] node8016;
	wire [4-1:0] node8019;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8026;
	wire [4-1:0] node8029;
	wire [4-1:0] node8031;
	wire [4-1:0] node8034;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8039;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8050;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8055;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8067;
	wire [4-1:0] node8070;
	wire [4-1:0] node8071;
	wire [4-1:0] node8072;
	wire [4-1:0] node8074;
	wire [4-1:0] node8077;
	wire [4-1:0] node8079;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8087;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8092;
	wire [4-1:0] node8093;
	wire [4-1:0] node8094;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8104;
	wire [4-1:0] node8106;
	wire [4-1:0] node8109;
	wire [4-1:0] node8110;
	wire [4-1:0] node8113;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8123;
	wire [4-1:0] node8124;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8129;
	wire [4-1:0] node8132;
	wire [4-1:0] node8133;
	wire [4-1:0] node8136;
	wire [4-1:0] node8139;
	wire [4-1:0] node8140;
	wire [4-1:0] node8143;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8154;
	wire [4-1:0] node8155;
	wire [4-1:0] node8158;
	wire [4-1:0] node8161;
	wire [4-1:0] node8162;
	wire [4-1:0] node8164;
	wire [4-1:0] node8167;
	wire [4-1:0] node8170;
	wire [4-1:0] node8172;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8177;
	wire [4-1:0] node8178;
	wire [4-1:0] node8179;
	wire [4-1:0] node8181;
	wire [4-1:0] node8184;
	wire [4-1:0] node8185;
	wire [4-1:0] node8187;
	wire [4-1:0] node8191;
	wire [4-1:0] node8192;
	wire [4-1:0] node8193;
	wire [4-1:0] node8196;
	wire [4-1:0] node8198;
	wire [4-1:0] node8201;
	wire [4-1:0] node8202;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8213;
	wire [4-1:0] node8214;
	wire [4-1:0] node8217;
	wire [4-1:0] node8218;
	wire [4-1:0] node8222;
	wire [4-1:0] node8223;
	wire [4-1:0] node8224;
	wire [4-1:0] node8226;
	wire [4-1:0] node8229;
	wire [4-1:0] node8231;
	wire [4-1:0] node8234;
	wire [4-1:0] node8236;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8243;
	wire [4-1:0] node8244;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8253;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8257;
	wire [4-1:0] node8260;
	wire [4-1:0] node8263;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8268;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8275;
	wire [4-1:0] node8276;
	wire [4-1:0] node8277;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8282;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8290;
	wire [4-1:0] node8291;
	wire [4-1:0] node8293;
	wire [4-1:0] node8295;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8302;
	wire [4-1:0] node8305;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8310;
	wire [4-1:0] node8313;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8318;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8325;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8332;
	wire [4-1:0] node8333;
	wire [4-1:0] node8337;
	wire [4-1:0] node8339;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8346;
	wire [4-1:0] node8349;
	wire [4-1:0] node8350;
	wire [4-1:0] node8354;
	wire [4-1:0] node8355;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8361;
	wire [4-1:0] node8362;
	wire [4-1:0] node8363;
	wire [4-1:0] node8364;
	wire [4-1:0] node8367;
	wire [4-1:0] node8370;
	wire [4-1:0] node8371;
	wire [4-1:0] node8372;
	wire [4-1:0] node8375;
	wire [4-1:0] node8379;
	wire [4-1:0] node8380;
	wire [4-1:0] node8381;
	wire [4-1:0] node8384;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8394;
	wire [4-1:0] node8395;
	wire [4-1:0] node8396;
	wire [4-1:0] node8397;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8405;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8416;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8421;
	wire [4-1:0] node8422;
	wire [4-1:0] node8423;
	wire [4-1:0] node8427;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8432;
	wire [4-1:0] node8435;
	wire [4-1:0] node8438;
	wire [4-1:0] node8439;
	wire [4-1:0] node8442;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8447;
	wire [4-1:0] node8448;
	wire [4-1:0] node8451;
	wire [4-1:0] node8454;
	wire [4-1:0] node8455;
	wire [4-1:0] node8456;
	wire [4-1:0] node8460;
	wire [4-1:0] node8461;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8471;
	wire [4-1:0] node8474;
	wire [4-1:0] node8475;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8483;
	wire [4-1:0] node8486;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8494;
	wire [4-1:0] node8496;
	wire [4-1:0] node8499;
	wire [4-1:0] node8500;
	wire [4-1:0] node8503;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8509;
	wire [4-1:0] node8512;
	wire [4-1:0] node8513;
	wire [4-1:0] node8516;
	wire [4-1:0] node8517;
	wire [4-1:0] node8521;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8524;
	wire [4-1:0] node8525;
	wire [4-1:0] node8527;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8539;
	wire [4-1:0] node8542;
	wire [4-1:0] node8543;
	wire [4-1:0] node8545;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8555;
	wire [4-1:0] node8557;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8565;
	wire [4-1:0] node8566;
	wire [4-1:0] node8568;
	wire [4-1:0] node8571;
	wire [4-1:0] node8572;
	wire [4-1:0] node8576;
	wire [4-1:0] node8577;
	wire [4-1:0] node8578;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8583;
	wire [4-1:0] node8586;
	wire [4-1:0] node8587;
	wire [4-1:0] node8591;
	wire [4-1:0] node8592;
	wire [4-1:0] node8594;
	wire [4-1:0] node8597;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8603;
	wire [4-1:0] node8605;
	wire [4-1:0] node8607;
	wire [4-1:0] node8610;
	wire [4-1:0] node8611;
	wire [4-1:0] node8615;
	wire [4-1:0] node8616;
	wire [4-1:0] node8617;
	wire [4-1:0] node8618;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8623;
	wire [4-1:0] node8624;
	wire [4-1:0] node8628;
	wire [4-1:0] node8630;
	wire [4-1:0] node8633;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8641;
	wire [4-1:0] node8642;
	wire [4-1:0] node8647;
	wire [4-1:0] node8648;
	wire [4-1:0] node8649;
	wire [4-1:0] node8650;
	wire [4-1:0] node8651;
	wire [4-1:0] node8653;
	wire [4-1:0] node8656;
	wire [4-1:0] node8657;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8664;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8680;
	wire [4-1:0] node8681;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8690;
	wire [4-1:0] node8691;
	wire [4-1:0] node8693;
	wire [4-1:0] node8696;
	wire [4-1:0] node8697;
	wire [4-1:0] node8699;
	wire [4-1:0] node8702;
	wire [4-1:0] node8704;
	wire [4-1:0] node8707;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8713;
	wire [4-1:0] node8716;
	wire [4-1:0] node8718;
	wire [4-1:0] node8721;
	wire [4-1:0] node8723;
	wire [4-1:0] node8724;
	wire [4-1:0] node8726;
	wire [4-1:0] node8729;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8736;
	wire [4-1:0] node8737;
	wire [4-1:0] node8738;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8744;
	wire [4-1:0] node8746;
	wire [4-1:0] node8748;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8754;
	wire [4-1:0] node8757;
	wire [4-1:0] node8759;
	wire [4-1:0] node8761;
	wire [4-1:0] node8764;
	wire [4-1:0] node8765;
	wire [4-1:0] node8766;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8772;
	wire [4-1:0] node8776;
	wire [4-1:0] node8779;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8783;
	wire [4-1:0] node8786;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8792;
	wire [4-1:0] node8793;
	wire [4-1:0] node8797;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8811;
	wire [4-1:0] node8812;
	wire [4-1:0] node8813;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8819;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8828;
	wire [4-1:0] node8829;
	wire [4-1:0] node8831;
	wire [4-1:0] node8835;
	wire [4-1:0] node8837;
	wire [4-1:0] node8839;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8845;
	wire [4-1:0] node8848;
	wire [4-1:0] node8850;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8855;
	wire [4-1:0] node8856;
	wire [4-1:0] node8859;
	wire [4-1:0] node8861;
	wire [4-1:0] node8864;
	wire [4-1:0] node8866;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8872;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8880;
	wire [4-1:0] node8881;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8890;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8904;
	wire [4-1:0] node8907;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8919;
	wire [4-1:0] node8921;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8928;
	wire [4-1:0] node8931;
	wire [4-1:0] node8933;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8940;
	wire [4-1:0] node8942;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8950;
	wire [4-1:0] node8951;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8955;
	wire [4-1:0] node8956;
	wire [4-1:0] node8959;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8969;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8984;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8996;
	wire [4-1:0] node8998;
	wire [4-1:0] node9001;
	wire [4-1:0] node9002;
	wire [4-1:0] node9003;
	wire [4-1:0] node9006;
	wire [4-1:0] node9007;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9016;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9028;
	wire [4-1:0] node9029;
	wire [4-1:0] node9031;
	wire [4-1:0] node9034;
	wire [4-1:0] node9036;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9044;
	wire [4-1:0] node9046;
	wire [4-1:0] node9049;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9059;
	wire [4-1:0] node9062;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9069;
	wire [4-1:0] node9072;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9078;
	wire [4-1:0] node9079;
	wire [4-1:0] node9082;
	wire [4-1:0] node9085;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9091;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9100;
	wire [4-1:0] node9102;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9108;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9121;
	wire [4-1:0] node9124;
	wire [4-1:0] node9127;
	wire [4-1:0] node9128;
	wire [4-1:0] node9129;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9135;
	wire [4-1:0] node9136;
	wire [4-1:0] node9140;
	wire [4-1:0] node9141;
	wire [4-1:0] node9143;
	wire [4-1:0] node9148;
	wire [4-1:0] node9149;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9152;
	wire [4-1:0] node9153;
	wire [4-1:0] node9155;
	wire [4-1:0] node9158;
	wire [4-1:0] node9160;
	wire [4-1:0] node9163;
	wire [4-1:0] node9164;
	wire [4-1:0] node9168;
	wire [4-1:0] node9169;
	wire [4-1:0] node9170;
	wire [4-1:0] node9171;
	wire [4-1:0] node9172;
	wire [4-1:0] node9175;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9182;
	wire [4-1:0] node9185;
	wire [4-1:0] node9186;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9197;
	wire [4-1:0] node9200;
	wire [4-1:0] node9201;
	wire [4-1:0] node9204;
	wire [4-1:0] node9206;
	wire [4-1:0] node9209;
	wire [4-1:0] node9210;
	wire [4-1:0] node9211;
	wire [4-1:0] node9212;
	wire [4-1:0] node9213;
	wire [4-1:0] node9216;
	wire [4-1:0] node9220;
	wire [4-1:0] node9221;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9229;
	wire [4-1:0] node9230;
	wire [4-1:0] node9231;
	wire [4-1:0] node9232;
	wire [4-1:0] node9235;
	wire [4-1:0] node9236;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9247;
	wire [4-1:0] node9248;
	wire [4-1:0] node9249;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9260;
	wire [4-1:0] node9263;
	wire [4-1:0] node9264;
	wire [4-1:0] node9268;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9271;
	wire [4-1:0] node9272;
	wire [4-1:0] node9274;
	wire [4-1:0] node9277;
	wire [4-1:0] node9279;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9288;
	wire [4-1:0] node9290;
	wire [4-1:0] node9293;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9298;
	wire [4-1:0] node9302;
	wire [4-1:0] node9303;
	wire [4-1:0] node9307;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9318;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9325;
	wire [4-1:0] node9326;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9336;
	wire [4-1:0] node9339;
	wire [4-1:0] node9340;
	wire [4-1:0] node9342;
	wire [4-1:0] node9343;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9353;
	wire [4-1:0] node9354;
	wire [4-1:0] node9355;
	wire [4-1:0] node9356;
	wire [4-1:0] node9357;
	wire [4-1:0] node9358;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9362;
	wire [4-1:0] node9365;
	wire [4-1:0] node9368;
	wire [4-1:0] node9369;
	wire [4-1:0] node9371;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9379;
	wire [4-1:0] node9380;
	wire [4-1:0] node9385;
	wire [4-1:0] node9386;
	wire [4-1:0] node9389;
	wire [4-1:0] node9390;
	wire [4-1:0] node9393;
	wire [4-1:0] node9396;
	wire [4-1:0] node9397;
	wire [4-1:0] node9398;
	wire [4-1:0] node9399;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9415;
	wire [4-1:0] node9416;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9424;
	wire [4-1:0] node9427;
	wire [4-1:0] node9428;
	wire [4-1:0] node9429;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9437;
	wire [4-1:0] node9438;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9449;
	wire [4-1:0] node9450;
	wire [4-1:0] node9454;
	wire [4-1:0] node9455;
	wire [4-1:0] node9456;
	wire [4-1:0] node9459;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9466;
	wire [4-1:0] node9469;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9477;
	wire [4-1:0] node9478;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9486;
	wire [4-1:0] node9489;
	wire [4-1:0] node9491;
	wire [4-1:0] node9492;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9502;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9509;
	wire [4-1:0] node9510;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9518;
	wire [4-1:0] node9519;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9525;
	wire [4-1:0] node9527;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9534;
	wire [4-1:0] node9537;
	wire [4-1:0] node9538;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9552;
	wire [4-1:0] node9556;
	wire [4-1:0] node9557;
	wire [4-1:0] node9560;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9568;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9574;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9583;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9588;
	wire [4-1:0] node9591;
	wire [4-1:0] node9594;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9603;
	wire [4-1:0] node9604;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9610;
	wire [4-1:0] node9613;
	wire [4-1:0] node9614;
	wire [4-1:0] node9617;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9623;
	wire [4-1:0] node9626;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9633;
	wire [4-1:0] node9635;
	wire [4-1:0] node9636;
	wire [4-1:0] node9639;
	wire [4-1:0] node9642;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9647;
	wire [4-1:0] node9650;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9664;
	wire [4-1:0] node9667;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9678;
	wire [4-1:0] node9682;
	wire [4-1:0] node9686;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9690;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9700;
	wire [4-1:0] node9702;
	wire [4-1:0] node9704;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9709;
	wire [4-1:0] node9711;
	wire [4-1:0] node9712;
	wire [4-1:0] node9713;
	wire [4-1:0] node9714;
	wire [4-1:0] node9717;
	wire [4-1:0] node9720;
	wire [4-1:0] node9721;
	wire [4-1:0] node9724;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9732;
	wire [4-1:0] node9733;
	wire [4-1:0] node9734;
	wire [4-1:0] node9736;
	wire [4-1:0] node9739;
	wire [4-1:0] node9740;
	wire [4-1:0] node9743;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9751;
	wire [4-1:0] node9754;
	wire [4-1:0] node9756;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9770;
	wire [4-1:0] node9774;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9777;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9786;
	wire [4-1:0] node9789;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9795;
	wire [4-1:0] node9798;
	wire [4-1:0] node9801;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9807;
	wire [4-1:0] node9810;
	wire [4-1:0] node9811;
	wire [4-1:0] node9814;
	wire [4-1:0] node9817;
	wire [4-1:0] node9819;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9824;
	wire [4-1:0] node9826;
	wire [4-1:0] node9827;
	wire [4-1:0] node9830;
	wire [4-1:0] node9833;
	wire [4-1:0] node9834;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9841;
	wire [4-1:0] node9844;
	wire [4-1:0] node9845;
	wire [4-1:0] node9846;
	wire [4-1:0] node9847;
	wire [4-1:0] node9851;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9858;
	wire [4-1:0] node9859;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9868;
	wire [4-1:0] node9872;
	wire [4-1:0] node9875;
	wire [4-1:0] node9876;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9883;
	wire [4-1:0] node9886;
	wire [4-1:0] node9887;
	wire [4-1:0] node9888;
	wire [4-1:0] node9891;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9897;
	wire [4-1:0] node9900;
	wire [4-1:0] node9901;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9910;
	wire [4-1:0] node9913;
	wire [4-1:0] node9914;
	wire [4-1:0] node9918;
	wire [4-1:0] node9919;
	wire [4-1:0] node9920;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9928;
	wire [4-1:0] node9931;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9935;
	wire [4-1:0] node9938;
	wire [4-1:0] node9940;
	wire [4-1:0] node9943;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9953;
	wire [4-1:0] node9954;
	wire [4-1:0] node9955;
	wire [4-1:0] node9959;
	wire [4-1:0] node9960;
	wire [4-1:0] node9963;
	wire [4-1:0] node9966;
	wire [4-1:0] node9967;
	wire [4-1:0] node9969;
	wire [4-1:0] node9972;
	wire [4-1:0] node9973;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9980;
	wire [4-1:0] node9983;
	wire [4-1:0] node9984;
	wire [4-1:0] node9985;
	wire [4-1:0] node9989;
	wire [4-1:0] node9990;
	wire [4-1:0] node9994;
	wire [4-1:0] node9995;
	wire [4-1:0] node9996;
	wire [4-1:0] node9998;
	wire [4-1:0] node10001;
	wire [4-1:0] node10002;
	wire [4-1:0] node10004;
	wire [4-1:0] node10007;
	wire [4-1:0] node10009;
	wire [4-1:0] node10012;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10018;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10025;
	wire [4-1:0] node10028;
	wire [4-1:0] node10029;
	wire [4-1:0] node10031;
	wire [4-1:0] node10034;
	wire [4-1:0] node10035;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10043;
	wire [4-1:0] node10044;
	wire [4-1:0] node10045;
	wire [4-1:0] node10046;
	wire [4-1:0] node10047;
	wire [4-1:0] node10050;
	wire [4-1:0] node10051;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10058;
	wire [4-1:0] node10061;
	wire [4-1:0] node10062;
	wire [4-1:0] node10066;
	wire [4-1:0] node10067;
	wire [4-1:0] node10070;
	wire [4-1:0] node10072;
	wire [4-1:0] node10074;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10080;
	wire [4-1:0] node10084;
	wire [4-1:0] node10085;
	wire [4-1:0] node10086;
	wire [4-1:0] node10090;
	wire [4-1:0] node10093;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10096;
	wire [4-1:0] node10100;
	wire [4-1:0] node10102;
	wire [4-1:0] node10105;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10113;
	wire [4-1:0] node10118;
	wire [4-1:0] node10121;
	wire [4-1:0] node10122;
	wire [4-1:0] node10124;
	wire [4-1:0] node10125;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10132;
	wire [4-1:0] node10134;
	wire [4-1:0] node10137;
	wire [4-1:0] node10139;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10145;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10152;
	wire [4-1:0] node10155;
	wire [4-1:0] node10157;
	wire [4-1:0] node10160;
	wire [4-1:0] node10161;
	wire [4-1:0] node10163;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10169;
	wire [4-1:0] node10171;
	wire [4-1:0] node10175;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10183;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10191;
	wire [4-1:0] node10192;
	wire [4-1:0] node10195;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10204;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10209;
	wire [4-1:0] node10212;
	wire [4-1:0] node10213;
	wire [4-1:0] node10216;
	wire [4-1:0] node10219;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10222;
	wire [4-1:0] node10224;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10236;
	wire [4-1:0] node10238;
	wire [4-1:0] node10242;
	wire [4-1:0] node10243;
	wire [4-1:0] node10244;
	wire [4-1:0] node10245;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10253;
	wire [4-1:0] node10254;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10264;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10268;
	wire [4-1:0] node10271;
	wire [4-1:0] node10272;
	wire [4-1:0] node10275;
	wire [4-1:0] node10278;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10284;
	wire [4-1:0] node10285;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10291;
	wire [4-1:0] node10292;
	wire [4-1:0] node10294;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10307;
	wire [4-1:0] node10308;
	wire [4-1:0] node10309;
	wire [4-1:0] node10313;
	wire [4-1:0] node10314;
	wire [4-1:0] node10317;
	wire [4-1:0] node10320;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10323;
	wire [4-1:0] node10324;
	wire [4-1:0] node10328;
	wire [4-1:0] node10329;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10339;
	wire [4-1:0] node10341;
	wire [4-1:0] node10342;
	wire [4-1:0] node10346;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10349;
	wire [4-1:0] node10350;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10360;
	wire [4-1:0] node10363;
	wire [4-1:0] node10365;
	wire [4-1:0] node10368;
	wire [4-1:0] node10369;
	wire [4-1:0] node10370;
	wire [4-1:0] node10371;
	wire [4-1:0] node10375;
	wire [4-1:0] node10377;
	wire [4-1:0] node10380;
	wire [4-1:0] node10381;
	wire [4-1:0] node10385;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10389;
	wire [4-1:0] node10390;
	wire [4-1:0] node10392;
	wire [4-1:0] node10395;
	wire [4-1:0] node10397;
	wire [4-1:0] node10400;
	wire [4-1:0] node10401;
	wire [4-1:0] node10403;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10410;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10415;
	wire [4-1:0] node10416;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10431;
	wire [4-1:0] node10434;
	wire [4-1:0] node10435;
	wire [4-1:0] node10436;
	wire [4-1:0] node10437;
	wire [4-1:0] node10438;
	wire [4-1:0] node10441;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10448;
	wire [4-1:0] node10451;
	wire [4-1:0] node10452;
	wire [4-1:0] node10453;
	wire [4-1:0] node10456;
	wire [4-1:0] node10459;
	wire [4-1:0] node10460;
	wire [4-1:0] node10463;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10468;
	wire [4-1:0] node10470;
	wire [4-1:0] node10473;
	wire [4-1:0] node10475;
	wire [4-1:0] node10478;
	wire [4-1:0] node10479;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10486;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10491;
	wire [4-1:0] node10492;
	wire [4-1:0] node10494;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10502;
	wire [4-1:0] node10503;
	wire [4-1:0] node10504;
	wire [4-1:0] node10508;
	wire [4-1:0] node10509;
	wire [4-1:0] node10510;
	wire [4-1:0] node10513;
	wire [4-1:0] node10516;
	wire [4-1:0] node10518;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10524;
	wire [4-1:0] node10525;
	wire [4-1:0] node10526;
	wire [4-1:0] node10527;
	wire [4-1:0] node10529;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10535;
	wire [4-1:0] node10538;
	wire [4-1:0] node10540;
	wire [4-1:0] node10543;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10547;
	wire [4-1:0] node10550;
	wire [4-1:0] node10552;
	wire [4-1:0] node10555;
	wire [4-1:0] node10556;
	wire [4-1:0] node10558;
	wire [4-1:0] node10561;
	wire [4-1:0] node10563;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10570;
	wire [4-1:0] node10571;
	wire [4-1:0] node10574;
	wire [4-1:0] node10577;
	wire [4-1:0] node10578;
	wire [4-1:0] node10579;
	wire [4-1:0] node10582;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10592;
	wire [4-1:0] node10596;
	wire [4-1:0] node10597;
	wire [4-1:0] node10599;
	wire [4-1:0] node10602;
	wire [4-1:0] node10604;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10611;
	wire [4-1:0] node10612;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10620;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10630;
	wire [4-1:0] node10631;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10639;
	wire [4-1:0] node10642;
	wire [4-1:0] node10644;
	wire [4-1:0] node10648;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10651;
	wire [4-1:0] node10652;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10659;
	wire [4-1:0] node10660;
	wire [4-1:0] node10661;
	wire [4-1:0] node10664;
	wire [4-1:0] node10668;
	wire [4-1:0] node10670;
	wire [4-1:0] node10672;
	wire [4-1:0] node10673;
	wire [4-1:0] node10676;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10683;
	wire [4-1:0] node10684;
	wire [4-1:0] node10685;
	wire [4-1:0] node10687;
	wire [4-1:0] node10688;
	wire [4-1:0] node10690;
	wire [4-1:0] node10691;
	wire [4-1:0] node10692;
	wire [4-1:0] node10694;
	wire [4-1:0] node10696;
	wire [4-1:0] node10699;
	wire [4-1:0] node10701;
	wire [4-1:0] node10702;
	wire [4-1:0] node10703;
	wire [4-1:0] node10709;
	wire [4-1:0] node10710;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10716;
	wire [4-1:0] node10720;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10726;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10734;
	wire [4-1:0] node10737;
	wire [4-1:0] node10739;
	wire [4-1:0] node10742;
	wire [4-1:0] node10743;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10746;
	wire [4-1:0] node10750;
	wire [4-1:0] node10753;
	wire [4-1:0] node10754;
	wire [4-1:0] node10756;
	wire [4-1:0] node10759;
	wire [4-1:0] node10761;
	wire [4-1:0] node10764;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10770;
	wire [4-1:0] node10771;
	wire [4-1:0] node10775;
	wire [4-1:0] node10777;
	wire [4-1:0] node10778;
	wire [4-1:0] node10779;
	wire [4-1:0] node10780;
	wire [4-1:0] node10783;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10790;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10800;
	wire [4-1:0] node10801;
	wire [4-1:0] node10802;
	wire [4-1:0] node10803;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10807;
	wire [4-1:0] node10811;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10817;
	wire [4-1:0] node10820;
	wire [4-1:0] node10821;
	wire [4-1:0] node10822;
	wire [4-1:0] node10827;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10831;
	wire [4-1:0] node10832;
	wire [4-1:0] node10836;
	wire [4-1:0] node10837;
	wire [4-1:0] node10838;
	wire [4-1:0] node10842;
	wire [4-1:0] node10844;
	wire [4-1:0] node10847;
	wire [4-1:0] node10848;
	wire [4-1:0] node10850;
	wire [4-1:0] node10853;
	wire [4-1:0] node10855;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10861;
	wire [4-1:0] node10863;
	wire [4-1:0] node10866;
	wire [4-1:0] node10867;
	wire [4-1:0] node10871;
	wire [4-1:0] node10872;
	wire [4-1:0] node10873;
	wire [4-1:0] node10875;
	wire [4-1:0] node10878;
	wire [4-1:0] node10880;
	wire [4-1:0] node10883;
	wire [4-1:0] node10884;
	wire [4-1:0] node10886;
	wire [4-1:0] node10889;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10897;
	wire [4-1:0] node10900;
	wire [4-1:0] node10902;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10908;
	wire [4-1:0] node10911;
	wire [4-1:0] node10913;
	wire [4-1:0] node10916;
	wire [4-1:0] node10917;
	wire [4-1:0] node10918;
	wire [4-1:0] node10922;
	wire [4-1:0] node10923;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10930;
	wire [4-1:0] node10931;
	wire [4-1:0] node10932;
	wire [4-1:0] node10936;
	wire [4-1:0] node10938;
	wire [4-1:0] node10941;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10947;
	wire [4-1:0] node10949;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10954;
	wire [4-1:0] node10958;
	wire [4-1:0] node10960;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10966;
	wire [4-1:0] node10970;
	wire [4-1:0] node10972;
	wire [4-1:0] node10975;
	wire [4-1:0] node10976;
	wire [4-1:0] node10977;
	wire [4-1:0] node10978;
	wire [4-1:0] node10982;
	wire [4-1:0] node10983;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10990;
	wire [4-1:0] node10993;
	wire [4-1:0] node10995;
	wire [4-1:0] node10998;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11003;
	wire [4-1:0] node11004;
	wire [4-1:0] node11008;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11015;
	wire [4-1:0] node11019;
	wire [4-1:0] node11020;
	wire [4-1:0] node11021;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11032;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11047;
	wire [4-1:0] node11048;
	wire [4-1:0] node11049;
	wire [4-1:0] node11050;
	wire [4-1:0] node11051;
	wire [4-1:0] node11056;
	wire [4-1:0] node11057;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11063;
	wire [4-1:0] node11064;
	wire [4-1:0] node11067;
	wire [4-1:0] node11069;
	wire [4-1:0] node11072;
	wire [4-1:0] node11073;
	wire [4-1:0] node11077;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11086;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11093;
	wire [4-1:0] node11094;
	wire [4-1:0] node11095;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11113;
	wire [4-1:0] node11116;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11121;
	wire [4-1:0] node11122;
	wire [4-1:0] node11123;
	wire [4-1:0] node11127;
	wire [4-1:0] node11128;
	wire [4-1:0] node11132;
	wire [4-1:0] node11133;
	wire [4-1:0] node11134;
	wire [4-1:0] node11138;
	wire [4-1:0] node11141;
	wire [4-1:0] node11142;
	wire [4-1:0] node11143;
	wire [4-1:0] node11147;
	wire [4-1:0] node11149;
	wire [4-1:0] node11152;
	wire [4-1:0] node11153;
	wire [4-1:0] node11154;
	wire [4-1:0] node11155;
	wire [4-1:0] node11159;
	wire [4-1:0] node11161;
	wire [4-1:0] node11164;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11168;
	wire [4-1:0] node11171;
	wire [4-1:0] node11172;
	wire [4-1:0] node11176;
	wire [4-1:0] node11177;
	wire [4-1:0] node11179;
	wire [4-1:0] node11182;
	wire [4-1:0] node11184;
	wire [4-1:0] node11187;
	wire [4-1:0] node11189;
	wire [4-1:0] node11191;
	wire [4-1:0] node11192;
	wire [4-1:0] node11193;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11209;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11216;
	wire [4-1:0] node11217;
	wire [4-1:0] node11218;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11224;
	wire [4-1:0] node11226;
	wire [4-1:0] node11229;
	wire [4-1:0] node11230;
	wire [4-1:0] node11231;
	wire [4-1:0] node11233;
	wire [4-1:0] node11236;
	wire [4-1:0] node11238;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11246;
	wire [4-1:0] node11247;
	wire [4-1:0] node11248;
	wire [4-1:0] node11249;
	wire [4-1:0] node11252;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11258;
	wire [4-1:0] node11262;
	wire [4-1:0] node11263;
	wire [4-1:0] node11264;
	wire [4-1:0] node11268;
	wire [4-1:0] node11269;
	wire [4-1:0] node11273;
	wire [4-1:0] node11275;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11279;
	wire [4-1:0] node11280;
	wire [4-1:0] node11282;
	wire [4-1:0] node11286;
	wire [4-1:0] node11287;
	wire [4-1:0] node11291;
	wire [4-1:0] node11293;
	wire [4-1:0] node11294;
	wire [4-1:0] node11295;
	wire [4-1:0] node11299;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11307;
	wire [4-1:0] node11308;
	wire [4-1:0] node11309;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11313;
	wire [4-1:0] node11316;
	wire [4-1:0] node11317;
	wire [4-1:0] node11318;
	wire [4-1:0] node11322;
	wire [4-1:0] node11325;
	wire [4-1:0] node11327;
	wire [4-1:0] node11330;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11333;
	wire [4-1:0] node11334;
	wire [4-1:0] node11335;
	wire [4-1:0] node11339;
	wire [4-1:0] node11341;
	wire [4-1:0] node11344;
	wire [4-1:0] node11345;
	wire [4-1:0] node11348;
	wire [4-1:0] node11349;
	wire [4-1:0] node11353;
	wire [4-1:0] node11354;
	wire [4-1:0] node11355;
	wire [4-1:0] node11357;
	wire [4-1:0] node11360;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11367;
	wire [4-1:0] node11368;
	wire [4-1:0] node11372;
	wire [4-1:0] node11373;
	wire [4-1:0] node11374;
	wire [4-1:0] node11376;
	wire [4-1:0] node11379;
	wire [4-1:0] node11380;
	wire [4-1:0] node11383;
	wire [4-1:0] node11384;
	wire [4-1:0] node11388;
	wire [4-1:0] node11390;
	wire [4-1:0] node11393;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11400;
	wire [4-1:0] node11401;
	wire [4-1:0] node11402;
	wire [4-1:0] node11405;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11418;
	wire [4-1:0] node11421;
	wire [4-1:0] node11424;
	wire [4-1:0] node11427;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11436;
	wire [4-1:0] node11439;
	wire [4-1:0] node11441;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11448;
	wire [4-1:0] node11450;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11455;
	wire [4-1:0] node11456;
	wire [4-1:0] node11457;
	wire [4-1:0] node11458;
	wire [4-1:0] node11461;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11470;
	wire [4-1:0] node11473;
	wire [4-1:0] node11475;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11480;
	wire [4-1:0] node11482;
	wire [4-1:0] node11485;
	wire [4-1:0] node11488;
	wire [4-1:0] node11489;
	wire [4-1:0] node11490;
	wire [4-1:0] node11493;
	wire [4-1:0] node11496;
	wire [4-1:0] node11497;
	wire [4-1:0] node11500;
	wire [4-1:0] node11503;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11507;
	wire [4-1:0] node11508;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11516;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11525;
	wire [4-1:0] node11528;
	wire [4-1:0] node11529;
	wire [4-1:0] node11532;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11538;
	wire [4-1:0] node11541;
	wire [4-1:0] node11543;
	wire [4-1:0] node11546;
	wire [4-1:0] node11547;
	wire [4-1:0] node11548;
	wire [4-1:0] node11549;
	wire [4-1:0] node11550;
	wire [4-1:0] node11552;
	wire [4-1:0] node11553;
	wire [4-1:0] node11555;
	wire [4-1:0] node11559;
	wire [4-1:0] node11560;
	wire [4-1:0] node11564;
	wire [4-1:0] node11565;
	wire [4-1:0] node11566;
	wire [4-1:0] node11568;
	wire [4-1:0] node11571;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11576;
	wire [4-1:0] node11579;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11585;
	wire [4-1:0] node11586;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11594;
	wire [4-1:0] node11595;
	wire [4-1:0] node11599;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11607;
	wire [4-1:0] node11610;
	wire [4-1:0] node11611;
	wire [4-1:0] node11614;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11621;
	wire [4-1:0] node11622;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11632;
	wire [4-1:0] node11635;
	wire [4-1:0] node11638;
	wire [4-1:0] node11639;
	wire [4-1:0] node11642;
	wire [4-1:0] node11645;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11648;
	wire [4-1:0] node11652;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11661;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11670;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11679;
	wire [4-1:0] node11680;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11686;
	wire [4-1:0] node11687;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11696;
	wire [4-1:0] node11697;
	wire [4-1:0] node11699;
	wire [4-1:0] node11702;
	wire [4-1:0] node11704;
	wire [4-1:0] node11707;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11711;
	wire [4-1:0] node11712;
	wire [4-1:0] node11716;
	wire [4-1:0] node11717;
	wire [4-1:0] node11718;
	wire [4-1:0] node11721;
	wire [4-1:0] node11724;
	wire [4-1:0] node11727;
	wire [4-1:0] node11728;
	wire [4-1:0] node11730;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11740;
	wire [4-1:0] node11741;
	wire [4-1:0] node11742;
	wire [4-1:0] node11745;
	wire [4-1:0] node11746;
	wire [4-1:0] node11749;
	wire [4-1:0] node11752;
	wire [4-1:0] node11753;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11765;
	wire [4-1:0] node11768;
	wire [4-1:0] node11771;
	wire [4-1:0] node11772;
	wire [4-1:0] node11774;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11781;
	wire [4-1:0] node11784;
	wire [4-1:0] node11785;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11790;
	wire [4-1:0] node11793;
	wire [4-1:0] node11794;
	wire [4-1:0] node11798;
	wire [4-1:0] node11799;
	wire [4-1:0] node11801;
	wire [4-1:0] node11803;
	wire [4-1:0] node11806;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11812;
	wire [4-1:0] node11813;
	wire [4-1:0] node11816;
	wire [4-1:0] node11819;
	wire [4-1:0] node11820;
	wire [4-1:0] node11821;
	wire [4-1:0] node11822;
	wire [4-1:0] node11823;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11830;
	wire [4-1:0] node11833;
	wire [4-1:0] node11834;
	wire [4-1:0] node11835;
	wire [4-1:0] node11839;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11848;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11855;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11861;
	wire [4-1:0] node11865;
	wire [4-1:0] node11868;
	wire [4-1:0] node11869;
	wire [4-1:0] node11872;
	wire [4-1:0] node11875;
	wire [4-1:0] node11876;
	wire [4-1:0] node11877;
	wire [4-1:0] node11878;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11886;
	wire [4-1:0] node11887;
	wire [4-1:0] node11888;
	wire [4-1:0] node11891;
	wire [4-1:0] node11894;
	wire [4-1:0] node11895;
	wire [4-1:0] node11898;
	wire [4-1:0] node11901;
	wire [4-1:0] node11902;
	wire [4-1:0] node11903;
	wire [4-1:0] node11905;
	wire [4-1:0] node11908;
	wire [4-1:0] node11910;
	wire [4-1:0] node11913;
	wire [4-1:0] node11914;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11921;
	wire [4-1:0] node11922;
	wire [4-1:0] node11923;
	wire [4-1:0] node11927;
	wire [4-1:0] node11930;
	wire [4-1:0] node11931;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11936;
	wire [4-1:0] node11940;
	wire [4-1:0] node11943;
	wire [4-1:0] node11944;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11953;
	wire [4-1:0] node11954;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11958;
	wire [4-1:0] node11962;
	wire [4-1:0] node11963;
	wire [4-1:0] node11966;
	wire [4-1:0] node11967;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11974;
	wire [4-1:0] node11977;
	wire [4-1:0] node11978;
	wire [4-1:0] node11981;
	wire [4-1:0] node11984;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11989;
	wire [4-1:0] node11994;
	wire [4-1:0] node11995;
	wire [4-1:0] node11998;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12003;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12014;
	wire [4-1:0] node12018;
	wire [4-1:0] node12019;
	wire [4-1:0] node12020;
	wire [4-1:0] node12024;
	wire [4-1:0] node12025;
	wire [4-1:0] node12027;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12034;
	wire [4-1:0] node12037;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12043;
	wire [4-1:0] node12045;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12052;
	wire [4-1:0] node12055;
	wire [4-1:0] node12056;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12063;
	wire [4-1:0] node12064;
	wire [4-1:0] node12068;
	wire [4-1:0] node12070;
	wire [4-1:0] node12071;
	wire [4-1:0] node12074;
	wire [4-1:0] node12077;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12081;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12088;
	wire [4-1:0] node12091;
	wire [4-1:0] node12092;
	wire [4-1:0] node12093;
	wire [4-1:0] node12096;
	wire [4-1:0] node12099;
	wire [4-1:0] node12101;
	wire [4-1:0] node12104;
	wire [4-1:0] node12105;
	wire [4-1:0] node12106;
	wire [4-1:0] node12107;
	wire [4-1:0] node12108;
	wire [4-1:0] node12110;
	wire [4-1:0] node12113;
	wire [4-1:0] node12115;
	wire [4-1:0] node12118;
	wire [4-1:0] node12119;
	wire [4-1:0] node12120;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12130;
	wire [4-1:0] node12132;
	wire [4-1:0] node12135;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12144;
	wire [4-1:0] node12145;
	wire [4-1:0] node12148;
	wire [4-1:0] node12151;
	wire [4-1:0] node12153;
	wire [4-1:0] node12156;
	wire [4-1:0] node12157;
	wire [4-1:0] node12158;
	wire [4-1:0] node12159;
	wire [4-1:0] node12163;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12173;
	wire [4-1:0] node12174;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12181;
	wire [4-1:0] node12182;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12187;
	wire [4-1:0] node12190;
	wire [4-1:0] node12193;
	wire [4-1:0] node12196;
	wire [4-1:0] node12197;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12207;
	wire [4-1:0] node12211;
	wire [4-1:0] node12212;
	wire [4-1:0] node12216;
	wire [4-1:0] node12217;
	wire [4-1:0] node12218;
	wire [4-1:0] node12219;
	wire [4-1:0] node12223;
	wire [4-1:0] node12226;
	wire [4-1:0] node12227;
	wire [4-1:0] node12231;
	wire [4-1:0] node12232;
	wire [4-1:0] node12233;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12238;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12246;
	wire [4-1:0] node12247;
	wire [4-1:0] node12249;
	wire [4-1:0] node12252;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12262;
	wire [4-1:0] node12265;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12273;
	wire [4-1:0] node12275;
	wire [4-1:0] node12278;
	wire [4-1:0] node12279;
	wire [4-1:0] node12281;
	wire [4-1:0] node12284;
	wire [4-1:0] node12286;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12295;
	wire [4-1:0] node12296;
	wire [4-1:0] node12297;
	wire [4-1:0] node12298;
	wire [4-1:0] node12302;
	wire [4-1:0] node12303;
	wire [4-1:0] node12304;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12313;
	wire [4-1:0] node12316;
	wire [4-1:0] node12317;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12328;
	wire [4-1:0] node12329;
	wire [4-1:0] node12333;
	wire [4-1:0] node12334;
	wire [4-1:0] node12336;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12343;
	wire [4-1:0] node12346;
	wire [4-1:0] node12347;
	wire [4-1:0] node12351;
	wire [4-1:0] node12352;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12356;
	wire [4-1:0] node12359;
	wire [4-1:0] node12361;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12369;
	wire [4-1:0] node12371;
	wire [4-1:0] node12374;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12380;
	wire [4-1:0] node12383;
	wire [4-1:0] node12384;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12387;
	wire [4-1:0] node12391;
	wire [4-1:0] node12392;
	wire [4-1:0] node12396;
	wire [4-1:0] node12397;
	wire [4-1:0] node12400;
	wire [4-1:0] node12401;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12410;
	wire [4-1:0] node12413;
	wire [4-1:0] node12416;
	wire [4-1:0] node12417;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12421;
	wire [4-1:0] node12422;
	wire [4-1:0] node12423;
	wire [4-1:0] node12428;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12434;
	wire [4-1:0] node12436;
	wire [4-1:0] node12437;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12444;
	wire [4-1:0] node12447;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12453;
	wire [4-1:0] node12457;
	wire [4-1:0] node12458;
	wire [4-1:0] node12459;
	wire [4-1:0] node12461;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12469;
	wire [4-1:0] node12472;
	wire [4-1:0] node12473;
	wire [4-1:0] node12474;
	wire [4-1:0] node12475;
	wire [4-1:0] node12476;
	wire [4-1:0] node12479;
	wire [4-1:0] node12480;
	wire [4-1:0] node12484;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12489;
	wire [4-1:0] node12492;
	wire [4-1:0] node12493;
	wire [4-1:0] node12496;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12503;
	wire [4-1:0] node12507;
	wire [4-1:0] node12508;
	wire [4-1:0] node12510;
	wire [4-1:0] node12513;
	wire [4-1:0] node12514;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12520;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12531;
	wire [4-1:0] node12534;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12539;
	wire [4-1:0] node12540;
	wire [4-1:0] node12541;
	wire [4-1:0] node12542;
	wire [4-1:0] node12543;
	wire [4-1:0] node12544;
	wire [4-1:0] node12547;
	wire [4-1:0] node12550;
	wire [4-1:0] node12551;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12559;
	wire [4-1:0] node12562;
	wire [4-1:0] node12563;
	wire [4-1:0] node12564;
	wire [4-1:0] node12568;
	wire [4-1:0] node12569;
	wire [4-1:0] node12573;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12577;
	wire [4-1:0] node12581;
	wire [4-1:0] node12582;
	wire [4-1:0] node12586;
	wire [4-1:0] node12587;
	wire [4-1:0] node12589;
	wire [4-1:0] node12592;
	wire [4-1:0] node12594;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12600;
	wire [4-1:0] node12603;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12608;
	wire [4-1:0] node12609;
	wire [4-1:0] node12613;
	wire [4-1:0] node12614;
	wire [4-1:0] node12616;
	wire [4-1:0] node12619;
	wire [4-1:0] node12622;
	wire [4-1:0] node12623;
	wire [4-1:0] node12624;
	wire [4-1:0] node12625;
	wire [4-1:0] node12628;
	wire [4-1:0] node12629;
	wire [4-1:0] node12633;
	wire [4-1:0] node12634;
	wire [4-1:0] node12637;
	wire [4-1:0] node12640;
	wire [4-1:0] node12641;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12647;
	wire [4-1:0] node12648;
	wire [4-1:0] node12651;
	wire [4-1:0] node12654;
	wire [4-1:0] node12656;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12661;
	wire [4-1:0] node12662;
	wire [4-1:0] node12663;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12669;
	wire [4-1:0] node12672;
	wire [4-1:0] node12673;
	wire [4-1:0] node12676;
	wire [4-1:0] node12679;
	wire [4-1:0] node12680;
	wire [4-1:0] node12681;
	wire [4-1:0] node12683;
	wire [4-1:0] node12686;
	wire [4-1:0] node12689;
	wire [4-1:0] node12690;
	wire [4-1:0] node12694;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12698;
	wire [4-1:0] node12699;
	wire [4-1:0] node12703;
	wire [4-1:0] node12705;
	wire [4-1:0] node12707;
	wire [4-1:0] node12710;
	wire [4-1:0] node12711;
	wire [4-1:0] node12712;
	wire [4-1:0] node12713;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12722;
	wire [4-1:0] node12723;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12730;
	wire [4-1:0] node12731;
	wire [4-1:0] node12733;
	wire [4-1:0] node12736;
	wire [4-1:0] node12740;
	wire [4-1:0] node12741;
	wire [4-1:0] node12742;
	wire [4-1:0] node12744;
	wire [4-1:0] node12747;
	wire [4-1:0] node12748;
	wire [4-1:0] node12751;
	wire [4-1:0] node12754;
	wire [4-1:0] node12756;
	wire [4-1:0] node12757;
	wire [4-1:0] node12761;
	wire [4-1:0] node12762;
	wire [4-1:0] node12763;
	wire [4-1:0] node12765;
	wire [4-1:0] node12766;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12772;
	wire [4-1:0] node12778;
	wire [4-1:0] node12779;
	wire [4-1:0] node12780;
	wire [4-1:0] node12781;
	wire [4-1:0] node12782;
	wire [4-1:0] node12783;
	wire [4-1:0] node12784;
	wire [4-1:0] node12787;
	wire [4-1:0] node12790;
	wire [4-1:0] node12791;
	wire [4-1:0] node12794;
	wire [4-1:0] node12796;
	wire [4-1:0] node12799;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12805;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12810;
	wire [4-1:0] node12813;
	wire [4-1:0] node12816;
	wire [4-1:0] node12817;
	wire [4-1:0] node12820;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12827;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12832;
	wire [4-1:0] node12834;
	wire [4-1:0] node12837;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12844;
	wire [4-1:0] node12845;
	wire [4-1:0] node12846;
	wire [4-1:0] node12847;
	wire [4-1:0] node12850;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12855;
	wire [4-1:0] node12858;
	wire [4-1:0] node12861;
	wire [4-1:0] node12862;
	wire [4-1:0] node12865;
	wire [4-1:0] node12868;
	wire [4-1:0] node12869;
	wire [4-1:0] node12870;
	wire [4-1:0] node12874;
	wire [4-1:0] node12875;
	wire [4-1:0] node12878;
	wire [4-1:0] node12881;
	wire [4-1:0] node12882;
	wire [4-1:0] node12883;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12889;
	wire [4-1:0] node12892;
	wire [4-1:0] node12893;
	wire [4-1:0] node12894;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12899;
	wire [4-1:0] node12902;
	wire [4-1:0] node12903;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12909;
	wire [4-1:0] node12913;
	wire [4-1:0] node12914;
	wire [4-1:0] node12917;
	wire [4-1:0] node12920;
	wire [4-1:0] node12922;
	wire [4-1:0] node12925;
	wire [4-1:0] node12926;
	wire [4-1:0] node12927;
	wire [4-1:0] node12930;
	wire [4-1:0] node12931;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12949;
	wire [4-1:0] node12952;
	wire [4-1:0] node12953;
	wire [4-1:0] node12957;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12963;
	wire [4-1:0] node12964;
	wire [4-1:0] node12967;
	wire [4-1:0] node12970;
	wire [4-1:0] node12971;
	wire [4-1:0] node12972;
	wire [4-1:0] node12974;
	wire [4-1:0] node12977;
	wire [4-1:0] node12978;
	wire [4-1:0] node12981;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12988;
	wire [4-1:0] node12990;
	wire [4-1:0] node12993;
	wire [4-1:0] node12994;
	wire [4-1:0] node12995;
	wire [4-1:0] node12996;
	wire [4-1:0] node12998;
	wire [4-1:0] node13001;
	wire [4-1:0] node13004;
	wire [4-1:0] node13005;
	wire [4-1:0] node13006;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13015;
	wire [4-1:0] node13017;
	wire [4-1:0] node13018;
	wire [4-1:0] node13022;
	wire [4-1:0] node13023;
	wire [4-1:0] node13024;
	wire [4-1:0] node13025;
	wire [4-1:0] node13026;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13034;
	wire [4-1:0] node13035;
	wire [4-1:0] node13037;
	wire [4-1:0] node13040;
	wire [4-1:0] node13042;
	wire [4-1:0] node13045;
	wire [4-1:0] node13047;
	wire [4-1:0] node13048;
	wire [4-1:0] node13052;
	wire [4-1:0] node13053;
	wire [4-1:0] node13054;
	wire [4-1:0] node13055;
	wire [4-1:0] node13056;
	wire [4-1:0] node13060;
	wire [4-1:0] node13062;
	wire [4-1:0] node13066;
	wire [4-1:0] node13069;
	wire [4-1:0] node13071;
	wire [4-1:0] node13072;
	wire [4-1:0] node13073;
	wire [4-1:0] node13075;
	wire [4-1:0] node13076;
	wire [4-1:0] node13077;
	wire [4-1:0] node13079;
	wire [4-1:0] node13080;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13084;
	wire [4-1:0] node13088;
	wire [4-1:0] node13089;
	wire [4-1:0] node13093;
	wire [4-1:0] node13095;
	wire [4-1:0] node13096;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13102;
	wire [4-1:0] node13103;
	wire [4-1:0] node13105;
	wire [4-1:0] node13108;
	wire [4-1:0] node13110;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13119;
	wire [4-1:0] node13123;
	wire [4-1:0] node13125;
	wire [4-1:0] node13128;
	wire [4-1:0] node13129;
	wire [4-1:0] node13130;
	wire [4-1:0] node13132;
	wire [4-1:0] node13135;
	wire [4-1:0] node13136;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13148;
	wire [4-1:0] node13150;
	wire [4-1:0] node13151;
	wire [4-1:0] node13154;
	wire [4-1:0] node13157;
	wire [4-1:0] node13159;
	wire [4-1:0] node13161;
	wire [4-1:0] node13162;
	wire [4-1:0] node13163;
	wire [4-1:0] node13164;
	wire [4-1:0] node13168;
	wire [4-1:0] node13170;
	wire [4-1:0] node13171;
	wire [4-1:0] node13175;
	wire [4-1:0] node13177;
	wire [4-1:0] node13178;
	wire [4-1:0] node13182;
	wire [4-1:0] node13183;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;
	wire [4-1:0] node13190;
	wire [4-1:0] node13193;
	wire [4-1:0] node13195;
	wire [4-1:0] node13198;
	wire [4-1:0] node13199;
	wire [4-1:0] node13201;
	wire [4-1:0] node13205;
	wire [4-1:0] node13206;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13210;
	wire [4-1:0] node13213;
	wire [4-1:0] node13216;
	wire [4-1:0] node13218;
	wire [4-1:0] node13219;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13231;
	wire [4-1:0] node13232;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13238;
	wire [4-1:0] node13239;
	wire [4-1:0] node13241;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13251;
	wire [4-1:0] node13252;
	wire [4-1:0] node13254;
	wire [4-1:0] node13257;
	wire [4-1:0] node13258;
	wire [4-1:0] node13259;
	wire [4-1:0] node13262;
	wire [4-1:0] node13265;
	wire [4-1:0] node13266;
	wire [4-1:0] node13270;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13273;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13279;
	wire [4-1:0] node13282;
	wire [4-1:0] node13285;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13292;
	wire [4-1:0] node13296;
	wire [4-1:0] node13297;
	wire [4-1:0] node13299;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13306;
	wire [4-1:0] node13309;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13312;
	wire [4-1:0] node13313;
	wire [4-1:0] node13316;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13321;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13328;
	wire [4-1:0] node13332;
	wire [4-1:0] node13333;
	wire [4-1:0] node13334;
	wire [4-1:0] node13335;
	wire [4-1:0] node13336;
	wire [4-1:0] node13340;
	wire [4-1:0] node13343;
	wire [4-1:0] node13344;
	wire [4-1:0] node13347;
	wire [4-1:0] node13350;
	wire [4-1:0] node13351;
	wire [4-1:0] node13353;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13363;
	wire [4-1:0] node13364;
	wire [4-1:0] node13365;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13369;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13377;
	wire [4-1:0] node13378;
	wire [4-1:0] node13381;
	wire [4-1:0] node13384;
	wire [4-1:0] node13385;
	wire [4-1:0] node13386;
	wire [4-1:0] node13389;
	wire [4-1:0] node13392;
	wire [4-1:0] node13394;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13400;
	wire [4-1:0] node13402;
	wire [4-1:0] node13405;
	wire [4-1:0] node13408;
	wire [4-1:0] node13409;
	wire [4-1:0] node13410;
	wire [4-1:0] node13413;
	wire [4-1:0] node13416;
	wire [4-1:0] node13417;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13431;
	wire [4-1:0] node13432;
	wire [4-1:0] node13433;
	wire [4-1:0] node13435;
	wire [4-1:0] node13438;
	wire [4-1:0] node13439;
	wire [4-1:0] node13443;
	wire [4-1:0] node13444;
	wire [4-1:0] node13445;
	wire [4-1:0] node13446;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13454;
	wire [4-1:0] node13458;
	wire [4-1:0] node13459;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13466;
	wire [4-1:0] node13469;
	wire [4-1:0] node13471;
	wire [4-1:0] node13472;
	wire [4-1:0] node13476;
	wire [4-1:0] node13477;
	wire [4-1:0] node13478;
	wire [4-1:0] node13480;
	wire [4-1:0] node13483;
	wire [4-1:0] node13484;
	wire [4-1:0] node13488;
	wire [4-1:0] node13489;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13497;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13503;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13513;
	wire [4-1:0] node13515;
	wire [4-1:0] node13518;
	wire [4-1:0] node13519;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13524;
	wire [4-1:0] node13528;
	wire [4-1:0] node13529;
	wire [4-1:0] node13533;
	wire [4-1:0] node13534;
	wire [4-1:0] node13535;
	wire [4-1:0] node13537;
	wire [4-1:0] node13540;
	wire [4-1:0] node13542;
	wire [4-1:0] node13545;
	wire [4-1:0] node13546;
	wire [4-1:0] node13547;
	wire [4-1:0] node13548;
	wire [4-1:0] node13552;
	wire [4-1:0] node13554;
	wire [4-1:0] node13557;
	wire [4-1:0] node13559;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13564;
	wire [4-1:0] node13565;
	wire [4-1:0] node13567;
	wire [4-1:0] node13570;
	wire [4-1:0] node13571;
	wire [4-1:0] node13572;
	wire [4-1:0] node13575;
	wire [4-1:0] node13578;
	wire [4-1:0] node13580;
	wire [4-1:0] node13583;
	wire [4-1:0] node13584;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13589;
	wire [4-1:0] node13593;
	wire [4-1:0] node13594;
	wire [4-1:0] node13596;
	wire [4-1:0] node13599;
	wire [4-1:0] node13600;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13606;
	wire [4-1:0] node13607;
	wire [4-1:0] node13608;
	wire [4-1:0] node13611;
	wire [4-1:0] node13615;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13622;
	wire [4-1:0] node13623;
	wire [4-1:0] node13624;
	wire [4-1:0] node13628;
	wire [4-1:0] node13631;
	wire [4-1:0] node13633;
	wire [4-1:0] node13635;
	wire [4-1:0] node13636;
	wire [4-1:0] node13638;
	wire [4-1:0] node13639;
	wire [4-1:0] node13640;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13646;
	wire [4-1:0] node13648;
	wire [4-1:0] node13651;
	wire [4-1:0] node13653;
	wire [4-1:0] node13654;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13663;
	wire [4-1:0] node13664;
	wire [4-1:0] node13665;
	wire [4-1:0] node13668;
	wire [4-1:0] node13672;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13682;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13687;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13695;
	wire [4-1:0] node13696;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13704;
	wire [4-1:0] node13705;
	wire [4-1:0] node13709;
	wire [4-1:0] node13710;
	wire [4-1:0] node13714;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13718;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13727;
	wire [4-1:0] node13728;
	wire [4-1:0] node13729;
	wire [4-1:0] node13731;
	wire [4-1:0] node13733;
	wire [4-1:0] node13738;
	wire [4-1:0] node13739;
	wire [4-1:0] node13740;
	wire [4-1:0] node13741;
	wire [4-1:0] node13742;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13745;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13748;
	wire [4-1:0] node13749;
	wire [4-1:0] node13750;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13757;
	wire [4-1:0] node13760;
	wire [4-1:0] node13761;
	wire [4-1:0] node13765;
	wire [4-1:0] node13766;
	wire [4-1:0] node13767;
	wire [4-1:0] node13769;
	wire [4-1:0] node13772;
	wire [4-1:0] node13773;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13782;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13786;
	wire [4-1:0] node13789;
	wire [4-1:0] node13790;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13797;
	wire [4-1:0] node13801;
	wire [4-1:0] node13802;
	wire [4-1:0] node13803;
	wire [4-1:0] node13804;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13807;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13816;
	wire [4-1:0] node13818;
	wire [4-1:0] node13821;
	wire [4-1:0] node13822;
	wire [4-1:0] node13824;
	wire [4-1:0] node13825;
	wire [4-1:0] node13829;
	wire [4-1:0] node13831;
	wire [4-1:0] node13834;
	wire [4-1:0] node13835;
	wire [4-1:0] node13836;
	wire [4-1:0] node13838;
	wire [4-1:0] node13841;
	wire [4-1:0] node13843;
	wire [4-1:0] node13846;
	wire [4-1:0] node13847;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13860;
	wire [4-1:0] node13861;
	wire [4-1:0] node13862;
	wire [4-1:0] node13864;
	wire [4-1:0] node13868;
	wire [4-1:0] node13870;
	wire [4-1:0] node13872;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13878;
	wire [4-1:0] node13881;
	wire [4-1:0] node13882;
	wire [4-1:0] node13883;
	wire [4-1:0] node13887;
	wire [4-1:0] node13888;
	wire [4-1:0] node13892;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13903;
	wire [4-1:0] node13906;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13912;
	wire [4-1:0] node13914;
	wire [4-1:0] node13915;
	wire [4-1:0] node13917;
	wire [4-1:0] node13918;
	wire [4-1:0] node13922;
	wire [4-1:0] node13923;
	wire [4-1:0] node13927;
	wire [4-1:0] node13928;
	wire [4-1:0] node13930;
	wire [4-1:0] node13933;
	wire [4-1:0] node13934;
	wire [4-1:0] node13936;
	wire [4-1:0] node13939;
	wire [4-1:0] node13941;
	wire [4-1:0] node13944;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13957;
	wire [4-1:0] node13958;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13965;
	wire [4-1:0] node13967;
	wire [4-1:0] node13970;
	wire [4-1:0] node13972;
	wire [4-1:0] node13975;
	wire [4-1:0] node13977;
	wire [4-1:0] node13980;
	wire [4-1:0] node13981;
	wire [4-1:0] node13982;
	wire [4-1:0] node13984;
	wire [4-1:0] node13987;
	wire [4-1:0] node13988;
	wire [4-1:0] node13992;
	wire [4-1:0] node13994;
	wire [4-1:0] node13997;
	wire [4-1:0] node13998;
	wire [4-1:0] node13999;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14002;
	wire [4-1:0] node14003;
	wire [4-1:0] node14005;
	wire [4-1:0] node14009;
	wire [4-1:0] node14011;
	wire [4-1:0] node14014;
	wire [4-1:0] node14015;
	wire [4-1:0] node14016;
	wire [4-1:0] node14017;
	wire [4-1:0] node14019;
	wire [4-1:0] node14022;
	wire [4-1:0] node14023;
	wire [4-1:0] node14027;
	wire [4-1:0] node14029;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14034;
	wire [4-1:0] node14036;
	wire [4-1:0] node14040;
	wire [4-1:0] node14042;
	wire [4-1:0] node14045;
	wire [4-1:0] node14046;
	wire [4-1:0] node14047;
	wire [4-1:0] node14048;
	wire [4-1:0] node14052;
	wire [4-1:0] node14053;
	wire [4-1:0] node14056;
	wire [4-1:0] node14058;
	wire [4-1:0] node14061;
	wire [4-1:0] node14062;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14068;
	wire [4-1:0] node14069;
	wire [4-1:0] node14073;
	wire [4-1:0] node14075;
	wire [4-1:0] node14078;
	wire [4-1:0] node14079;
	wire [4-1:0] node14080;
	wire [4-1:0] node14081;
	wire [4-1:0] node14082;
	wire [4-1:0] node14083;
	wire [4-1:0] node14084;
	wire [4-1:0] node14088;
	wire [4-1:0] node14090;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14096;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14103;
	wire [4-1:0] node14105;
	wire [4-1:0] node14108;
	wire [4-1:0] node14110;
	wire [4-1:0] node14113;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14119;
	wire [4-1:0] node14120;
	wire [4-1:0] node14122;
	wire [4-1:0] node14125;
	wire [4-1:0] node14126;
	wire [4-1:0] node14130;
	wire [4-1:0] node14131;
	wire [4-1:0] node14132;
	wire [4-1:0] node14134;
	wire [4-1:0] node14137;
	wire [4-1:0] node14138;
	wire [4-1:0] node14141;
	wire [4-1:0] node14142;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14152;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14158;
	wire [4-1:0] node14159;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14166;
	wire [4-1:0] node14167;
	wire [4-1:0] node14169;
	wire [4-1:0] node14173;
	wire [4-1:0] node14174;
	wire [4-1:0] node14178;
	wire [4-1:0] node14179;
	wire [4-1:0] node14180;
	wire [4-1:0] node14181;
	wire [4-1:0] node14182;
	wire [4-1:0] node14186;
	wire [4-1:0] node14187;
	wire [4-1:0] node14191;
	wire [4-1:0] node14193;
	wire [4-1:0] node14196;
	wire [4-1:0] node14197;
	wire [4-1:0] node14198;
	wire [4-1:0] node14200;
	wire [4-1:0] node14204;
	wire [4-1:0] node14206;
	wire [4-1:0] node14209;
	wire [4-1:0] node14210;
	wire [4-1:0] node14211;
	wire [4-1:0] node14212;
	wire [4-1:0] node14216;
	wire [4-1:0] node14217;
	wire [4-1:0] node14219;
	wire [4-1:0] node14221;
	wire [4-1:0] node14224;
	wire [4-1:0] node14225;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14231;
	wire [4-1:0] node14232;
	wire [4-1:0] node14236;
	wire [4-1:0] node14238;
	wire [4-1:0] node14241;
	wire [4-1:0] node14243;
	wire [4-1:0] node14246;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14251;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14261;
	wire [4-1:0] node14262;
	wire [4-1:0] node14264;
	wire [4-1:0] node14267;
	wire [4-1:0] node14269;
	wire [4-1:0] node14272;
	wire [4-1:0] node14274;
	wire [4-1:0] node14276;
	wire [4-1:0] node14279;
	wire [4-1:0] node14280;
	wire [4-1:0] node14281;
	wire [4-1:0] node14282;
	wire [4-1:0] node14286;
	wire [4-1:0] node14287;
	wire [4-1:0] node14289;
	wire [4-1:0] node14292;
	wire [4-1:0] node14295;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14302;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14309;
	wire [4-1:0] node14313;
	wire [4-1:0] node14314;
	wire [4-1:0] node14315;
	wire [4-1:0] node14316;
	wire [4-1:0] node14317;
	wire [4-1:0] node14319;
	wire [4-1:0] node14322;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14334;
	wire [4-1:0] node14336;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14343;
	wire [4-1:0] node14346;
	wire [4-1:0] node14347;
	wire [4-1:0] node14348;
	wire [4-1:0] node14349;
	wire [4-1:0] node14350;
	wire [4-1:0] node14354;
	wire [4-1:0] node14357;
	wire [4-1:0] node14358;
	wire [4-1:0] node14359;
	wire [4-1:0] node14363;
	wire [4-1:0] node14365;
	wire [4-1:0] node14368;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14374;
	wire [4-1:0] node14376;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14381;
	wire [4-1:0] node14382;
	wire [4-1:0] node14384;
	wire [4-1:0] node14385;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14404;
	wire [4-1:0] node14409;
	wire [4-1:0] node14410;
	wire [4-1:0] node14411;
	wire [4-1:0] node14412;
	wire [4-1:0] node14416;
	wire [4-1:0] node14417;
	wire [4-1:0] node14419;
	wire [4-1:0] node14422;
	wire [4-1:0] node14425;
	wire [4-1:0] node14426;
	wire [4-1:0] node14427;
	wire [4-1:0] node14431;
	wire [4-1:0] node14432;
	wire [4-1:0] node14433;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14442;
	wire [4-1:0] node14443;
	wire [4-1:0] node14445;
	wire [4-1:0] node14446;
	wire [4-1:0] node14450;
	wire [4-1:0] node14452;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14463;
	wire [4-1:0] node14468;
	wire [4-1:0] node14469;
	wire [4-1:0] node14470;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14477;
	wire [4-1:0] node14480;
	wire [4-1:0] node14482;
	wire [4-1:0] node14485;
	wire [4-1:0] node14486;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14490;
	wire [4-1:0] node14493;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14499;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14505;
	wire [4-1:0] node14507;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14515;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14521;
	wire [4-1:0] node14522;
	wire [4-1:0] node14524;
	wire [4-1:0] node14527;
	wire [4-1:0] node14528;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14534;
	wire [4-1:0] node14535;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14539;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14547;
	wire [4-1:0] node14549;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14555;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14564;
	wire [4-1:0] node14566;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14572;
	wire [4-1:0] node14574;
	wire [4-1:0] node14577;
	wire [4-1:0] node14579;
	wire [4-1:0] node14582;
	wire [4-1:0] node14583;
	wire [4-1:0] node14587;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14593;
	wire [4-1:0] node14594;
	wire [4-1:0] node14596;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14602;
	wire [4-1:0] node14603;
	wire [4-1:0] node14604;
	wire [4-1:0] node14608;
	wire [4-1:0] node14610;
	wire [4-1:0] node14613;
	wire [4-1:0] node14615;
	wire [4-1:0] node14618;
	wire [4-1:0] node14619;
	wire [4-1:0] node14620;
	wire [4-1:0] node14621;
	wire [4-1:0] node14625;
	wire [4-1:0] node14626;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14636;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14640;
	wire [4-1:0] node14641;
	wire [4-1:0] node14642;
	wire [4-1:0] node14643;
	wire [4-1:0] node14644;
	wire [4-1:0] node14647;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14655;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14666;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14675;
	wire [4-1:0] node14676;
	wire [4-1:0] node14679;
	wire [4-1:0] node14682;
	wire [4-1:0] node14683;
	wire [4-1:0] node14686;
	wire [4-1:0] node14689;
	wire [4-1:0] node14690;
	wire [4-1:0] node14691;
	wire [4-1:0] node14693;
	wire [4-1:0] node14694;
	wire [4-1:0] node14698;
	wire [4-1:0] node14699;
	wire [4-1:0] node14700;
	wire [4-1:0] node14703;
	wire [4-1:0] node14707;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14710;
	wire [4-1:0] node14711;
	wire [4-1:0] node14715;
	wire [4-1:0] node14717;
	wire [4-1:0] node14720;
	wire [4-1:0] node14721;
	wire [4-1:0] node14723;
	wire [4-1:0] node14726;
	wire [4-1:0] node14729;
	wire [4-1:0] node14730;
	wire [4-1:0] node14732;
	wire [4-1:0] node14735;
	wire [4-1:0] node14736;
	wire [4-1:0] node14737;
	wire [4-1:0] node14740;
	wire [4-1:0] node14744;
	wire [4-1:0] node14745;
	wire [4-1:0] node14746;
	wire [4-1:0] node14747;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14751;
	wire [4-1:0] node14754;
	wire [4-1:0] node14755;
	wire [4-1:0] node14758;
	wire [4-1:0] node14761;
	wire [4-1:0] node14762;
	wire [4-1:0] node14764;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14771;
	wire [4-1:0] node14774;
	wire [4-1:0] node14776;
	wire [4-1:0] node14779;
	wire [4-1:0] node14780;
	wire [4-1:0] node14782;
	wire [4-1:0] node14784;
	wire [4-1:0] node14786;
	wire [4-1:0] node14789;
	wire [4-1:0] node14790;
	wire [4-1:0] node14791;
	wire [4-1:0] node14792;
	wire [4-1:0] node14795;
	wire [4-1:0] node14799;
	wire [4-1:0] node14801;
	wire [4-1:0] node14802;
	wire [4-1:0] node14805;
	wire [4-1:0] node14808;
	wire [4-1:0] node14809;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14813;
	wire [4-1:0] node14817;
	wire [4-1:0] node14818;
	wire [4-1:0] node14821;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14828;
	wire [4-1:0] node14829;
	wire [4-1:0] node14833;
	wire [4-1:0] node14834;
	wire [4-1:0] node14835;
	wire [4-1:0] node14838;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14845;
	wire [4-1:0] node14848;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14855;
	wire [4-1:0] node14856;
	wire [4-1:0] node14858;
	wire [4-1:0] node14861;
	wire [4-1:0] node14864;
	wire [4-1:0] node14866;
	wire [4-1:0] node14868;
	wire [4-1:0] node14871;
	wire [4-1:0] node14872;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14876;
	wire [4-1:0] node14878;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14884;
	wire [4-1:0] node14887;
	wire [4-1:0] node14888;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14895;
	wire [4-1:0] node14897;
	wire [4-1:0] node14900;
	wire [4-1:0] node14901;
	wire [4-1:0] node14902;
	wire [4-1:0] node14907;
	wire [4-1:0] node14908;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14912;
	wire [4-1:0] node14915;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14923;
	wire [4-1:0] node14924;
	wire [4-1:0] node14926;
	wire [4-1:0] node14927;
	wire [4-1:0] node14930;
	wire [4-1:0] node14934;
	wire [4-1:0] node14935;
	wire [4-1:0] node14936;
	wire [4-1:0] node14937;
	wire [4-1:0] node14938;
	wire [4-1:0] node14939;
	wire [4-1:0] node14942;
	wire [4-1:0] node14945;
	wire [4-1:0] node14946;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14955;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14958;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14965;
	wire [4-1:0] node14968;
	wire [4-1:0] node14971;
	wire [4-1:0] node14972;
	wire [4-1:0] node14975;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14980;
	wire [4-1:0] node14984;
	wire [4-1:0] node14985;
	wire [4-1:0] node14986;
	wire [4-1:0] node14988;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14995;
	wire [4-1:0] node14998;
	wire [4-1:0] node15000;
	wire [4-1:0] node15003;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15006;
	wire [4-1:0] node15007;
	wire [4-1:0] node15008;
	wire [4-1:0] node15012;
	wire [4-1:0] node15013;
	wire [4-1:0] node15015;
	wire [4-1:0] node15018;
	wire [4-1:0] node15019;
	wire [4-1:0] node15022;
	wire [4-1:0] node15025;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15028;
	wire [4-1:0] node15031;
	wire [4-1:0] node15034;
	wire [4-1:0] node15035;
	wire [4-1:0] node15038;
	wire [4-1:0] node15041;
	wire [4-1:0] node15042;
	wire [4-1:0] node15046;
	wire [4-1:0] node15047;
	wire [4-1:0] node15048;
	wire [4-1:0] node15049;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15055;
	wire [4-1:0] node15059;
	wire [4-1:0] node15060;
	wire [4-1:0] node15063;
	wire [4-1:0] node15066;
	wire [4-1:0] node15067;
	wire [4-1:0] node15068;
	wire [4-1:0] node15070;
	wire [4-1:0] node15073;
	wire [4-1:0] node15074;
	wire [4-1:0] node15077;
	wire [4-1:0] node15080;
	wire [4-1:0] node15082;
	wire [4-1:0] node15085;
	wire [4-1:0] node15086;
	wire [4-1:0] node15087;
	wire [4-1:0] node15089;
	wire [4-1:0] node15092;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15097;
	wire [4-1:0] node15100;
	wire [4-1:0] node15101;
	wire [4-1:0] node15103;
	wire [4-1:0] node15106;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15111;
	wire [4-1:0] node15112;
	wire [4-1:0] node15115;
	wire [4-1:0] node15118;
	wire [4-1:0] node15119;
	wire [4-1:0] node15122;
	wire [4-1:0] node15125;
	wire [4-1:0] node15127;
	wire [4-1:0] node15130;
	wire [4-1:0] node15131;
	wire [4-1:0] node15132;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15136;
	wire [4-1:0] node15137;
	wire [4-1:0] node15140;
	wire [4-1:0] node15143;
	wire [4-1:0] node15144;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15150;
	wire [4-1:0] node15153;
	wire [4-1:0] node15156;
	wire [4-1:0] node15158;
	wire [4-1:0] node15159;
	wire [4-1:0] node15162;
	wire [4-1:0] node15165;
	wire [4-1:0] node15166;
	wire [4-1:0] node15167;
	wire [4-1:0] node15168;
	wire [4-1:0] node15172;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15178;
	wire [4-1:0] node15182;
	wire [4-1:0] node15183;
	wire [4-1:0] node15184;
	wire [4-1:0] node15185;
	wire [4-1:0] node15186;
	wire [4-1:0] node15189;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15196;
	wire [4-1:0] node15199;
	wire [4-1:0] node15200;
	wire [4-1:0] node15201;
	wire [4-1:0] node15204;
	wire [4-1:0] node15207;
	wire [4-1:0] node15209;
	wire [4-1:0] node15212;
	wire [4-1:0] node15213;
	wire [4-1:0] node15214;
	wire [4-1:0] node15216;
	wire [4-1:0] node15220;
	wire [4-1:0] node15221;
	wire [4-1:0] node15222;
	wire [4-1:0] node15225;
	wire [4-1:0] node15228;
	wire [4-1:0] node15230;
	wire [4-1:0] node15231;
	wire [4-1:0] node15234;
	wire [4-1:0] node15237;
	wire [4-1:0] node15238;
	wire [4-1:0] node15239;
	wire [4-1:0] node15240;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15243;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15251;
	wire [4-1:0] node15254;
	wire [4-1:0] node15255;
	wire [4-1:0] node15258;
	wire [4-1:0] node15261;
	wire [4-1:0] node15262;
	wire [4-1:0] node15264;
	wire [4-1:0] node15267;
	wire [4-1:0] node15269;
	wire [4-1:0] node15272;
	wire [4-1:0] node15273;
	wire [4-1:0] node15275;
	wire [4-1:0] node15277;
	wire [4-1:0] node15280;
	wire [4-1:0] node15281;
	wire [4-1:0] node15283;
	wire [4-1:0] node15286;
	wire [4-1:0] node15289;
	wire [4-1:0] node15290;
	wire [4-1:0] node15291;
	wire [4-1:0] node15292;
	wire [4-1:0] node15294;
	wire [4-1:0] node15297;
	wire [4-1:0] node15300;
	wire [4-1:0] node15302;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15307;
	wire [4-1:0] node15308;
	wire [4-1:0] node15311;
	wire [4-1:0] node15315;
	wire [4-1:0] node15316;
	wire [4-1:0] node15319;
	wire [4-1:0] node15320;
	wire [4-1:0] node15324;
	wire [4-1:0] node15325;
	wire [4-1:0] node15326;
	wire [4-1:0] node15327;
	wire [4-1:0] node15328;
	wire [4-1:0] node15330;
	wire [4-1:0] node15331;
	wire [4-1:0] node15334;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15341;
	wire [4-1:0] node15343;
	wire [4-1:0] node15346;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15351;
	wire [4-1:0] node15353;
	wire [4-1:0] node15357;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15360;
	wire [4-1:0] node15362;
	wire [4-1:0] node15363;
	wire [4-1:0] node15366;
	wire [4-1:0] node15369;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15377;
	wire [4-1:0] node15380;
	wire [4-1:0] node15381;
	wire [4-1:0] node15383;
	wire [4-1:0] node15386;
	wire [4-1:0] node15387;
	wire [4-1:0] node15391;
	wire [4-1:0] node15392;
	wire [4-1:0] node15394;
	wire [4-1:0] node15397;
	wire [4-1:0] node15398;
	wire [4-1:0] node15400;
	wire [4-1:0] node15404;
	wire [4-1:0] node15405;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15409;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15416;
	wire [4-1:0] node15419;
	wire [4-1:0] node15420;
	wire [4-1:0] node15422;
	wire [4-1:0] node15425;
	wire [4-1:0] node15426;
	wire [4-1:0] node15429;
	wire [4-1:0] node15432;
	wire [4-1:0] node15433;
	wire [4-1:0] node15435;
	wire [4-1:0] node15436;
	wire [4-1:0] node15440;
	wire [4-1:0] node15442;
	wire [4-1:0] node15445;
	wire [4-1:0] node15446;
	wire [4-1:0] node15447;
	wire [4-1:0] node15448;
	wire [4-1:0] node15449;
	wire [4-1:0] node15450;
	wire [4-1:0] node15451;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15455;
	wire [4-1:0] node15460;
	wire [4-1:0] node15461;
	wire [4-1:0] node15463;
	wire [4-1:0] node15466;
	wire [4-1:0] node15467;
	wire [4-1:0] node15469;
	wire [4-1:0] node15472;
	wire [4-1:0] node15473;
	wire [4-1:0] node15477;
	wire [4-1:0] node15478;
	wire [4-1:0] node15480;
	wire [4-1:0] node15482;
	wire [4-1:0] node15484;
	wire [4-1:0] node15488;
	wire [4-1:0] node15489;
	wire [4-1:0] node15490;
	wire [4-1:0] node15492;
	wire [4-1:0] node15495;
	wire [4-1:0] node15496;
	wire [4-1:0] node15497;
	wire [4-1:0] node15501;
	wire [4-1:0] node15503;
	wire [4-1:0] node15506;
	wire [4-1:0] node15507;
	wire [4-1:0] node15508;
	wire [4-1:0] node15510;
	wire [4-1:0] node15513;
	wire [4-1:0] node15515;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15532;
	wire [4-1:0] node15534;
	wire [4-1:0] node15537;
	wire [4-1:0] node15538;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15545;
	wire [4-1:0] node15548;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15553;
	wire [4-1:0] node15556;
	wire [4-1:0] node15557;
	wire [4-1:0] node15561;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15564;
	wire [4-1:0] node15566;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15574;
	wire [4-1:0] node15576;
	wire [4-1:0] node15579;
	wire [4-1:0] node15580;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15584;
	wire [4-1:0] node15587;
	wire [4-1:0] node15588;
	wire [4-1:0] node15592;
	wire [4-1:0] node15594;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15600;
	wire [4-1:0] node15603;
	wire [4-1:0] node15604;
	wire [4-1:0] node15605;
	wire [4-1:0] node15609;
	wire [4-1:0] node15612;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15615;
	wire [4-1:0] node15616;
	wire [4-1:0] node15617;
	wire [4-1:0] node15619;
	wire [4-1:0] node15622;
	wire [4-1:0] node15623;
	wire [4-1:0] node15627;
	wire [4-1:0] node15628;
	wire [4-1:0] node15629;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15638;
	wire [4-1:0] node15639;
	wire [4-1:0] node15640;
	wire [4-1:0] node15644;
	wire [4-1:0] node15645;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15651;
	wire [4-1:0] node15653;
	wire [4-1:0] node15656;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15665;
	wire [4-1:0] node15669;
	wire [4-1:0] node15670;
	wire [4-1:0] node15671;
	wire [4-1:0] node15675;
	wire [4-1:0] node15676;
	wire [4-1:0] node15680;
	wire [4-1:0] node15681;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15685;
	wire [4-1:0] node15687;
	wire [4-1:0] node15690;
	wire [4-1:0] node15691;
	wire [4-1:0] node15695;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15705;
	wire [4-1:0] node15708;
	wire [4-1:0] node15709;
	wire [4-1:0] node15712;
	wire [4-1:0] node15715;
	wire [4-1:0] node15716;
	wire [4-1:0] node15717;
	wire [4-1:0] node15719;
	wire [4-1:0] node15722;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15728;
	wire [4-1:0] node15731;
	wire [4-1:0] node15732;
	wire [4-1:0] node15734;
	wire [4-1:0] node15737;
	wire [4-1:0] node15738;
	wire [4-1:0] node15742;
	wire [4-1:0] node15743;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15746;
	wire [4-1:0] node15749;
	wire [4-1:0] node15751;
	wire [4-1:0] node15754;
	wire [4-1:0] node15756;
	wire [4-1:0] node15758;
	wire [4-1:0] node15761;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15767;
	wire [4-1:0] node15768;
	wire [4-1:0] node15772;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15776;
	wire [4-1:0] node15779;
	wire [4-1:0] node15782;
	wire [4-1:0] node15783;
	wire [4-1:0] node15785;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15794;
	wire [4-1:0] node15796;
	wire [4-1:0] node15800;
	wire [4-1:0] node15801;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15805;
	wire [4-1:0] node15806;
	wire [4-1:0] node15807;
	wire [4-1:0] node15809;
	wire [4-1:0] node15810;
	wire [4-1:0] node15811;
	wire [4-1:0] node15816;
	wire [4-1:0] node15817;
	wire [4-1:0] node15819;
	wire [4-1:0] node15822;
	wire [4-1:0] node15823;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15829;
	wire [4-1:0] node15830;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15839;
	wire [4-1:0] node15840;
	wire [4-1:0] node15844;
	wire [4-1:0] node15845;
	wire [4-1:0] node15846;
	wire [4-1:0] node15847;
	wire [4-1:0] node15848;
	wire [4-1:0] node15851;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15859;
	wire [4-1:0] node15863;
	wire [4-1:0] node15864;
	wire [4-1:0] node15865;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15873;
	wire [4-1:0] node15875;
	wire [4-1:0] node15878;
	wire [4-1:0] node15880;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15886;
	wire [4-1:0] node15890;
	wire [4-1:0] node15891;
	wire [4-1:0] node15893;
	wire [4-1:0] node15894;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15903;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15906;
	wire [4-1:0] node15907;
	wire [4-1:0] node15910;
	wire [4-1:0] node15911;
	wire [4-1:0] node15913;
	wire [4-1:0] node15916;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15925;
	wire [4-1:0] node15928;
	wire [4-1:0] node15929;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15936;
	wire [4-1:0] node15939;
	wire [4-1:0] node15940;
	wire [4-1:0] node15944;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15953;
	wire [4-1:0] node15956;
	wire [4-1:0] node15957;
	wire [4-1:0] node15960;
	wire [4-1:0] node15961;
	wire [4-1:0] node15963;
	wire [4-1:0] node15966;
	wire [4-1:0] node15967;
	wire [4-1:0] node15971;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15975;
	wire [4-1:0] node15978;
	wire [4-1:0] node15979;
	wire [4-1:0] node15980;
	wire [4-1:0] node15983;
	wire [4-1:0] node15987;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15997;
	wire [4-1:0] node15998;
	wire [4-1:0] node16002;
	wire [4-1:0] node16003;
	wire [4-1:0] node16004;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16009;
	wire [4-1:0] node16013;
	wire [4-1:0] node16016;
	wire [4-1:0] node16018;
	wire [4-1:0] node16021;
	wire [4-1:0] node16022;
	wire [4-1:0] node16023;
	wire [4-1:0] node16026;
	wire [4-1:0] node16029;
	wire [4-1:0] node16032;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16041;
	wire [4-1:0] node16044;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16048;
	wire [4-1:0] node16052;
	wire [4-1:0] node16055;
	wire [4-1:0] node16056;
	wire [4-1:0] node16057;
	wire [4-1:0] node16058;
	wire [4-1:0] node16059;
	wire [4-1:0] node16063;
	wire [4-1:0] node16064;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16070;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16081;
	wire [4-1:0] node16082;
	wire [4-1:0] node16083;
	wire [4-1:0] node16087;
	wire [4-1:0] node16089;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16097;
	wire [4-1:0] node16098;
	wire [4-1:0] node16099;
	wire [4-1:0] node16102;
	wire [4-1:0] node16105;
	wire [4-1:0] node16106;
	wire [4-1:0] node16110;
	wire [4-1:0] node16111;
	wire [4-1:0] node16112;
	wire [4-1:0] node16113;
	wire [4-1:0] node16114;
	wire [4-1:0] node16115;
	wire [4-1:0] node16119;
	wire [4-1:0] node16120;
	wire [4-1:0] node16122;
	wire [4-1:0] node16125;
	wire [4-1:0] node16126;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16132;
	wire [4-1:0] node16136;
	wire [4-1:0] node16137;
	wire [4-1:0] node16138;
	wire [4-1:0] node16142;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16149;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16157;
	wire [4-1:0] node16160;
	wire [4-1:0] node16161;
	wire [4-1:0] node16165;
	wire [4-1:0] node16166;
	wire [4-1:0] node16168;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16177;
	wire [4-1:0] node16178;
	wire [4-1:0] node16179;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16182;
	wire [4-1:0] node16183;
	wire [4-1:0] node16184;
	wire [4-1:0] node16185;
	wire [4-1:0] node16189;
	wire [4-1:0] node16191;
	wire [4-1:0] node16194;
	wire [4-1:0] node16195;
	wire [4-1:0] node16196;
	wire [4-1:0] node16200;
	wire [4-1:0] node16201;
	wire [4-1:0] node16204;
	wire [4-1:0] node16207;
	wire [4-1:0] node16209;
	wire [4-1:0] node16210;
	wire [4-1:0] node16213;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16225;
	wire [4-1:0] node16226;
	wire [4-1:0] node16228;
	wire [4-1:0] node16231;
	wire [4-1:0] node16232;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16246;
	wire [4-1:0] node16249;
	wire [4-1:0] node16250;
	wire [4-1:0] node16251;
	wire [4-1:0] node16252;
	wire [4-1:0] node16253;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16266;
	wire [4-1:0] node16267;
	wire [4-1:0] node16268;
	wire [4-1:0] node16269;
	wire [4-1:0] node16273;
	wire [4-1:0] node16274;
	wire [4-1:0] node16277;
	wire [4-1:0] node16280;
	wire [4-1:0] node16281;
	wire [4-1:0] node16285;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16288;
	wire [4-1:0] node16291;
	wire [4-1:0] node16294;
	wire [4-1:0] node16297;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16303;
	wire [4-1:0] node16304;
	wire [4-1:0] node16307;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16313;
	wire [4-1:0] node16314;
	wire [4-1:0] node16316;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16324;
	wire [4-1:0] node16325;
	wire [4-1:0] node16327;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16333;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16344;
	wire [4-1:0] node16346;
	wire [4-1:0] node16349;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16356;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16360;
	wire [4-1:0] node16361;
	wire [4-1:0] node16365;
	wire [4-1:0] node16368;
	wire [4-1:0] node16370;
	wire [4-1:0] node16373;
	wire [4-1:0] node16374;
	wire [4-1:0] node16375;
	wire [4-1:0] node16376;
	wire [4-1:0] node16380;
	wire [4-1:0] node16381;
	wire [4-1:0] node16384;
	wire [4-1:0] node16387;
	wire [4-1:0] node16390;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16396;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16402;
	wire [4-1:0] node16406;
	wire [4-1:0] node16408;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16415;
	wire [4-1:0] node16416;
	wire [4-1:0] node16419;
	wire [4-1:0] node16421;
	wire [4-1:0] node16424;
	wire [4-1:0] node16425;
	wire [4-1:0] node16426;
	wire [4-1:0] node16429;
	wire [4-1:0] node16430;
	wire [4-1:0] node16434;
	wire [4-1:0] node16436;
	wire [4-1:0] node16438;
	wire [4-1:0] node16441;
	wire [4-1:0] node16442;
	wire [4-1:0] node16443;
	wire [4-1:0] node16444;
	wire [4-1:0] node16446;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16454;
	wire [4-1:0] node16455;
	wire [4-1:0] node16456;
	wire [4-1:0] node16460;
	wire [4-1:0] node16463;
	wire [4-1:0] node16464;
	wire [4-1:0] node16465;
	wire [4-1:0] node16468;
	wire [4-1:0] node16471;
	wire [4-1:0] node16473;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16479;
	wire [4-1:0] node16480;
	wire [4-1:0] node16481;
	wire [4-1:0] node16484;
	wire [4-1:0] node16488;
	wire [4-1:0] node16489;
	wire [4-1:0] node16491;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16499;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16507;
	wire [4-1:0] node16509;
	wire [4-1:0] node16512;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16515;
	wire [4-1:0] node16519;
	wire [4-1:0] node16521;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16526;
	wire [4-1:0] node16527;
	wire [4-1:0] node16530;
	wire [4-1:0] node16534;
	wire [4-1:0] node16536;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16541;
	wire [4-1:0] node16542;
	wire [4-1:0] node16543;
	wire [4-1:0] node16547;
	wire [4-1:0] node16548;
	wire [4-1:0] node16550;
	wire [4-1:0] node16553;
	wire [4-1:0] node16554;
	wire [4-1:0] node16557;
	wire [4-1:0] node16560;
	wire [4-1:0] node16561;
	wire [4-1:0] node16562;
	wire [4-1:0] node16564;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16571;
	wire [4-1:0] node16574;
	wire [4-1:0] node16575;
	wire [4-1:0] node16576;
	wire [4-1:0] node16579;
	wire [4-1:0] node16582;
	wire [4-1:0] node16584;
	wire [4-1:0] node16587;
	wire [4-1:0] node16588;
	wire [4-1:0] node16589;
	wire [4-1:0] node16591;
	wire [4-1:0] node16594;
	wire [4-1:0] node16595;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16603;
	wire [4-1:0] node16604;
	wire [4-1:0] node16605;
	wire [4-1:0] node16606;
	wire [4-1:0] node16608;
	wire [4-1:0] node16609;
	wire [4-1:0] node16610;
	wire [4-1:0] node16613;
	wire [4-1:0] node16616;
	wire [4-1:0] node16619;
	wire [4-1:0] node16620;
	wire [4-1:0] node16621;
	wire [4-1:0] node16622;
	wire [4-1:0] node16627;
	wire [4-1:0] node16628;
	wire [4-1:0] node16630;
	wire [4-1:0] node16633;
	wire [4-1:0] node16634;
	wire [4-1:0] node16637;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16644;
	wire [4-1:0] node16645;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16659;
	wire [4-1:0] node16660;
	wire [4-1:0] node16661;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16669;
	wire [4-1:0] node16672;
	wire [4-1:0] node16673;
	wire [4-1:0] node16675;
	wire [4-1:0] node16679;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16682;
	wire [4-1:0] node16683;
	wire [4-1:0] node16684;
	wire [4-1:0] node16689;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16699;
	wire [4-1:0] node16703;
	wire [4-1:0] node16706;
	wire [4-1:0] node16707;
	wire [4-1:0] node16711;
	wire [4-1:0] node16712;
	wire [4-1:0] node16713;
	wire [4-1:0] node16714;
	wire [4-1:0] node16717;
	wire [4-1:0] node16720;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16731;
	wire [4-1:0] node16734;
	wire [4-1:0] node16737;
	wire [4-1:0] node16740;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16745;
	wire [4-1:0] node16747;
	wire [4-1:0] node16750;
	wire [4-1:0] node16753;
	wire [4-1:0] node16754;
	wire [4-1:0] node16755;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16766;
	wire [4-1:0] node16767;
	wire [4-1:0] node16769;
	wire [4-1:0] node16772;
	wire [4-1:0] node16774;
	wire [4-1:0] node16776;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16781;
	wire [4-1:0] node16782;
	wire [4-1:0] node16783;
	wire [4-1:0] node16787;
	wire [4-1:0] node16789;
	wire [4-1:0] node16792;
	wire [4-1:0] node16793;
	wire [4-1:0] node16794;
	wire [4-1:0] node16797;
	wire [4-1:0] node16800;
	wire [4-1:0] node16803;
	wire [4-1:0] node16804;
	wire [4-1:0] node16806;
	wire [4-1:0] node16807;
	wire [4-1:0] node16810;
	wire [4-1:0] node16813;
	wire [4-1:0] node16814;
	wire [4-1:0] node16817;
	wire [4-1:0] node16818;
	wire [4-1:0] node16821;
	wire [4-1:0] node16824;
	wire [4-1:0] node16825;
	wire [4-1:0] node16826;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16836;
	wire [4-1:0] node16838;
	wire [4-1:0] node16841;
	wire [4-1:0] node16842;
	wire [4-1:0] node16844;
	wire [4-1:0] node16847;
	wire [4-1:0] node16850;
	wire [4-1:0] node16851;
	wire [4-1:0] node16852;
	wire [4-1:0] node16853;
	wire [4-1:0] node16857;
	wire [4-1:0] node16858;
	wire [4-1:0] node16861;
	wire [4-1:0] node16862;
	wire [4-1:0] node16865;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16870;
	wire [4-1:0] node16871;
	wire [4-1:0] node16875;
	wire [4-1:0] node16877;
	wire [4-1:0] node16880;
	wire [4-1:0] node16881;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16890;
	wire [4-1:0] node16892;
	wire [4-1:0] node16895;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16901;
	wire [4-1:0] node16903;
	wire [4-1:0] node16906;
	wire [4-1:0] node16907;
	wire [4-1:0] node16911;
	wire [4-1:0] node16912;
	wire [4-1:0] node16913;
	wire [4-1:0] node16915;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16928;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16936;
	wire [4-1:0] node16937;
	wire [4-1:0] node16938;
	wire [4-1:0] node16939;
	wire [4-1:0] node16940;
	wire [4-1:0] node16944;
	wire [4-1:0] node16945;
	wire [4-1:0] node16949;
	wire [4-1:0] node16950;
	wire [4-1:0] node16951;
	wire [4-1:0] node16954;
	wire [4-1:0] node16957;
	wire [4-1:0] node16959;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16966;
	wire [4-1:0] node16969;
	wire [4-1:0] node16970;
	wire [4-1:0] node16973;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16978;
	wire [4-1:0] node16981;
	wire [4-1:0] node16984;
	wire [4-1:0] node16985;
	wire [4-1:0] node16988;
	wire [4-1:0] node16991;
	wire [4-1:0] node16992;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16995;
	wire [4-1:0] node16996;
	wire [4-1:0] node17000;
	wire [4-1:0] node17002;
	wire [4-1:0] node17005;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17010;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17015;
	wire [4-1:0] node17018;
	wire [4-1:0] node17022;
	wire [4-1:0] node17024;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17030;
	wire [4-1:0] node17031;
	wire [4-1:0] node17034;
	wire [4-1:0] node17037;
	wire [4-1:0] node17038;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17042;
	wire [4-1:0] node17045;
	wire [4-1:0] node17047;
	wire [4-1:0] node17050;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17058;
	wire [4-1:0] node17059;
	wire [4-1:0] node17060;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17063;
	wire [4-1:0] node17064;
	wire [4-1:0] node17066;
	wire [4-1:0] node17069;
	wire [4-1:0] node17070;
	wire [4-1:0] node17072;
	wire [4-1:0] node17075;
	wire [4-1:0] node17078;
	wire [4-1:0] node17079;
	wire [4-1:0] node17081;
	wire [4-1:0] node17083;
	wire [4-1:0] node17086;
	wire [4-1:0] node17088;
	wire [4-1:0] node17091;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17095;
	wire [4-1:0] node17098;
	wire [4-1:0] node17101;
	wire [4-1:0] node17103;
	wire [4-1:0] node17106;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17113;
	wire [4-1:0] node17114;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17121;
	wire [4-1:0] node17124;
	wire [4-1:0] node17125;
	wire [4-1:0] node17126;
	wire [4-1:0] node17127;
	wire [4-1:0] node17128;
	wire [4-1:0] node17129;
	wire [4-1:0] node17133;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17141;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17144;
	wire [4-1:0] node17148;
	wire [4-1:0] node17151;
	wire [4-1:0] node17152;
	wire [4-1:0] node17153;
	wire [4-1:0] node17156;
	wire [4-1:0] node17160;
	wire [4-1:0] node17161;
	wire [4-1:0] node17162;
	wire [4-1:0] node17163;
	wire [4-1:0] node17164;
	wire [4-1:0] node17167;
	wire [4-1:0] node17170;
	wire [4-1:0] node17171;
	wire [4-1:0] node17174;
	wire [4-1:0] node17177;
	wire [4-1:0] node17178;
	wire [4-1:0] node17179;
	wire [4-1:0] node17182;
	wire [4-1:0] node17185;
	wire [4-1:0] node17187;
	wire [4-1:0] node17190;
	wire [4-1:0] node17191;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17198;
	wire [4-1:0] node17200;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17207;
	wire [4-1:0] node17209;
	wire [4-1:0] node17212;
	wire [4-1:0] node17213;
	wire [4-1:0] node17215;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17223;
	wire [4-1:0] node17224;
	wire [4-1:0] node17226;
	wire [4-1:0] node17227;
	wire [4-1:0] node17230;
	wire [4-1:0] node17233;
	wire [4-1:0] node17234;
	wire [4-1:0] node17236;
	wire [4-1:0] node17240;
	wire [4-1:0] node17241;
	wire [4-1:0] node17242;
	wire [4-1:0] node17243;
	wire [4-1:0] node17244;
	wire [4-1:0] node17248;
	wire [4-1:0] node17250;
	wire [4-1:0] node17253;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17262;
	wire [4-1:0] node17265;
	wire [4-1:0] node17267;
	wire [4-1:0] node17270;
	wire [4-1:0] node17271;
	wire [4-1:0] node17273;
	wire [4-1:0] node17277;
	wire [4-1:0] node17278;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17285;
	wire [4-1:0] node17286;
	wire [4-1:0] node17287;
	wire [4-1:0] node17290;
	wire [4-1:0] node17293;
	wire [4-1:0] node17294;
	wire [4-1:0] node17297;
	wire [4-1:0] node17300;
	wire [4-1:0] node17301;
	wire [4-1:0] node17302;
	wire [4-1:0] node17306;
	wire [4-1:0] node17307;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17314;
	wire [4-1:0] node17315;
	wire [4-1:0] node17316;
	wire [4-1:0] node17317;
	wire [4-1:0] node17319;
	wire [4-1:0] node17320;
	wire [4-1:0] node17324;
	wire [4-1:0] node17325;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17333;
	wire [4-1:0] node17337;
	wire [4-1:0] node17340;
	wire [4-1:0] node17341;
	wire [4-1:0] node17342;
	wire [4-1:0] node17343;
	wire [4-1:0] node17344;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17353;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17360;
	wire [4-1:0] node17361;
	wire [4-1:0] node17362;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17373;
	wire [4-1:0] node17374;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17378;
	wire [4-1:0] node17380;
	wire [4-1:0] node17383;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17389;
	wire [4-1:0] node17391;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17397;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17403;
	wire [4-1:0] node17408;
	wire [4-1:0] node17409;
	wire [4-1:0] node17410;
	wire [4-1:0] node17411;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17415;
	wire [4-1:0] node17419;
	wire [4-1:0] node17420;
	wire [4-1:0] node17422;
	wire [4-1:0] node17425;
	wire [4-1:0] node17426;
	wire [4-1:0] node17429;
	wire [4-1:0] node17432;
	wire [4-1:0] node17433;
	wire [4-1:0] node17434;
	wire [4-1:0] node17436;
	wire [4-1:0] node17439;
	wire [4-1:0] node17440;
	wire [4-1:0] node17443;
	wire [4-1:0] node17446;
	wire [4-1:0] node17447;
	wire [4-1:0] node17449;
	wire [4-1:0] node17452;
	wire [4-1:0] node17454;
	wire [4-1:0] node17459;
	wire [4-1:0] node17460;
	wire [4-1:0] node17461;
	wire [4-1:0] node17462;
	wire [4-1:0] node17464;
	wire [4-1:0] node17465;
	wire [4-1:0] node17466;
	wire [4-1:0] node17467;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17470;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17478;
	wire [4-1:0] node17479;
	wire [4-1:0] node17481;
	wire [4-1:0] node17483;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17498;
	wire [4-1:0] node17500;
	wire [4-1:0] node17503;
	wire [4-1:0] node17505;
	wire [4-1:0] node17508;
	wire [4-1:0] node17509;
	wire [4-1:0] node17510;
	wire [4-1:0] node17511;
	wire [4-1:0] node17512;
	wire [4-1:0] node17514;
	wire [4-1:0] node17518;
	wire [4-1:0] node17520;
	wire [4-1:0] node17523;
	wire [4-1:0] node17524;
	wire [4-1:0] node17525;
	wire [4-1:0] node17527;
	wire [4-1:0] node17530;
	wire [4-1:0] node17532;
	wire [4-1:0] node17535;
	wire [4-1:0] node17537;
	wire [4-1:0] node17540;
	wire [4-1:0] node17541;
	wire [4-1:0] node17542;
	wire [4-1:0] node17544;
	wire [4-1:0] node17548;
	wire [4-1:0] node17550;
	wire [4-1:0] node17553;
	wire [4-1:0] node17555;
	wire [4-1:0] node17556;
	wire [4-1:0] node17557;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17561;
	wire [4-1:0] node17566;
	wire [4-1:0] node17567;
	wire [4-1:0] node17568;
	wire [4-1:0] node17571;
	wire [4-1:0] node17572;
	wire [4-1:0] node17576;
	wire [4-1:0] node17578;
	wire [4-1:0] node17580;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17585;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17592;
	wire [4-1:0] node17594;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17599;
	wire [4-1:0] node17603;
	wire [4-1:0] node17605;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17611;
	wire [4-1:0] node17612;
	wire [4-1:0] node17613;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17616;
	wire [4-1:0] node17618;
	wire [4-1:0] node17619;
	wire [4-1:0] node17622;
	wire [4-1:0] node17625;
	wire [4-1:0] node17626;
	wire [4-1:0] node17629;
	wire [4-1:0] node17630;
	wire [4-1:0] node17634;
	wire [4-1:0] node17636;
	wire [4-1:0] node17637;
	wire [4-1:0] node17641;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17644;
	wire [4-1:0] node17648;
	wire [4-1:0] node17649;
	wire [4-1:0] node17653;
	wire [4-1:0] node17654;
	wire [4-1:0] node17655;
	wire [4-1:0] node17656;
	wire [4-1:0] node17660;
	wire [4-1:0] node17662;
	wire [4-1:0] node17665;
	wire [4-1:0] node17666;
	wire [4-1:0] node17669;
	wire [4-1:0] node17671;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17676;
	wire [4-1:0] node17677;
	wire [4-1:0] node17678;
	wire [4-1:0] node17682;
	wire [4-1:0] node17684;
	wire [4-1:0] node17687;
	wire [4-1:0] node17688;
	wire [4-1:0] node17689;
	wire [4-1:0] node17690;
	wire [4-1:0] node17694;
	wire [4-1:0] node17695;
	wire [4-1:0] node17699;
	wire [4-1:0] node17700;
	wire [4-1:0] node17704;
	wire [4-1:0] node17705;
	wire [4-1:0] node17706;
	wire [4-1:0] node17708;
	wire [4-1:0] node17711;
	wire [4-1:0] node17712;
	wire [4-1:0] node17716;
	wire [4-1:0] node17717;
	wire [4-1:0] node17718;
	wire [4-1:0] node17721;
	wire [4-1:0] node17723;
	wire [4-1:0] node17726;
	wire [4-1:0] node17727;
	wire [4-1:0] node17730;
	wire [4-1:0] node17731;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17738;
	wire [4-1:0] node17739;
	wire [4-1:0] node17741;
	wire [4-1:0] node17744;
	wire [4-1:0] node17746;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17751;
	wire [4-1:0] node17755;
	wire [4-1:0] node17757;
	wire [4-1:0] node17760;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17766;
	wire [4-1:0] node17768;
	wire [4-1:0] node17771;
	wire [4-1:0] node17772;
	wire [4-1:0] node17773;
	wire [4-1:0] node17775;
	wire [4-1:0] node17778;
	wire [4-1:0] node17779;
	wire [4-1:0] node17783;
	wire [4-1:0] node17784;
	wire [4-1:0] node17785;
	wire [4-1:0] node17786;
	wire [4-1:0] node17790;
	wire [4-1:0] node17791;
	wire [4-1:0] node17795;
	wire [4-1:0] node17796;
	wire [4-1:0] node17798;
	wire [4-1:0] node17801;
	wire [4-1:0] node17803;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17808;
	wire [4-1:0] node17809;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17813;
	wire [4-1:0] node17816;
	wire [4-1:0] node17817;
	wire [4-1:0] node17821;
	wire [4-1:0] node17822;
	wire [4-1:0] node17825;
	wire [4-1:0] node17827;
	wire [4-1:0] node17830;
	wire [4-1:0] node17831;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17838;
	wire [4-1:0] node17841;
	wire [4-1:0] node17842;
	wire [4-1:0] node17843;
	wire [4-1:0] node17844;
	wire [4-1:0] node17846;
	wire [4-1:0] node17850;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17856;
	wire [4-1:0] node17857;
	wire [4-1:0] node17861;
	wire [4-1:0] node17862;
	wire [4-1:0] node17863;
	wire [4-1:0] node17867;
	wire [4-1:0] node17869;
	wire [4-1:0] node17872;
	wire [4-1:0] node17873;
	wire [4-1:0] node17874;
	wire [4-1:0] node17875;
	wire [4-1:0] node17876;
	wire [4-1:0] node17877;
	wire [4-1:0] node17881;
	wire [4-1:0] node17883;
	wire [4-1:0] node17886;
	wire [4-1:0] node17887;
	wire [4-1:0] node17888;
	wire [4-1:0] node17889;
	wire [4-1:0] node17893;
	wire [4-1:0] node17894;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17900;
	wire [4-1:0] node17904;
	wire [4-1:0] node17906;
	wire [4-1:0] node17909;
	wire [4-1:0] node17910;
	wire [4-1:0] node17911;
	wire [4-1:0] node17912;
	wire [4-1:0] node17916;
	wire [4-1:0] node17918;
	wire [4-1:0] node17921;
	wire [4-1:0] node17922;
	wire [4-1:0] node17923;
	wire [4-1:0] node17925;
	wire [4-1:0] node17928;
	wire [4-1:0] node17929;
	wire [4-1:0] node17933;
	wire [4-1:0] node17935;
	wire [4-1:0] node17937;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17943;
	wire [4-1:0] node17945;
	wire [4-1:0] node17948;
	wire [4-1:0] node17949;
	wire [4-1:0] node17953;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17960;
	wire [4-1:0] node17961;
	wire [4-1:0] node17965;
	wire [4-1:0] node17966;
	wire [4-1:0] node17968;
	wire [4-1:0] node17971;
	wire [4-1:0] node17973;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17978;
	wire [4-1:0] node17979;
	wire [4-1:0] node17982;
	wire [4-1:0] node17983;
	wire [4-1:0] node17987;
	wire [4-1:0] node17988;
	wire [4-1:0] node17989;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17998;
	wire [4-1:0] node17999;
	wire [4-1:0] node18000;
	wire [4-1:0] node18004;
	wire [4-1:0] node18006;
	wire [4-1:0] node18009;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18023;
	wire [4-1:0] node18024;
	wire [4-1:0] node18026;
	wire [4-1:0] node18029;
	wire [4-1:0] node18031;
	wire [4-1:0] node18034;
	wire [4-1:0] node18036;
	wire [4-1:0] node18038;
	wire [4-1:0] node18040;
	wire [4-1:0] node18043;
	wire [4-1:0] node18044;
	wire [4-1:0] node18045;
	wire [4-1:0] node18047;
	wire [4-1:0] node18050;
	wire [4-1:0] node18051;
	wire [4-1:0] node18054;
	wire [4-1:0] node18057;
	wire [4-1:0] node18058;
	wire [4-1:0] node18059;
	wire [4-1:0] node18061;
	wire [4-1:0] node18065;
	wire [4-1:0] node18067;
	wire [4-1:0] node18068;
	wire [4-1:0] node18073;
	wire [4-1:0] node18074;
	wire [4-1:0] node18075;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18079;
	wire [4-1:0] node18080;
	wire [4-1:0] node18084;
	wire [4-1:0] node18085;
	wire [4-1:0] node18089;
	wire [4-1:0] node18090;
	wire [4-1:0] node18092;
	wire [4-1:0] node18093;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18101;
	wire [4-1:0] node18102;
	wire [4-1:0] node18106;
	wire [4-1:0] node18107;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18114;
	wire [4-1:0] node18116;
	wire [4-1:0] node18117;
	wire [4-1:0] node18121;
	wire [4-1:0] node18123;
	wire [4-1:0] node18126;
	wire [4-1:0] node18127;
	wire [4-1:0] node18129;
	wire [4-1:0] node18132;
	wire [4-1:0] node18135;
	wire [4-1:0] node18136;
	wire [4-1:0] node18137;
	wire [4-1:0] node18139;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18148;
	wire [4-1:0] node18149;
	wire [4-1:0] node18150;
	wire [4-1:0] node18151;
	wire [4-1:0] node18152;
	wire [4-1:0] node18153;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18156;
	wire [4-1:0] node18157;
	wire [4-1:0] node18159;
	wire [4-1:0] node18162;
	wire [4-1:0] node18164;
	wire [4-1:0] node18167;
	wire [4-1:0] node18168;
	wire [4-1:0] node18169;
	wire [4-1:0] node18172;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18179;
	wire [4-1:0] node18182;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18186;
	wire [4-1:0] node18189;
	wire [4-1:0] node18190;
	wire [4-1:0] node18193;
	wire [4-1:0] node18196;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18202;
	wire [4-1:0] node18203;
	wire [4-1:0] node18207;
	wire [4-1:0] node18208;
	wire [4-1:0] node18209;
	wire [4-1:0] node18210;
	wire [4-1:0] node18211;
	wire [4-1:0] node18214;
	wire [4-1:0] node18217;
	wire [4-1:0] node18218;
	wire [4-1:0] node18221;
	wire [4-1:0] node18224;
	wire [4-1:0] node18225;
	wire [4-1:0] node18227;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18234;
	wire [4-1:0] node18237;
	wire [4-1:0] node18238;
	wire [4-1:0] node18239;
	wire [4-1:0] node18240;
	wire [4-1:0] node18243;
	wire [4-1:0] node18246;
	wire [4-1:0] node18247;
	wire [4-1:0] node18250;
	wire [4-1:0] node18253;
	wire [4-1:0] node18254;
	wire [4-1:0] node18255;
	wire [4-1:0] node18258;
	wire [4-1:0] node18261;
	wire [4-1:0] node18262;
	wire [4-1:0] node18266;
	wire [4-1:0] node18267;
	wire [4-1:0] node18268;
	wire [4-1:0] node18269;
	wire [4-1:0] node18270;
	wire [4-1:0] node18273;
	wire [4-1:0] node18276;
	wire [4-1:0] node18277;
	wire [4-1:0] node18279;
	wire [4-1:0] node18282;
	wire [4-1:0] node18285;
	wire [4-1:0] node18286;
	wire [4-1:0] node18287;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18296;
	wire [4-1:0] node18299;
	wire [4-1:0] node18300;
	wire [4-1:0] node18304;
	wire [4-1:0] node18305;
	wire [4-1:0] node18306;
	wire [4-1:0] node18307;
	wire [4-1:0] node18311;
	wire [4-1:0] node18312;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18318;
	wire [4-1:0] node18321;
	wire [4-1:0] node18324;
	wire [4-1:0] node18326;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18333;
	wire [4-1:0] node18334;
	wire [4-1:0] node18338;
	wire [4-1:0] node18339;
	wire [4-1:0] node18343;
	wire [4-1:0] node18344;
	wire [4-1:0] node18346;
	wire [4-1:0] node18349;
	wire [4-1:0] node18350;
	wire [4-1:0] node18352;
	wire [4-1:0] node18355;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18364;
	wire [4-1:0] node18366;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18373;
	wire [4-1:0] node18374;
	wire [4-1:0] node18375;
	wire [4-1:0] node18376;
	wire [4-1:0] node18378;
	wire [4-1:0] node18381;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18388;
	wire [4-1:0] node18391;
	wire [4-1:0] node18392;
	wire [4-1:0] node18393;
	wire [4-1:0] node18395;
	wire [4-1:0] node18398;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18404;
	wire [4-1:0] node18405;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18413;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18419;
	wire [4-1:0] node18420;
	wire [4-1:0] node18421;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18427;
	wire [4-1:0] node18429;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18435;
	wire [4-1:0] node18438;
	wire [4-1:0] node18439;
	wire [4-1:0] node18443;
	wire [4-1:0] node18444;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18450;
	wire [4-1:0] node18451;
	wire [4-1:0] node18454;
	wire [4-1:0] node18457;
	wire [4-1:0] node18458;
	wire [4-1:0] node18459;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18474;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18482;
	wire [4-1:0] node18485;
	wire [4-1:0] node18486;
	wire [4-1:0] node18490;
	wire [4-1:0] node18491;
	wire [4-1:0] node18492;
	wire [4-1:0] node18493;
	wire [4-1:0] node18496;
	wire [4-1:0] node18499;
	wire [4-1:0] node18500;
	wire [4-1:0] node18503;
	wire [4-1:0] node18506;
	wire [4-1:0] node18507;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18514;
	wire [4-1:0] node18517;
	wire [4-1:0] node18518;
	wire [4-1:0] node18519;
	wire [4-1:0] node18520;
	wire [4-1:0] node18523;
	wire [4-1:0] node18524;
	wire [4-1:0] node18528;
	wire [4-1:0] node18529;
	wire [4-1:0] node18530;
	wire [4-1:0] node18533;
	wire [4-1:0] node18534;
	wire [4-1:0] node18538;
	wire [4-1:0] node18539;
	wire [4-1:0] node18541;
	wire [4-1:0] node18544;
	wire [4-1:0] node18546;
	wire [4-1:0] node18549;
	wire [4-1:0] node18550;
	wire [4-1:0] node18551;
	wire [4-1:0] node18552;
	wire [4-1:0] node18555;
	wire [4-1:0] node18558;
	wire [4-1:0] node18559;
	wire [4-1:0] node18562;
	wire [4-1:0] node18563;
	wire [4-1:0] node18567;
	wire [4-1:0] node18568;
	wire [4-1:0] node18569;
	wire [4-1:0] node18570;
	wire [4-1:0] node18573;
	wire [4-1:0] node18577;
	wire [4-1:0] node18578;
	wire [4-1:0] node18580;
	wire [4-1:0] node18583;
	wire [4-1:0] node18586;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18589;
	wire [4-1:0] node18590;
	wire [4-1:0] node18591;
	wire [4-1:0] node18594;
	wire [4-1:0] node18597;
	wire [4-1:0] node18598;
	wire [4-1:0] node18601;
	wire [4-1:0] node18604;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18609;
	wire [4-1:0] node18612;
	wire [4-1:0] node18613;
	wire [4-1:0] node18616;
	wire [4-1:0] node18619;
	wire [4-1:0] node18620;
	wire [4-1:0] node18621;
	wire [4-1:0] node18623;
	wire [4-1:0] node18625;
	wire [4-1:0] node18628;
	wire [4-1:0] node18631;
	wire [4-1:0] node18632;
	wire [4-1:0] node18634;
	wire [4-1:0] node18635;
	wire [4-1:0] node18639;
	wire [4-1:0] node18640;
	wire [4-1:0] node18641;
	wire [4-1:0] node18645;
	wire [4-1:0] node18646;
	wire [4-1:0] node18649;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18654;
	wire [4-1:0] node18655;
	wire [4-1:0] node18656;
	wire [4-1:0] node18657;
	wire [4-1:0] node18661;
	wire [4-1:0] node18662;
	wire [4-1:0] node18666;
	wire [4-1:0] node18668;
	wire [4-1:0] node18669;
	wire [4-1:0] node18672;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18679;
	wire [4-1:0] node18682;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18691;
	wire [4-1:0] node18694;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18706;
	wire [4-1:0] node18707;
	wire [4-1:0] node18708;
	wire [4-1:0] node18711;
	wire [4-1:0] node18713;
	wire [4-1:0] node18716;
	wire [4-1:0] node18717;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18726;
	wire [4-1:0] node18727;
	wire [4-1:0] node18729;
	wire [4-1:0] node18733;
	wire [4-1:0] node18734;
	wire [4-1:0] node18735;
	wire [4-1:0] node18739;
	wire [4-1:0] node18740;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18748;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18756;
	wire [4-1:0] node18757;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18765;
	wire [4-1:0] node18766;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18771;
	wire [4-1:0] node18772;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18778;
	wire [4-1:0] node18779;
	wire [4-1:0] node18782;
	wire [4-1:0] node18785;
	wire [4-1:0] node18786;
	wire [4-1:0] node18790;
	wire [4-1:0] node18791;
	wire [4-1:0] node18792;
	wire [4-1:0] node18796;
	wire [4-1:0] node18798;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18803;
	wire [4-1:0] node18804;
	wire [4-1:0] node18807;
	wire [4-1:0] node18810;
	wire [4-1:0] node18811;
	wire [4-1:0] node18814;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18819;
	wire [4-1:0] node18822;
	wire [4-1:0] node18826;
	wire [4-1:0] node18827;
	wire [4-1:0] node18828;
	wire [4-1:0] node18829;
	wire [4-1:0] node18830;
	wire [4-1:0] node18832;
	wire [4-1:0] node18835;
	wire [4-1:0] node18837;
	wire [4-1:0] node18840;
	wire [4-1:0] node18841;
	wire [4-1:0] node18843;
	wire [4-1:0] node18846;
	wire [4-1:0] node18847;
	wire [4-1:0] node18850;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18859;
	wire [4-1:0] node18861;
	wire [4-1:0] node18862;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18870;
	wire [4-1:0] node18873;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18879;
	wire [4-1:0] node18881;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18886;
	wire [4-1:0] node18888;
	wire [4-1:0] node18891;
	wire [4-1:0] node18893;
	wire [4-1:0] node18896;
	wire [4-1:0] node18897;
	wire [4-1:0] node18900;
	wire [4-1:0] node18901;
	wire [4-1:0] node18904;
	wire [4-1:0] node18907;
	wire [4-1:0] node18908;
	wire [4-1:0] node18909;
	wire [4-1:0] node18910;
	wire [4-1:0] node18911;
	wire [4-1:0] node18912;
	wire [4-1:0] node18913;
	wire [4-1:0] node18916;
	wire [4-1:0] node18919;
	wire [4-1:0] node18921;
	wire [4-1:0] node18924;
	wire [4-1:0] node18925;
	wire [4-1:0] node18926;
	wire [4-1:0] node18928;
	wire [4-1:0] node18931;
	wire [4-1:0] node18932;
	wire [4-1:0] node18935;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18943;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18948;
	wire [4-1:0] node18949;
	wire [4-1:0] node18953;
	wire [4-1:0] node18954;
	wire [4-1:0] node18955;
	wire [4-1:0] node18958;
	wire [4-1:0] node18961;
	wire [4-1:0] node18962;
	wire [4-1:0] node18965;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18970;
	wire [4-1:0] node18971;
	wire [4-1:0] node18973;
	wire [4-1:0] node18976;
	wire [4-1:0] node18977;
	wire [4-1:0] node18981;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18984;
	wire [4-1:0] node18987;
	wire [4-1:0] node18990;
	wire [4-1:0] node18991;
	wire [4-1:0] node18994;
	wire [4-1:0] node18997;
	wire [4-1:0] node18999;
	wire [4-1:0] node19002;
	wire [4-1:0] node19003;
	wire [4-1:0] node19004;
	wire [4-1:0] node19005;
	wire [4-1:0] node19008;
	wire [4-1:0] node19011;
	wire [4-1:0] node19012;
	wire [4-1:0] node19015;
	wire [4-1:0] node19018;
	wire [4-1:0] node19019;
	wire [4-1:0] node19020;
	wire [4-1:0] node19024;
	wire [4-1:0] node19025;
	wire [4-1:0] node19028;
	wire [4-1:0] node19031;
	wire [4-1:0] node19032;
	wire [4-1:0] node19033;
	wire [4-1:0] node19034;
	wire [4-1:0] node19035;
	wire [4-1:0] node19036;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19044;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19052;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19056;
	wire [4-1:0] node19059;
	wire [4-1:0] node19062;
	wire [4-1:0] node19063;
	wire [4-1:0] node19064;
	wire [4-1:0] node19068;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19075;
	wire [4-1:0] node19078;
	wire [4-1:0] node19079;
	wire [4-1:0] node19080;
	wire [4-1:0] node19083;
	wire [4-1:0] node19086;
	wire [4-1:0] node19087;
	wire [4-1:0] node19088;
	wire [4-1:0] node19091;
	wire [4-1:0] node19094;
	wire [4-1:0] node19095;
	wire [4-1:0] node19099;
	wire [4-1:0] node19100;
	wire [4-1:0] node19104;
	wire [4-1:0] node19105;
	wire [4-1:0] node19106;
	wire [4-1:0] node19107;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19113;
	wire [4-1:0] node19117;
	wire [4-1:0] node19120;
	wire [4-1:0] node19121;
	wire [4-1:0] node19124;
	wire [4-1:0] node19125;
	wire [4-1:0] node19129;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19132;
	wire [4-1:0] node19136;
	wire [4-1:0] node19138;
	wire [4-1:0] node19141;
	wire [4-1:0] node19142;
	wire [4-1:0] node19143;
	wire [4-1:0] node19146;
	wire [4-1:0] node19149;
	wire [4-1:0] node19151;
	wire [4-1:0] node19154;
	wire [4-1:0] node19155;
	wire [4-1:0] node19156;
	wire [4-1:0] node19159;
	wire [4-1:0] node19160;
	wire [4-1:0] node19161;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19169;
	wire [4-1:0] node19173;
	wire [4-1:0] node19176;
	wire [4-1:0] node19177;
	wire [4-1:0] node19180;
	wire [4-1:0] node19181;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19187;
	wire [4-1:0] node19188;
	wire [4-1:0] node19189;
	wire [4-1:0] node19193;
	wire [4-1:0] node19195;
	wire [4-1:0] node19198;
	wire [4-1:0] node19200;
	wire [4-1:0] node19201;
	wire [4-1:0] node19205;
	wire [4-1:0] node19206;
	wire [4-1:0] node19207;
	wire [4-1:0] node19208;
	wire [4-1:0] node19211;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19219;
	wire [4-1:0] node19223;
	wire [4-1:0] node19224;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19229;
	wire [4-1:0] node19232;
	wire [4-1:0] node19235;
	wire [4-1:0] node19236;
	wire [4-1:0] node19238;
	wire [4-1:0] node19241;
	wire [4-1:0] node19244;
	wire [4-1:0] node19245;
	wire [4-1:0] node19246;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19252;
	wire [4-1:0] node19255;
	wire [4-1:0] node19256;
	wire [4-1:0] node19260;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19269;
	wire [4-1:0] node19270;
	wire [4-1:0] node19273;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19281;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19284;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19291;
	wire [4-1:0] node19294;
	wire [4-1:0] node19297;
	wire [4-1:0] node19298;
	wire [4-1:0] node19301;
	wire [4-1:0] node19304;
	wire [4-1:0] node19305;
	wire [4-1:0] node19306;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19316;
	wire [4-1:0] node19319;
	wire [4-1:0] node19320;
	wire [4-1:0] node19321;
	wire [4-1:0] node19325;
	wire [4-1:0] node19328;
	wire [4-1:0] node19329;
	wire [4-1:0] node19331;
	wire [4-1:0] node19334;
	wire [4-1:0] node19336;
	wire [4-1:0] node19339;
	wire [4-1:0] node19340;
	wire [4-1:0] node19341;
	wire [4-1:0] node19342;
	wire [4-1:0] node19343;
	wire [4-1:0] node19344;
	wire [4-1:0] node19345;
	wire [4-1:0] node19347;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19354;
	wire [4-1:0] node19358;
	wire [4-1:0] node19359;
	wire [4-1:0] node19361;
	wire [4-1:0] node19364;
	wire [4-1:0] node19367;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19373;
	wire [4-1:0] node19374;
	wire [4-1:0] node19378;
	wire [4-1:0] node19379;
	wire [4-1:0] node19382;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19388;
	wire [4-1:0] node19392;
	wire [4-1:0] node19393;
	wire [4-1:0] node19394;
	wire [4-1:0] node19395;
	wire [4-1:0] node19397;
	wire [4-1:0] node19399;
	wire [4-1:0] node19402;
	wire [4-1:0] node19404;
	wire [4-1:0] node19406;
	wire [4-1:0] node19409;
	wire [4-1:0] node19410;
	wire [4-1:0] node19411;
	wire [4-1:0] node19413;
	wire [4-1:0] node19416;
	wire [4-1:0] node19419;
	wire [4-1:0] node19421;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19429;
	wire [4-1:0] node19432;
	wire [4-1:0] node19436;
	wire [4-1:0] node19437;
	wire [4-1:0] node19438;
	wire [4-1:0] node19439;
	wire [4-1:0] node19442;
	wire [4-1:0] node19445;
	wire [4-1:0] node19448;
	wire [4-1:0] node19449;
	wire [4-1:0] node19450;
	wire [4-1:0] node19453;
	wire [4-1:0] node19457;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19461;
	wire [4-1:0] node19462;
	wire [4-1:0] node19463;
	wire [4-1:0] node19467;
	wire [4-1:0] node19468;
	wire [4-1:0] node19471;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19478;
	wire [4-1:0] node19481;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19486;
	wire [4-1:0] node19487;
	wire [4-1:0] node19492;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19496;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19504;
	wire [4-1:0] node19505;
	wire [4-1:0] node19506;
	wire [4-1:0] node19508;
	wire [4-1:0] node19511;
	wire [4-1:0] node19514;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19524;
	wire [4-1:0] node19525;
	wire [4-1:0] node19529;
	wire [4-1:0] node19530;
	wire [4-1:0] node19534;
	wire [4-1:0] node19535;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19541;
	wire [4-1:0] node19543;
	wire [4-1:0] node19546;
	wire [4-1:0] node19547;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19556;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19559;
	wire [4-1:0] node19560;
	wire [4-1:0] node19565;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19572;
	wire [4-1:0] node19573;
	wire [4-1:0] node19575;
	wire [4-1:0] node19576;
	wire [4-1:0] node19580;
	wire [4-1:0] node19581;
	wire [4-1:0] node19582;
	wire [4-1:0] node19585;
	wire [4-1:0] node19588;
	wire [4-1:0] node19590;
	wire [4-1:0] node19593;
	wire [4-1:0] node19594;
	wire [4-1:0] node19595;
	wire [4-1:0] node19598;
	wire [4-1:0] node19600;
	wire [4-1:0] node19603;
	wire [4-1:0] node19604;
	wire [4-1:0] node19605;
	wire [4-1:0] node19606;
	wire [4-1:0] node19611;
	wire [4-1:0] node19612;
	wire [4-1:0] node19614;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19620;
	wire [4-1:0] node19621;
	wire [4-1:0] node19622;
	wire [4-1:0] node19625;
	wire [4-1:0] node19626;
	wire [4-1:0] node19629;
	wire [4-1:0] node19632;
	wire [4-1:0] node19633;
	wire [4-1:0] node19634;
	wire [4-1:0] node19638;
	wire [4-1:0] node19641;
	wire [4-1:0] node19642;
	wire [4-1:0] node19643;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19654;
	wire [4-1:0] node19655;
	wire [4-1:0] node19656;
	wire [4-1:0] node19657;
	wire [4-1:0] node19660;
	wire [4-1:0] node19663;
	wire [4-1:0] node19665;
	wire [4-1:0] node19668;
	wire [4-1:0] node19669;
	wire [4-1:0] node19670;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19678;
	wire [4-1:0] node19681;
	wire [4-1:0] node19682;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19686;
	wire [4-1:0] node19689;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19697;
	wire [4-1:0] node19700;
	wire [4-1:0] node19701;
	wire [4-1:0] node19704;
	wire [4-1:0] node19707;
	wire [4-1:0] node19708;
	wire [4-1:0] node19709;
	wire [4-1:0] node19712;
	wire [4-1:0] node19715;
	wire [4-1:0] node19716;
	wire [4-1:0] node19717;
	wire [4-1:0] node19721;
	wire [4-1:0] node19724;
	wire [4-1:0] node19725;
	wire [4-1:0] node19726;
	wire [4-1:0] node19728;
	wire [4-1:0] node19731;
	wire [4-1:0] node19733;
	wire [4-1:0] node19736;
	wire [4-1:0] node19737;
	wire [4-1:0] node19740;
	wire [4-1:0] node19741;
	wire [4-1:0] node19742;
	wire [4-1:0] node19747;
	wire [4-1:0] node19748;
	wire [4-1:0] node19749;
	wire [4-1:0] node19750;
	wire [4-1:0] node19751;
	wire [4-1:0] node19755;
	wire [4-1:0] node19757;
	wire [4-1:0] node19759;
	wire [4-1:0] node19762;
	wire [4-1:0] node19763;
	wire [4-1:0] node19764;
	wire [4-1:0] node19767;
	wire [4-1:0] node19770;
	wire [4-1:0] node19771;
	wire [4-1:0] node19774;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19779;
	wire [4-1:0] node19781;
	wire [4-1:0] node19783;
	wire [4-1:0] node19786;
	wire [4-1:0] node19787;
	wire [4-1:0] node19789;
	wire [4-1:0] node19792;
	wire [4-1:0] node19794;
	wire [4-1:0] node19798;
	wire [4-1:0] node19799;
	wire [4-1:0] node19800;
	wire [4-1:0] node19801;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19804;
	wire [4-1:0] node19807;
	wire [4-1:0] node19809;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19815;
	wire [4-1:0] node19818;
	wire [4-1:0] node19820;
	wire [4-1:0] node19823;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19826;
	wire [4-1:0] node19830;
	wire [4-1:0] node19831;
	wire [4-1:0] node19835;
	wire [4-1:0] node19836;
	wire [4-1:0] node19838;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19845;
	wire [4-1:0] node19848;
	wire [4-1:0] node19849;
	wire [4-1:0] node19851;
	wire [4-1:0] node19852;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19859;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19864;
	wire [4-1:0] node19867;
	wire [4-1:0] node19868;
	wire [4-1:0] node19871;
	wire [4-1:0] node19874;
	wire [4-1:0] node19876;
	wire [4-1:0] node19878;
	wire [4-1:0] node19881;
	wire [4-1:0] node19882;
	wire [4-1:0] node19883;
	wire [4-1:0] node19884;
	wire [4-1:0] node19888;
	wire [4-1:0] node19889;
	wire [4-1:0] node19892;
	wire [4-1:0] node19896;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19899;
	wire [4-1:0] node19900;
	wire [4-1:0] node19901;
	wire [4-1:0] node19904;
	wire [4-1:0] node19906;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19912;
	wire [4-1:0] node19915;
	wire [4-1:0] node19918;
	wire [4-1:0] node19919;
	wire [4-1:0] node19921;
	wire [4-1:0] node19924;
	wire [4-1:0] node19925;
	wire [4-1:0] node19928;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19933;
	wire [4-1:0] node19935;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19942;
	wire [4-1:0] node19946;
	wire [4-1:0] node19948;
	wire [4-1:0] node19949;
	wire [4-1:0] node19950;
	wire [4-1:0] node19951;
	wire [4-1:0] node19952;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19963;
	wire [4-1:0] node19965;
	wire [4-1:0] node19966;
	wire [4-1:0] node19968;
	wire [4-1:0] node19969;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19975;
	wire [4-1:0] node19976;
	wire [4-1:0] node19977;
	wire [4-1:0] node19982;
	wire [4-1:0] node19983;
	wire [4-1:0] node19984;
	wire [4-1:0] node19985;
	wire [4-1:0] node19989;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node19999;
	wire [4-1:0] node20000;
	wire [4-1:0] node20003;
	wire [4-1:0] node20005;
	wire [4-1:0] node20008;
	wire [4-1:0] node20010;
	wire [4-1:0] node20013;
	wire [4-1:0] node20014;
	wire [4-1:0] node20015;
	wire [4-1:0] node20016;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20025;
	wire [4-1:0] node20027;
	wire [4-1:0] node20031;
	wire [4-1:0] node20032;
	wire [4-1:0] node20033;
	wire [4-1:0] node20034;
	wire [4-1:0] node20035;
	wire [4-1:0] node20036;
	wire [4-1:0] node20038;
	wire [4-1:0] node20042;
	wire [4-1:0] node20044;
	wire [4-1:0] node20047;
	wire [4-1:0] node20048;
	wire [4-1:0] node20049;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20056;
	wire [4-1:0] node20057;
	wire [4-1:0] node20061;
	wire [4-1:0] node20062;
	wire [4-1:0] node20066;
	wire [4-1:0] node20067;
	wire [4-1:0] node20071;
	wire [4-1:0] node20072;
	wire [4-1:0] node20073;
	wire [4-1:0] node20075;
	wire [4-1:0] node20078;
	wire [4-1:0] node20079;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20085;
	wire [4-1:0] node20086;
	wire [4-1:0] node20087;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20097;
	wire [4-1:0] node20098;
	wire [4-1:0] node20099;
	wire [4-1:0] node20103;
	wire [4-1:0] node20105;
	wire [4-1:0] node20109;
	wire [4-1:0] node20110;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20113;
	wire [4-1:0] node20114;
	wire [4-1:0] node20115;
	wire [4-1:0] node20116;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20123;
	wire [4-1:0] node20126;
	wire [4-1:0] node20127;
	wire [4-1:0] node20129;
	wire [4-1:0] node20132;
	wire [4-1:0] node20133;
	wire [4-1:0] node20137;
	wire [4-1:0] node20138;
	wire [4-1:0] node20139;
	wire [4-1:0] node20140;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20148;
	wire [4-1:0] node20149;
	wire [4-1:0] node20150;
	wire [4-1:0] node20153;
	wire [4-1:0] node20156;
	wire [4-1:0] node20159;
	wire [4-1:0] node20160;
	wire [4-1:0] node20161;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20167;
	wire [4-1:0] node20170;
	wire [4-1:0] node20173;
	wire [4-1:0] node20176;
	wire [4-1:0] node20177;
	wire [4-1:0] node20178;
	wire [4-1:0] node20179;
	wire [4-1:0] node20181;
	wire [4-1:0] node20184;
	wire [4-1:0] node20187;
	wire [4-1:0] node20188;
	wire [4-1:0] node20189;
	wire [4-1:0] node20192;
	wire [4-1:0] node20193;
	wire [4-1:0] node20197;
	wire [4-1:0] node20198;
	wire [4-1:0] node20202;
	wire [4-1:0] node20203;
	wire [4-1:0] node20204;
	wire [4-1:0] node20206;
	wire [4-1:0] node20210;
	wire [4-1:0] node20211;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20218;
	wire [4-1:0] node20221;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20227;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20235;
	wire [4-1:0] node20238;
	wire [4-1:0] node20239;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20245;
	wire [4-1:0] node20246;
	wire [4-1:0] node20249;
	wire [4-1:0] node20252;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20259;
	wire [4-1:0] node20260;
	wire [4-1:0] node20262;
	wire [4-1:0] node20265;
	wire [4-1:0] node20267;
	wire [4-1:0] node20270;
	wire [4-1:0] node20271;
	wire [4-1:0] node20272;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20279;
	wire [4-1:0] node20280;
	wire [4-1:0] node20281;
	wire [4-1:0] node20284;
	wire [4-1:0] node20287;
	wire [4-1:0] node20289;
	wire [4-1:0] node20292;
	wire [4-1:0] node20293;
	wire [4-1:0] node20295;
	wire [4-1:0] node20297;
	wire [4-1:0] node20300;
	wire [4-1:0] node20302;
	wire [4-1:0] node20303;
	wire [4-1:0] node20307;
	wire [4-1:0] node20308;
	wire [4-1:0] node20309;
	wire [4-1:0] node20310;
	wire [4-1:0] node20311;
	wire [4-1:0] node20314;
	wire [4-1:0] node20317;
	wire [4-1:0] node20318;
	wire [4-1:0] node20321;
	wire [4-1:0] node20324;
	wire [4-1:0] node20325;
	wire [4-1:0] node20327;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20336;
	wire [4-1:0] node20339;
	wire [4-1:0] node20340;
	wire [4-1:0] node20344;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20347;
	wire [4-1:0] node20348;
	wire [4-1:0] node20349;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20356;
	wire [4-1:0] node20359;
	wire [4-1:0] node20360;
	wire [4-1:0] node20362;
	wire [4-1:0] node20363;
	wire [4-1:0] node20366;
	wire [4-1:0] node20369;
	wire [4-1:0] node20370;
	wire [4-1:0] node20372;
	wire [4-1:0] node20375;
	wire [4-1:0] node20378;
	wire [4-1:0] node20379;
	wire [4-1:0] node20380;
	wire [4-1:0] node20381;
	wire [4-1:0] node20382;
	wire [4-1:0] node20386;
	wire [4-1:0] node20388;
	wire [4-1:0] node20391;
	wire [4-1:0] node20393;
	wire [4-1:0] node20394;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20402;
	wire [4-1:0] node20405;
	wire [4-1:0] node20407;
	wire [4-1:0] node20410;
	wire [4-1:0] node20411;
	wire [4-1:0] node20413;
	wire [4-1:0] node20416;
	wire [4-1:0] node20419;
	wire [4-1:0] node20420;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20423;
	wire [4-1:0] node20427;
	wire [4-1:0] node20428;
	wire [4-1:0] node20429;
	wire [4-1:0] node20432;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20439;
	wire [4-1:0] node20442;
	wire [4-1:0] node20444;
	wire [4-1:0] node20445;
	wire [4-1:0] node20446;
	wire [4-1:0] node20450;
	wire [4-1:0] node20451;
	wire [4-1:0] node20455;
	wire [4-1:0] node20456;
	wire [4-1:0] node20457;
	wire [4-1:0] node20458;
	wire [4-1:0] node20463;
	wire [4-1:0] node20464;
	wire [4-1:0] node20466;
	wire [4-1:0] node20470;
	wire [4-1:0] node20471;
	wire [4-1:0] node20472;
	wire [4-1:0] node20473;
	wire [4-1:0] node20474;
	wire [4-1:0] node20475;
	wire [4-1:0] node20477;
	wire [4-1:0] node20480;
	wire [4-1:0] node20481;
	wire [4-1:0] node20484;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20493;
	wire [4-1:0] node20494;
	wire [4-1:0] node20497;
	wire [4-1:0] node20500;
	wire [4-1:0] node20501;
	wire [4-1:0] node20502;
	wire [4-1:0] node20504;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20511;
	wire [4-1:0] node20514;
	wire [4-1:0] node20515;
	wire [4-1:0] node20517;
	wire [4-1:0] node20520;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20527;
	wire [4-1:0] node20531;
	wire [4-1:0] node20533;
	wire [4-1:0] node20536;
	wire [4-1:0] node20537;
	wire [4-1:0] node20538;
	wire [4-1:0] node20541;
	wire [4-1:0] node20545;
	wire [4-1:0] node20546;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20556;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20565;
	wire [4-1:0] node20566;
	wire [4-1:0] node20567;
	wire [4-1:0] node20573;
	wire [4-1:0] node20575;
	wire [4-1:0] node20576;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20582;
	wire [4-1:0] node20584;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20590;
	wire [4-1:0] node20593;
	wire [4-1:0] node20595;
	wire [4-1:0] node20598;
	wire [4-1:0] node20600;
	wire [4-1:0] node20602;
	wire [4-1:0] node20604;
	wire [4-1:0] node20607;
	wire [4-1:0] node20608;
	wire [4-1:0] node20609;
	wire [4-1:0] node20611;
	wire [4-1:0] node20613;
	wire [4-1:0] node20616;
	wire [4-1:0] node20618;
	wire [4-1:0] node20619;
	wire [4-1:0] node20623;
	wire [4-1:0] node20624;
	wire [4-1:0] node20625;
	wire [4-1:0] node20629;
	wire [4-1:0] node20630;
	wire [4-1:0] node20631;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20639;
	wire [4-1:0] node20640;
	wire [4-1:0] node20641;
	wire [4-1:0] node20642;
	wire [4-1:0] node20643;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20654;
	wire [4-1:0] node20655;
	wire [4-1:0] node20659;
	wire [4-1:0] node20662;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20665;
	wire [4-1:0] node20667;
	wire [4-1:0] node20670;
	wire [4-1:0] node20672;
	wire [4-1:0] node20675;
	wire [4-1:0] node20676;
	wire [4-1:0] node20677;
	wire [4-1:0] node20680;
	wire [4-1:0] node20683;
	wire [4-1:0] node20685;
	wire [4-1:0] node20688;
	wire [4-1:0] node20690;
	wire [4-1:0] node20692;
	wire [4-1:0] node20695;
	wire [4-1:0] node20696;
	wire [4-1:0] node20697;
	wire [4-1:0] node20698;
	wire [4-1:0] node20700;
	wire [4-1:0] node20701;
	wire [4-1:0] node20704;
	wire [4-1:0] node20707;
	wire [4-1:0] node20708;
	wire [4-1:0] node20710;
	wire [4-1:0] node20713;
	wire [4-1:0] node20714;
	wire [4-1:0] node20717;
	wire [4-1:0] node20720;
	wire [4-1:0] node20721;
	wire [4-1:0] node20722;
	wire [4-1:0] node20723;
	wire [4-1:0] node20727;
	wire [4-1:0] node20731;
	wire [4-1:0] node20732;
	wire [4-1:0] node20734;
	wire [4-1:0] node20735;
	wire [4-1:0] node20740;
	wire [4-1:0] node20741;
	wire [4-1:0] node20742;
	wire [4-1:0] node20743;
	wire [4-1:0] node20744;
	wire [4-1:0] node20745;
	wire [4-1:0] node20746;
	wire [4-1:0] node20747;
	wire [4-1:0] node20748;
	wire [4-1:0] node20750;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20754;
	wire [4-1:0] node20755;
	wire [4-1:0] node20760;
	wire [4-1:0] node20761;
	wire [4-1:0] node20762;
	wire [4-1:0] node20764;
	wire [4-1:0] node20767;
	wire [4-1:0] node20769;
	wire [4-1:0] node20772;
	wire [4-1:0] node20774;
	wire [4-1:0] node20775;
	wire [4-1:0] node20780;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20783;
	wire [4-1:0] node20784;
	wire [4-1:0] node20785;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20792;
	wire [4-1:0] node20795;
	wire [4-1:0] node20797;
	wire [4-1:0] node20800;
	wire [4-1:0] node20801;
	wire [4-1:0] node20802;
	wire [4-1:0] node20804;
	wire [4-1:0] node20807;
	wire [4-1:0] node20808;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20817;
	wire [4-1:0] node20818;
	wire [4-1:0] node20819;
	wire [4-1:0] node20821;
	wire [4-1:0] node20824;
	wire [4-1:0] node20825;
	wire [4-1:0] node20829;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20833;
	wire [4-1:0] node20836;
	wire [4-1:0] node20838;
	wire [4-1:0] node20841;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20847;
	wire [4-1:0] node20849;
	wire [4-1:0] node20852;
	wire [4-1:0] node20854;
	wire [4-1:0] node20855;
	wire [4-1:0] node20856;
	wire [4-1:0] node20860;
	wire [4-1:0] node20861;
	wire [4-1:0] node20862;
	wire [4-1:0] node20865;
	wire [4-1:0] node20866;
	wire [4-1:0] node20870;
	wire [4-1:0] node20872;
	wire [4-1:0] node20873;
	wire [4-1:0] node20877;
	wire [4-1:0] node20878;
	wire [4-1:0] node20879;
	wire [4-1:0] node20880;
	wire [4-1:0] node20881;
	wire [4-1:0] node20883;
	wire [4-1:0] node20886;
	wire [4-1:0] node20887;
	wire [4-1:0] node20889;
	wire [4-1:0] node20892;
	wire [4-1:0] node20893;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20899;
	wire [4-1:0] node20901;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20907;
	wire [4-1:0] node20910;
	wire [4-1:0] node20912;
	wire [4-1:0] node20915;
	wire [4-1:0] node20917;
	wire [4-1:0] node20920;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20923;
	wire [4-1:0] node20925;
	wire [4-1:0] node20928;
	wire [4-1:0] node20929;
	wire [4-1:0] node20930;
	wire [4-1:0] node20934;
	wire [4-1:0] node20937;
	wire [4-1:0] node20938;
	wire [4-1:0] node20940;
	wire [4-1:0] node20943;
	wire [4-1:0] node20945;
	wire [4-1:0] node20946;
	wire [4-1:0] node20950;
	wire [4-1:0] node20951;
	wire [4-1:0] node20952;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20959;
	wire [4-1:0] node20962;
	wire [4-1:0] node20963;
	wire [4-1:0] node20967;
	wire [4-1:0] node20968;
	wire [4-1:0] node20969;
	wire [4-1:0] node20970;
	wire [4-1:0] node20971;
	wire [4-1:0] node20972;
	wire [4-1:0] node20974;
	wire [4-1:0] node20977;
	wire [4-1:0] node20978;
	wire [4-1:0] node20982;
	wire [4-1:0] node20983;
	wire [4-1:0] node20985;
	wire [4-1:0] node20988;
	wire [4-1:0] node20990;
	wire [4-1:0] node20993;
	wire [4-1:0] node20994;
	wire [4-1:0] node20996;
	wire [4-1:0] node20999;
	wire [4-1:0] node21001;
	wire [4-1:0] node21004;
	wire [4-1:0] node21005;
	wire [4-1:0] node21006;
	wire [4-1:0] node21007;
	wire [4-1:0] node21008;
	wire [4-1:0] node21012;
	wire [4-1:0] node21015;
	wire [4-1:0] node21016;
	wire [4-1:0] node21017;
	wire [4-1:0] node21021;
	wire [4-1:0] node21022;
	wire [4-1:0] node21026;
	wire [4-1:0] node21027;
	wire [4-1:0] node21029;
	wire [4-1:0] node21032;
	wire [4-1:0] node21033;
	wire [4-1:0] node21037;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21040;
	wire [4-1:0] node21041;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21050;
	wire [4-1:0] node21051;
	wire [4-1:0] node21052;
	wire [4-1:0] node21053;
	wire [4-1:0] node21057;
	wire [4-1:0] node21059;
	wire [4-1:0] node21062;
	wire [4-1:0] node21064;
	wire [4-1:0] node21067;
	wire [4-1:0] node21068;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21074;
	wire [4-1:0] node21076;
	wire [4-1:0] node21079;
	wire [4-1:0] node21080;
	wire [4-1:0] node21081;
	wire [4-1:0] node21085;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21091;
	wire [4-1:0] node21092;
	wire [4-1:0] node21097;
	wire [4-1:0] node21098;
	wire [4-1:0] node21099;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21105;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21111;
	wire [4-1:0] node21114;
	wire [4-1:0] node21115;
	wire [4-1:0] node21119;
	wire [4-1:0] node21120;
	wire [4-1:0] node21121;
	wire [4-1:0] node21123;
	wire [4-1:0] node21126;
	wire [4-1:0] node21127;
	wire [4-1:0] node21128;
	wire [4-1:0] node21132;
	wire [4-1:0] node21133;
	wire [4-1:0] node21137;
	wire [4-1:0] node21139;
	wire [4-1:0] node21142;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21146;
	wire [4-1:0] node21149;
	wire [4-1:0] node21150;
	wire [4-1:0] node21152;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21160;
	wire [4-1:0] node21161;
	wire [4-1:0] node21162;
	wire [4-1:0] node21164;
	wire [4-1:0] node21168;
	wire [4-1:0] node21169;
	wire [4-1:0] node21171;
	wire [4-1:0] node21174;
	wire [4-1:0] node21175;
	wire [4-1:0] node21177;
	wire [4-1:0] node21180;
	wire [4-1:0] node21183;
	wire [4-1:0] node21184;
	wire [4-1:0] node21185;
	wire [4-1:0] node21186;
	wire [4-1:0] node21187;
	wire [4-1:0] node21189;
	wire [4-1:0] node21190;
	wire [4-1:0] node21194;
	wire [4-1:0] node21196;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21211;
	wire [4-1:0] node21213;
	wire [4-1:0] node21216;
	wire [4-1:0] node21217;
	wire [4-1:0] node21218;
	wire [4-1:0] node21219;
	wire [4-1:0] node21223;
	wire [4-1:0] node21224;
	wire [4-1:0] node21228;
	wire [4-1:0] node21229;
	wire [4-1:0] node21230;
	wire [4-1:0] node21232;
	wire [4-1:0] node21235;
	wire [4-1:0] node21238;
	wire [4-1:0] node21239;
	wire [4-1:0] node21243;
	wire [4-1:0] node21244;
	wire [4-1:0] node21245;
	wire [4-1:0] node21246;
	wire [4-1:0] node21247;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21254;
	wire [4-1:0] node21258;
	wire [4-1:0] node21259;
	wire [4-1:0] node21260;
	wire [4-1:0] node21262;
	wire [4-1:0] node21265;
	wire [4-1:0] node21266;
	wire [4-1:0] node21270;
	wire [4-1:0] node21272;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21280;
	wire [4-1:0] node21283;
	wire [4-1:0] node21285;
	wire [4-1:0] node21289;
	wire [4-1:0] node21290;
	wire [4-1:0] node21291;
	wire [4-1:0] node21295;
	wire [4-1:0] node21296;
	wire [4-1:0] node21299;
	wire [4-1:0] node21300;
	wire [4-1:0] node21304;
	wire [4-1:0] node21305;
	wire [4-1:0] node21306;
	wire [4-1:0] node21308;
	wire [4-1:0] node21309;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21314;
	wire [4-1:0] node21318;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21325;
	wire [4-1:0] node21327;
	wire [4-1:0] node21330;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21337;
	wire [4-1:0] node21338;
	wire [4-1:0] node21339;
	wire [4-1:0] node21340;
	wire [4-1:0] node21342;
	wire [4-1:0] node21345;
	wire [4-1:0] node21346;
	wire [4-1:0] node21348;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21356;
	wire [4-1:0] node21357;
	wire [4-1:0] node21359;
	wire [4-1:0] node21362;
	wire [4-1:0] node21364;
	wire [4-1:0] node21366;
	wire [4-1:0] node21369;
	wire [4-1:0] node21370;
	wire [4-1:0] node21371;
	wire [4-1:0] node21372;
	wire [4-1:0] node21373;
	wire [4-1:0] node21377;
	wire [4-1:0] node21380;
	wire [4-1:0] node21381;
	wire [4-1:0] node21384;
	wire [4-1:0] node21386;
	wire [4-1:0] node21389;
	wire [4-1:0] node21390;
	wire [4-1:0] node21391;
	wire [4-1:0] node21395;
	wire [4-1:0] node21397;
	wire [4-1:0] node21400;
	wire [4-1:0] node21402;
	wire [4-1:0] node21404;
	wire [4-1:0] node21405;
	wire [4-1:0] node21407;
	wire [4-1:0] node21410;
	wire [4-1:0] node21411;
	wire [4-1:0] node21412;
	wire [4-1:0] node21416;
	wire [4-1:0] node21418;
	wire [4-1:0] node21421;
	wire [4-1:0] node21422;
	wire [4-1:0] node21423;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21428;
	wire [4-1:0] node21431;
	wire [4-1:0] node21433;
	wire [4-1:0] node21436;
	wire [4-1:0] node21438;
	wire [4-1:0] node21441;
	wire [4-1:0] node21442;
	wire [4-1:0] node21443;
	wire [4-1:0] node21444;
	wire [4-1:0] node21448;
	wire [4-1:0] node21449;
	wire [4-1:0] node21450;
	wire [4-1:0] node21454;
	wire [4-1:0] node21455;
	wire [4-1:0] node21459;
	wire [4-1:0] node21460;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21466;
	wire [4-1:0] node21467;
	wire [4-1:0] node21469;
	wire [4-1:0] node21472;
	wire [4-1:0] node21473;
	wire [4-1:0] node21475;
	wire [4-1:0] node21478;
	wire [4-1:0] node21479;
	wire [4-1:0] node21483;
	wire [4-1:0] node21484;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21491;
	wire [4-1:0] node21493;
	wire [4-1:0] node21496;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21500;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21506;
	wire [4-1:0] node21509;
	wire [4-1:0] node21510;
	wire [4-1:0] node21514;
	wire [4-1:0] node21515;
	wire [4-1:0] node21516;
	wire [4-1:0] node21520;
	wire [4-1:0] node21521;
	wire [4-1:0] node21522;
	wire [4-1:0] node21526;
	wire [4-1:0] node21527;
	wire [4-1:0] node21531;
	wire [4-1:0] node21532;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21535;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21543;
	wire [4-1:0] node21546;
	wire [4-1:0] node21547;
	wire [4-1:0] node21551;
	wire [4-1:0] node21552;
	wire [4-1:0] node21553;
	wire [4-1:0] node21555;
	wire [4-1:0] node21559;
	wire [4-1:0] node21561;
	wire [4-1:0] node21563;
	wire [4-1:0] node21566;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21569;
	wire [4-1:0] node21573;
	wire [4-1:0] node21574;
	wire [4-1:0] node21575;
	wire [4-1:0] node21579;
	wire [4-1:0] node21580;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21587;
	wire [4-1:0] node21590;
	wire [4-1:0] node21591;
	wire [4-1:0] node21592;
	wire [4-1:0] node21596;
	wire [4-1:0] node21597;
	wire [4-1:0] node21601;
	wire [4-1:0] node21602;
	wire [4-1:0] node21603;
	wire [4-1:0] node21604;
	wire [4-1:0] node21605;
	wire [4-1:0] node21609;
	wire [4-1:0] node21610;
	wire [4-1:0] node21614;
	wire [4-1:0] node21616;
	wire [4-1:0] node21619;
	wire [4-1:0] node21620;
	wire [4-1:0] node21621;
	wire [4-1:0] node21623;
	wire [4-1:0] node21626;
	wire [4-1:0] node21628;
	wire [4-1:0] node21631;
	wire [4-1:0] node21633;
	wire [4-1:0] node21637;
	wire [4-1:0] node21638;
	wire [4-1:0] node21639;
	wire [4-1:0] node21640;
	wire [4-1:0] node21641;
	wire [4-1:0] node21642;
	wire [4-1:0] node21643;
	wire [4-1:0] node21644;
	wire [4-1:0] node21645;
	wire [4-1:0] node21646;
	wire [4-1:0] node21649;
	wire [4-1:0] node21652;
	wire [4-1:0] node21653;
	wire [4-1:0] node21654;
	wire [4-1:0] node21658;
	wire [4-1:0] node21659;
	wire [4-1:0] node21662;
	wire [4-1:0] node21665;
	wire [4-1:0] node21666;
	wire [4-1:0] node21667;
	wire [4-1:0] node21668;
	wire [4-1:0] node21671;
	wire [4-1:0] node21674;
	wire [4-1:0] node21675;
	wire [4-1:0] node21678;
	wire [4-1:0] node21681;
	wire [4-1:0] node21682;
	wire [4-1:0] node21685;
	wire [4-1:0] node21688;
	wire [4-1:0] node21689;
	wire [4-1:0] node21690;
	wire [4-1:0] node21691;
	wire [4-1:0] node21692;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21701;
	wire [4-1:0] node21702;
	wire [4-1:0] node21703;
	wire [4-1:0] node21705;
	wire [4-1:0] node21708;
	wire [4-1:0] node21709;
	wire [4-1:0] node21713;
	wire [4-1:0] node21714;
	wire [4-1:0] node21716;
	wire [4-1:0] node21720;
	wire [4-1:0] node21721;
	wire [4-1:0] node21722;
	wire [4-1:0] node21725;
	wire [4-1:0] node21726;
	wire [4-1:0] node21730;
	wire [4-1:0] node21731;
	wire [4-1:0] node21732;
	wire [4-1:0] node21735;
	wire [4-1:0] node21737;
	wire [4-1:0] node21740;
	wire [4-1:0] node21741;
	wire [4-1:0] node21744;
	wire [4-1:0] node21747;
	wire [4-1:0] node21748;
	wire [4-1:0] node21749;
	wire [4-1:0] node21750;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21756;
	wire [4-1:0] node21758;
	wire [4-1:0] node21761;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21769;
	wire [4-1:0] node21770;
	wire [4-1:0] node21774;
	wire [4-1:0] node21775;
	wire [4-1:0] node21776;
	wire [4-1:0] node21780;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21785;
	wire [4-1:0] node21786;
	wire [4-1:0] node21787;
	wire [4-1:0] node21788;
	wire [4-1:0] node21791;
	wire [4-1:0] node21794;
	wire [4-1:0] node21795;
	wire [4-1:0] node21798;
	wire [4-1:0] node21801;
	wire [4-1:0] node21802;
	wire [4-1:0] node21805;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21810;
	wire [4-1:0] node21811;
	wire [4-1:0] node21815;
	wire [4-1:0] node21816;
	wire [4-1:0] node21819;
	wire [4-1:0] node21822;
	wire [4-1:0] node21823;
	wire [4-1:0] node21824;
	wire [4-1:0] node21827;
	wire [4-1:0] node21830;
	wire [4-1:0] node21832;
	wire [4-1:0] node21835;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21838;
	wire [4-1:0] node21840;
	wire [4-1:0] node21843;
	wire [4-1:0] node21846;
	wire [4-1:0] node21847;
	wire [4-1:0] node21848;
	wire [4-1:0] node21851;
	wire [4-1:0] node21854;
	wire [4-1:0] node21855;
	wire [4-1:0] node21858;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21867;
	wire [4-1:0] node21870;
	wire [4-1:0] node21871;
	wire [4-1:0] node21874;
	wire [4-1:0] node21877;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21882;
	wire [4-1:0] node21885;
	wire [4-1:0] node21886;
	wire [4-1:0] node21889;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21898;
	wire [4-1:0] node21901;
	wire [4-1:0] node21902;
	wire [4-1:0] node21903;
	wire [4-1:0] node21907;
	wire [4-1:0] node21909;
	wire [4-1:0] node21912;
	wire [4-1:0] node21913;
	wire [4-1:0] node21914;
	wire [4-1:0] node21915;
	wire [4-1:0] node21919;
	wire [4-1:0] node21920;
	wire [4-1:0] node21923;
	wire [4-1:0] node21925;
	wire [4-1:0] node21928;
	wire [4-1:0] node21929;
	wire [4-1:0] node21933;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21941;
	wire [4-1:0] node21943;
	wire [4-1:0] node21946;
	wire [4-1:0] node21947;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21954;
	wire [4-1:0] node21955;
	wire [4-1:0] node21956;
	wire [4-1:0] node21960;
	wire [4-1:0] node21962;
	wire [4-1:0] node21965;
	wire [4-1:0] node21966;
	wire [4-1:0] node21967;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21973;
	wire [4-1:0] node21974;
	wire [4-1:0] node21978;
	wire [4-1:0] node21979;
	wire [4-1:0] node21981;
	wire [4-1:0] node21984;
	wire [4-1:0] node21986;
	wire [4-1:0] node21989;
	wire [4-1:0] node21990;
	wire [4-1:0] node21991;
	wire [4-1:0] node21994;
	wire [4-1:0] node21996;
	wire [4-1:0] node21999;
	wire [4-1:0] node22000;
	wire [4-1:0] node22002;
	wire [4-1:0] node22005;
	wire [4-1:0] node22007;
	wire [4-1:0] node22010;
	wire [4-1:0] node22011;
	wire [4-1:0] node22012;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22021;
	wire [4-1:0] node22022;
	wire [4-1:0] node22025;
	wire [4-1:0] node22028;
	wire [4-1:0] node22029;
	wire [4-1:0] node22032;
	wire [4-1:0] node22033;
	wire [4-1:0] node22037;
	wire [4-1:0] node22038;
	wire [4-1:0] node22039;
	wire [4-1:0] node22041;
	wire [4-1:0] node22044;
	wire [4-1:0] node22045;
	wire [4-1:0] node22049;
	wire [4-1:0] node22050;
	wire [4-1:0] node22051;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22059;
	wire [4-1:0] node22060;
	wire [4-1:0] node22062;
	wire [4-1:0] node22065;
	wire [4-1:0] node22066;
	wire [4-1:0] node22069;
	wire [4-1:0] node22072;
	wire [4-1:0] node22073;
	wire [4-1:0] node22074;
	wire [4-1:0] node22075;
	wire [4-1:0] node22076;
	wire [4-1:0] node22080;
	wire [4-1:0] node22081;
	wire [4-1:0] node22085;
	wire [4-1:0] node22086;
	wire [4-1:0] node22087;
	wire [4-1:0] node22090;
	wire [4-1:0] node22093;
	wire [4-1:0] node22096;
	wire [4-1:0] node22097;
	wire [4-1:0] node22099;
	wire [4-1:0] node22102;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22109;
	wire [4-1:0] node22110;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22115;
	wire [4-1:0] node22116;
	wire [4-1:0] node22117;
	wire [4-1:0] node22122;
	wire [4-1:0] node22123;
	wire [4-1:0] node22124;
	wire [4-1:0] node22127;
	wire [4-1:0] node22128;
	wire [4-1:0] node22132;
	wire [4-1:0] node22133;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22141;
	wire [4-1:0] node22142;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22146;
	wire [4-1:0] node22149;
	wire [4-1:0] node22150;
	wire [4-1:0] node22154;
	wire [4-1:0] node22155;
	wire [4-1:0] node22156;
	wire [4-1:0] node22159;
	wire [4-1:0] node22162;
	wire [4-1:0] node22164;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22169;
	wire [4-1:0] node22170;
	wire [4-1:0] node22173;
	wire [4-1:0] node22176;
	wire [4-1:0] node22178;
	wire [4-1:0] node22181;
	wire [4-1:0] node22182;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22190;
	wire [4-1:0] node22191;
	wire [4-1:0] node22192;
	wire [4-1:0] node22193;
	wire [4-1:0] node22194;
	wire [4-1:0] node22195;
	wire [4-1:0] node22196;
	wire [4-1:0] node22199;
	wire [4-1:0] node22202;
	wire [4-1:0] node22203;
	wire [4-1:0] node22206;
	wire [4-1:0] node22209;
	wire [4-1:0] node22210;
	wire [4-1:0] node22214;
	wire [4-1:0] node22215;
	wire [4-1:0] node22216;
	wire [4-1:0] node22217;
	wire [4-1:0] node22220;
	wire [4-1:0] node22223;
	wire [4-1:0] node22224;
	wire [4-1:0] node22227;
	wire [4-1:0] node22230;
	wire [4-1:0] node22231;
	wire [4-1:0] node22234;
	wire [4-1:0] node22237;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22242;
	wire [4-1:0] node22245;
	wire [4-1:0] node22247;
	wire [4-1:0] node22250;
	wire [4-1:0] node22251;
	wire [4-1:0] node22252;
	wire [4-1:0] node22253;
	wire [4-1:0] node22254;
	wire [4-1:0] node22255;
	wire [4-1:0] node22259;
	wire [4-1:0] node22260;
	wire [4-1:0] node22263;
	wire [4-1:0] node22266;
	wire [4-1:0] node22267;
	wire [4-1:0] node22268;
	wire [4-1:0] node22271;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22278;
	wire [4-1:0] node22281;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22286;
	wire [4-1:0] node22289;
	wire [4-1:0] node22291;
	wire [4-1:0] node22294;
	wire [4-1:0] node22295;
	wire [4-1:0] node22296;
	wire [4-1:0] node22297;
	wire [4-1:0] node22300;
	wire [4-1:0] node22303;
	wire [4-1:0] node22304;
	wire [4-1:0] node22308;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22313;
	wire [4-1:0] node22316;
	wire [4-1:0] node22317;
	wire [4-1:0] node22318;
	wire [4-1:0] node22322;
	wire [4-1:0] node22324;
	wire [4-1:0] node22327;
	wire [4-1:0] node22328;
	wire [4-1:0] node22329;
	wire [4-1:0] node22330;
	wire [4-1:0] node22331;
	wire [4-1:0] node22332;
	wire [4-1:0] node22335;
	wire [4-1:0] node22336;
	wire [4-1:0] node22339;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22346;
	wire [4-1:0] node22349;
	wire [4-1:0] node22350;
	wire [4-1:0] node22352;
	wire [4-1:0] node22355;
	wire [4-1:0] node22356;
	wire [4-1:0] node22359;
	wire [4-1:0] node22361;
	wire [4-1:0] node22364;
	wire [4-1:0] node22365;
	wire [4-1:0] node22366;
	wire [4-1:0] node22367;
	wire [4-1:0] node22371;
	wire [4-1:0] node22372;
	wire [4-1:0] node22373;
	wire [4-1:0] node22376;
	wire [4-1:0] node22380;
	wire [4-1:0] node22381;
	wire [4-1:0] node22382;
	wire [4-1:0] node22384;
	wire [4-1:0] node22387;
	wire [4-1:0] node22388;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22395;
	wire [4-1:0] node22398;
	wire [4-1:0] node22399;
	wire [4-1:0] node22402;
	wire [4-1:0] node22405;
	wire [4-1:0] node22406;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22409;
	wire [4-1:0] node22412;
	wire [4-1:0] node22415;
	wire [4-1:0] node22416;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22423;
	wire [4-1:0] node22426;
	wire [4-1:0] node22427;
	wire [4-1:0] node22430;
	wire [4-1:0] node22433;
	wire [4-1:0] node22434;
	wire [4-1:0] node22436;
	wire [4-1:0] node22437;
	wire [4-1:0] node22441;
	wire [4-1:0] node22442;
	wire [4-1:0] node22446;
	wire [4-1:0] node22447;
	wire [4-1:0] node22448;
	wire [4-1:0] node22449;
	wire [4-1:0] node22451;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22456;
	wire [4-1:0] node22457;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22464;
	wire [4-1:0] node22466;
	wire [4-1:0] node22470;
	wire [4-1:0] node22472;
	wire [4-1:0] node22473;
	wire [4-1:0] node22478;
	wire [4-1:0] node22479;
	wire [4-1:0] node22480;
	wire [4-1:0] node22481;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22488;
	wire [4-1:0] node22490;
	wire [4-1:0] node22493;
	wire [4-1:0] node22494;
	wire [4-1:0] node22498;
	wire [4-1:0] node22499;
	wire [4-1:0] node22500;
	wire [4-1:0] node22502;
	wire [4-1:0] node22506;
	wire [4-1:0] node22508;
	wire [4-1:0] node22511;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22514;
	wire [4-1:0] node22518;
	wire [4-1:0] node22519;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22525;
	wire [4-1:0] node22526;
	wire [4-1:0] node22530;
	wire [4-1:0] node22533;
	wire [4-1:0] node22534;
	wire [4-1:0] node22537;
	wire [4-1:0] node22540;
	wire [4-1:0] node22542;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22546;
	wire [4-1:0] node22548;
	wire [4-1:0] node22551;
	wire [4-1:0] node22552;
	wire [4-1:0] node22553;
	wire [4-1:0] node22557;
	wire [4-1:0] node22559;
	wire [4-1:0] node22562;
	wire [4-1:0] node22564;
	wire [4-1:0] node22566;
	wire [4-1:0] node22569;
	wire [4-1:0] node22570;
	wire [4-1:0] node22571;
	wire [4-1:0] node22572;
	wire [4-1:0] node22573;
	wire [4-1:0] node22574;
	wire [4-1:0] node22576;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22584;
	wire [4-1:0] node22585;
	wire [4-1:0] node22586;
	wire [4-1:0] node22588;
	wire [4-1:0] node22591;
	wire [4-1:0] node22592;
	wire [4-1:0] node22596;
	wire [4-1:0] node22597;
	wire [4-1:0] node22600;
	wire [4-1:0] node22603;
	wire [4-1:0] node22604;
	wire [4-1:0] node22605;
	wire [4-1:0] node22607;
	wire [4-1:0] node22610;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22617;
	wire [4-1:0] node22621;
	wire [4-1:0] node22622;
	wire [4-1:0] node22623;
	wire [4-1:0] node22627;
	wire [4-1:0] node22629;
	wire [4-1:0] node22632;
	wire [4-1:0] node22633;
	wire [4-1:0] node22634;
	wire [4-1:0] node22635;
	wire [4-1:0] node22637;
	wire [4-1:0] node22638;
	wire [4-1:0] node22642;
	wire [4-1:0] node22644;
	wire [4-1:0] node22645;
	wire [4-1:0] node22649;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22655;
	wire [4-1:0] node22656;
	wire [4-1:0] node22660;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22664;
	wire [4-1:0] node22667;
	wire [4-1:0] node22668;
	wire [4-1:0] node22672;
	wire [4-1:0] node22673;
	wire [4-1:0] node22674;
	wire [4-1:0] node22675;
	wire [4-1:0] node22679;
	wire [4-1:0] node22680;
	wire [4-1:0] node22684;
	wire [4-1:0] node22685;
	wire [4-1:0] node22688;
	wire [4-1:0] node22689;
	wire [4-1:0] node22693;
	wire [4-1:0] node22694;
	wire [4-1:0] node22695;
	wire [4-1:0] node22696;
	wire [4-1:0] node22697;
	wire [4-1:0] node22700;
	wire [4-1:0] node22701;
	wire [4-1:0] node22705;
	wire [4-1:0] node22706;
	wire [4-1:0] node22707;
	wire [4-1:0] node22711;
	wire [4-1:0] node22713;
	wire [4-1:0] node22716;
	wire [4-1:0] node22717;
	wire [4-1:0] node22718;
	wire [4-1:0] node22722;
	wire [4-1:0] node22724;
	wire [4-1:0] node22725;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22731;
	wire [4-1:0] node22732;
	wire [4-1:0] node22734;
	wire [4-1:0] node22737;
	wire [4-1:0] node22738;
	wire [4-1:0] node22741;
	wire [4-1:0] node22744;
	wire [4-1:0] node22745;
	wire [4-1:0] node22746;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22753;
	wire [4-1:0] node22757;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22763;
	wire [4-1:0] node22764;
	wire [4-1:0] node22765;
	wire [4-1:0] node22769;
	wire [4-1:0] node22770;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22777;
	wire [4-1:0] node22778;
	wire [4-1:0] node22779;
	wire [4-1:0] node22780;
	wire [4-1:0] node22781;
	wire [4-1:0] node22782;
	wire [4-1:0] node22783;
	wire [4-1:0] node22784;
	wire [4-1:0] node22787;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22793;
	wire [4-1:0] node22796;
	wire [4-1:0] node22798;
	wire [4-1:0] node22801;
	wire [4-1:0] node22802;
	wire [4-1:0] node22803;
	wire [4-1:0] node22805;
	wire [4-1:0] node22808;
	wire [4-1:0] node22811;
	wire [4-1:0] node22813;
	wire [4-1:0] node22816;
	wire [4-1:0] node22817;
	wire [4-1:0] node22818;
	wire [4-1:0] node22820;
	wire [4-1:0] node22823;
	wire [4-1:0] node22825;
	wire [4-1:0] node22828;
	wire [4-1:0] node22829;
	wire [4-1:0] node22830;
	wire [4-1:0] node22832;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22839;
	wire [4-1:0] node22843;
	wire [4-1:0] node22844;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22849;
	wire [4-1:0] node22852;
	wire [4-1:0] node22855;
	wire [4-1:0] node22856;
	wire [4-1:0] node22858;
	wire [4-1:0] node22861;
	wire [4-1:0] node22863;
	wire [4-1:0] node22866;
	wire [4-1:0] node22867;
	wire [4-1:0] node22869;
	wire [4-1:0] node22872;
	wire [4-1:0] node22874;
	wire [4-1:0] node22877;
	wire [4-1:0] node22878;
	wire [4-1:0] node22879;
	wire [4-1:0] node22880;
	wire [4-1:0] node22883;
	wire [4-1:0] node22886;
	wire [4-1:0] node22887;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22894;
	wire [4-1:0] node22897;
	wire [4-1:0] node22900;
	wire [4-1:0] node22901;
	wire [4-1:0] node22902;
	wire [4-1:0] node22903;
	wire [4-1:0] node22905;
	wire [4-1:0] node22908;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22914;
	wire [4-1:0] node22915;
	wire [4-1:0] node22919;
	wire [4-1:0] node22920;
	wire [4-1:0] node22921;
	wire [4-1:0] node22922;
	wire [4-1:0] node22923;
	wire [4-1:0] node22927;
	wire [4-1:0] node22930;
	wire [4-1:0] node22931;
	wire [4-1:0] node22935;
	wire [4-1:0] node22936;
	wire [4-1:0] node22939;
	wire [4-1:0] node22942;
	wire [4-1:0] node22943;
	wire [4-1:0] node22944;
	wire [4-1:0] node22945;
	wire [4-1:0] node22946;
	wire [4-1:0] node22947;
	wire [4-1:0] node22951;
	wire [4-1:0] node22954;
	wire [4-1:0] node22955;
	wire [4-1:0] node22956;
	wire [4-1:0] node22960;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22966;
	wire [4-1:0] node22970;
	wire [4-1:0] node22971;
	wire [4-1:0] node22972;
	wire [4-1:0] node22973;
	wire [4-1:0] node22974;
	wire [4-1:0] node22978;
	wire [4-1:0] node22981;
	wire [4-1:0] node22983;
	wire [4-1:0] node22986;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22993;
	wire [4-1:0] node22994;
	wire [4-1:0] node22995;
	wire [4-1:0] node22996;
	wire [4-1:0] node22997;
	wire [4-1:0] node22999;
	wire [4-1:0] node23002;
	wire [4-1:0] node23003;
	wire [4-1:0] node23004;
	wire [4-1:0] node23005;
	wire [4-1:0] node23009;
	wire [4-1:0] node23011;
	wire [4-1:0] node23014;
	wire [4-1:0] node23016;
	wire [4-1:0] node23019;
	wire [4-1:0] node23020;
	wire [4-1:0] node23021;
	wire [4-1:0] node23022;
	wire [4-1:0] node23025;
	wire [4-1:0] node23028;
	wire [4-1:0] node23029;
	wire [4-1:0] node23030;
	wire [4-1:0] node23034;
	wire [4-1:0] node23035;
	wire [4-1:0] node23039;
	wire [4-1:0] node23040;
	wire [4-1:0] node23041;
	wire [4-1:0] node23045;
	wire [4-1:0] node23047;
	wire [4-1:0] node23050;
	wire [4-1:0] node23051;
	wire [4-1:0] node23052;
	wire [4-1:0] node23053;
	wire [4-1:0] node23054;
	wire [4-1:0] node23058;
	wire [4-1:0] node23059;
	wire [4-1:0] node23063;
	wire [4-1:0] node23064;
	wire [4-1:0] node23066;
	wire [4-1:0] node23069;
	wire [4-1:0] node23070;
	wire [4-1:0] node23074;
	wire [4-1:0] node23075;
	wire [4-1:0] node23076;
	wire [4-1:0] node23077;
	wire [4-1:0] node23081;
	wire [4-1:0] node23082;
	wire [4-1:0] node23084;
	wire [4-1:0] node23087;
	wire [4-1:0] node23089;
	wire [4-1:0] node23092;
	wire [4-1:0] node23093;
	wire [4-1:0] node23094;
	wire [4-1:0] node23098;
	wire [4-1:0] node23099;
	wire [4-1:0] node23101;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23109;
	wire [4-1:0] node23110;
	wire [4-1:0] node23112;
	wire [4-1:0] node23113;
	wire [4-1:0] node23114;
	wire [4-1:0] node23116;
	wire [4-1:0] node23118;
	wire [4-1:0] node23121;
	wire [4-1:0] node23122;
	wire [4-1:0] node23124;
	wire [4-1:0] node23127;
	wire [4-1:0] node23128;
	wire [4-1:0] node23132;
	wire [4-1:0] node23134;
	wire [4-1:0] node23136;
	wire [4-1:0] node23140;
	wire [4-1:0] node23141;
	wire [4-1:0] node23142;
	wire [4-1:0] node23143;
	wire [4-1:0] node23144;
	wire [4-1:0] node23145;
	wire [4-1:0] node23146;
	wire [4-1:0] node23149;
	wire [4-1:0] node23150;
	wire [4-1:0] node23152;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23161;
	wire [4-1:0] node23162;
	wire [4-1:0] node23165;
	wire [4-1:0] node23168;
	wire [4-1:0] node23169;
	wire [4-1:0] node23170;
	wire [4-1:0] node23173;
	wire [4-1:0] node23177;
	wire [4-1:0] node23178;
	wire [4-1:0] node23179;
	wire [4-1:0] node23181;
	wire [4-1:0] node23182;
	wire [4-1:0] node23187;
	wire [4-1:0] node23188;
	wire [4-1:0] node23189;
	wire [4-1:0] node23191;
	wire [4-1:0] node23195;
	wire [4-1:0] node23196;
	wire [4-1:0] node23198;
	wire [4-1:0] node23202;
	wire [4-1:0] node23203;
	wire [4-1:0] node23204;
	wire [4-1:0] node23205;
	wire [4-1:0] node23209;
	wire [4-1:0] node23210;
	wire [4-1:0] node23211;
	wire [4-1:0] node23212;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23221;
	wire [4-1:0] node23222;
	wire [4-1:0] node23226;
	wire [4-1:0] node23227;
	wire [4-1:0] node23228;
	wire [4-1:0] node23229;
	wire [4-1:0] node23230;
	wire [4-1:0] node23234;
	wire [4-1:0] node23237;
	wire [4-1:0] node23238;
	wire [4-1:0] node23241;
	wire [4-1:0] node23244;
	wire [4-1:0] node23245;
	wire [4-1:0] node23246;
	wire [4-1:0] node23249;
	wire [4-1:0] node23252;
	wire [4-1:0] node23254;
	wire [4-1:0] node23257;
	wire [4-1:0] node23258;
	wire [4-1:0] node23259;
	wire [4-1:0] node23260;
	wire [4-1:0] node23261;
	wire [4-1:0] node23262;
	wire [4-1:0] node23263;
	wire [4-1:0] node23267;
	wire [4-1:0] node23269;
	wire [4-1:0] node23272;
	wire [4-1:0] node23273;
	wire [4-1:0] node23276;
	wire [4-1:0] node23279;
	wire [4-1:0] node23280;
	wire [4-1:0] node23281;
	wire [4-1:0] node23282;
	wire [4-1:0] node23285;
	wire [4-1:0] node23288;
	wire [4-1:0] node23289;
	wire [4-1:0] node23292;
	wire [4-1:0] node23295;
	wire [4-1:0] node23296;
	wire [4-1:0] node23297;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23304;
	wire [4-1:0] node23305;
	wire [4-1:0] node23307;
	wire [4-1:0] node23310;
	wire [4-1:0] node23313;
	wire [4-1:0] node23314;
	wire [4-1:0] node23315;
	wire [4-1:0] node23318;
	wire [4-1:0] node23321;
	wire [4-1:0] node23323;
	wire [4-1:0] node23326;
	wire [4-1:0] node23327;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23333;
	wire [4-1:0] node23334;
	wire [4-1:0] node23337;
	wire [4-1:0] node23340;
	wire [4-1:0] node23341;
	wire [4-1:0] node23342;
	wire [4-1:0] node23345;
	wire [4-1:0] node23348;
	wire [4-1:0] node23349;
	wire [4-1:0] node23352;
	wire [4-1:0] node23355;
	wire [4-1:0] node23356;
	wire [4-1:0] node23357;
	wire [4-1:0] node23358;
	wire [4-1:0] node23359;
	wire [4-1:0] node23360;
	wire [4-1:0] node23364;
	wire [4-1:0] node23367;
	wire [4-1:0] node23368;
	wire [4-1:0] node23370;
	wire [4-1:0] node23373;
	wire [4-1:0] node23374;
	wire [4-1:0] node23377;
	wire [4-1:0] node23380;
	wire [4-1:0] node23381;
	wire [4-1:0] node23382;
	wire [4-1:0] node23386;
	wire [4-1:0] node23387;
	wire [4-1:0] node23390;
	wire [4-1:0] node23393;
	wire [4-1:0] node23395;
	wire [4-1:0] node23397;
	wire [4-1:0] node23398;
	wire [4-1:0] node23399;
	wire [4-1:0] node23402;
	wire [4-1:0] node23405;
	wire [4-1:0] node23406;
	wire [4-1:0] node23410;
	wire [4-1:0] node23411;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23414;
	wire [4-1:0] node23415;
	wire [4-1:0] node23417;
	wire [4-1:0] node23420;
	wire [4-1:0] node23421;
	wire [4-1:0] node23425;
	wire [4-1:0] node23426;
	wire [4-1:0] node23427;
	wire [4-1:0] node23430;
	wire [4-1:0] node23433;
	wire [4-1:0] node23435;
	wire [4-1:0] node23438;
	wire [4-1:0] node23439;
	wire [4-1:0] node23440;
	wire [4-1:0] node23441;
	wire [4-1:0] node23445;
	wire [4-1:0] node23446;
	wire [4-1:0] node23450;
	wire [4-1:0] node23451;
	wire [4-1:0] node23452;
	wire [4-1:0] node23456;
	wire [4-1:0] node23458;
	wire [4-1:0] node23461;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23464;
	wire [4-1:0] node23467;
	wire [4-1:0] node23468;
	wire [4-1:0] node23472;
	wire [4-1:0] node23473;
	wire [4-1:0] node23474;
	wire [4-1:0] node23477;
	wire [4-1:0] node23481;
	wire [4-1:0] node23482;
	wire [4-1:0] node23483;
	wire [4-1:0] node23485;
	wire [4-1:0] node23488;
	wire [4-1:0] node23491;
	wire [4-1:0] node23493;
	wire [4-1:0] node23494;
	wire [4-1:0] node23498;
	wire [4-1:0] node23499;
	wire [4-1:0] node23500;
	wire [4-1:0] node23502;
	wire [4-1:0] node23503;
	wire [4-1:0] node23506;
	wire [4-1:0] node23507;
	wire [4-1:0] node23511;
	wire [4-1:0] node23512;
	wire [4-1:0] node23513;
	wire [4-1:0] node23515;
	wire [4-1:0] node23518;
	wire [4-1:0] node23519;
	wire [4-1:0] node23522;
	wire [4-1:0] node23525;
	wire [4-1:0] node23526;
	wire [4-1:0] node23527;
	wire [4-1:0] node23530;
	wire [4-1:0] node23533;
	wire [4-1:0] node23535;
	wire [4-1:0] node23538;
	wire [4-1:0] node23539;
	wire [4-1:0] node23540;
	wire [4-1:0] node23542;
	wire [4-1:0] node23545;
	wire [4-1:0] node23546;
	wire [4-1:0] node23549;
	wire [4-1:0] node23553;
	wire [4-1:0] node23554;
	wire [4-1:0] node23555;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23559;
	wire [4-1:0] node23560;
	wire [4-1:0] node23561;
	wire [4-1:0] node23562;
	wire [4-1:0] node23566;
	wire [4-1:0] node23567;
	wire [4-1:0] node23570;
	wire [4-1:0] node23573;
	wire [4-1:0] node23574;
	wire [4-1:0] node23575;
	wire [4-1:0] node23578;
	wire [4-1:0] node23581;
	wire [4-1:0] node23583;
	wire [4-1:0] node23586;
	wire [4-1:0] node23587;
	wire [4-1:0] node23589;
	wire [4-1:0] node23591;
	wire [4-1:0] node23594;
	wire [4-1:0] node23595;
	wire [4-1:0] node23596;
	wire [4-1:0] node23599;
	wire [4-1:0] node23602;
	wire [4-1:0] node23603;
	wire [4-1:0] node23607;
	wire [4-1:0] node23608;
	wire [4-1:0] node23609;
	wire [4-1:0] node23610;
	wire [4-1:0] node23614;
	wire [4-1:0] node23615;
	wire [4-1:0] node23616;
	wire [4-1:0] node23620;
	wire [4-1:0] node23621;
	wire [4-1:0] node23625;
	wire [4-1:0] node23626;
	wire [4-1:0] node23628;
	wire [4-1:0] node23631;
	wire [4-1:0] node23632;
	wire [4-1:0] node23634;
	wire [4-1:0] node23637;
	wire [4-1:0] node23640;
	wire [4-1:0] node23641;
	wire [4-1:0] node23642;
	wire [4-1:0] node23643;
	wire [4-1:0] node23645;
	wire [4-1:0] node23648;
	wire [4-1:0] node23649;
	wire [4-1:0] node23650;
	wire [4-1:0] node23654;
	wire [4-1:0] node23657;
	wire [4-1:0] node23658;
	wire [4-1:0] node23660;
	wire [4-1:0] node23663;
	wire [4-1:0] node23665;
	wire [4-1:0] node23668;
	wire [4-1:0] node23669;
	wire [4-1:0] node23670;
	wire [4-1:0] node23671;
	wire [4-1:0] node23674;
	wire [4-1:0] node23677;
	wire [4-1:0] node23678;
	wire [4-1:0] node23680;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23686;
	wire [4-1:0] node23689;
	wire [4-1:0] node23690;
	wire [4-1:0] node23694;
	wire [4-1:0] node23695;
	wire [4-1:0] node23697;
	wire [4-1:0] node23700;
	wire [4-1:0] node23702;
	wire [4-1:0] node23705;
	wire [4-1:0] node23706;
	wire [4-1:0] node23707;
	wire [4-1:0] node23708;
	wire [4-1:0] node23709;
	wire [4-1:0] node23710;
	wire [4-1:0] node23713;
	wire [4-1:0] node23716;
	wire [4-1:0] node23717;
	wire [4-1:0] node23718;
	wire [4-1:0] node23723;
	wire [4-1:0] node23724;
	wire [4-1:0] node23727;
	wire [4-1:0] node23728;
	wire [4-1:0] node23729;
	wire [4-1:0] node23733;
	wire [4-1:0] node23734;
	wire [4-1:0] node23738;
	wire [4-1:0] node23739;
	wire [4-1:0] node23740;
	wire [4-1:0] node23741;
	wire [4-1:0] node23742;
	wire [4-1:0] node23745;
	wire [4-1:0] node23748;
	wire [4-1:0] node23750;
	wire [4-1:0] node23753;
	wire [4-1:0] node23754;
	wire [4-1:0] node23755;
	wire [4-1:0] node23758;
	wire [4-1:0] node23761;
	wire [4-1:0] node23764;
	wire [4-1:0] node23765;
	wire [4-1:0] node23766;
	wire [4-1:0] node23770;
	wire [4-1:0] node23771;
	wire [4-1:0] node23772;
	wire [4-1:0] node23775;
	wire [4-1:0] node23778;
	wire [4-1:0] node23780;
	wire [4-1:0] node23783;
	wire [4-1:0] node23784;
	wire [4-1:0] node23785;
	wire [4-1:0] node23786;
	wire [4-1:0] node23788;
	wire [4-1:0] node23790;
	wire [4-1:0] node23793;
	wire [4-1:0] node23795;
	wire [4-1:0] node23796;
	wire [4-1:0] node23799;
	wire [4-1:0] node23802;
	wire [4-1:0] node23803;
	wire [4-1:0] node23804;
	wire [4-1:0] node23805;
	wire [4-1:0] node23809;
	wire [4-1:0] node23810;
	wire [4-1:0] node23814;
	wire [4-1:0] node23815;
	wire [4-1:0] node23816;
	wire [4-1:0] node23821;
	wire [4-1:0] node23822;
	wire [4-1:0] node23823;
	wire [4-1:0] node23824;
	wire [4-1:0] node23828;
	wire [4-1:0] node23829;
	wire [4-1:0] node23831;
	wire [4-1:0] node23835;
	wire [4-1:0] node23836;
	wire [4-1:0] node23837;
	wire [4-1:0] node23839;
	wire [4-1:0] node23842;
	wire [4-1:0] node23845;
	wire [4-1:0] node23846;
	wire [4-1:0] node23848;
	wire [4-1:0] node23851;
	wire [4-1:0] node23852;
	wire [4-1:0] node23855;
	wire [4-1:0] node23858;
	wire [4-1:0] node23859;
	wire [4-1:0] node23860;
	wire [4-1:0] node23861;
	wire [4-1:0] node23862;
	wire [4-1:0] node23863;
	wire [4-1:0] node23865;
	wire [4-1:0] node23868;
	wire [4-1:0] node23869;
	wire [4-1:0] node23873;
	wire [4-1:0] node23874;
	wire [4-1:0] node23875;
	wire [4-1:0] node23878;
	wire [4-1:0] node23881;
	wire [4-1:0] node23883;
	wire [4-1:0] node23886;
	wire [4-1:0] node23887;
	wire [4-1:0] node23888;
	wire [4-1:0] node23891;
	wire [4-1:0] node23892;
	wire [4-1:0] node23895;
	wire [4-1:0] node23898;
	wire [4-1:0] node23899;
	wire [4-1:0] node23901;
	wire [4-1:0] node23904;
	wire [4-1:0] node23905;
	wire [4-1:0] node23908;
	wire [4-1:0] node23911;
	wire [4-1:0] node23912;
	wire [4-1:0] node23913;
	wire [4-1:0] node23914;
	wire [4-1:0] node23916;
	wire [4-1:0] node23917;
	wire [4-1:0] node23920;
	wire [4-1:0] node23923;
	wire [4-1:0] node23924;
	wire [4-1:0] node23928;
	wire [4-1:0] node23929;
	wire [4-1:0] node23930;
	wire [4-1:0] node23933;
	wire [4-1:0] node23936;
	wire [4-1:0] node23937;
	wire [4-1:0] node23938;
	wire [4-1:0] node23942;
	wire [4-1:0] node23943;
	wire [4-1:0] node23947;
	wire [4-1:0] node23948;
	wire [4-1:0] node23949;
	wire [4-1:0] node23950;
	wire [4-1:0] node23954;
	wire [4-1:0] node23956;
	wire [4-1:0] node23959;
	wire [4-1:0] node23960;
	wire [4-1:0] node23961;
	wire [4-1:0] node23964;
	wire [4-1:0] node23967;
	wire [4-1:0] node23969;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23977;
	wire [4-1:0] node23979;
	wire [4-1:0] node23982;
	wire [4-1:0] node23983;
	wire [4-1:0] node23984;
	wire [4-1:0] node23988;
	wire [4-1:0] node23990;
	wire [4-1:0] node23993;
	wire [4-1:0] node23994;
	wire [4-1:0] node23995;
	wire [4-1:0] node23997;
	wire [4-1:0] node24001;
	wire [4-1:0] node24002;
	wire [4-1:0] node24005;
	wire [4-1:0] node24006;
	wire [4-1:0] node24010;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24013;
	wire [4-1:0] node24014;
	wire [4-1:0] node24017;
	wire [4-1:0] node24020;
	wire [4-1:0] node24021;
	wire [4-1:0] node24024;
	wire [4-1:0] node24027;
	wire [4-1:0] node24029;
	wire [4-1:0] node24033;
	wire [4-1:0] node24034;
	wire [4-1:0] node24035;
	wire [4-1:0] node24036;
	wire [4-1:0] node24037;
	wire [4-1:0] node24038;
	wire [4-1:0] node24039;
	wire [4-1:0] node24040;
	wire [4-1:0] node24042;
	wire [4-1:0] node24045;
	wire [4-1:0] node24047;
	wire [4-1:0] node24050;
	wire [4-1:0] node24051;
	wire [4-1:0] node24052;
	wire [4-1:0] node24055;
	wire [4-1:0] node24058;
	wire [4-1:0] node24060;
	wire [4-1:0] node24063;
	wire [4-1:0] node24064;
	wire [4-1:0] node24065;
	wire [4-1:0] node24068;
	wire [4-1:0] node24071;
	wire [4-1:0] node24072;
	wire [4-1:0] node24073;
	wire [4-1:0] node24078;
	wire [4-1:0] node24079;
	wire [4-1:0] node24080;
	wire [4-1:0] node24083;
	wire [4-1:0] node24084;
	wire [4-1:0] node24085;
	wire [4-1:0] node24089;
	wire [4-1:0] node24090;
	wire [4-1:0] node24094;
	wire [4-1:0] node24095;
	wire [4-1:0] node24096;
	wire [4-1:0] node24097;
	wire [4-1:0] node24100;
	wire [4-1:0] node24103;
	wire [4-1:0] node24105;
	wire [4-1:0] node24108;
	wire [4-1:0] node24110;
	wire [4-1:0] node24113;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24116;
	wire [4-1:0] node24117;
	wire [4-1:0] node24118;
	wire [4-1:0] node24121;
	wire [4-1:0] node24124;
	wire [4-1:0] node24125;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24133;
	wire [4-1:0] node24136;
	wire [4-1:0] node24137;
	wire [4-1:0] node24138;
	wire [4-1:0] node24139;
	wire [4-1:0] node24143;
	wire [4-1:0] node24145;
	wire [4-1:0] node24148;
	wire [4-1:0] node24149;
	wire [4-1:0] node24152;
	wire [4-1:0] node24155;
	wire [4-1:0] node24156;
	wire [4-1:0] node24157;
	wire [4-1:0] node24159;
	wire [4-1:0] node24162;
	wire [4-1:0] node24163;
	wire [4-1:0] node24166;
	wire [4-1:0] node24169;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24175;
	wire [4-1:0] node24177;
	wire [4-1:0] node24180;
	wire [4-1:0] node24181;
	wire [4-1:0] node24182;
	wire [4-1:0] node24183;
	wire [4-1:0] node24184;
	wire [4-1:0] node24185;
	wire [4-1:0] node24187;
	wire [4-1:0] node24191;
	wire [4-1:0] node24194;
	wire [4-1:0] node24195;
	wire [4-1:0] node24197;
	wire [4-1:0] node24198;
	wire [4-1:0] node24202;
	wire [4-1:0] node24203;
	wire [4-1:0] node24204;
	wire [4-1:0] node24207;
	wire [4-1:0] node24210;
	wire [4-1:0] node24212;
	wire [4-1:0] node24215;
	wire [4-1:0] node24216;
	wire [4-1:0] node24217;
	wire [4-1:0] node24219;
	wire [4-1:0] node24220;
	wire [4-1:0] node24224;
	wire [4-1:0] node24225;
	wire [4-1:0] node24228;
	wire [4-1:0] node24230;
	wire [4-1:0] node24233;
	wire [4-1:0] node24234;
	wire [4-1:0] node24235;
	wire [4-1:0] node24239;
	wire [4-1:0] node24240;
	wire [4-1:0] node24244;
	wire [4-1:0] node24245;
	wire [4-1:0] node24246;
	wire [4-1:0] node24247;
	wire [4-1:0] node24249;
	wire [4-1:0] node24250;
	wire [4-1:0] node24254;
	wire [4-1:0] node24255;
	wire [4-1:0] node24257;
	wire [4-1:0] node24260;
	wire [4-1:0] node24262;
	wire [4-1:0] node24265;
	wire [4-1:0] node24266;
	wire [4-1:0] node24267;
	wire [4-1:0] node24269;
	wire [4-1:0] node24272;
	wire [4-1:0] node24274;
	wire [4-1:0] node24277;
	wire [4-1:0] node24279;
	wire [4-1:0] node24281;
	wire [4-1:0] node24285;
	wire [4-1:0] node24286;
	wire [4-1:0] node24287;
	wire [4-1:0] node24288;
	wire [4-1:0] node24289;
	wire [4-1:0] node24290;
	wire [4-1:0] node24291;
	wire [4-1:0] node24292;
	wire [4-1:0] node24295;
	wire [4-1:0] node24299;
	wire [4-1:0] node24301;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24307;
	wire [4-1:0] node24310;
	wire [4-1:0] node24312;
	wire [4-1:0] node24313;
	wire [4-1:0] node24317;
	wire [4-1:0] node24318;
	wire [4-1:0] node24319;
	wire [4-1:0] node24321;
	wire [4-1:0] node24324;
	wire [4-1:0] node24326;
	wire [4-1:0] node24327;
	wire [4-1:0] node24331;
	wire [4-1:0] node24332;
	wire [4-1:0] node24333;
	wire [4-1:0] node24334;
	wire [4-1:0] node24339;
	wire [4-1:0] node24340;
	wire [4-1:0] node24344;
	wire [4-1:0] node24345;
	wire [4-1:0] node24346;
	wire [4-1:0] node24347;
	wire [4-1:0] node24348;
	wire [4-1:0] node24349;
	wire [4-1:0] node24353;
	wire [4-1:0] node24354;
	wire [4-1:0] node24357;
	wire [4-1:0] node24360;
	wire [4-1:0] node24361;
	wire [4-1:0] node24363;
	wire [4-1:0] node24366;
	wire [4-1:0] node24367;
	wire [4-1:0] node24371;
	wire [4-1:0] node24372;
	wire [4-1:0] node24373;
	wire [4-1:0] node24375;
	wire [4-1:0] node24379;
	wire [4-1:0] node24380;
	wire [4-1:0] node24381;
	wire [4-1:0] node24385;
	wire [4-1:0] node24387;
	wire [4-1:0] node24391;
	wire [4-1:0] node24392;
	wire [4-1:0] node24393;
	wire [4-1:0] node24394;
	wire [4-1:0] node24395;
	wire [4-1:0] node24396;
	wire [4-1:0] node24398;
	wire [4-1:0] node24401;
	wire [4-1:0] node24403;
	wire [4-1:0] node24406;
	wire [4-1:0] node24407;
	wire [4-1:0] node24408;
	wire [4-1:0] node24413;
	wire [4-1:0] node24414;
	wire [4-1:0] node24415;
	wire [4-1:0] node24419;
	wire [4-1:0] node24420;
	wire [4-1:0] node24423;
	wire [4-1:0] node24428;
	wire [4-1:0] node24429;
	wire [4-1:0] node24430;
	wire [4-1:0] node24431;
	wire [4-1:0] node24432;
	wire [4-1:0] node24434;
	wire [4-1:0] node24435;
	wire [4-1:0] node24436;
	wire [4-1:0] node24438;
	wire [4-1:0] node24439;
	wire [4-1:0] node24440;
	wire [4-1:0] node24441;
	wire [4-1:0] node24442;
	wire [4-1:0] node24447;
	wire [4-1:0] node24448;
	wire [4-1:0] node24451;
	wire [4-1:0] node24452;
	wire [4-1:0] node24456;
	wire [4-1:0] node24458;
	wire [4-1:0] node24460;
	wire [4-1:0] node24462;
	wire [4-1:0] node24465;
	wire [4-1:0] node24466;
	wire [4-1:0] node24467;
	wire [4-1:0] node24468;
	wire [4-1:0] node24469;
	wire [4-1:0] node24473;
	wire [4-1:0] node24474;
	wire [4-1:0] node24476;
	wire [4-1:0] node24480;
	wire [4-1:0] node24481;
	wire [4-1:0] node24484;
	wire [4-1:0] node24485;
	wire [4-1:0] node24489;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24493;
	wire [4-1:0] node24494;
	wire [4-1:0] node24498;
	wire [4-1:0] node24499;
	wire [4-1:0] node24501;
	wire [4-1:0] node24504;
	wire [4-1:0] node24506;
	wire [4-1:0] node24509;
	wire [4-1:0] node24510;
	wire [4-1:0] node24511;
	wire [4-1:0] node24515;
	wire [4-1:0] node24517;
	wire [4-1:0] node24520;
	wire [4-1:0] node24522;
	wire [4-1:0] node24524;
	wire [4-1:0] node24525;
	wire [4-1:0] node24526;
	wire [4-1:0] node24528;
	wire [4-1:0] node24529;
	wire [4-1:0] node24534;
	wire [4-1:0] node24535;
	wire [4-1:0] node24536;
	wire [4-1:0] node24538;
	wire [4-1:0] node24541;
	wire [4-1:0] node24542;
	wire [4-1:0] node24546;
	wire [4-1:0] node24548;
	wire [4-1:0] node24550;
	wire [4-1:0] node24553;
	wire [4-1:0] node24554;
	wire [4-1:0] node24555;
	wire [4-1:0] node24556;
	wire [4-1:0] node24557;
	wire [4-1:0] node24558;
	wire [4-1:0] node24560;
	wire [4-1:0] node24563;
	wire [4-1:0] node24564;
	wire [4-1:0] node24566;
	wire [4-1:0] node24570;
	wire [4-1:0] node24571;
	wire [4-1:0] node24572;
	wire [4-1:0] node24573;
	wire [4-1:0] node24575;
	wire [4-1:0] node24579;
	wire [4-1:0] node24581;
	wire [4-1:0] node24584;
	wire [4-1:0] node24585;
	wire [4-1:0] node24587;
	wire [4-1:0] node24589;
	wire [4-1:0] node24592;
	wire [4-1:0] node24593;
	wire [4-1:0] node24597;
	wire [4-1:0] node24598;
	wire [4-1:0] node24599;
	wire [4-1:0] node24600;
	wire [4-1:0] node24604;
	wire [4-1:0] node24605;
	wire [4-1:0] node24606;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24615;
	wire [4-1:0] node24616;
	wire [4-1:0] node24617;
	wire [4-1:0] node24619;
	wire [4-1:0] node24622;
	wire [4-1:0] node24624;
	wire [4-1:0] node24626;
	wire [4-1:0] node24629;
	wire [4-1:0] node24630;
	wire [4-1:0] node24632;
	wire [4-1:0] node24634;
	wire [4-1:0] node24637;
	wire [4-1:0] node24639;
	wire [4-1:0] node24642;
	wire [4-1:0] node24643;
	wire [4-1:0] node24644;
	wire [4-1:0] node24645;
	wire [4-1:0] node24646;
	wire [4-1:0] node24647;
	wire [4-1:0] node24651;
	wire [4-1:0] node24652;
	wire [4-1:0] node24656;
	wire [4-1:0] node24657;
	wire [4-1:0] node24658;
	wire [4-1:0] node24662;
	wire [4-1:0] node24664;
	wire [4-1:0] node24667;
	wire [4-1:0] node24668;
	wire [4-1:0] node24670;
	wire [4-1:0] node24673;
	wire [4-1:0] node24675;
	wire [4-1:0] node24678;
	wire [4-1:0] node24679;
	wire [4-1:0] node24680;
	wire [4-1:0] node24681;
	wire [4-1:0] node24683;
	wire [4-1:0] node24686;
	wire [4-1:0] node24687;
	wire [4-1:0] node24691;
	wire [4-1:0] node24692;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24698;
	wire [4-1:0] node24700;
	wire [4-1:0] node24703;
	wire [4-1:0] node24704;
	wire [4-1:0] node24706;
	wire [4-1:0] node24709;
	wire [4-1:0] node24712;
	wire [4-1:0] node24713;
	wire [4-1:0] node24714;
	wire [4-1:0] node24715;
	wire [4-1:0] node24716;
	wire [4-1:0] node24720;
	wire [4-1:0] node24722;
	wire [4-1:0] node24725;
	wire [4-1:0] node24726;
	wire [4-1:0] node24727;
	wire [4-1:0] node24731;
	wire [4-1:0] node24732;
	wire [4-1:0] node24736;
	wire [4-1:0] node24737;
	wire [4-1:0] node24738;
	wire [4-1:0] node24742;
	wire [4-1:0] node24744;
	wire [4-1:0] node24747;
	wire [4-1:0] node24748;
	wire [4-1:0] node24749;
	wire [4-1:0] node24750;
	wire [4-1:0] node24751;
	wire [4-1:0] node24752;
	wire [4-1:0] node24753;
	wire [4-1:0] node24754;
	wire [4-1:0] node24759;
	wire [4-1:0] node24760;
	wire [4-1:0] node24762;
	wire [4-1:0] node24765;
	wire [4-1:0] node24768;
	wire [4-1:0] node24769;
	wire [4-1:0] node24771;
	wire [4-1:0] node24774;
	wire [4-1:0] node24776;
	wire [4-1:0] node24779;
	wire [4-1:0] node24780;
	wire [4-1:0] node24781;
	wire [4-1:0] node24782;
	wire [4-1:0] node24783;
	wire [4-1:0] node24788;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24795;
	wire [4-1:0] node24796;
	wire [4-1:0] node24797;
	wire [4-1:0] node24801;
	wire [4-1:0] node24802;
	wire [4-1:0] node24806;
	wire [4-1:0] node24807;
	wire [4-1:0] node24808;
	wire [4-1:0] node24809;
	wire [4-1:0] node24810;
	wire [4-1:0] node24811;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24820;
	wire [4-1:0] node24821;
	wire [4-1:0] node24822;
	wire [4-1:0] node24826;
	wire [4-1:0] node24827;
	wire [4-1:0] node24831;
	wire [4-1:0] node24832;
	wire [4-1:0] node24834;
	wire [4-1:0] node24837;
	wire [4-1:0] node24838;
	wire [4-1:0] node24842;
	wire [4-1:0] node24843;
	wire [4-1:0] node24844;
	wire [4-1:0] node24845;
	wire [4-1:0] node24847;
	wire [4-1:0] node24850;
	wire [4-1:0] node24852;
	wire [4-1:0] node24855;
	wire [4-1:0] node24856;
	wire [4-1:0] node24857;
	wire [4-1:0] node24861;
	wire [4-1:0] node24862;
	wire [4-1:0] node24866;
	wire [4-1:0] node24867;
	wire [4-1:0] node24869;
	wire [4-1:0] node24872;
	wire [4-1:0] node24873;
	wire [4-1:0] node24877;
	wire [4-1:0] node24878;
	wire [4-1:0] node24879;
	wire [4-1:0] node24880;
	wire [4-1:0] node24881;
	wire [4-1:0] node24882;
	wire [4-1:0] node24886;
	wire [4-1:0] node24888;
	wire [4-1:0] node24891;
	wire [4-1:0] node24892;
	wire [4-1:0] node24896;
	wire [4-1:0] node24897;
	wire [4-1:0] node24898;
	wire [4-1:0] node24899;
	wire [4-1:0] node24903;
	wire [4-1:0] node24905;
	wire [4-1:0] node24908;
	wire [4-1:0] node24910;
	wire [4-1:0] node24913;
	wire [4-1:0] node24914;
	wire [4-1:0] node24915;
	wire [4-1:0] node24917;
	wire [4-1:0] node24920;
	wire [4-1:0] node24922;
	wire [4-1:0] node24925;
	wire [4-1:0] node24926;
	wire [4-1:0] node24927;
	wire [4-1:0] node24928;
	wire [4-1:0] node24932;
	wire [4-1:0] node24934;
	wire [4-1:0] node24937;
	wire [4-1:0] node24938;
	wire [4-1:0] node24939;
	wire [4-1:0] node24943;
	wire [4-1:0] node24945;
	wire [4-1:0] node24948;
	wire [4-1:0] node24950;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24954;
	wire [4-1:0] node24956;
	wire [4-1:0] node24957;
	wire [4-1:0] node24959;
	wire [4-1:0] node24961;
	wire [4-1:0] node24964;
	wire [4-1:0] node24965;
	wire [4-1:0] node24966;
	wire [4-1:0] node24970;
	wire [4-1:0] node24972;
	wire [4-1:0] node24974;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24980;
	wire [4-1:0] node24981;
	wire [4-1:0] node24982;
	wire [4-1:0] node24983;
	wire [4-1:0] node24985;
	wire [4-1:0] node24988;
	wire [4-1:0] node24989;
	wire [4-1:0] node24993;
	wire [4-1:0] node24994;
	wire [4-1:0] node24995;
	wire [4-1:0] node24999;
	wire [4-1:0] node25000;
	wire [4-1:0] node25004;
	wire [4-1:0] node25005;
	wire [4-1:0] node25007;
	wire [4-1:0] node25010;
	wire [4-1:0] node25011;
	wire [4-1:0] node25015;
	wire [4-1:0] node25016;
	wire [4-1:0] node25017;
	wire [4-1:0] node25018;
	wire [4-1:0] node25020;
	wire [4-1:0] node25023;
	wire [4-1:0] node25024;
	wire [4-1:0] node25028;
	wire [4-1:0] node25030;
	wire [4-1:0] node25031;
	wire [4-1:0] node25035;
	wire [4-1:0] node25036;
	wire [4-1:0] node25037;
	wire [4-1:0] node25041;
	wire [4-1:0] node25042;
	wire [4-1:0] node25046;
	wire [4-1:0] node25048;
	wire [4-1:0] node25049;
	wire [4-1:0] node25050;
	wire [4-1:0] node25052;
	wire [4-1:0] node25053;
	wire [4-1:0] node25058;
	wire [4-1:0] node25059;
	wire [4-1:0] node25060;
	wire [4-1:0] node25062;
	wire [4-1:0] node25065;
	wire [4-1:0] node25067;
	wire [4-1:0] node25070;
	wire [4-1:0] node25072;
	wire [4-1:0] node25073;
	wire [4-1:0] node25077;
	wire [4-1:0] node25078;
	wire [4-1:0] node25079;
	wire [4-1:0] node25080;
	wire [4-1:0] node25081;
	wire [4-1:0] node25082;
	wire [4-1:0] node25083;
	wire [4-1:0] node25084;
	wire [4-1:0] node25085;
	wire [4-1:0] node25089;
	wire [4-1:0] node25091;
	wire [4-1:0] node25092;
	wire [4-1:0] node25094;
	wire [4-1:0] node25098;
	wire [4-1:0] node25099;
	wire [4-1:0] node25103;
	wire [4-1:0] node25104;
	wire [4-1:0] node25105;
	wire [4-1:0] node25106;
	wire [4-1:0] node25108;
	wire [4-1:0] node25112;
	wire [4-1:0] node25113;
	wire [4-1:0] node25115;
	wire [4-1:0] node25116;
	wire [4-1:0] node25120;
	wire [4-1:0] node25122;
	wire [4-1:0] node25123;
	wire [4-1:0] node25127;
	wire [4-1:0] node25128;
	wire [4-1:0] node25129;
	wire [4-1:0] node25130;
	wire [4-1:0] node25132;
	wire [4-1:0] node25135;
	wire [4-1:0] node25138;
	wire [4-1:0] node25142;
	wire [4-1:0] node25143;
	wire [4-1:0] node25144;
	wire [4-1:0] node25145;
	wire [4-1:0] node25146;
	wire [4-1:0] node25150;
	wire [4-1:0] node25151;
	wire [4-1:0] node25153;
	wire [4-1:0] node25157;
	wire [4-1:0] node25158;
	wire [4-1:0] node25159;
	wire [4-1:0] node25161;
	wire [4-1:0] node25164;
	wire [4-1:0] node25165;
	wire [4-1:0] node25168;
	wire [4-1:0] node25169;
	wire [4-1:0] node25173;
	wire [4-1:0] node25174;
	wire [4-1:0] node25175;
	wire [4-1:0] node25179;
	wire [4-1:0] node25180;
	wire [4-1:0] node25184;
	wire [4-1:0] node25185;
	wire [4-1:0] node25186;
	wire [4-1:0] node25187;
	wire [4-1:0] node25188;
	wire [4-1:0] node25192;
	wire [4-1:0] node25194;
	wire [4-1:0] node25197;
	wire [4-1:0] node25199;
	wire [4-1:0] node25202;
	wire [4-1:0] node25203;
	wire [4-1:0] node25204;
	wire [4-1:0] node25205;
	wire [4-1:0] node25209;
	wire [4-1:0] node25210;
	wire [4-1:0] node25211;
	wire [4-1:0] node25214;
	wire [4-1:0] node25217;
	wire [4-1:0] node25218;
	wire [4-1:0] node25222;
	wire [4-1:0] node25223;
	wire [4-1:0] node25224;
	wire [4-1:0] node25227;
	wire [4-1:0] node25228;
	wire [4-1:0] node25232;
	wire [4-1:0] node25234;
	wire [4-1:0] node25237;
	wire [4-1:0] node25238;
	wire [4-1:0] node25239;
	wire [4-1:0] node25240;
	wire [4-1:0] node25241;
	wire [4-1:0] node25243;
	wire [4-1:0] node25246;
	wire [4-1:0] node25248;
	wire [4-1:0] node25251;
	wire [4-1:0] node25252;
	wire [4-1:0] node25253;
	wire [4-1:0] node25254;
	wire [4-1:0] node25258;
	wire [4-1:0] node25259;
	wire [4-1:0] node25263;
	wire [4-1:0] node25264;
	wire [4-1:0] node25266;
	wire [4-1:0] node25269;
	wire [4-1:0] node25270;
	wire [4-1:0] node25274;
	wire [4-1:0] node25275;
	wire [4-1:0] node25276;
	wire [4-1:0] node25278;
	wire [4-1:0] node25281;
	wire [4-1:0] node25282;
	wire [4-1:0] node25283;
	wire [4-1:0] node25287;
	wire [4-1:0] node25288;
	wire [4-1:0] node25292;
	wire [4-1:0] node25293;
	wire [4-1:0] node25294;
	wire [4-1:0] node25295;
	wire [4-1:0] node25299;
	wire [4-1:0] node25301;
	wire [4-1:0] node25304;
	wire [4-1:0] node25306;
	wire [4-1:0] node25309;
	wire [4-1:0] node25310;
	wire [4-1:0] node25311;
	wire [4-1:0] node25312;
	wire [4-1:0] node25314;
	wire [4-1:0] node25317;
	wire [4-1:0] node25319;
	wire [4-1:0] node25320;
	wire [4-1:0] node25322;
	wire [4-1:0] node25326;
	wire [4-1:0] node25327;
	wire [4-1:0] node25328;
	wire [4-1:0] node25329;
	wire [4-1:0] node25330;
	wire [4-1:0] node25333;
	wire [4-1:0] node25336;
	wire [4-1:0] node25337;
	wire [4-1:0] node25340;
	wire [4-1:0] node25343;
	wire [4-1:0] node25344;
	wire [4-1:0] node25345;
	wire [4-1:0] node25349;
	wire [4-1:0] node25350;
	wire [4-1:0] node25354;
	wire [4-1:0] node25355;
	wire [4-1:0] node25356;
	wire [4-1:0] node25359;
	wire [4-1:0] node25360;
	wire [4-1:0] node25364;
	wire [4-1:0] node25365;
	wire [4-1:0] node25366;
	wire [4-1:0] node25369;
	wire [4-1:0] node25372;
	wire [4-1:0] node25373;
	wire [4-1:0] node25376;
	wire [4-1:0] node25379;
	wire [4-1:0] node25380;
	wire [4-1:0] node25381;
	wire [4-1:0] node25382;
	wire [4-1:0] node25383;
	wire [4-1:0] node25387;
	wire [4-1:0] node25388;
	wire [4-1:0] node25392;
	wire [4-1:0] node25393;
	wire [4-1:0] node25395;
	wire [4-1:0] node25398;
	wire [4-1:0] node25399;
	wire [4-1:0] node25403;
	wire [4-1:0] node25404;
	wire [4-1:0] node25405;
	wire [4-1:0] node25408;
	wire [4-1:0] node25409;
	wire [4-1:0] node25413;
	wire [4-1:0] node25414;
	wire [4-1:0] node25415;
	wire [4-1:0] node25418;
	wire [4-1:0] node25421;
	wire [4-1:0] node25422;
	wire [4-1:0] node25425;
	wire [4-1:0] node25428;
	wire [4-1:0] node25429;
	wire [4-1:0] node25430;
	wire [4-1:0] node25431;
	wire [4-1:0] node25432;
	wire [4-1:0] node25433;
	wire [4-1:0] node25434;
	wire [4-1:0] node25436;
	wire [4-1:0] node25439;
	wire [4-1:0] node25440;
	wire [4-1:0] node25444;
	wire [4-1:0] node25445;
	wire [4-1:0] node25449;
	wire [4-1:0] node25450;
	wire [4-1:0] node25451;
	wire [4-1:0] node25453;
	wire [4-1:0] node25454;
	wire [4-1:0] node25458;
	wire [4-1:0] node25459;
	wire [4-1:0] node25460;
	wire [4-1:0] node25463;
	wire [4-1:0] node25466;
	wire [4-1:0] node25467;
	wire [4-1:0] node25471;
	wire [4-1:0] node25472;
	wire [4-1:0] node25473;
	wire [4-1:0] node25477;
	wire [4-1:0] node25478;
	wire [4-1:0] node25482;
	wire [4-1:0] node25483;
	wire [4-1:0] node25484;
	wire [4-1:0] node25485;
	wire [4-1:0] node25486;
	wire [4-1:0] node25487;
	wire [4-1:0] node25490;
	wire [4-1:0] node25493;
	wire [4-1:0] node25494;
	wire [4-1:0] node25497;
	wire [4-1:0] node25500;
	wire [4-1:0] node25501;
	wire [4-1:0] node25502;
	wire [4-1:0] node25505;
	wire [4-1:0] node25508;
	wire [4-1:0] node25509;
	wire [4-1:0] node25513;
	wire [4-1:0] node25514;
	wire [4-1:0] node25515;
	wire [4-1:0] node25516;
	wire [4-1:0] node25519;
	wire [4-1:0] node25522;
	wire [4-1:0] node25525;
	wire [4-1:0] node25526;
	wire [4-1:0] node25528;
	wire [4-1:0] node25531;
	wire [4-1:0] node25534;
	wire [4-1:0] node25535;
	wire [4-1:0] node25536;
	wire [4-1:0] node25538;
	wire [4-1:0] node25541;
	wire [4-1:0] node25542;
	wire [4-1:0] node25544;
	wire [4-1:0] node25547;
	wire [4-1:0] node25549;
	wire [4-1:0] node25552;
	wire [4-1:0] node25553;
	wire [4-1:0] node25554;
	wire [4-1:0] node25555;
	wire [4-1:0] node25558;
	wire [4-1:0] node25561;
	wire [4-1:0] node25562;
	wire [4-1:0] node25565;
	wire [4-1:0] node25568;
	wire [4-1:0] node25569;
	wire [4-1:0] node25570;
	wire [4-1:0] node25574;
	wire [4-1:0] node25575;
	wire [4-1:0] node25578;
	wire [4-1:0] node25581;
	wire [4-1:0] node25582;
	wire [4-1:0] node25583;
	wire [4-1:0] node25584;
	wire [4-1:0] node25585;
	wire [4-1:0] node25586;
	wire [4-1:0] node25589;
	wire [4-1:0] node25592;
	wire [4-1:0] node25593;
	wire [4-1:0] node25596;
	wire [4-1:0] node25598;
	wire [4-1:0] node25601;
	wire [4-1:0] node25602;
	wire [4-1:0] node25603;
	wire [4-1:0] node25604;
	wire [4-1:0] node25608;
	wire [4-1:0] node25610;
	wire [4-1:0] node25613;
	wire [4-1:0] node25614;
	wire [4-1:0] node25617;
	wire [4-1:0] node25620;
	wire [4-1:0] node25621;
	wire [4-1:0] node25622;
	wire [4-1:0] node25624;
	wire [4-1:0] node25627;
	wire [4-1:0] node25630;
	wire [4-1:0] node25631;
	wire [4-1:0] node25633;
	wire [4-1:0] node25636;
	wire [4-1:0] node25639;
	wire [4-1:0] node25640;
	wire [4-1:0] node25641;
	wire [4-1:0] node25642;
	wire [4-1:0] node25644;
	wire [4-1:0] node25646;
	wire [4-1:0] node25649;
	wire [4-1:0] node25651;
	wire [4-1:0] node25654;
	wire [4-1:0] node25655;
	wire [4-1:0] node25656;
	wire [4-1:0] node25657;
	wire [4-1:0] node25662;
	wire [4-1:0] node25664;
	wire [4-1:0] node25667;
	wire [4-1:0] node25668;
	wire [4-1:0] node25669;
	wire [4-1:0] node25670;
	wire [4-1:0] node25671;
	wire [4-1:0] node25675;
	wire [4-1:0] node25676;
	wire [4-1:0] node25679;
	wire [4-1:0] node25682;
	wire [4-1:0] node25683;
	wire [4-1:0] node25685;
	wire [4-1:0] node25689;
	wire [4-1:0] node25690;
	wire [4-1:0] node25692;
	wire [4-1:0] node25693;
	wire [4-1:0] node25696;
	wire [4-1:0] node25699;
	wire [4-1:0] node25700;
	wire [4-1:0] node25701;
	wire [4-1:0] node25705;
	wire [4-1:0] node25708;
	wire [4-1:0] node25709;
	wire [4-1:0] node25710;
	wire [4-1:0] node25711;
	wire [4-1:0] node25712;
	wire [4-1:0] node25713;
	wire [4-1:0] node25716;
	wire [4-1:0] node25719;
	wire [4-1:0] node25720;
	wire [4-1:0] node25721;
	wire [4-1:0] node25725;
	wire [4-1:0] node25726;
	wire [4-1:0] node25729;
	wire [4-1:0] node25732;
	wire [4-1:0] node25733;
	wire [4-1:0] node25736;
	wire [4-1:0] node25737;
	wire [4-1:0] node25741;
	wire [4-1:0] node25742;
	wire [4-1:0] node25743;
	wire [4-1:0] node25745;
	wire [4-1:0] node25748;
	wire [4-1:0] node25749;
	wire [4-1:0] node25751;
	wire [4-1:0] node25755;
	wire [4-1:0] node25756;
	wire [4-1:0] node25757;
	wire [4-1:0] node25758;
	wire [4-1:0] node25761;
	wire [4-1:0] node25764;
	wire [4-1:0] node25765;
	wire [4-1:0] node25769;
	wire [4-1:0] node25770;
	wire [4-1:0] node25772;
	wire [4-1:0] node25775;
	wire [4-1:0] node25778;
	wire [4-1:0] node25779;
	wire [4-1:0] node25780;
	wire [4-1:0] node25782;
	wire [4-1:0] node25783;
	wire [4-1:0] node25787;
	wire [4-1:0] node25788;
	wire [4-1:0] node25789;
	wire [4-1:0] node25792;
	wire [4-1:0] node25795;
	wire [4-1:0] node25797;
	wire [4-1:0] node25800;
	wire [4-1:0] node25801;
	wire [4-1:0] node25802;
	wire [4-1:0] node25803;
	wire [4-1:0] node25807;
	wire [4-1:0] node25808;
	wire [4-1:0] node25811;
	wire [4-1:0] node25814;
	wire [4-1:0] node25815;
	wire [4-1:0] node25819;
	wire [4-1:0] node25820;
	wire [4-1:0] node25821;
	wire [4-1:0] node25822;
	wire [4-1:0] node25823;
	wire [4-1:0] node25824;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25830;
	wire [4-1:0] node25833;
	wire [4-1:0] node25835;
	wire [4-1:0] node25838;
	wire [4-1:0] node25839;
	wire [4-1:0] node25840;
	wire [4-1:0] node25841;
	wire [4-1:0] node25845;
	wire [4-1:0] node25847;
	wire [4-1:0] node25850;
	wire [4-1:0] node25851;
	wire [4-1:0] node25852;
	wire [4-1:0] node25855;
	wire [4-1:0] node25859;
	wire [4-1:0] node25860;
	wire [4-1:0] node25861;
	wire [4-1:0] node25862;
	wire [4-1:0] node25863;
	wire [4-1:0] node25867;
	wire [4-1:0] node25869;
	wire [4-1:0] node25872;
	wire [4-1:0] node25873;
	wire [4-1:0] node25876;
	wire [4-1:0] node25878;
	wire [4-1:0] node25881;
	wire [4-1:0] node25882;
	wire [4-1:0] node25885;
	wire [4-1:0] node25886;
	wire [4-1:0] node25890;
	wire [4-1:0] node25891;
	wire [4-1:0] node25892;
	wire [4-1:0] node25893;
	wire [4-1:0] node25894;
	wire [4-1:0] node25896;
	wire [4-1:0] node25899;
	wire [4-1:0] node25900;
	wire [4-1:0] node25903;
	wire [4-1:0] node25906;
	wire [4-1:0] node25907;
	wire [4-1:0] node25910;
	wire [4-1:0] node25911;
	wire [4-1:0] node25914;
	wire [4-1:0] node25917;
	wire [4-1:0] node25918;
	wire [4-1:0] node25919;
	wire [4-1:0] node25920;
	wire [4-1:0] node25924;
	wire [4-1:0] node25925;
	wire [4-1:0] node25929;
	wire [4-1:0] node25931;
	wire [4-1:0] node25934;
	wire [4-1:0] node25935;
	wire [4-1:0] node25936;
	wire [4-1:0] node25938;
	wire [4-1:0] node25941;
	wire [4-1:0] node25942;
	wire [4-1:0] node25944;
	wire [4-1:0] node25947;
	wire [4-1:0] node25948;
	wire [4-1:0] node25951;
	wire [4-1:0] node25954;
	wire [4-1:0] node25955;
	wire [4-1:0] node25957;
	wire [4-1:0] node25959;
	wire [4-1:0] node25962;
	wire [4-1:0] node25963;
	wire [4-1:0] node25967;
	wire [4-1:0] node25968;
	wire [4-1:0] node25969;
	wire [4-1:0] node25970;
	wire [4-1:0] node25972;
	wire [4-1:0] node25975;
	wire [4-1:0] node25976;
	wire [4-1:0] node25977;
	wire [4-1:0] node25981;
	wire [4-1:0] node25982;
	wire [4-1:0] node25986;
	wire [4-1:0] node25987;
	wire [4-1:0] node25988;
	wire [4-1:0] node25992;
	wire [4-1:0] node25993;
	wire [4-1:0] node25994;
	wire [4-1:0] node25997;
	wire [4-1:0] node26000;
	wire [4-1:0] node26001;
	wire [4-1:0] node26005;
	wire [4-1:0] node26006;
	wire [4-1:0] node26007;
	wire [4-1:0] node26008;
	wire [4-1:0] node26009;
	wire [4-1:0] node26010;
	wire [4-1:0] node26014;
	wire [4-1:0] node26017;
	wire [4-1:0] node26018;
	wire [4-1:0] node26019;
	wire [4-1:0] node26022;
	wire [4-1:0] node26025;
	wire [4-1:0] node26028;
	wire [4-1:0] node26029;
	wire [4-1:0] node26030;
	wire [4-1:0] node26034;
	wire [4-1:0] node26035;
	wire [4-1:0] node26036;
	wire [4-1:0] node26040;
	wire [4-1:0] node26043;
	wire [4-1:0] node26044;
	wire [4-1:0] node26045;
	wire [4-1:0] node26047;
	wire [4-1:0] node26050;
	wire [4-1:0] node26051;
	wire [4-1:0] node26054;
	wire [4-1:0] node26057;
	wire [4-1:0] node26058;
	wire [4-1:0] node26059;
	wire [4-1:0] node26062;
	wire [4-1:0] node26065;
	wire [4-1:0] node26066;
	wire [4-1:0] node26069;
	wire [4-1:0] node26071;
	wire [4-1:0] node26074;
	wire [4-1:0] node26075;
	wire [4-1:0] node26076;
	wire [4-1:0] node26077;
	wire [4-1:0] node26078;
	wire [4-1:0] node26079;
	wire [4-1:0] node26082;
	wire [4-1:0] node26085;
	wire [4-1:0] node26086;
	wire [4-1:0] node26087;
	wire [4-1:0] node26091;
	wire [4-1:0] node26094;
	wire [4-1:0] node26095;
	wire [4-1:0] node26096;
	wire [4-1:0] node26098;
	wire [4-1:0] node26101;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26106;
	wire [4-1:0] node26109;
	wire [4-1:0] node26112;
	wire [4-1:0] node26113;
	wire [4-1:0] node26116;
	wire [4-1:0] node26119;
	wire [4-1:0] node26120;
	wire [4-1:0] node26121;
	wire [4-1:0] node26122;
	wire [4-1:0] node26124;
	wire [4-1:0] node26127;
	wire [4-1:0] node26128;
	wire [4-1:0] node26132;
	wire [4-1:0] node26133;
	wire [4-1:0] node26134;
	wire [4-1:0] node26137;
	wire [4-1:0] node26141;
	wire [4-1:0] node26142;
	wire [4-1:0] node26144;
	wire [4-1:0] node26145;
	wire [4-1:0] node26149;
	wire [4-1:0] node26150;
	wire [4-1:0] node26152;
	wire [4-1:0] node26155;
	wire [4-1:0] node26158;
	wire [4-1:0] node26159;
	wire [4-1:0] node26160;
	wire [4-1:0] node26161;
	wire [4-1:0] node26162;
	wire [4-1:0] node26164;
	wire [4-1:0] node26167;
	wire [4-1:0] node26169;
	wire [4-1:0] node26172;
	wire [4-1:0] node26173;
	wire [4-1:0] node26176;
	wire [4-1:0] node26179;
	wire [4-1:0] node26180;
	wire [4-1:0] node26182;
	wire [4-1:0] node26185;
	wire [4-1:0] node26186;
	wire [4-1:0] node26188;
	wire [4-1:0] node26192;
	wire [4-1:0] node26193;
	wire [4-1:0] node26194;
	wire [4-1:0] node26195;
	wire [4-1:0] node26197;
	wire [4-1:0] node26200;
	wire [4-1:0] node26203;
	wire [4-1:0] node26204;
	wire [4-1:0] node26205;
	wire [4-1:0] node26208;
	wire [4-1:0] node26211;
	wire [4-1:0] node26212;
	wire [4-1:0] node26213;
	wire [4-1:0] node26216;
	wire [4-1:0] node26220;
	wire [4-1:0] node26221;
	wire [4-1:0] node26223;
	wire [4-1:0] node26227;
	wire [4-1:0] node26228;
	wire [4-1:0] node26229;
	wire [4-1:0] node26230;
	wire [4-1:0] node26231;
	wire [4-1:0] node26232;
	wire [4-1:0] node26233;
	wire [4-1:0] node26235;
	wire [4-1:0] node26238;
	wire [4-1:0] node26240;
	wire [4-1:0] node26241;
	wire [4-1:0] node26245;
	wire [4-1:0] node26246;
	wire [4-1:0] node26247;
	wire [4-1:0] node26248;
	wire [4-1:0] node26252;
	wire [4-1:0] node26253;
	wire [4-1:0] node26257;
	wire [4-1:0] node26258;
	wire [4-1:0] node26260;
	wire [4-1:0] node26263;
	wire [4-1:0] node26264;
	wire [4-1:0] node26268;
	wire [4-1:0] node26269;
	wire [4-1:0] node26270;
	wire [4-1:0] node26271;
	wire [4-1:0] node26272;
	wire [4-1:0] node26275;
	wire [4-1:0] node26278;
	wire [4-1:0] node26279;
	wire [4-1:0] node26283;
	wire [4-1:0] node26284;
	wire [4-1:0] node26285;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26292;
	wire [4-1:0] node26295;
	wire [4-1:0] node26296;
	wire [4-1:0] node26300;
	wire [4-1:0] node26302;
	wire [4-1:0] node26305;
	wire [4-1:0] node26306;
	wire [4-1:0] node26307;
	wire [4-1:0] node26308;
	wire [4-1:0] node26310;
	wire [4-1:0] node26311;
	wire [4-1:0] node26314;
	wire [4-1:0] node26317;
	wire [4-1:0] node26318;
	wire [4-1:0] node26319;
	wire [4-1:0] node26322;
	wire [4-1:0] node26325;
	wire [4-1:0] node26328;
	wire [4-1:0] node26329;
	wire [4-1:0] node26330;
	wire [4-1:0] node26331;
	wire [4-1:0] node26335;
	wire [4-1:0] node26336;
	wire [4-1:0] node26340;
	wire [4-1:0] node26341;
	wire [4-1:0] node26342;
	wire [4-1:0] node26346;
	wire [4-1:0] node26349;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26354;
	wire [4-1:0] node26356;
	wire [4-1:0] node26359;
	wire [4-1:0] node26360;
	wire [4-1:0] node26361;
	wire [4-1:0] node26365;
	wire [4-1:0] node26366;
	wire [4-1:0] node26367;
	wire [4-1:0] node26371;
	wire [4-1:0] node26374;
	wire [4-1:0] node26375;
	wire [4-1:0] node26376;
	wire [4-1:0] node26377;
	wire [4-1:0] node26378;
	wire [4-1:0] node26379;
	wire [4-1:0] node26383;
	wire [4-1:0] node26386;
	wire [4-1:0] node26387;
	wire [4-1:0] node26389;
	wire [4-1:0] node26391;
	wire [4-1:0] node26394;
	wire [4-1:0] node26395;
	wire [4-1:0] node26399;
	wire [4-1:0] node26400;
	wire [4-1:0] node26402;
	wire [4-1:0] node26403;
	wire [4-1:0] node26406;
	wire [4-1:0] node26409;
	wire [4-1:0] node26410;
	wire [4-1:0] node26412;
	wire [4-1:0] node26415;
	wire [4-1:0] node26416;
	wire [4-1:0] node26420;
	wire [4-1:0] node26421;
	wire [4-1:0] node26422;
	wire [4-1:0] node26423;
	wire [4-1:0] node26426;
	wire [4-1:0] node26427;
	wire [4-1:0] node26431;
	wire [4-1:0] node26432;
	wire [4-1:0] node26434;
	wire [4-1:0] node26435;
	wire [4-1:0] node26440;
	wire [4-1:0] node26441;
	wire [4-1:0] node26443;
	wire [4-1:0] node26447;
	wire [4-1:0] node26448;
	wire [4-1:0] node26449;
	wire [4-1:0] node26450;
	wire [4-1:0] node26451;
	wire [4-1:0] node26452;
	wire [4-1:0] node26454;
	wire [4-1:0] node26455;
	wire [4-1:0] node26459;
	wire [4-1:0] node26460;
	wire [4-1:0] node26461;
	wire [4-1:0] node26465;
	wire [4-1:0] node26466;
	wire [4-1:0] node26470;
	wire [4-1:0] node26471;
	wire [4-1:0] node26472;
	wire [4-1:0] node26473;
	wire [4-1:0] node26476;
	wire [4-1:0] node26480;
	wire [4-1:0] node26481;
	wire [4-1:0] node26485;
	wire [4-1:0] node26486;
	wire [4-1:0] node26487;
	wire [4-1:0] node26488;
	wire [4-1:0] node26492;
	wire [4-1:0] node26493;
	wire [4-1:0] node26496;
	wire [4-1:0] node26499;
	wire [4-1:0] node26500;
	wire [4-1:0] node26501;
	wire [4-1:0] node26502;
	wire [4-1:0] node26506;
	wire [4-1:0] node26509;
	wire [4-1:0] node26510;
	wire [4-1:0] node26511;
	wire [4-1:0] node26515;
	wire [4-1:0] node26517;
	wire [4-1:0] node26520;
	wire [4-1:0] node26521;
	wire [4-1:0] node26522;
	wire [4-1:0] node26523;
	wire [4-1:0] node26524;
	wire [4-1:0] node26525;
	wire [4-1:0] node26528;
	wire [4-1:0] node26533;
	wire [4-1:0] node26534;
	wire [4-1:0] node26535;
	wire [4-1:0] node26536;
	wire [4-1:0] node26539;
	wire [4-1:0] node26542;
	wire [4-1:0] node26544;
	wire [4-1:0] node26547;
	wire [4-1:0] node26548;
	wire [4-1:0] node26552;
	wire [4-1:0] node26553;
	wire [4-1:0] node26554;
	wire [4-1:0] node26555;
	wire [4-1:0] node26556;
	wire [4-1:0] node26560;
	wire [4-1:0] node26562;
	wire [4-1:0] node26565;
	wire [4-1:0] node26566;
	wire [4-1:0] node26567;
	wire [4-1:0] node26571;
	wire [4-1:0] node26573;
	wire [4-1:0] node26577;
	wire [4-1:0] node26578;
	wire [4-1:0] node26579;
	wire [4-1:0] node26580;
	wire [4-1:0] node26581;
	wire [4-1:0] node26582;
	wire [4-1:0] node26584;
	wire [4-1:0] node26587;
	wire [4-1:0] node26590;
	wire [4-1:0] node26591;
	wire [4-1:0] node26592;
	wire [4-1:0] node26596;
	wire [4-1:0] node26598;
	wire [4-1:0] node26601;
	wire [4-1:0] node26602;
	wire [4-1:0] node26603;
	wire [4-1:0] node26604;
	wire [4-1:0] node26607;
	wire [4-1:0] node26611;
	wire [4-1:0] node26612;
	wire [4-1:0] node26613;
	wire [4-1:0] node26616;
	wire [4-1:0] node26620;
	wire [4-1:0] node26621;
	wire [4-1:0] node26622;
	wire [4-1:0] node26623;
	wire [4-1:0] node26627;
	wire [4-1:0] node26629;
	wire [4-1:0] node26633;
	wire [4-1:0] node26634;
	wire [4-1:0] node26635;
	wire [4-1:0] node26636;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26641;
	wire [4-1:0] node26645;
	wire [4-1:0] node26647;
	wire [4-1:0] node26649;
	wire [4-1:0] node26654;
	wire [4-1:0] node26656;
	wire [4-1:0] node26657;
	wire [4-1:0] node26658;
	wire [4-1:0] node26660;
	wire [4-1:0] node26661;
	wire [4-1:0] node26662;
	wire [4-1:0] node26664;
	wire [4-1:0] node26665;
	wire [4-1:0] node26667;
	wire [4-1:0] node26668;
	wire [4-1:0] node26669;
	wire [4-1:0] node26673;
	wire [4-1:0] node26675;
	wire [4-1:0] node26679;
	wire [4-1:0] node26680;
	wire [4-1:0] node26681;
	wire [4-1:0] node26682;
	wire [4-1:0] node26684;
	wire [4-1:0] node26687;
	wire [4-1:0] node26688;
	wire [4-1:0] node26689;
	wire [4-1:0] node26694;
	wire [4-1:0] node26695;
	wire [4-1:0] node26696;
	wire [4-1:0] node26699;
	wire [4-1:0] node26701;
	wire [4-1:0] node26704;
	wire [4-1:0] node26705;
	wire [4-1:0] node26709;
	wire [4-1:0] node26710;
	wire [4-1:0] node26711;
	wire [4-1:0] node26713;
	wire [4-1:0] node26716;
	wire [4-1:0] node26717;
	wire [4-1:0] node26721;
	wire [4-1:0] node26722;
	wire [4-1:0] node26723;
	wire [4-1:0] node26724;
	wire [4-1:0] node26728;
	wire [4-1:0] node26731;
	wire [4-1:0] node26732;
	wire [4-1:0] node26735;
	wire [4-1:0] node26737;
	wire [4-1:0] node26740;
	wire [4-1:0] node26742;
	wire [4-1:0] node26744;
	wire [4-1:0] node26745;
	wire [4-1:0] node26747;
	wire [4-1:0] node26748;
	wire [4-1:0] node26750;
	wire [4-1:0] node26753;
	wire [4-1:0] node26754;
	wire [4-1:0] node26759;
	wire [4-1:0] node26760;
	wire [4-1:0] node26761;
	wire [4-1:0] node26762;
	wire [4-1:0] node26763;
	wire [4-1:0] node26764;
	wire [4-1:0] node26765;
	wire [4-1:0] node26768;
	wire [4-1:0] node26769;
	wire [4-1:0] node26773;
	wire [4-1:0] node26774;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26780;
	wire [4-1:0] node26782;
	wire [4-1:0] node26785;
	wire [4-1:0] node26786;
	wire [4-1:0] node26790;
	wire [4-1:0] node26791;
	wire [4-1:0] node26792;
	wire [4-1:0] node26794;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26802;
	wire [4-1:0] node26803;
	wire [4-1:0] node26807;
	wire [4-1:0] node26808;
	wire [4-1:0] node26809;
	wire [4-1:0] node26810;
	wire [4-1:0] node26811;
	wire [4-1:0] node26813;
	wire [4-1:0] node26816;
	wire [4-1:0] node26817;
	wire [4-1:0] node26821;
	wire [4-1:0] node26822;
	wire [4-1:0] node26823;
	wire [4-1:0] node26827;
	wire [4-1:0] node26829;
	wire [4-1:0] node26832;
	wire [4-1:0] node26833;
	wire [4-1:0] node26834;
	wire [4-1:0] node26836;
	wire [4-1:0] node26839;
	wire [4-1:0] node26840;
	wire [4-1:0] node26844;
	wire [4-1:0] node26845;
	wire [4-1:0] node26847;
	wire [4-1:0] node26851;
	wire [4-1:0] node26852;
	wire [4-1:0] node26853;
	wire [4-1:0] node26855;
	wire [4-1:0] node26857;
	wire [4-1:0] node26861;
	wire [4-1:0] node26862;
	wire [4-1:0] node26863;
	wire [4-1:0] node26865;
	wire [4-1:0] node26869;
	wire [4-1:0] node26871;
	wire [4-1:0] node26872;
	wire [4-1:0] node26876;
	wire [4-1:0] node26877;
	wire [4-1:0] node26878;
	wire [4-1:0] node26879;
	wire [4-1:0] node26881;
	wire [4-1:0] node26882;
	wire [4-1:0] node26884;
	wire [4-1:0] node26887;
	wire [4-1:0] node26890;
	wire [4-1:0] node26891;
	wire [4-1:0] node26894;
	wire [4-1:0] node26895;
	wire [4-1:0] node26898;
	wire [4-1:0] node26901;
	wire [4-1:0] node26902;
	wire [4-1:0] node26903;
	wire [4-1:0] node26904;
	wire [4-1:0] node26906;
	wire [4-1:0] node26910;
	wire [4-1:0] node26912;
	wire [4-1:0] node26915;
	wire [4-1:0] node26916;
	wire [4-1:0] node26917;
	wire [4-1:0] node26921;
	wire [4-1:0] node26922;
	wire [4-1:0] node26926;
	wire [4-1:0] node26927;
	wire [4-1:0] node26928;
	wire [4-1:0] node26929;
	wire [4-1:0] node26930;
	wire [4-1:0] node26931;
	wire [4-1:0] node26935;
	wire [4-1:0] node26936;
	wire [4-1:0] node26940;
	wire [4-1:0] node26941;
	wire [4-1:0] node26945;
	wire [4-1:0] node26946;
	wire [4-1:0] node26947;
	wire [4-1:0] node26950;
	wire [4-1:0] node26952;
	wire [4-1:0] node26955;
	wire [4-1:0] node26957;
	wire [4-1:0] node26960;
	wire [4-1:0] node26961;
	wire [4-1:0] node26962;
	wire [4-1:0] node26963;
	wire [4-1:0] node26966;
	wire [4-1:0] node26968;
	wire [4-1:0] node26971;
	wire [4-1:0] node26973;
	wire [4-1:0] node26976;
	wire [4-1:0] node26977;
	wire [4-1:0] node26978;
	wire [4-1:0] node26980;
	wire [4-1:0] node26983;
	wire [4-1:0] node26984;
	wire [4-1:0] node26987;
	wire [4-1:0] node26991;
	wire [4-1:0] node26992;
	wire [4-1:0] node26993;
	wire [4-1:0] node26994;
	wire [4-1:0] node26995;
	wire [4-1:0] node26996;
	wire [4-1:0] node26998;
	wire [4-1:0] node26999;
	wire [4-1:0] node27002;
	wire [4-1:0] node27005;
	wire [4-1:0] node27006;
	wire [4-1:0] node27007;
	wire [4-1:0] node27010;
	wire [4-1:0] node27013;
	wire [4-1:0] node27014;
	wire [4-1:0] node27018;
	wire [4-1:0] node27019;
	wire [4-1:0] node27020;
	wire [4-1:0] node27024;
	wire [4-1:0] node27025;
	wire [4-1:0] node27027;
	wire [4-1:0] node27031;
	wire [4-1:0] node27032;
	wire [4-1:0] node27033;
	wire [4-1:0] node27035;
	wire [4-1:0] node27038;
	wire [4-1:0] node27039;
	wire [4-1:0] node27041;
	wire [4-1:0] node27044;
	wire [4-1:0] node27045;
	wire [4-1:0] node27049;
	wire [4-1:0] node27051;
	wire [4-1:0] node27052;
	wire [4-1:0] node27053;
	wire [4-1:0] node27058;
	wire [4-1:0] node27059;
	wire [4-1:0] node27060;
	wire [4-1:0] node27061;
	wire [4-1:0] node27062;
	wire [4-1:0] node27064;
	wire [4-1:0] node27067;
	wire [4-1:0] node27070;
	wire [4-1:0] node27071;
	wire [4-1:0] node27073;
	wire [4-1:0] node27076;
	wire [4-1:0] node27079;
	wire [4-1:0] node27080;
	wire [4-1:0] node27081;
	wire [4-1:0] node27083;
	wire [4-1:0] node27086;
	wire [4-1:0] node27087;
	wire [4-1:0] node27090;
	wire [4-1:0] node27093;
	wire [4-1:0] node27094;
	wire [4-1:0] node27095;
	wire [4-1:0] node27098;
	wire [4-1:0] node27101;
	wire [4-1:0] node27102;
	wire [4-1:0] node27105;
	wire [4-1:0] node27108;
	wire [4-1:0] node27109;
	wire [4-1:0] node27110;
	wire [4-1:0] node27113;
	wire [4-1:0] node27115;
	wire [4-1:0] node27116;
	wire [4-1:0] node27121;
	wire [4-1:0] node27122;
	wire [4-1:0] node27123;
	wire [4-1:0] node27124;
	wire [4-1:0] node27125;
	wire [4-1:0] node27126;
	wire [4-1:0] node27129;
	wire [4-1:0] node27132;
	wire [4-1:0] node27134;
	wire [4-1:0] node27137;
	wire [4-1:0] node27139;
	wire [4-1:0] node27142;
	wire [4-1:0] node27143;
	wire [4-1:0] node27144;
	wire [4-1:0] node27145;
	wire [4-1:0] node27149;
	wire [4-1:0] node27150;
	wire [4-1:0] node27154;
	wire [4-1:0] node27155;
	wire [4-1:0] node27159;
	wire [4-1:0] node27160;
	wire [4-1:0] node27161;
	wire [4-1:0] node27162;
	wire [4-1:0] node27163;
	wire [4-1:0] node27166;
	wire [4-1:0] node27170;
	wire [4-1:0] node27172;
	wire [4-1:0] node27173;
	wire [4-1:0] node27177;
	wire [4-1:0] node27178;
	wire [4-1:0] node27179;
	wire [4-1:0] node27184;
	wire [4-1:0] node27186;
	wire [4-1:0] node27188;
	wire [4-1:0] node27189;
	wire [4-1:0] node27190;
	wire [4-1:0] node27192;
	wire [4-1:0] node27194;
	wire [4-1:0] node27195;
	wire [4-1:0] node27196;
	wire [4-1:0] node27198;
	wire [4-1:0] node27201;
	wire [4-1:0] node27202;
	wire [4-1:0] node27207;
	wire [4-1:0] node27208;
	wire [4-1:0] node27209;
	wire [4-1:0] node27210;
	wire [4-1:0] node27212;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27217;
	wire [4-1:0] node27221;
	wire [4-1:0] node27224;
	wire [4-1:0] node27225;
	wire [4-1:0] node27226;
	wire [4-1:0] node27227;
	wire [4-1:0] node27231;
	wire [4-1:0] node27232;
	wire [4-1:0] node27236;
	wire [4-1:0] node27237;
	wire [4-1:0] node27238;
	wire [4-1:0] node27241;
	wire [4-1:0] node27245;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27248;
	wire [4-1:0] node27249;
	wire [4-1:0] node27252;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27261;
	wire [4-1:0] node27262;
	wire [4-1:0] node27263;
	wire [4-1:0] node27268;
	wire [4-1:0] node27270;
	wire [4-1:0] node27272;
	wire [4-1:0] node27273;
	wire [4-1:0] node27275;
	wire [4-1:0] node27276;
	wire [4-1:0] node27277;

	assign outp = (inp[8]) ? node13738 : node1;
		assign node1 = (inp[9]) ? node6813 : node2;
			assign node2 = (inp[6]) ? node1474 : node3;
				assign node3 = (inp[15]) ? node809 : node4;
					assign node4 = (inp[0]) ? 4'b1101 : node5;
						assign node5 = (inp[5]) ? node349 : node6;
							assign node6 = (inp[2]) ? 4'b1111 : node7;
								assign node7 = (inp[3]) ? node135 : node8;
									assign node8 = (inp[4]) ? node60 : node9;
										assign node9 = (inp[7]) ? 4'b1111 : node10;
											assign node10 = (inp[13]) ? node34 : node11;
												assign node11 = (inp[12]) ? node23 : node12;
													assign node12 = (inp[1]) ? node18 : node13;
														assign node13 = (inp[14]) ? node15 : 4'b0000;
															assign node15 = (inp[11]) ? 4'b0000 : 4'b1111;
														assign node18 = (inp[14]) ? node20 : 4'b0001;
															assign node20 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node23 = (inp[10]) ? node25 : 4'b1111;
														assign node25 = (inp[1]) ? node29 : node26;
															assign node26 = (inp[14]) ? 4'b1111 : 4'b0000;
															assign node29 = (inp[14]) ? node31 : 4'b0001;
																assign node31 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node34 = (inp[12]) ? node46 : node35;
													assign node35 = (inp[1]) ? node41 : node36;
														assign node36 = (inp[14]) ? node38 : 4'b1000;
															assign node38 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node41 = (inp[11]) ? 4'b1001 : node42;
															assign node42 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node46 = (inp[10]) ? node54 : node47;
														assign node47 = (inp[1]) ? node49 : 4'b0000;
															assign node49 = (inp[14]) ? node51 : 4'b0001;
																assign node51 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node54 = (inp[11]) ? 4'b1001 : node55;
															assign node55 = (inp[14]) ? 4'b0001 : 4'b1000;
										assign node60 = (inp[13]) ? node100 : node61;
											assign node61 = (inp[10]) ? node87 : node62;
												assign node62 = (inp[12]) ? node76 : node63;
													assign node63 = (inp[1]) ? node71 : node64;
														assign node64 = (inp[11]) ? 4'b0000 : node65;
															assign node65 = (inp[14]) ? node67 : 4'b0000;
																assign node67 = (inp[7]) ? 4'b1111 : 4'b1001;
														assign node71 = (inp[11]) ? 4'b0001 : node72;
															assign node72 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node76 = (inp[7]) ? 4'b1111 : node77;
														assign node77 = (inp[14]) ? node79 : 4'b1001;
															assign node79 = (inp[1]) ? node83 : node80;
																assign node80 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node83 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node87 = (inp[1]) ? node95 : node88;
													assign node88 = (inp[14]) ? node90 : 4'b0000;
														assign node90 = (inp[11]) ? 4'b0000 : node91;
															assign node91 = (inp[12]) ? 4'b1111 : 4'b0001;
													assign node95 = (inp[11]) ? 4'b0001 : node96;
														assign node96 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node100 = (inp[1]) ? node118 : node101;
												assign node101 = (inp[14]) ? node107 : node102;
													assign node102 = (inp[12]) ? node104 : 4'b1000;
														assign node104 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node107 = (inp[11]) ? node113 : node108;
														assign node108 = (inp[12]) ? 4'b0001 : node109;
															assign node109 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node113 = (inp[12]) ? node115 : 4'b1000;
															assign node115 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node118 = (inp[14]) ? node124 : node119;
													assign node119 = (inp[10]) ? 4'b1001 : node120;
														assign node120 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node124 = (inp[11]) ? node130 : node125;
														assign node125 = (inp[12]) ? node127 : 4'b1000;
															assign node127 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node130 = (inp[12]) ? node132 : 4'b1001;
															assign node132 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node135 = (inp[4]) ? node267 : node136;
										assign node136 = (inp[7]) ? node198 : node137;
											assign node137 = (inp[1]) ? node167 : node138;
												assign node138 = (inp[14]) ? node150 : node139;
													assign node139 = (inp[13]) ? node145 : node140;
														assign node140 = (inp[12]) ? node142 : 4'b0100;
															assign node142 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node145 = (inp[10]) ? 4'b1100 : node146;
															assign node146 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node150 = (inp[11]) ? node160 : node151;
														assign node151 = (inp[13]) ? node157 : node152;
															assign node152 = (inp[10]) ? node154 : 4'b1001;
																assign node154 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node157 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node160 = (inp[13]) ? 4'b1100 : node161;
															assign node161 = (inp[10]) ? 4'b0100 : node162;
																assign node162 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node167 = (inp[13]) ? node185 : node168;
													assign node168 = (inp[12]) ? node174 : node169;
														assign node169 = (inp[11]) ? 4'b0101 : node170;
															assign node170 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node174 = (inp[10]) ? node180 : node175;
															assign node175 = (inp[14]) ? node177 : 4'b1001;
																assign node177 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node180 = (inp[14]) ? node182 : 4'b0101;
																assign node182 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node185 = (inp[12]) ? node191 : node186;
														assign node186 = (inp[11]) ? 4'b1101 : node187;
															assign node187 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node191 = (inp[10]) ? node193 : 4'b0101;
															assign node193 = (inp[14]) ? node195 : 4'b1101;
																assign node195 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node198 = (inp[1]) ? node232 : node199;
												assign node199 = (inp[11]) ? node221 : node200;
													assign node200 = (inp[14]) ? node210 : node201;
														assign node201 = (inp[13]) ? node207 : node202;
															assign node202 = (inp[12]) ? node204 : 4'b0000;
																assign node204 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node207 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node210 = (inp[13]) ? node216 : node211;
															assign node211 = (inp[12]) ? 4'b1001 : node212;
																assign node212 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node216 = (inp[12]) ? 4'b0001 : node217;
																assign node217 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node221 = (inp[13]) ? node227 : node222;
														assign node222 = (inp[12]) ? node224 : 4'b0000;
															assign node224 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node227 = (inp[10]) ? 4'b1000 : node228;
															assign node228 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node232 = (inp[14]) ? node244 : node233;
													assign node233 = (inp[13]) ? node239 : node234;
														assign node234 = (inp[10]) ? 4'b0001 : node235;
															assign node235 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node239 = (inp[12]) ? node241 : 4'b1001;
															assign node241 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node244 = (inp[11]) ? node256 : node245;
														assign node245 = (inp[13]) ? node251 : node246;
															assign node246 = (inp[10]) ? 4'b0000 : node247;
																assign node247 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node251 = (inp[10]) ? 4'b1000 : node252;
																assign node252 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node256 = (inp[13]) ? node262 : node257;
															assign node257 = (inp[12]) ? node259 : 4'b0001;
																assign node259 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node262 = (inp[10]) ? 4'b1001 : node263;
																assign node263 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node267 = (inp[1]) ? node307 : node268;
											assign node268 = (inp[11]) ? node294 : node269;
												assign node269 = (inp[14]) ? node277 : node270;
													assign node270 = (inp[13]) ? node272 : 4'b0100;
														assign node272 = (inp[10]) ? 4'b1100 : node273;
															assign node273 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node277 = (inp[13]) ? node289 : node278;
														assign node278 = (inp[7]) ? node284 : node279;
															assign node279 = (inp[12]) ? 4'b1101 : node280;
																assign node280 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node284 = (inp[10]) ? node286 : 4'b1001;
																assign node286 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node289 = (inp[12]) ? 4'b0101 : node290;
															assign node290 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node294 = (inp[13]) ? node302 : node295;
													assign node295 = (inp[10]) ? 4'b0100 : node296;
														assign node296 = (inp[12]) ? node298 : 4'b0100;
															assign node298 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node302 = (inp[10]) ? 4'b1100 : node303;
														assign node303 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node307 = (inp[13]) ? node331 : node308;
												assign node308 = (inp[12]) ? node314 : node309;
													assign node309 = (inp[14]) ? node311 : 4'b0101;
														assign node311 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node314 = (inp[10]) ? node326 : node315;
														assign node315 = (inp[7]) ? node321 : node316;
															assign node316 = (inp[14]) ? node318 : 4'b1101;
																assign node318 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node321 = (inp[14]) ? node323 : 4'b1001;
																assign node323 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node326 = (inp[14]) ? node328 : 4'b0101;
															assign node328 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node331 = (inp[11]) ? node343 : node332;
													assign node332 = (inp[14]) ? node338 : node333;
														assign node333 = (inp[12]) ? node335 : 4'b1101;
															assign node335 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node338 = (inp[10]) ? 4'b1100 : node339;
															assign node339 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node343 = (inp[12]) ? node345 : 4'b1101;
														assign node345 = (inp[10]) ? 4'b1101 : 4'b0101;
							assign node349 = (inp[1]) ? node595 : node350;
								assign node350 = (inp[11]) ? node516 : node351;
									assign node351 = (inp[14]) ? node431 : node352;
										assign node352 = (inp[13]) ? node398 : node353;
											assign node353 = (inp[10]) ? node385 : node354;
												assign node354 = (inp[12]) ? node368 : node355;
													assign node355 = (inp[3]) ? node363 : node356;
														assign node356 = (inp[7]) ? node358 : 4'b0000;
															assign node358 = (inp[4]) ? 4'b0000 : node359;
																assign node359 = (inp[2]) ? 4'b1111 : 4'b0100;
														assign node363 = (inp[4]) ? 4'b0100 : node364;
															assign node364 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node368 = (inp[3]) ? node380 : node369;
														assign node369 = (inp[2]) ? node375 : node370;
															assign node370 = (inp[4]) ? node372 : 4'b1100;
																assign node372 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node375 = (inp[4]) ? node377 : 4'b1111;
																assign node377 = (inp[7]) ? 4'b1111 : 4'b1000;
														assign node380 = (inp[4]) ? node382 : 4'b1000;
															assign node382 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node385 = (inp[3]) ? node393 : node386;
													assign node386 = (inp[4]) ? 4'b0000 : node387;
														assign node387 = (inp[7]) ? node389 : 4'b0000;
															assign node389 = (inp[2]) ? 4'b1111 : 4'b0100;
													assign node393 = (inp[4]) ? 4'b0100 : node394;
														assign node394 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node398 = (inp[3]) ? node418 : node399;
												assign node399 = (inp[4]) ? node413 : node400;
													assign node400 = (inp[7]) ? node406 : node401;
														assign node401 = (inp[10]) ? 4'b1000 : node402;
															assign node402 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node406 = (inp[2]) ? 4'b1111 : node407;
															assign node407 = (inp[10]) ? 4'b1100 : node408;
																assign node408 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node413 = (inp[12]) ? node415 : 4'b1000;
														assign node415 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node418 = (inp[4]) ? node426 : node419;
													assign node419 = (inp[7]) ? node421 : 4'b1100;
														assign node421 = (inp[10]) ? 4'b1000 : node422;
															assign node422 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node426 = (inp[10]) ? 4'b1100 : node427;
														assign node427 = (inp[12]) ? 4'b0100 : 4'b1100;
										assign node431 = (inp[13]) ? node477 : node432;
											assign node432 = (inp[10]) ? node450 : node433;
												assign node433 = (inp[3]) ? node445 : node434;
													assign node434 = (inp[2]) ? node440 : node435;
														assign node435 = (inp[7]) ? 4'b1101 : node436;
															assign node436 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node440 = (inp[4]) ? node442 : 4'b1111;
															assign node442 = (inp[7]) ? 4'b1111 : 4'b1001;
													assign node445 = (inp[4]) ? node447 : 4'b1001;
														assign node447 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node450 = (inp[12]) ? node466 : node451;
													assign node451 = (inp[3]) ? node459 : node452;
														assign node452 = (inp[7]) ? node454 : 4'b0001;
															assign node454 = (inp[4]) ? 4'b0001 : node455;
																assign node455 = (inp[2]) ? 4'b1111 : 4'b0101;
														assign node459 = (inp[2]) ? node461 : 4'b0101;
															assign node461 = (inp[4]) ? 4'b0101 : node462;
																assign node462 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node466 = (inp[3]) ? node474 : node467;
														assign node467 = (inp[7]) ? node471 : node468;
															assign node468 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node471 = (inp[2]) ? 4'b1111 : 4'b1101;
														assign node474 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node477 = (inp[12]) ? node503 : node478;
												assign node478 = (inp[10]) ? node490 : node479;
													assign node479 = (inp[3]) ? node485 : node480;
														assign node480 = (inp[7]) ? node482 : 4'b0001;
															assign node482 = (inp[2]) ? 4'b1111 : 4'b0101;
														assign node485 = (inp[7]) ? node487 : 4'b0101;
															assign node487 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node490 = (inp[3]) ? node498 : node491;
														assign node491 = (inp[7]) ? node493 : 4'b1001;
															assign node493 = (inp[4]) ? 4'b1001 : node494;
																assign node494 = (inp[2]) ? 4'b1111 : 4'b1101;
														assign node498 = (inp[7]) ? node500 : 4'b1101;
															assign node500 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node503 = (inp[3]) ? node511 : node504;
													assign node504 = (inp[7]) ? node506 : 4'b0001;
														assign node506 = (inp[4]) ? 4'b0001 : node507;
															assign node507 = (inp[2]) ? 4'b1111 : 4'b0101;
													assign node511 = (inp[7]) ? node513 : 4'b0101;
														assign node513 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node516 = (inp[3]) ? node560 : node517;
										assign node517 = (inp[4]) ? node545 : node518;
											assign node518 = (inp[7]) ? node532 : node519;
												assign node519 = (inp[13]) ? node527 : node520;
													assign node520 = (inp[10]) ? 4'b0000 : node521;
														assign node521 = (inp[12]) ? node523 : 4'b0000;
															assign node523 = (inp[2]) ? 4'b1111 : 4'b1100;
													assign node527 = (inp[12]) ? node529 : 4'b1000;
														assign node529 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node532 = (inp[2]) ? 4'b1111 : node533;
													assign node533 = (inp[13]) ? node539 : node534;
														assign node534 = (inp[10]) ? 4'b0100 : node535;
															assign node535 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node539 = (inp[10]) ? 4'b1100 : node540;
															assign node540 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node545 = (inp[13]) ? node555 : node546;
												assign node546 = (inp[10]) ? 4'b0000 : node547;
													assign node547 = (inp[12]) ? node549 : 4'b0000;
														assign node549 = (inp[7]) ? node551 : 4'b1000;
															assign node551 = (inp[2]) ? 4'b1111 : 4'b1100;
												assign node555 = (inp[10]) ? 4'b1000 : node556;
													assign node556 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node560 = (inp[13]) ? node578 : node561;
											assign node561 = (inp[12]) ? node567 : node562;
												assign node562 = (inp[7]) ? node564 : 4'b0100;
													assign node564 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node567 = (inp[10]) ? node573 : node568;
													assign node568 = (inp[7]) ? 4'b1000 : node569;
														assign node569 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node573 = (inp[7]) ? node575 : 4'b0100;
														assign node575 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node578 = (inp[10]) ? node590 : node579;
												assign node579 = (inp[12]) ? node585 : node580;
													assign node580 = (inp[7]) ? node582 : 4'b1100;
														assign node582 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node585 = (inp[7]) ? node587 : 4'b0100;
														assign node587 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node590 = (inp[7]) ? node592 : 4'b1100;
													assign node592 = (inp[4]) ? 4'b1100 : 4'b1000;
								assign node595 = (inp[13]) ? node709 : node596;
									assign node596 = (inp[10]) ? node672 : node597;
										assign node597 = (inp[12]) ? node635 : node598;
											assign node598 = (inp[3]) ? node618 : node599;
												assign node599 = (inp[4]) ? node613 : node600;
													assign node600 = (inp[7]) ? node606 : node601;
														assign node601 = (inp[11]) ? 4'b0001 : node602;
															assign node602 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node606 = (inp[2]) ? 4'b1111 : node607;
															assign node607 = (inp[11]) ? 4'b0101 : node608;
																assign node608 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node613 = (inp[11]) ? 4'b0001 : node614;
														assign node614 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node618 = (inp[7]) ? node624 : node619;
													assign node619 = (inp[11]) ? 4'b0101 : node620;
														assign node620 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node624 = (inp[4]) ? node630 : node625;
														assign node625 = (inp[11]) ? 4'b0001 : node626;
															assign node626 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node630 = (inp[11]) ? 4'b0101 : node631;
															assign node631 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node635 = (inp[3]) ? node655 : node636;
												assign node636 = (inp[2]) ? node646 : node637;
													assign node637 = (inp[14]) ? node643 : node638;
														assign node638 = (inp[7]) ? 4'b1101 : node639;
															assign node639 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node643 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node646 = (inp[4]) ? node648 : 4'b1111;
														assign node648 = (inp[7]) ? 4'b1111 : node649;
															assign node649 = (inp[14]) ? node651 : 4'b1001;
																assign node651 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node655 = (inp[14]) ? node661 : node656;
													assign node656 = (inp[4]) ? node658 : 4'b1001;
														assign node658 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node661 = (inp[11]) ? node667 : node662;
														assign node662 = (inp[4]) ? node664 : 4'b1000;
															assign node664 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node667 = (inp[7]) ? 4'b1001 : node668;
															assign node668 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node672 = (inp[3]) ? node692 : node673;
											assign node673 = (inp[7]) ? node679 : node674;
												assign node674 = (inp[11]) ? 4'b0001 : node675;
													assign node675 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node679 = (inp[4]) ? node687 : node680;
													assign node680 = (inp[2]) ? 4'b1111 : node681;
														assign node681 = (inp[11]) ? 4'b0101 : node682;
															assign node682 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node687 = (inp[14]) ? node689 : 4'b0001;
														assign node689 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node692 = (inp[7]) ? node698 : node693;
												assign node693 = (inp[14]) ? node695 : 4'b0101;
													assign node695 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node698 = (inp[4]) ? node704 : node699;
													assign node699 = (inp[14]) ? node701 : 4'b0001;
														assign node701 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node704 = (inp[11]) ? 4'b0101 : node705;
														assign node705 = (inp[14]) ? 4'b0100 : 4'b0101;
									assign node709 = (inp[3]) ? node755 : node710;
										assign node710 = (inp[7]) ? node728 : node711;
											assign node711 = (inp[10]) ? node723 : node712;
												assign node712 = (inp[12]) ? node718 : node713;
													assign node713 = (inp[14]) ? node715 : 4'b1001;
														assign node715 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node718 = (inp[11]) ? 4'b0001 : node719;
														assign node719 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node723 = (inp[14]) ? node725 : 4'b1001;
													assign node725 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node728 = (inp[4]) ? node740 : node729;
												assign node729 = (inp[2]) ? 4'b1111 : node730;
													assign node730 = (inp[10]) ? node734 : node731;
														assign node731 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node734 = (inp[14]) ? node736 : 4'b1101;
															assign node736 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node740 = (inp[14]) ? node746 : node741;
													assign node741 = (inp[10]) ? 4'b1001 : node742;
														assign node742 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node746 = (inp[11]) ? node752 : node747;
														assign node747 = (inp[12]) ? node749 : 4'b1000;
															assign node749 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node752 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node755 = (inp[7]) ? node773 : node756;
											assign node756 = (inp[12]) ? node762 : node757;
												assign node757 = (inp[14]) ? node759 : 4'b1101;
													assign node759 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node762 = (inp[10]) ? node768 : node763;
													assign node763 = (inp[11]) ? 4'b0101 : node764;
														assign node764 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node768 = (inp[11]) ? 4'b1101 : node769;
														assign node769 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node773 = (inp[4]) ? node791 : node774;
												assign node774 = (inp[12]) ? node780 : node775;
													assign node775 = (inp[14]) ? node777 : 4'b1001;
														assign node777 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node780 = (inp[10]) ? node786 : node781;
														assign node781 = (inp[14]) ? node783 : 4'b0001;
															assign node783 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node786 = (inp[11]) ? 4'b1001 : node787;
															assign node787 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node791 = (inp[12]) ? node797 : node792;
													assign node792 = (inp[11]) ? 4'b1101 : node793;
														assign node793 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node797 = (inp[10]) ? node803 : node798;
														assign node798 = (inp[11]) ? 4'b0101 : node799;
															assign node799 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node803 = (inp[11]) ? 4'b1101 : node804;
															assign node804 = (inp[14]) ? 4'b1100 : 4'b1101;
					assign node809 = (inp[0]) ? 4'b1001 : node810;
						assign node810 = (inp[5]) ? node956 : node811;
							assign node811 = (inp[3]) ? node813 : 4'b1011;
								assign node813 = (inp[2]) ? 4'b1011 : node814;
									assign node814 = (inp[7]) ? node898 : node815;
										assign node815 = (inp[1]) ? node861 : node816;
											assign node816 = (inp[14]) ? node830 : node817;
												assign node817 = (inp[13]) ? node825 : node818;
													assign node818 = (inp[10]) ? 4'b0000 : node819;
														assign node819 = (inp[12]) ? node821 : 4'b0000;
															assign node821 = (inp[4]) ? 4'b1000 : 4'b1011;
													assign node825 = (inp[12]) ? node827 : 4'b1000;
														assign node827 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node830 = (inp[11]) ? node848 : node831;
													assign node831 = (inp[13]) ? node843 : node832;
														assign node832 = (inp[4]) ? node838 : node833;
															assign node833 = (inp[10]) ? node835 : 4'b1011;
																assign node835 = (inp[12]) ? 4'b1011 : 4'b0001;
															assign node838 = (inp[12]) ? 4'b1001 : node839;
																assign node839 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node843 = (inp[12]) ? 4'b0001 : node844;
															assign node844 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node848 = (inp[13]) ? node856 : node849;
														assign node849 = (inp[12]) ? node851 : 4'b0000;
															assign node851 = (inp[4]) ? node853 : 4'b1011;
																assign node853 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node856 = (inp[12]) ? node858 : 4'b1000;
															assign node858 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node861 = (inp[13]) ? node881 : node862;
												assign node862 = (inp[12]) ? node868 : node863;
													assign node863 = (inp[14]) ? node865 : 4'b0001;
														assign node865 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node868 = (inp[10]) ? node876 : node869;
														assign node869 = (inp[4]) ? node871 : 4'b1011;
															assign node871 = (inp[14]) ? node873 : 4'b1001;
																assign node873 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node876 = (inp[14]) ? node878 : 4'b0001;
															assign node878 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node881 = (inp[11]) ? node893 : node882;
													assign node882 = (inp[14]) ? node888 : node883;
														assign node883 = (inp[10]) ? 4'b1001 : node884;
															assign node884 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node888 = (inp[10]) ? 4'b1000 : node889;
															assign node889 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node893 = (inp[12]) ? node895 : 4'b1001;
														assign node895 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node898 = (inp[4]) ? node900 : 4'b1011;
											assign node900 = (inp[13]) ? node926 : node901;
												assign node901 = (inp[12]) ? node915 : node902;
													assign node902 = (inp[1]) ? node910 : node903;
														assign node903 = (inp[11]) ? 4'b0000 : node904;
															assign node904 = (inp[14]) ? node906 : 4'b0000;
																assign node906 = (inp[10]) ? 4'b0001 : 4'b1011;
														assign node910 = (inp[14]) ? node912 : 4'b0001;
															assign node912 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node915 = (inp[10]) ? node917 : 4'b1011;
														assign node917 = (inp[1]) ? node921 : node918;
															assign node918 = (inp[14]) ? 4'b1011 : 4'b0000;
															assign node921 = (inp[11]) ? 4'b0001 : node922;
																assign node922 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node926 = (inp[10]) ? node946 : node927;
													assign node927 = (inp[12]) ? node937 : node928;
														assign node928 = (inp[1]) ? node932 : node929;
															assign node929 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node932 = (inp[14]) ? node934 : 4'b1001;
																assign node934 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node937 = (inp[11]) ? 4'b0001 : node938;
															assign node938 = (inp[14]) ? node942 : node939;
																assign node939 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node942 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node946 = (inp[1]) ? node952 : node947;
														assign node947 = (inp[11]) ? 4'b1000 : node948;
															assign node948 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node952 = (inp[14]) ? 4'b1000 : 4'b1001;
							assign node956 = (inp[2]) ? node1334 : node957;
								assign node957 = (inp[1]) ? node1159 : node958;
									assign node958 = (inp[11]) ? node1088 : node959;
										assign node959 = (inp[14]) ? node1021 : node960;
											assign node960 = (inp[13]) ? node988 : node961;
												assign node961 = (inp[10]) ? node977 : node962;
													assign node962 = (inp[12]) ? node970 : node963;
														assign node963 = (inp[3]) ? 4'b0000 : node964;
															assign node964 = (inp[4]) ? 4'b0100 : node965;
																assign node965 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node970 = (inp[3]) ? 4'b1100 : node971;
															assign node971 = (inp[7]) ? 4'b1000 : node972;
																assign node972 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node977 = (inp[3]) ? node983 : node978;
														assign node978 = (inp[7]) ? node980 : 4'b0100;
															assign node980 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node983 = (inp[4]) ? 4'b0000 : node984;
															assign node984 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node988 = (inp[12]) ? node1000 : node989;
													assign node989 = (inp[3]) ? node995 : node990;
														assign node990 = (inp[7]) ? node992 : 4'b1100;
															assign node992 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node995 = (inp[4]) ? 4'b1000 : node996;
															assign node996 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node1000 = (inp[10]) ? node1012 : node1001;
														assign node1001 = (inp[3]) ? node1007 : node1002;
															assign node1002 = (inp[7]) ? node1004 : 4'b0100;
																assign node1004 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node1007 = (inp[7]) ? node1009 : 4'b0000;
																assign node1009 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1012 = (inp[7]) ? node1014 : 4'b1100;
															assign node1014 = (inp[4]) ? node1018 : node1015;
																assign node1015 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node1018 = (inp[3]) ? 4'b1000 : 4'b1100;
											assign node1021 = (inp[13]) ? node1055 : node1022;
												assign node1022 = (inp[10]) ? node1034 : node1023;
													assign node1023 = (inp[3]) ? node1029 : node1024;
														assign node1024 = (inp[7]) ? 4'b1001 : node1025;
															assign node1025 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node1029 = (inp[7]) ? 4'b1101 : node1030;
															assign node1030 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node1034 = (inp[12]) ? node1046 : node1035;
														assign node1035 = (inp[3]) ? node1041 : node1036;
															assign node1036 = (inp[4]) ? 4'b0101 : node1037;
																assign node1037 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node1041 = (inp[4]) ? 4'b0001 : node1042;
																assign node1042 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node1046 = (inp[3]) ? node1052 : node1047;
															assign node1047 = (inp[7]) ? 4'b1001 : node1048;
																assign node1048 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node1052 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node1055 = (inp[10]) ? node1067 : node1056;
													assign node1056 = (inp[3]) ? node1062 : node1057;
														assign node1057 = (inp[7]) ? node1059 : 4'b0101;
															assign node1059 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node1062 = (inp[4]) ? 4'b0001 : node1063;
															assign node1063 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node1067 = (inp[12]) ? node1079 : node1068;
														assign node1068 = (inp[3]) ? node1074 : node1069;
															assign node1069 = (inp[4]) ? 4'b1101 : node1070;
																assign node1070 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node1074 = (inp[4]) ? 4'b1001 : node1075;
																assign node1075 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1079 = (inp[3]) ? node1083 : node1080;
															assign node1080 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node1083 = (inp[4]) ? 4'b0001 : node1084;
																assign node1084 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node1088 = (inp[13]) ? node1124 : node1089;
											assign node1089 = (inp[10]) ? node1113 : node1090;
												assign node1090 = (inp[12]) ? node1102 : node1091;
													assign node1091 = (inp[3]) ? node1097 : node1092;
														assign node1092 = (inp[4]) ? 4'b0100 : node1093;
															assign node1093 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1097 = (inp[4]) ? 4'b0000 : node1098;
															assign node1098 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1102 = (inp[3]) ? node1108 : node1103;
														assign node1103 = (inp[7]) ? 4'b1000 : node1104;
															assign node1104 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1108 = (inp[7]) ? 4'b1100 : node1109;
															assign node1109 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node1113 = (inp[3]) ? node1119 : node1114;
													assign node1114 = (inp[4]) ? 4'b0100 : node1115;
														assign node1115 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node1119 = (inp[4]) ? 4'b0000 : node1120;
														assign node1120 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node1124 = (inp[12]) ? node1136 : node1125;
												assign node1125 = (inp[3]) ? node1131 : node1126;
													assign node1126 = (inp[4]) ? 4'b1100 : node1127;
														assign node1127 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node1131 = (inp[7]) ? node1133 : 4'b1000;
														assign node1133 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node1136 = (inp[10]) ? node1148 : node1137;
													assign node1137 = (inp[3]) ? node1143 : node1138;
														assign node1138 = (inp[4]) ? 4'b0100 : node1139;
															assign node1139 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1143 = (inp[4]) ? 4'b0000 : node1144;
															assign node1144 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1148 = (inp[3]) ? node1154 : node1149;
														assign node1149 = (inp[4]) ? 4'b1100 : node1150;
															assign node1150 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node1154 = (inp[4]) ? 4'b1000 : node1155;
															assign node1155 = (inp[7]) ? 4'b1100 : 4'b1000;
									assign node1159 = (inp[14]) ? node1219 : node1160;
										assign node1160 = (inp[13]) ? node1192 : node1161;
											assign node1161 = (inp[10]) ? node1181 : node1162;
												assign node1162 = (inp[12]) ? node1170 : node1163;
													assign node1163 = (inp[3]) ? node1165 : 4'b0101;
														assign node1165 = (inp[4]) ? 4'b0001 : node1166;
															assign node1166 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node1170 = (inp[3]) ? node1176 : node1171;
														assign node1171 = (inp[4]) ? node1173 : 4'b1001;
															assign node1173 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1176 = (inp[4]) ? node1178 : 4'b1101;
															assign node1178 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node1181 = (inp[3]) ? node1187 : node1182;
													assign node1182 = (inp[4]) ? 4'b0101 : node1183;
														assign node1183 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1187 = (inp[7]) ? node1189 : 4'b0001;
														assign node1189 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node1192 = (inp[3]) ? node1206 : node1193;
												assign node1193 = (inp[4]) ? node1201 : node1194;
													assign node1194 = (inp[7]) ? node1196 : 4'b1101;
														assign node1196 = (inp[12]) ? node1198 : 4'b1001;
															assign node1198 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node1201 = (inp[10]) ? 4'b1101 : node1202;
														assign node1202 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node1206 = (inp[7]) ? node1212 : node1207;
													assign node1207 = (inp[10]) ? 4'b1001 : node1208;
														assign node1208 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1212 = (inp[4]) ? node1214 : 4'b1101;
														assign node1214 = (inp[10]) ? 4'b1001 : node1215;
															assign node1215 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node1219 = (inp[11]) ? node1277 : node1220;
											assign node1220 = (inp[13]) ? node1252 : node1221;
												assign node1221 = (inp[12]) ? node1233 : node1222;
													assign node1222 = (inp[3]) ? node1228 : node1223;
														assign node1223 = (inp[4]) ? 4'b0100 : node1224;
															assign node1224 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node1228 = (inp[4]) ? 4'b0000 : node1229;
															assign node1229 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node1233 = (inp[10]) ? node1245 : node1234;
														assign node1234 = (inp[3]) ? node1240 : node1235;
															assign node1235 = (inp[4]) ? node1237 : 4'b1000;
																assign node1237 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node1240 = (inp[7]) ? 4'b1100 : node1241;
																assign node1241 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node1245 = (inp[3]) ? node1249 : node1246;
															assign node1246 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node1249 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node1252 = (inp[3]) ? node1266 : node1253;
													assign node1253 = (inp[12]) ? node1259 : node1254;
														assign node1254 = (inp[7]) ? node1256 : 4'b1100;
															assign node1256 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1259 = (inp[10]) ? 4'b1100 : node1260;
															assign node1260 = (inp[7]) ? node1262 : 4'b0100;
																assign node1262 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node1266 = (inp[10]) ? node1272 : node1267;
														assign node1267 = (inp[12]) ? 4'b0000 : node1268;
															assign node1268 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node1272 = (inp[4]) ? 4'b1000 : node1273;
															assign node1273 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node1277 = (inp[3]) ? node1301 : node1278;
												assign node1278 = (inp[13]) ? node1290 : node1279;
													assign node1279 = (inp[10]) ? 4'b0101 : node1280;
														assign node1280 = (inp[12]) ? node1284 : node1281;
															assign node1281 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node1284 = (inp[4]) ? node1286 : 4'b1001;
																assign node1286 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node1290 = (inp[10]) ? node1296 : node1291;
														assign node1291 = (inp[12]) ? 4'b0101 : node1292;
															assign node1292 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1296 = (inp[7]) ? node1298 : 4'b1101;
															assign node1298 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node1301 = (inp[4]) ? node1321 : node1302;
													assign node1302 = (inp[7]) ? node1312 : node1303;
														assign node1303 = (inp[13]) ? node1307 : node1304;
															assign node1304 = (inp[10]) ? 4'b0001 : 4'b1101;
															assign node1307 = (inp[10]) ? 4'b1001 : node1308;
																assign node1308 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node1312 = (inp[12]) ? node1314 : 4'b1101;
															assign node1314 = (inp[13]) ? node1318 : node1315;
																assign node1315 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node1318 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node1321 = (inp[13]) ? node1329 : node1322;
														assign node1322 = (inp[12]) ? node1324 : 4'b0001;
															assign node1324 = (inp[10]) ? 4'b0001 : node1325;
																assign node1325 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node1329 = (inp[10]) ? 4'b1001 : node1330;
															assign node1330 = (inp[12]) ? 4'b0001 : 4'b1001;
								assign node1334 = (inp[3]) ? node1336 : 4'b1011;
									assign node1336 = (inp[7]) ? node1418 : node1337;
										assign node1337 = (inp[1]) ? node1383 : node1338;
											assign node1338 = (inp[11]) ? node1370 : node1339;
												assign node1339 = (inp[14]) ? node1353 : node1340;
													assign node1340 = (inp[13]) ? node1348 : node1341;
														assign node1341 = (inp[10]) ? 4'b0000 : node1342;
															assign node1342 = (inp[12]) ? node1344 : 4'b0000;
																assign node1344 = (inp[4]) ? 4'b1000 : 4'b1011;
														assign node1348 = (inp[10]) ? 4'b1000 : node1349;
															assign node1349 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node1353 = (inp[13]) ? node1365 : node1354;
														assign node1354 = (inp[4]) ? node1360 : node1355;
															assign node1355 = (inp[10]) ? node1357 : 4'b1011;
																assign node1357 = (inp[12]) ? 4'b1011 : 4'b0001;
															assign node1360 = (inp[12]) ? 4'b1001 : node1361;
																assign node1361 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node1365 = (inp[12]) ? 4'b0001 : node1366;
															assign node1366 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node1370 = (inp[13]) ? node1378 : node1371;
													assign node1371 = (inp[10]) ? 4'b0000 : node1372;
														assign node1372 = (inp[12]) ? node1374 : 4'b0000;
															assign node1374 = (inp[4]) ? 4'b1000 : 4'b1011;
													assign node1378 = (inp[12]) ? node1380 : 4'b1000;
														assign node1380 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node1383 = (inp[13]) ? node1401 : node1384;
												assign node1384 = (inp[12]) ? node1390 : node1385;
													assign node1385 = (inp[14]) ? node1387 : 4'b0001;
														assign node1387 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1390 = (inp[10]) ? node1398 : node1391;
														assign node1391 = (inp[4]) ? node1393 : 4'b1011;
															assign node1393 = (inp[11]) ? 4'b1001 : node1394;
																assign node1394 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1398 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node1401 = (inp[14]) ? node1407 : node1402;
													assign node1402 = (inp[10]) ? 4'b1001 : node1403;
														assign node1403 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node1407 = (inp[11]) ? node1413 : node1408;
														assign node1408 = (inp[12]) ? node1410 : 4'b1000;
															assign node1410 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node1413 = (inp[10]) ? 4'b1001 : node1414;
															assign node1414 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node1418 = (inp[4]) ? node1420 : 4'b1011;
											assign node1420 = (inp[13]) ? node1442 : node1421;
												assign node1421 = (inp[10]) ? node1435 : node1422;
													assign node1422 = (inp[12]) ? 4'b1011 : node1423;
														assign node1423 = (inp[1]) ? node1429 : node1424;
															assign node1424 = (inp[14]) ? node1426 : 4'b0000;
																assign node1426 = (inp[11]) ? 4'b0000 : 4'b1011;
															assign node1429 = (inp[14]) ? node1431 : 4'b0001;
																assign node1431 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node1435 = (inp[1]) ? node1437 : 4'b0000;
														assign node1437 = (inp[14]) ? node1439 : 4'b0001;
															assign node1439 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node1442 = (inp[1]) ? node1460 : node1443;
													assign node1443 = (inp[10]) ? node1455 : node1444;
														assign node1444 = (inp[12]) ? node1450 : node1445;
															assign node1445 = (inp[11]) ? 4'b1000 : node1446;
																assign node1446 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node1450 = (inp[11]) ? 4'b0000 : node1451;
																assign node1451 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node1455 = (inp[14]) ? node1457 : 4'b1000;
															assign node1457 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node1460 = (inp[12]) ? node1466 : node1461;
														assign node1461 = (inp[11]) ? 4'b1001 : node1462;
															assign node1462 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node1466 = (inp[10]) ? 4'b1001 : node1467;
															assign node1467 = (inp[14]) ? node1469 : 4'b0001;
																assign node1469 = (inp[11]) ? 4'b0001 : 4'b0000;
				assign node1474 = (inp[5]) ? node3638 : node1475;
					assign node1475 = (inp[0]) ? node3161 : node1476;
						assign node1476 = (inp[11]) ? node2532 : node1477;
							assign node1477 = (inp[10]) ? node2027 : node1478;
								assign node1478 = (inp[12]) ? node1708 : node1479;
									assign node1479 = (inp[3]) ? node1611 : node1480;
										assign node1480 = (inp[2]) ? node1534 : node1481;
											assign node1481 = (inp[15]) ? node1497 : node1482;
												assign node1482 = (inp[4]) ? node1492 : node1483;
													assign node1483 = (inp[7]) ? node1485 : 4'b0000;
														assign node1485 = (inp[13]) ? 4'b0000 : node1486;
															assign node1486 = (inp[14]) ? node1488 : 4'b0100;
																assign node1488 = (inp[1]) ? 4'b0100 : 4'b1101;
													assign node1492 = (inp[7]) ? node1494 : 4'b0100;
														assign node1494 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node1497 = (inp[4]) ? node1523 : node1498;
													assign node1498 = (inp[7]) ? node1510 : node1499;
														assign node1499 = (inp[13]) ? node1505 : node1500;
															assign node1500 = (inp[14]) ? 4'b1001 : node1501;
																assign node1501 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node1505 = (inp[1]) ? node1507 : 4'b1100;
																assign node1507 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node1510 = (inp[13]) ? node1516 : node1511;
															assign node1511 = (inp[1]) ? node1513 : 4'b1001;
																assign node1513 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node1516 = (inp[1]) ? node1520 : node1517;
																assign node1517 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node1520 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node1523 = (inp[7]) ? node1525 : 4'b0000;
														assign node1525 = (inp[13]) ? 4'b0000 : node1526;
															assign node1526 = (inp[14]) ? node1530 : node1527;
																assign node1527 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node1530 = (inp[1]) ? 4'b0100 : 4'b1001;
											assign node1534 = (inp[13]) ? node1570 : node1535;
												assign node1535 = (inp[1]) ? node1551 : node1536;
													assign node1536 = (inp[14]) ? node1544 : node1537;
														assign node1537 = (inp[15]) ? 4'b0100 : node1538;
															assign node1538 = (inp[7]) ? node1540 : 4'b0000;
																assign node1540 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1544 = (inp[15]) ? node1546 : 4'b1101;
															assign node1546 = (inp[7]) ? 4'b1001 : node1547;
																assign node1547 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node1551 = (inp[14]) ? node1559 : node1552;
														assign node1552 = (inp[15]) ? 4'b0101 : node1553;
															assign node1553 = (inp[7]) ? node1555 : 4'b0001;
																assign node1555 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1559 = (inp[15]) ? node1565 : node1560;
															assign node1560 = (inp[4]) ? 4'b0000 : node1561;
																assign node1561 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node1565 = (inp[4]) ? 4'b0100 : node1566;
																assign node1566 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node1570 = (inp[1]) ? node1590 : node1571;
													assign node1571 = (inp[14]) ? node1579 : node1572;
														assign node1572 = (inp[15]) ? node1574 : 4'b1000;
															assign node1574 = (inp[7]) ? node1576 : 4'b1100;
																assign node1576 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1579 = (inp[15]) ? node1585 : node1580;
															assign node1580 = (inp[7]) ? node1582 : 4'b0001;
																assign node1582 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node1585 = (inp[4]) ? 4'b0101 : node1586;
																assign node1586 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node1590 = (inp[14]) ? node1600 : node1591;
														assign node1591 = (inp[4]) ? node1597 : node1592;
															assign node1592 = (inp[7]) ? node1594 : 4'b1001;
																assign node1594 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node1597 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node1600 = (inp[15]) ? node1606 : node1601;
															assign node1601 = (inp[4]) ? 4'b1000 : node1602;
																assign node1602 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1606 = (inp[7]) ? node1608 : 4'b1100;
																assign node1608 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node1611 = (inp[15]) ? node1653 : node1612;
											assign node1612 = (inp[4]) ? node1626 : node1613;
												assign node1613 = (inp[7]) ? node1615 : 4'b0000;
													assign node1615 = (inp[2]) ? node1619 : node1616;
														assign node1616 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node1619 = (inp[13]) ? 4'b0000 : node1620;
															assign node1620 = (inp[14]) ? node1622 : 4'b0000;
																assign node1622 = (inp[1]) ? 4'b0000 : 4'b1001;
												assign node1626 = (inp[2]) ? node1648 : node1627;
													assign node1627 = (inp[13]) ? node1635 : node1628;
														assign node1628 = (inp[1]) ? node1632 : node1629;
															assign node1629 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node1632 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node1635 = (inp[7]) ? node1641 : node1636;
															assign node1636 = (inp[14]) ? node1638 : 4'b0100;
																assign node1638 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node1641 = (inp[14]) ? node1645 : node1642;
																assign node1642 = (inp[1]) ? 4'b0100 : 4'b1001;
																assign node1645 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node1648 = (inp[13]) ? 4'b0100 : node1649;
														assign node1649 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node1653 = (inp[4]) ? node1687 : node1654;
												assign node1654 = (inp[2]) ? node1660 : node1655;
													assign node1655 = (inp[7]) ? node1657 : 4'b0100;
														assign node1657 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node1660 = (inp[7]) ? node1674 : node1661;
														assign node1661 = (inp[13]) ? node1669 : node1662;
															assign node1662 = (inp[14]) ? node1666 : node1663;
																assign node1663 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node1666 = (inp[1]) ? 4'b0000 : 4'b1101;
															assign node1669 = (inp[1]) ? 4'b1000 : node1670;
																assign node1670 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node1674 = (inp[13]) ? node1682 : node1675;
															assign node1675 = (inp[14]) ? node1679 : node1676;
																assign node1676 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node1679 = (inp[1]) ? 4'b0100 : 4'b1101;
															assign node1682 = (inp[14]) ? 4'b0101 : node1683;
																assign node1683 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node1687 = (inp[13]) ? node1699 : node1688;
													assign node1688 = (inp[7]) ? node1690 : 4'b0000;
														assign node1690 = (inp[2]) ? node1692 : 4'b0100;
															assign node1692 = (inp[1]) ? node1696 : node1693;
																assign node1693 = (inp[14]) ? 4'b1101 : 4'b0000;
																assign node1696 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node1699 = (inp[2]) ? 4'b0000 : node1700;
														assign node1700 = (inp[7]) ? 4'b0000 : node1701;
															assign node1701 = (inp[1]) ? 4'b1001 : node1702;
																assign node1702 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node1708 = (inp[13]) ? node1850 : node1709;
										assign node1709 = (inp[1]) ? node1775 : node1710;
											assign node1710 = (inp[14]) ? node1742 : node1711;
												assign node1711 = (inp[4]) ? node1723 : node1712;
													assign node1712 = (inp[15]) ? node1718 : node1713;
														assign node1713 = (inp[3]) ? node1715 : 4'b1100;
															assign node1715 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node1718 = (inp[3]) ? node1720 : 4'b1000;
															assign node1720 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node1723 = (inp[15]) ? node1735 : node1724;
														assign node1724 = (inp[3]) ? node1730 : node1725;
															assign node1725 = (inp[2]) ? node1727 : 4'b1000;
																assign node1727 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1730 = (inp[7]) ? 4'b1000 : node1731;
																assign node1731 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node1735 = (inp[2]) ? 4'b1000 : node1736;
															assign node1736 = (inp[3]) ? 4'b1100 : node1737;
																assign node1737 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node1742 = (inp[3]) ? node1760 : node1743;
													assign node1743 = (inp[2]) ? node1751 : node1744;
														assign node1744 = (inp[4]) ? node1748 : node1745;
															assign node1745 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node1748 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node1751 = (inp[15]) ? node1757 : node1752;
															assign node1752 = (inp[7]) ? 4'b1101 : node1753;
																assign node1753 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node1757 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node1760 = (inp[2]) ? node1768 : node1761;
														assign node1761 = (inp[15]) ? node1765 : node1762;
															assign node1762 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node1765 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1768 = (inp[15]) ? node1772 : node1769;
															assign node1769 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node1772 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node1775 = (inp[2]) ? node1809 : node1776;
												assign node1776 = (inp[3]) ? node1794 : node1777;
													assign node1777 = (inp[7]) ? node1785 : node1778;
														assign node1778 = (inp[15]) ? node1782 : node1779;
															assign node1779 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node1782 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node1785 = (inp[4]) ? node1791 : node1786;
															assign node1786 = (inp[14]) ? 4'b1100 : node1787;
																assign node1787 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node1791 = (inp[15]) ? 4'b1001 : 4'b0000;
													assign node1794 = (inp[4]) ? node1802 : node1795;
														assign node1795 = (inp[7]) ? node1799 : node1796;
															assign node1796 = (inp[15]) ? 4'b0100 : 4'b0000;
															assign node1799 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1802 = (inp[15]) ? node1806 : node1803;
															assign node1803 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node1806 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node1809 = (inp[14]) ? node1829 : node1810;
													assign node1810 = (inp[3]) ? node1822 : node1811;
														assign node1811 = (inp[15]) ? node1817 : node1812;
															assign node1812 = (inp[4]) ? node1814 : 4'b1101;
																assign node1814 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node1817 = (inp[4]) ? node1819 : 4'b1001;
																assign node1819 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node1822 = (inp[4]) ? node1824 : 4'b1101;
															assign node1824 = (inp[7]) ? 4'b0000 : node1825;
																assign node1825 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node1829 = (inp[3]) ? node1841 : node1830;
														assign node1830 = (inp[15]) ? node1836 : node1831;
															assign node1831 = (inp[4]) ? node1833 : 4'b1100;
																assign node1833 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node1836 = (inp[7]) ? 4'b1000 : node1837;
																assign node1837 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node1841 = (inp[7]) ? 4'b1100 : node1842;
															assign node1842 = (inp[4]) ? node1846 : node1843;
																assign node1843 = (inp[15]) ? 4'b1100 : 4'b0000;
																assign node1846 = (inp[15]) ? 4'b0000 : 4'b0100;
										assign node1850 = (inp[1]) ? node1946 : node1851;
											assign node1851 = (inp[14]) ? node1899 : node1852;
												assign node1852 = (inp[2]) ? node1876 : node1853;
													assign node1853 = (inp[7]) ? node1869 : node1854;
														assign node1854 = (inp[3]) ? node1862 : node1855;
															assign node1855 = (inp[15]) ? node1859 : node1856;
																assign node1856 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node1859 = (inp[4]) ? 4'b1000 : 4'b0100;
															assign node1862 = (inp[4]) ? node1866 : node1863;
																assign node1863 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node1866 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node1869 = (inp[3]) ? 4'b1100 : node1870;
															assign node1870 = (inp[15]) ? 4'b0100 : node1871;
																assign node1871 = (inp[4]) ? 4'b1000 : 4'b0100;
													assign node1876 = (inp[3]) ? node1886 : node1877;
														assign node1877 = (inp[15]) ? node1883 : node1878;
															assign node1878 = (inp[7]) ? node1880 : 4'b0000;
																assign node1880 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node1883 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node1886 = (inp[15]) ? node1892 : node1887;
															assign node1887 = (inp[4]) ? node1889 : 4'b1000;
																assign node1889 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node1892 = (inp[4]) ? node1896 : node1893;
																assign node1893 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node1896 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node1899 = (inp[2]) ? node1925 : node1900;
													assign node1900 = (inp[3]) ? node1914 : node1901;
														assign node1901 = (inp[15]) ? node1907 : node1902;
															assign node1902 = (inp[4]) ? node1904 : 4'b1000;
																assign node1904 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node1907 = (inp[4]) ? node1911 : node1908;
																assign node1908 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node1911 = (inp[7]) ? 4'b0101 : 4'b1000;
														assign node1914 = (inp[15]) ? node1918 : node1915;
															assign node1915 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node1918 = (inp[4]) ? node1922 : node1919;
																assign node1919 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node1922 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node1925 = (inp[3]) ? node1933 : node1926;
														assign node1926 = (inp[15]) ? 4'b0101 : node1927;
															assign node1927 = (inp[7]) ? node1929 : 4'b0001;
																assign node1929 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1933 = (inp[15]) ? node1941 : node1934;
															assign node1934 = (inp[7]) ? node1938 : node1935;
																assign node1935 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node1938 = (inp[4]) ? 4'b1000 : 4'b0001;
															assign node1941 = (inp[4]) ? 4'b0001 : node1942;
																assign node1942 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node1946 = (inp[14]) ? node1988 : node1947;
												assign node1947 = (inp[3]) ? node1969 : node1948;
													assign node1948 = (inp[2]) ? node1960 : node1949;
														assign node1949 = (inp[7]) ? node1953 : node1950;
															assign node1950 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node1953 = (inp[4]) ? node1957 : node1954;
																assign node1954 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node1957 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node1960 = (inp[15]) ? node1966 : node1961;
															assign node1961 = (inp[7]) ? node1963 : 4'b0001;
																assign node1963 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node1966 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node1969 = (inp[2]) ? node1979 : node1970;
														assign node1970 = (inp[15]) ? node1976 : node1971;
															assign node1971 = (inp[4]) ? node1973 : 4'b0000;
																assign node1973 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node1976 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1979 = (inp[4]) ? node1985 : node1980;
															assign node1980 = (inp[15]) ? node1982 : 4'b0000;
																assign node1982 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node1985 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node1988 = (inp[4]) ? node2004 : node1989;
													assign node1989 = (inp[15]) ? node1995 : node1990;
														assign node1990 = (inp[2]) ? node1992 : 4'b0000;
															assign node1992 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node1995 = (inp[3]) ? node1999 : node1996;
															assign node1996 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node1999 = (inp[7]) ? 4'b0100 : node2000;
																assign node2000 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node2004 = (inp[2]) ? node2016 : node2005;
														assign node2005 = (inp[3]) ? node2009 : node2006;
															assign node2006 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node2009 = (inp[15]) ? node2013 : node2010;
																assign node2010 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node2013 = (inp[7]) ? 4'b0000 : 4'b1001;
														assign node2016 = (inp[7]) ? node2022 : node2017;
															assign node2017 = (inp[3]) ? node2019 : 4'b0000;
																assign node2019 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node2022 = (inp[3]) ? 4'b0100 : node2023;
																assign node2023 = (inp[15]) ? 4'b0100 : 4'b0000;
								assign node2027 = (inp[13]) ? node2305 : node2028;
									assign node2028 = (inp[3]) ? node2172 : node2029;
										assign node2029 = (inp[2]) ? node2101 : node2030;
											assign node2030 = (inp[15]) ? node2062 : node2031;
												assign node2031 = (inp[7]) ? node2045 : node2032;
													assign node2032 = (inp[4]) ? node2038 : node2033;
														assign node2033 = (inp[12]) ? node2035 : 4'b1000;
															assign node2035 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node2038 = (inp[14]) ? 4'b1100 : node2039;
															assign node2039 = (inp[1]) ? 4'b1100 : node2040;
																assign node2040 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2045 = (inp[4]) ? node2057 : node2046;
														assign node2046 = (inp[12]) ? node2052 : node2047;
															assign node2047 = (inp[1]) ? node2049 : 4'b0101;
																assign node2049 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node2052 = (inp[1]) ? 4'b0100 : node2053;
																assign node2053 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node2057 = (inp[1]) ? 4'b1000 : node2058;
															assign node2058 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2062 = (inp[4]) ? node2088 : node2063;
													assign node2063 = (inp[7]) ? node2079 : node2064;
														assign node2064 = (inp[12]) ? node2072 : node2065;
															assign node2065 = (inp[1]) ? node2069 : node2066;
																assign node2066 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node2069 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node2072 = (inp[14]) ? node2076 : node2073;
																assign node2073 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node2076 = (inp[1]) ? 4'b0100 : 4'b1001;
														assign node2079 = (inp[14]) ? node2083 : node2080;
															assign node2080 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2083 = (inp[1]) ? 4'b0000 : node2084;
																assign node2084 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2088 = (inp[7]) ? node2094 : node2089;
														assign node2089 = (inp[12]) ? node2091 : 4'b1000;
															assign node2091 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node2094 = (inp[14]) ? node2098 : node2095;
															assign node2095 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2098 = (inp[1]) ? 4'b0100 : 4'b1001;
											assign node2101 = (inp[15]) ? node2137 : node2102;
												assign node2102 = (inp[7]) ? node2114 : node2103;
													assign node2103 = (inp[1]) ? node2111 : node2104;
														assign node2104 = (inp[14]) ? node2106 : 4'b0000;
															assign node2106 = (inp[12]) ? node2108 : 4'b0001;
																assign node2108 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node2111 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node2114 = (inp[4]) ? node2128 : node2115;
														assign node2115 = (inp[12]) ? node2123 : node2116;
															assign node2116 = (inp[1]) ? node2120 : node2117;
																assign node2117 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node2120 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node2123 = (inp[1]) ? node2125 : 4'b1101;
																assign node2125 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node2128 = (inp[14]) ? node2132 : node2129;
															assign node2129 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2132 = (inp[1]) ? 4'b0000 : node2133;
																assign node2133 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node2137 = (inp[4]) ? node2161 : node2138;
													assign node2138 = (inp[7]) ? node2152 : node2139;
														assign node2139 = (inp[12]) ? node2147 : node2140;
															assign node2140 = (inp[1]) ? node2144 : node2141;
																assign node2141 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node2144 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node2147 = (inp[1]) ? 4'b0100 : node2148;
																assign node2148 = (inp[14]) ? 4'b1001 : 4'b0100;
														assign node2152 = (inp[14]) ? node2156 : node2153;
															assign node2153 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2156 = (inp[1]) ? 4'b0000 : node2157;
																assign node2157 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node2161 = (inp[14]) ? node2165 : node2162;
														assign node2162 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node2165 = (inp[12]) ? node2169 : node2166;
															assign node2166 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node2169 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node2172 = (inp[2]) ? node2240 : node2173;
											assign node2173 = (inp[4]) ? node2211 : node2174;
												assign node2174 = (inp[1]) ? node2190 : node2175;
													assign node2175 = (inp[12]) ? node2183 : node2176;
														assign node2176 = (inp[7]) ? node2180 : node2177;
															assign node2177 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node2180 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node2183 = (inp[15]) ? node2187 : node2184;
															assign node2184 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node2187 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node2190 = (inp[12]) ? node2204 : node2191;
														assign node2191 = (inp[14]) ? node2199 : node2192;
															assign node2192 = (inp[15]) ? node2196 : node2193;
																assign node2193 = (inp[7]) ? 4'b1100 : 4'b1000;
																assign node2196 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node2199 = (inp[15]) ? 4'b1000 : node2200;
																assign node2200 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node2204 = (inp[7]) ? node2208 : node2205;
															assign node2205 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node2208 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node2211 = (inp[15]) ? node2225 : node2212;
													assign node2212 = (inp[1]) ? node2216 : node2213;
														assign node2213 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node2216 = (inp[14]) ? node2220 : node2217;
															assign node2217 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node2220 = (inp[12]) ? 4'b1001 : node2221;
																assign node2221 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2225 = (inp[7]) ? node2235 : node2226;
														assign node2226 = (inp[12]) ? node2230 : node2227;
															assign node2227 = (inp[1]) ? 4'b0001 : 4'b1000;
															assign node2230 = (inp[14]) ? node2232 : 4'b0000;
																assign node2232 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node2235 = (inp[1]) ? 4'b1100 : node2236;
															assign node2236 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node2240 = (inp[15]) ? node2268 : node2241;
												assign node2241 = (inp[7]) ? node2253 : node2242;
													assign node2242 = (inp[4]) ? node2248 : node2243;
														assign node2243 = (inp[1]) ? 4'b1000 : node2244;
															assign node2244 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2248 = (inp[1]) ? 4'b1100 : node2249;
															assign node2249 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2253 = (inp[4]) ? node2263 : node2254;
														assign node2254 = (inp[14]) ? node2258 : node2255;
															assign node2255 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2258 = (inp[1]) ? 4'b0000 : node2259;
																assign node2259 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node2263 = (inp[1]) ? 4'b1000 : node2264;
															assign node2264 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node2268 = (inp[7]) ? node2284 : node2269;
													assign node2269 = (inp[4]) ? node2279 : node2270;
														assign node2270 = (inp[14]) ? node2274 : node2271;
															assign node2271 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2274 = (inp[12]) ? 4'b1101 : node2275;
																assign node2275 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node2279 = (inp[12]) ? node2281 : 4'b1000;
															assign node2281 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node2284 = (inp[4]) ? node2296 : node2285;
														assign node2285 = (inp[12]) ? node2291 : node2286;
															assign node2286 = (inp[1]) ? node2288 : 4'b0100;
																assign node2288 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node2291 = (inp[14]) ? 4'b1101 : node2292;
																assign node2292 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node2296 = (inp[14]) ? node2300 : node2297;
															assign node2297 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node2300 = (inp[12]) ? 4'b1101 : node2301;
																assign node2301 = (inp[1]) ? 4'b0000 : 4'b0001;
									assign node2305 = (inp[1]) ? node2443 : node2306;
										assign node2306 = (inp[12]) ? node2376 : node2307;
											assign node2307 = (inp[2]) ? node2337 : node2308;
												assign node2308 = (inp[3]) ? node2320 : node2309;
													assign node2309 = (inp[15]) ? node2313 : node2310;
														assign node2310 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2313 = (inp[4]) ? 4'b1000 : node2314;
															assign node2314 = (inp[7]) ? node2316 : 4'b1100;
																assign node2316 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node2320 = (inp[14]) ? node2328 : node2321;
														assign node2321 = (inp[4]) ? node2325 : node2322;
															assign node2322 = (inp[15]) ? 4'b1100 : 4'b0001;
															assign node2325 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node2328 = (inp[4]) ? node2334 : node2329;
															assign node2329 = (inp[15]) ? 4'b1100 : node2330;
																assign node2330 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node2334 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node2337 = (inp[14]) ? node2363 : node2338;
													assign node2338 = (inp[4]) ? node2348 : node2339;
														assign node2339 = (inp[15]) ? node2341 : 4'b1000;
															assign node2341 = (inp[3]) ? node2345 : node2342;
																assign node2342 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node2345 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node2348 = (inp[7]) ? node2356 : node2349;
															assign node2349 = (inp[3]) ? node2353 : node2350;
																assign node2350 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node2353 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node2356 = (inp[15]) ? node2360 : node2357;
																assign node2357 = (inp[3]) ? 4'b1100 : 4'b1000;
																assign node2360 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node2363 = (inp[3]) ? node2369 : node2364;
														assign node2364 = (inp[15]) ? node2366 : 4'b1001;
															assign node2366 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node2369 = (inp[4]) ? node2373 : node2370;
															assign node2370 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node2373 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node2376 = (inp[14]) ? node2414 : node2377;
												assign node2377 = (inp[2]) ? node2395 : node2378;
													assign node2378 = (inp[3]) ? node2388 : node2379;
														assign node2379 = (inp[4]) ? node2385 : node2380;
															assign node2380 = (inp[15]) ? node2382 : 4'b0000;
																assign node2382 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node2385 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node2388 = (inp[4]) ? node2392 : node2389;
															assign node2389 = (inp[15]) ? 4'b0100 : 4'b0001;
															assign node2392 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node2395 = (inp[3]) ? node2405 : node2396;
														assign node2396 = (inp[7]) ? node2398 : 4'b1000;
															assign node2398 = (inp[15]) ? node2402 : node2399;
																assign node2399 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node2402 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node2405 = (inp[15]) ? node2409 : node2406;
															assign node2406 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node2409 = (inp[4]) ? 4'b0000 : node2410;
																assign node2410 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node2414 = (inp[3]) ? node2432 : node2415;
													assign node2415 = (inp[2]) ? node2425 : node2416;
														assign node2416 = (inp[4]) ? node2422 : node2417;
															assign node2417 = (inp[15]) ? node2419 : 4'b0000;
																assign node2419 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node2422 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node2425 = (inp[15]) ? node2427 : 4'b0001;
															assign node2427 = (inp[4]) ? 4'b0101 : node2428;
																assign node2428 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node2432 = (inp[4]) ? node2440 : node2433;
														assign node2433 = (inp[15]) ? node2435 : 4'b0000;
															assign node2435 = (inp[2]) ? node2437 : 4'b0100;
																assign node2437 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node2440 = (inp[15]) ? 4'b0000 : 4'b0100;
										assign node2443 = (inp[14]) ? node2477 : node2444;
											assign node2444 = (inp[2]) ? node2456 : node2445;
												assign node2445 = (inp[15]) ? node2449 : node2446;
													assign node2446 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2449 = (inp[4]) ? 4'b1000 : node2450;
														assign node2450 = (inp[3]) ? 4'b1100 : node2451;
															assign node2451 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2456 = (inp[3]) ? node2468 : node2457;
													assign node2457 = (inp[15]) ? node2463 : node2458;
														assign node2458 = (inp[4]) ? 4'b1001 : node2459;
															assign node2459 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node2463 = (inp[7]) ? node2465 : 4'b1101;
															assign node2465 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node2468 = (inp[4]) ? node2474 : node2469;
														assign node2469 = (inp[15]) ? node2471 : 4'b1000;
															assign node2471 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node2474 = (inp[15]) ? 4'b1000 : 4'b1100;
											assign node2477 = (inp[3]) ? node2509 : node2478;
												assign node2478 = (inp[7]) ? node2490 : node2479;
													assign node2479 = (inp[15]) ? node2485 : node2480;
														assign node2480 = (inp[4]) ? node2482 : 4'b1000;
															assign node2482 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node2485 = (inp[2]) ? 4'b1100 : node2486;
															assign node2486 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node2490 = (inp[2]) ? node2496 : node2491;
														assign node2491 = (inp[4]) ? node2493 : 4'b1000;
															assign node2493 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node2496 = (inp[12]) ? node2504 : node2497;
															assign node2497 = (inp[4]) ? node2501 : node2498;
																assign node2498 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node2501 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node2504 = (inp[15]) ? 4'b1000 : node2505;
																assign node2505 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node2509 = (inp[2]) ? node2523 : node2510;
													assign node2510 = (inp[4]) ? node2518 : node2511;
														assign node2511 = (inp[15]) ? 4'b1100 : node2512;
															assign node2512 = (inp[7]) ? 4'b1000 : node2513;
																assign node2513 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2518 = (inp[15]) ? node2520 : 4'b1101;
															assign node2520 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2523 = (inp[4]) ? node2529 : node2524;
														assign node2524 = (inp[15]) ? node2526 : 4'b1000;
															assign node2526 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node2529 = (inp[15]) ? 4'b1000 : 4'b1100;
							assign node2532 = (inp[1]) ? node2902 : node2533;
								assign node2533 = (inp[3]) ? node2703 : node2534;
									assign node2534 = (inp[2]) ? node2632 : node2535;
										assign node2535 = (inp[15]) ? node2585 : node2536;
											assign node2536 = (inp[4]) ? node2560 : node2537;
												assign node2537 = (inp[13]) ? node2551 : node2538;
													assign node2538 = (inp[7]) ? node2546 : node2539;
														assign node2539 = (inp[12]) ? node2543 : node2540;
															assign node2540 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2543 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node2546 = (inp[10]) ? 4'b0100 : node2547;
															assign node2547 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node2551 = (inp[10]) ? node2557 : node2552;
														assign node2552 = (inp[12]) ? node2554 : 4'b0001;
															assign node2554 = (inp[7]) ? 4'b0100 : 4'b1001;
														assign node2557 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node2560 = (inp[13]) ? node2576 : node2561;
													assign node2561 = (inp[7]) ? node2569 : node2562;
														assign node2562 = (inp[12]) ? node2566 : node2563;
															assign node2563 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node2566 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node2569 = (inp[12]) ? node2573 : node2570;
															assign node2570 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2573 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node2576 = (inp[12]) ? node2580 : node2577;
														assign node2577 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node2580 = (inp[10]) ? 4'b0101 : node2581;
															assign node2581 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node2585 = (inp[4]) ? node2609 : node2586;
												assign node2586 = (inp[7]) ? node2598 : node2587;
													assign node2587 = (inp[13]) ? node2593 : node2588;
														assign node2588 = (inp[12]) ? node2590 : 4'b0100;
															assign node2590 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node2593 = (inp[10]) ? 4'b1100 : node2594;
															assign node2594 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2598 = (inp[13]) ? node2604 : node2599;
														assign node2599 = (inp[12]) ? node2601 : 4'b0000;
															assign node2601 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node2604 = (inp[12]) ? node2606 : 4'b1000;
															assign node2606 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node2609 = (inp[13]) ? node2623 : node2610;
													assign node2610 = (inp[7]) ? node2618 : node2611;
														assign node2611 = (inp[10]) ? node2615 : node2612;
															assign node2612 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node2615 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2618 = (inp[12]) ? node2620 : 4'b0100;
															assign node2620 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node2623 = (inp[12]) ? node2627 : node2624;
														assign node2624 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node2627 = (inp[10]) ? 4'b0001 : node2628;
															assign node2628 = (inp[7]) ? 4'b0100 : 4'b1001;
										assign node2632 = (inp[13]) ? node2668 : node2633;
											assign node2633 = (inp[12]) ? node2645 : node2634;
												assign node2634 = (inp[15]) ? node2640 : node2635;
													assign node2635 = (inp[4]) ? 4'b0000 : node2636;
														assign node2636 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2640 = (inp[7]) ? node2642 : 4'b0100;
														assign node2642 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node2645 = (inp[10]) ? node2657 : node2646;
													assign node2646 = (inp[15]) ? node2652 : node2647;
														assign node2647 = (inp[7]) ? 4'b1100 : node2648;
															assign node2648 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node2652 = (inp[4]) ? node2654 : 4'b1000;
															assign node2654 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node2657 = (inp[15]) ? node2663 : node2658;
														assign node2658 = (inp[4]) ? 4'b0000 : node2659;
															assign node2659 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node2663 = (inp[4]) ? 4'b0100 : node2664;
															assign node2664 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node2668 = (inp[15]) ? node2686 : node2669;
												assign node2669 = (inp[10]) ? node2681 : node2670;
													assign node2670 = (inp[12]) ? node2676 : node2671;
														assign node2671 = (inp[7]) ? node2673 : 4'b1000;
															assign node2673 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node2676 = (inp[4]) ? 4'b0000 : node2677;
															assign node2677 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node2681 = (inp[4]) ? 4'b1000 : node2682;
														assign node2682 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node2686 = (inp[12]) ? node2692 : node2687;
													assign node2687 = (inp[7]) ? node2689 : 4'b1100;
														assign node2689 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node2692 = (inp[10]) ? node2698 : node2693;
														assign node2693 = (inp[7]) ? node2695 : 4'b0100;
															assign node2695 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node2698 = (inp[7]) ? node2700 : 4'b1100;
															assign node2700 = (inp[4]) ? 4'b1100 : 4'b1000;
									assign node2703 = (inp[13]) ? node2811 : node2704;
										assign node2704 = (inp[2]) ? node2756 : node2705;
											assign node2705 = (inp[4]) ? node2731 : node2706;
												assign node2706 = (inp[12]) ? node2720 : node2707;
													assign node2707 = (inp[10]) ? node2713 : node2708;
														assign node2708 = (inp[15]) ? node2710 : 4'b0001;
															assign node2710 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node2713 = (inp[7]) ? node2717 : node2714;
															assign node2714 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node2717 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node2720 = (inp[10]) ? node2724 : node2721;
														assign node2721 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node2724 = (inp[7]) ? node2728 : node2725;
															assign node2725 = (inp[15]) ? 4'b0101 : 4'b0001;
															assign node2728 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node2731 = (inp[15]) ? node2741 : node2732;
													assign node2732 = (inp[12]) ? node2738 : node2733;
														assign node2733 = (inp[10]) ? node2735 : 4'b0000;
															assign node2735 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node2738 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node2741 = (inp[7]) ? node2749 : node2742;
														assign node2742 = (inp[10]) ? node2746 : node2743;
															assign node2743 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node2746 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node2749 = (inp[10]) ? node2753 : node2750;
															assign node2750 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node2753 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node2756 = (inp[15]) ? node2786 : node2757;
												assign node2757 = (inp[4]) ? node2771 : node2758;
													assign node2758 = (inp[7]) ? node2766 : node2759;
														assign node2759 = (inp[12]) ? node2763 : node2760;
															assign node2760 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2763 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node2766 = (inp[12]) ? node2768 : 4'b0000;
															assign node2768 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node2771 = (inp[7]) ? node2779 : node2772;
														assign node2772 = (inp[12]) ? node2776 : node2773;
															assign node2773 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node2776 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node2779 = (inp[10]) ? node2783 : node2780;
															assign node2780 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node2783 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node2786 = (inp[7]) ? node2800 : node2787;
													assign node2787 = (inp[4]) ? node2793 : node2788;
														assign node2788 = (inp[10]) ? 4'b0000 : node2789;
															assign node2789 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node2793 = (inp[10]) ? node2797 : node2794;
															assign node2794 = (inp[12]) ? 4'b1000 : 4'b0001;
															assign node2797 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2800 = (inp[4]) ? node2806 : node2801;
														assign node2801 = (inp[12]) ? node2803 : 4'b0100;
															assign node2803 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node2806 = (inp[10]) ? 4'b0000 : node2807;
															assign node2807 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node2811 = (inp[2]) ? node2855 : node2812;
											assign node2812 = (inp[4]) ? node2838 : node2813;
												assign node2813 = (inp[15]) ? node2829 : node2814;
													assign node2814 = (inp[7]) ? node2822 : node2815;
														assign node2815 = (inp[10]) ? node2819 : node2816;
															assign node2816 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node2819 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2822 = (inp[12]) ? node2826 : node2823;
															assign node2823 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node2826 = (inp[10]) ? 4'b0001 : 4'b1101;
													assign node2829 = (inp[12]) ? node2833 : node2830;
														assign node2830 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node2833 = (inp[10]) ? 4'b0101 : node2834;
															assign node2834 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2838 = (inp[15]) ? node2846 : node2839;
													assign node2839 = (inp[10]) ? node2843 : node2840;
														assign node2840 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node2843 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node2846 = (inp[10]) ? node2852 : node2847;
														assign node2847 = (inp[7]) ? node2849 : 4'b1000;
															assign node2849 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node2852 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node2855 = (inp[15]) ? node2881 : node2856;
												assign node2856 = (inp[4]) ? node2872 : node2857;
													assign node2857 = (inp[7]) ? node2865 : node2858;
														assign node2858 = (inp[10]) ? node2862 : node2859;
															assign node2859 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node2862 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node2865 = (inp[10]) ? node2869 : node2866;
															assign node2866 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node2869 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2872 = (inp[12]) ? node2876 : node2873;
														assign node2873 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node2876 = (inp[10]) ? 4'b0101 : node2877;
															assign node2877 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node2881 = (inp[4]) ? node2893 : node2882;
													assign node2882 = (inp[7]) ? node2888 : node2883;
														assign node2883 = (inp[10]) ? 4'b1000 : node2884;
															assign node2884 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node2888 = (inp[12]) ? node2890 : 4'b1100;
															assign node2890 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node2893 = (inp[12]) ? node2897 : node2894;
														assign node2894 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node2897 = (inp[10]) ? 4'b0001 : node2898;
															assign node2898 = (inp[7]) ? 4'b0000 : 4'b1001;
								assign node2902 = (inp[10]) ? node3054 : node2903;
									assign node2903 = (inp[3]) ? node2993 : node2904;
										assign node2904 = (inp[2]) ? node2944 : node2905;
											assign node2905 = (inp[15]) ? node2919 : node2906;
												assign node2906 = (inp[4]) ? node2914 : node2907;
													assign node2907 = (inp[13]) ? 4'b0001 : node2908;
														assign node2908 = (inp[7]) ? node2910 : 4'b0001;
															assign node2910 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node2914 = (inp[13]) ? 4'b0101 : node2915;
														assign node2915 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node2919 = (inp[4]) ? node2933 : node2920;
													assign node2920 = (inp[7]) ? node2926 : node2921;
														assign node2921 = (inp[13]) ? node2923 : 4'b1001;
															assign node2923 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node2926 = (inp[12]) ? node2930 : node2927;
															assign node2927 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node2930 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node2933 = (inp[12]) ? node2939 : node2934;
														assign node2934 = (inp[7]) ? node2936 : 4'b0001;
															assign node2936 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node2939 = (inp[13]) ? 4'b0001 : node2940;
															assign node2940 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node2944 = (inp[15]) ? node2968 : node2945;
												assign node2945 = (inp[7]) ? node2955 : node2946;
													assign node2946 = (inp[12]) ? node2950 : node2947;
														assign node2947 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node2950 = (inp[13]) ? 4'b0001 : node2951;
															assign node2951 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node2955 = (inp[4]) ? node2963 : node2956;
														assign node2956 = (inp[12]) ? node2960 : node2957;
															assign node2957 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node2960 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node2963 = (inp[12]) ? 4'b1101 : node2964;
															assign node2964 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node2968 = (inp[4]) ? node2984 : node2969;
													assign node2969 = (inp[7]) ? node2977 : node2970;
														assign node2970 = (inp[12]) ? node2974 : node2971;
															assign node2971 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node2974 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node2977 = (inp[13]) ? node2981 : node2978;
															assign node2978 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node2981 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node2984 = (inp[12]) ? node2988 : node2985;
														assign node2985 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node2988 = (inp[13]) ? 4'b0101 : node2989;
															assign node2989 = (inp[7]) ? 4'b1001 : 4'b1101;
										assign node2993 = (inp[15]) ? node3017 : node2994;
											assign node2994 = (inp[4]) ? node3002 : node2995;
												assign node2995 = (inp[7]) ? node2997 : 4'b0001;
													assign node2997 = (inp[13]) ? 4'b0001 : node2998;
														assign node2998 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node3002 = (inp[13]) ? node3010 : node3003;
													assign node3003 = (inp[2]) ? node3007 : node3004;
														assign node3004 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3007 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3010 = (inp[12]) ? node3012 : 4'b0101;
														assign node3012 = (inp[2]) ? 4'b0101 : node3013;
															assign node3013 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node3017 = (inp[4]) ? node3039 : node3018;
												assign node3018 = (inp[2]) ? node3024 : node3019;
													assign node3019 = (inp[7]) ? node3021 : 4'b0101;
														assign node3021 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node3024 = (inp[7]) ? node3032 : node3025;
														assign node3025 = (inp[12]) ? node3029 : node3026;
															assign node3026 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node3029 = (inp[13]) ? 4'b0001 : 4'b1101;
														assign node3032 = (inp[13]) ? node3036 : node3033;
															assign node3033 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node3036 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node3039 = (inp[13]) ? node3047 : node3040;
													assign node3040 = (inp[7]) ? node3042 : 4'b0001;
														assign node3042 = (inp[2]) ? node3044 : 4'b0101;
															assign node3044 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node3047 = (inp[2]) ? 4'b0001 : node3048;
														assign node3048 = (inp[12]) ? node3050 : 4'b0001;
															assign node3050 = (inp[7]) ? 4'b0001 : 4'b1001;
									assign node3054 = (inp[13]) ? node3112 : node3055;
										assign node3055 = (inp[2]) ? node3085 : node3056;
											assign node3056 = (inp[7]) ? node3070 : node3057;
												assign node3057 = (inp[4]) ? node3063 : node3058;
													assign node3058 = (inp[15]) ? node3060 : 4'b1001;
														assign node3060 = (inp[3]) ? 4'b1101 : 4'b0101;
													assign node3063 = (inp[15]) ? node3067 : node3064;
														assign node3064 = (inp[3]) ? 4'b0101 : 4'b1101;
														assign node3067 = (inp[3]) ? 4'b0001 : 4'b1001;
												assign node3070 = (inp[3]) ? node3078 : node3071;
													assign node3071 = (inp[4]) ? node3075 : node3072;
														assign node3072 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node3075 = (inp[15]) ? 4'b0101 : 4'b1001;
													assign node3078 = (inp[15]) ? node3082 : node3079;
														assign node3079 = (inp[4]) ? 4'b0001 : 4'b1101;
														assign node3082 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node3085 = (inp[3]) ? node3097 : node3086;
												assign node3086 = (inp[15]) ? node3092 : node3087;
													assign node3087 = (inp[7]) ? node3089 : 4'b0001;
														assign node3089 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node3092 = (inp[4]) ? 4'b0101 : node3093;
														assign node3093 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node3097 = (inp[7]) ? node3105 : node3098;
													assign node3098 = (inp[4]) ? node3102 : node3099;
														assign node3099 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node3102 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node3105 = (inp[15]) ? node3109 : node3106;
														assign node3106 = (inp[4]) ? 4'b1001 : 4'b0001;
														assign node3109 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node3112 = (inp[4]) ? node3150 : node3113;
											assign node3113 = (inp[15]) ? node3121 : node3114;
												assign node3114 = (inp[2]) ? node3116 : 4'b1001;
													assign node3116 = (inp[7]) ? node3118 : 4'b1001;
														assign node3118 = (inp[3]) ? 4'b1001 : 4'b1101;
												assign node3121 = (inp[2]) ? node3127 : node3122;
													assign node3122 = (inp[3]) ? 4'b1101 : node3123;
														assign node3123 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node3127 = (inp[14]) ? node3143 : node3128;
														assign node3128 = (inp[12]) ? node3136 : node3129;
															assign node3129 = (inp[3]) ? node3133 : node3130;
																assign node3130 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node3133 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node3136 = (inp[3]) ? node3140 : node3137;
																assign node3137 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node3140 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node3143 = (inp[3]) ? node3147 : node3144;
															assign node3144 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node3147 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node3150 = (inp[15]) ? node3156 : node3151;
												assign node3151 = (inp[3]) ? 4'b1101 : node3152;
													assign node3152 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node3156 = (inp[2]) ? node3158 : 4'b1001;
													assign node3158 = (inp[3]) ? 4'b1001 : 4'b1101;
						assign node3161 = (inp[15]) ? node3499 : node3162;
							assign node3162 = (inp[2]) ? 4'b1101 : node3163;
								assign node3163 = (inp[1]) ? node3333 : node3164;
									assign node3164 = (inp[3]) ? node3240 : node3165;
										assign node3165 = (inp[7]) ? node3207 : node3166;
											assign node3166 = (inp[14]) ? node3180 : node3167;
												assign node3167 = (inp[13]) ? node3175 : node3168;
													assign node3168 = (inp[12]) ? node3170 : 4'b0000;
														assign node3170 = (inp[10]) ? 4'b0000 : node3171;
															assign node3171 = (inp[4]) ? 4'b1000 : 4'b1101;
													assign node3175 = (inp[10]) ? 4'b1000 : node3176;
														assign node3176 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3180 = (inp[11]) ? node3194 : node3181;
													assign node3181 = (inp[13]) ? node3189 : node3182;
														assign node3182 = (inp[10]) ? node3186 : node3183;
															assign node3183 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node3186 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3189 = (inp[12]) ? 4'b0001 : node3190;
															assign node3190 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3194 = (inp[13]) ? node3202 : node3195;
														assign node3195 = (inp[12]) ? node3197 : 4'b0000;
															assign node3197 = (inp[10]) ? 4'b0000 : node3198;
																assign node3198 = (inp[4]) ? 4'b1000 : 4'b1101;
														assign node3202 = (inp[12]) ? node3204 : 4'b1000;
															assign node3204 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node3207 = (inp[4]) ? node3209 : 4'b1101;
												assign node3209 = (inp[11]) ? node3229 : node3210;
													assign node3210 = (inp[14]) ? node3218 : node3211;
														assign node3211 = (inp[13]) ? 4'b1000 : node3212;
															assign node3212 = (inp[12]) ? node3214 : 4'b0000;
																assign node3214 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node3218 = (inp[13]) ? node3224 : node3219;
															assign node3219 = (inp[10]) ? node3221 : 4'b1101;
																assign node3221 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node3224 = (inp[10]) ? node3226 : 4'b0001;
																assign node3226 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3229 = (inp[13]) ? node3235 : node3230;
														assign node3230 = (inp[10]) ? 4'b0000 : node3231;
															assign node3231 = (inp[12]) ? 4'b1101 : 4'b0000;
														assign node3235 = (inp[10]) ? 4'b1000 : node3236;
															assign node3236 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node3240 = (inp[7]) ? node3280 : node3241;
											assign node3241 = (inp[14]) ? node3255 : node3242;
												assign node3242 = (inp[13]) ? node3250 : node3243;
													assign node3243 = (inp[10]) ? 4'b0100 : node3244;
														assign node3244 = (inp[12]) ? node3246 : 4'b0100;
															assign node3246 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node3250 = (inp[10]) ? 4'b1100 : node3251;
														assign node3251 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node3255 = (inp[11]) ? node3267 : node3256;
													assign node3256 = (inp[13]) ? node3262 : node3257;
														assign node3257 = (inp[4]) ? 4'b1101 : node3258;
															assign node3258 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node3262 = (inp[12]) ? 4'b0101 : node3263;
															assign node3263 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node3267 = (inp[13]) ? node3275 : node3268;
														assign node3268 = (inp[12]) ? node3270 : 4'b0100;
															assign node3270 = (inp[4]) ? node3272 : 4'b1000;
																assign node3272 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node3275 = (inp[10]) ? 4'b1100 : node3276;
															assign node3276 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node3280 = (inp[4]) ? node3312 : node3281;
												assign node3281 = (inp[11]) ? node3301 : node3282;
													assign node3282 = (inp[14]) ? node3294 : node3283;
														assign node3283 = (inp[13]) ? node3289 : node3284;
															assign node3284 = (inp[12]) ? node3286 : 4'b0000;
																assign node3286 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node3289 = (inp[12]) ? node3291 : 4'b1000;
																assign node3291 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3294 = (inp[13]) ? node3296 : 4'b1001;
															assign node3296 = (inp[10]) ? node3298 : 4'b0001;
																assign node3298 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3301 = (inp[13]) ? node3307 : node3302;
														assign node3302 = (inp[12]) ? node3304 : 4'b0000;
															assign node3304 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node3307 = (inp[12]) ? node3309 : 4'b1000;
															assign node3309 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node3312 = (inp[13]) ? node3328 : node3313;
													assign node3313 = (inp[12]) ? node3321 : node3314;
														assign node3314 = (inp[14]) ? node3316 : 4'b0100;
															assign node3316 = (inp[11]) ? 4'b0100 : node3317;
																assign node3317 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node3321 = (inp[14]) ? node3325 : node3322;
															assign node3322 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node3325 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3328 = (inp[12]) ? node3330 : 4'b1100;
														assign node3330 = (inp[10]) ? 4'b1100 : 4'b0100;
									assign node3333 = (inp[13]) ? node3419 : node3334;
										assign node3334 = (inp[12]) ? node3366 : node3335;
											assign node3335 = (inp[3]) ? node3349 : node3336;
												assign node3336 = (inp[7]) ? node3342 : node3337;
													assign node3337 = (inp[14]) ? node3339 : 4'b0001;
														assign node3339 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3342 = (inp[4]) ? node3344 : 4'b1101;
														assign node3344 = (inp[14]) ? node3346 : 4'b0001;
															assign node3346 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node3349 = (inp[7]) ? node3355 : node3350;
													assign node3350 = (inp[14]) ? node3352 : 4'b0101;
														assign node3352 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node3355 = (inp[4]) ? node3361 : node3356;
														assign node3356 = (inp[11]) ? 4'b0001 : node3357;
															assign node3357 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node3361 = (inp[14]) ? node3363 : 4'b0101;
															assign node3363 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node3366 = (inp[10]) ? node3390 : node3367;
												assign node3367 = (inp[3]) ? node3377 : node3368;
													assign node3368 = (inp[4]) ? node3370 : 4'b1101;
														assign node3370 = (inp[7]) ? 4'b1101 : node3371;
															assign node3371 = (inp[14]) ? node3373 : 4'b1001;
																assign node3373 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node3377 = (inp[11]) ? node3385 : node3378;
														assign node3378 = (inp[14]) ? node3380 : 4'b1001;
															assign node3380 = (inp[7]) ? 4'b1000 : node3381;
																assign node3381 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node3385 = (inp[4]) ? node3387 : 4'b1001;
															assign node3387 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node3390 = (inp[3]) ? node3400 : node3391;
													assign node3391 = (inp[4]) ? node3395 : node3392;
														assign node3392 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node3395 = (inp[14]) ? node3397 : 4'b0001;
															assign node3397 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3400 = (inp[7]) ? node3408 : node3401;
														assign node3401 = (inp[4]) ? 4'b0101 : node3402;
															assign node3402 = (inp[14]) ? node3404 : 4'b0101;
																assign node3404 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node3408 = (inp[4]) ? node3414 : node3409;
															assign node3409 = (inp[11]) ? 4'b0001 : node3410;
																assign node3410 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node3414 = (inp[11]) ? 4'b0101 : node3415;
																assign node3415 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node3419 = (inp[3]) ? node3453 : node3420;
											assign node3420 = (inp[7]) ? node3438 : node3421;
												assign node3421 = (inp[14]) ? node3427 : node3422;
													assign node3422 = (inp[12]) ? node3424 : 4'b1001;
														assign node3424 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3427 = (inp[11]) ? node3433 : node3428;
														assign node3428 = (inp[12]) ? node3430 : 4'b1000;
															assign node3430 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3433 = (inp[12]) ? node3435 : 4'b1001;
															assign node3435 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node3438 = (inp[4]) ? node3440 : 4'b1101;
													assign node3440 = (inp[12]) ? node3446 : node3441;
														assign node3441 = (inp[11]) ? 4'b1001 : node3442;
															assign node3442 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3446 = (inp[10]) ? 4'b1001 : node3447;
															assign node3447 = (inp[11]) ? 4'b0001 : node3448;
																assign node3448 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node3453 = (inp[10]) ? node3481 : node3454;
												assign node3454 = (inp[12]) ? node3468 : node3455;
													assign node3455 = (inp[7]) ? node3457 : 4'b1101;
														assign node3457 = (inp[4]) ? node3463 : node3458;
															assign node3458 = (inp[11]) ? 4'b1001 : node3459;
																assign node3459 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node3463 = (inp[14]) ? node3465 : 4'b1101;
																assign node3465 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node3468 = (inp[4]) ? node3476 : node3469;
														assign node3469 = (inp[7]) ? node3471 : 4'b0101;
															assign node3471 = (inp[14]) ? node3473 : 4'b0001;
																assign node3473 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node3476 = (inp[14]) ? node3478 : 4'b0101;
															assign node3478 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node3481 = (inp[11]) ? node3493 : node3482;
													assign node3482 = (inp[14]) ? node3488 : node3483;
														assign node3483 = (inp[4]) ? 4'b1101 : node3484;
															assign node3484 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node3488 = (inp[4]) ? 4'b1100 : node3489;
															assign node3489 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node3493 = (inp[7]) ? node3495 : 4'b1101;
														assign node3495 = (inp[4]) ? 4'b1101 : 4'b1001;
							assign node3499 = (inp[3]) ? node3501 : 4'b1001;
								assign node3501 = (inp[2]) ? 4'b1001 : node3502;
									assign node3502 = (inp[4]) ? node3566 : node3503;
										assign node3503 = (inp[7]) ? 4'b1001 : node3504;
											assign node3504 = (inp[1]) ? node3534 : node3505;
												assign node3505 = (inp[11]) ? node3523 : node3506;
													assign node3506 = (inp[14]) ? node3514 : node3507;
														assign node3507 = (inp[13]) ? 4'b1000 : node3508;
															assign node3508 = (inp[10]) ? 4'b0000 : node3509;
																assign node3509 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node3514 = (inp[13]) ? node3520 : node3515;
															assign node3515 = (inp[10]) ? node3517 : 4'b1001;
																assign node3517 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node3520 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node3523 = (inp[13]) ? node3529 : node3524;
														assign node3524 = (inp[12]) ? node3526 : 4'b0000;
															assign node3526 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node3529 = (inp[10]) ? 4'b1000 : node3530;
															assign node3530 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node3534 = (inp[11]) ? node3554 : node3535;
													assign node3535 = (inp[14]) ? node3543 : node3536;
														assign node3536 = (inp[13]) ? node3540 : node3537;
															assign node3537 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node3540 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3543 = (inp[13]) ? node3549 : node3544;
															assign node3544 = (inp[12]) ? node3546 : 4'b0000;
																assign node3546 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node3549 = (inp[12]) ? node3551 : 4'b1000;
																assign node3551 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node3554 = (inp[13]) ? node3560 : node3555;
														assign node3555 = (inp[10]) ? 4'b0001 : node3556;
															assign node3556 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node3560 = (inp[12]) ? node3562 : 4'b1001;
															assign node3562 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node3566 = (inp[1]) ? node3604 : node3567;
											assign node3567 = (inp[14]) ? node3581 : node3568;
												assign node3568 = (inp[13]) ? node3576 : node3569;
													assign node3569 = (inp[10]) ? 4'b0000 : node3570;
														assign node3570 = (inp[12]) ? node3572 : 4'b0000;
															assign node3572 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3576 = (inp[10]) ? 4'b1000 : node3577;
														assign node3577 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node3581 = (inp[11]) ? node3593 : node3582;
													assign node3582 = (inp[13]) ? node3588 : node3583;
														assign node3583 = (inp[12]) ? 4'b1001 : node3584;
															assign node3584 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node3588 = (inp[10]) ? node3590 : 4'b0001;
															assign node3590 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3593 = (inp[13]) ? node3599 : node3594;
														assign node3594 = (inp[12]) ? node3596 : 4'b0000;
															assign node3596 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node3599 = (inp[12]) ? node3601 : 4'b1000;
															assign node3601 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node3604 = (inp[13]) ? node3620 : node3605;
												assign node3605 = (inp[14]) ? node3611 : node3606;
													assign node3606 = (inp[10]) ? 4'b0001 : node3607;
														assign node3607 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node3611 = (inp[11]) ? 4'b0001 : node3612;
														assign node3612 = (inp[12]) ? node3614 : 4'b0000;
															assign node3614 = (inp[10]) ? 4'b0000 : node3615;
																assign node3615 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node3620 = (inp[10]) ? node3632 : node3621;
													assign node3621 = (inp[12]) ? node3627 : node3622;
														assign node3622 = (inp[11]) ? 4'b1001 : node3623;
															assign node3623 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3627 = (inp[14]) ? node3629 : 4'b0001;
															assign node3629 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node3632 = (inp[11]) ? 4'b1001 : node3633;
														assign node3633 = (inp[14]) ? 4'b1000 : 4'b1001;
					assign node3638 = (inp[3]) ? node5158 : node3639;
						assign node3639 = (inp[2]) ? node4567 : node3640;
							assign node3640 = (inp[11]) ? node4196 : node3641;
								assign node3641 = (inp[0]) ? node3913 : node3642;
									assign node3642 = (inp[4]) ? node3782 : node3643;
										assign node3643 = (inp[15]) ? node3709 : node3644;
											assign node3644 = (inp[10]) ? node3684 : node3645;
												assign node3645 = (inp[13]) ? node3669 : node3646;
													assign node3646 = (inp[7]) ? node3656 : node3647;
														assign node3647 = (inp[1]) ? node3653 : node3648;
															assign node3648 = (inp[12]) ? node3650 : 4'b0001;
																assign node3650 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node3653 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3656 = (inp[1]) ? node3664 : node3657;
															assign node3657 = (inp[12]) ? node3661 : node3658;
																assign node3658 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node3661 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node3664 = (inp[14]) ? 4'b0101 : node3665;
																assign node3665 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node3669 = (inp[7]) ? node3677 : node3670;
														assign node3670 = (inp[12]) ? node3674 : node3671;
															assign node3671 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node3674 = (inp[1]) ? 4'b0101 : 4'b1001;
														assign node3677 = (inp[12]) ? node3681 : node3678;
															assign node3678 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node3681 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node3684 = (inp[13]) ? node3694 : node3685;
													assign node3685 = (inp[12]) ? node3689 : node3686;
														assign node3686 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node3689 = (inp[1]) ? 4'b0001 : node3690;
															assign node3690 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node3694 = (inp[12]) ? node3700 : node3695;
														assign node3695 = (inp[1]) ? node3697 : 4'b0101;
															assign node3697 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node3700 = (inp[1]) ? node3704 : node3701;
															assign node3701 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node3704 = (inp[7]) ? 4'b0101 : node3705;
																assign node3705 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node3709 = (inp[13]) ? node3749 : node3710;
												assign node3710 = (inp[7]) ? node3730 : node3711;
													assign node3711 = (inp[1]) ? node3719 : node3712;
														assign node3712 = (inp[14]) ? node3716 : node3713;
															assign node3713 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node3716 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node3719 = (inp[14]) ? node3725 : node3720;
															assign node3720 = (inp[10]) ? 4'b0100 : node3721;
																assign node3721 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node3725 = (inp[10]) ? node3727 : 4'b0101;
																assign node3727 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node3730 = (inp[1]) ? node3738 : node3731;
														assign node3731 = (inp[14]) ? node3733 : 4'b1001;
															assign node3733 = (inp[12]) ? 4'b1000 : node3734;
																assign node3734 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node3738 = (inp[14]) ? node3744 : node3739;
															assign node3739 = (inp[10]) ? 4'b0100 : node3740;
																assign node3740 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node3744 = (inp[10]) ? node3746 : 4'b0001;
																assign node3746 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node3749 = (inp[7]) ? node3759 : node3750;
													assign node3750 = (inp[12]) ? node3754 : node3751;
														assign node3751 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node3754 = (inp[1]) ? 4'b0001 : node3755;
															assign node3755 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node3759 = (inp[10]) ? node3773 : node3760;
														assign node3760 = (inp[14]) ? node3768 : node3761;
															assign node3761 = (inp[1]) ? node3765 : node3762;
																assign node3762 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node3765 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node3768 = (inp[1]) ? 4'b1101 : node3769;
																assign node3769 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node3773 = (inp[12]) ? node3777 : node3774;
															assign node3774 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node3777 = (inp[1]) ? 4'b0001 : node3778;
																assign node3778 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node3782 = (inp[13]) ? node3858 : node3783;
											assign node3783 = (inp[15]) ? node3819 : node3784;
												assign node3784 = (inp[1]) ? node3802 : node3785;
													assign node3785 = (inp[14]) ? node3793 : node3786;
														assign node3786 = (inp[10]) ? node3788 : 4'b0000;
															assign node3788 = (inp[7]) ? node3790 : 4'b1100;
																assign node3790 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node3793 = (inp[12]) ? node3795 : 4'b0001;
															assign node3795 = (inp[10]) ? node3799 : node3796;
																assign node3796 = (inp[7]) ? 4'b1101 : 4'b1001;
																assign node3799 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node3802 = (inp[14]) ? node3810 : node3803;
														assign node3803 = (inp[10]) ? node3805 : 4'b1001;
															assign node3805 = (inp[7]) ? node3807 : 4'b0000;
																assign node3807 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node3810 = (inp[10]) ? node3812 : 4'b1000;
															assign node3812 = (inp[12]) ? node3816 : node3813;
																assign node3813 = (inp[7]) ? 4'b0100 : 4'b1000;
																assign node3816 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node3819 = (inp[10]) ? node3837 : node3820;
													assign node3820 = (inp[7]) ? node3828 : node3821;
														assign node3821 = (inp[1]) ? node3825 : node3822;
															assign node3822 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node3825 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node3828 = (inp[14]) ? 4'b0001 : node3829;
															assign node3829 = (inp[1]) ? node3833 : node3830;
																assign node3830 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node3833 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node3837 = (inp[7]) ? node3849 : node3838;
														assign node3838 = (inp[1]) ? node3844 : node3839;
															assign node3839 = (inp[14]) ? 4'b0001 : node3840;
																assign node3840 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node3844 = (inp[12]) ? node3846 : 4'b0001;
																assign node3846 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node3849 = (inp[12]) ? node3855 : node3850;
															assign node3850 = (inp[1]) ? node3852 : 4'b0101;
																assign node3852 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node3855 = (inp[1]) ? 4'b0101 : 4'b1001;
											assign node3858 = (inp[10]) ? node3888 : node3859;
												assign node3859 = (inp[15]) ? node3869 : node3860;
													assign node3860 = (inp[12]) ? node3866 : node3861;
														assign node3861 = (inp[7]) ? 4'b0000 : node3862;
															assign node3862 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node3866 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node3869 = (inp[1]) ? node3875 : node3870;
														assign node3870 = (inp[14]) ? node3872 : 4'b1000;
															assign node3872 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3875 = (inp[14]) ? node3883 : node3876;
															assign node3876 = (inp[12]) ? node3880 : node3877;
																assign node3877 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node3880 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node3883 = (inp[7]) ? 4'b0000 : node3884;
																assign node3884 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node3888 = (inp[1]) ? node3902 : node3889;
													assign node3889 = (inp[7]) ? node3897 : node3890;
														assign node3890 = (inp[14]) ? 4'b1000 : node3891;
															assign node3891 = (inp[15]) ? 4'b1000 : node3892;
																assign node3892 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node3897 = (inp[15]) ? node3899 : 4'b1000;
															assign node3899 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node3902 = (inp[12]) ? node3908 : node3903;
														assign node3903 = (inp[14]) ? node3905 : 4'b1000;
															assign node3905 = (inp[15]) ? 4'b1000 : 4'b0001;
														assign node3908 = (inp[15]) ? 4'b0000 : node3909;
															assign node3909 = (inp[14]) ? 4'b0001 : 4'b0000;
									assign node3913 = (inp[13]) ? node4095 : node3914;
										assign node3914 = (inp[12]) ? node4006 : node3915;
											assign node3915 = (inp[10]) ? node3961 : node3916;
												assign node3916 = (inp[4]) ? node3946 : node3917;
													assign node3917 = (inp[1]) ? node3931 : node3918;
														assign node3918 = (inp[14]) ? node3924 : node3919;
															assign node3919 = (inp[15]) ? node3921 : 4'b0000;
																assign node3921 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node3924 = (inp[7]) ? node3928 : node3925;
																assign node3925 = (inp[15]) ? 4'b1001 : 4'b0000;
																assign node3928 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node3931 = (inp[14]) ? node3939 : node3932;
															assign node3932 = (inp[7]) ? node3936 : node3933;
																assign node3933 = (inp[15]) ? 4'b0101 : 4'b0000;
																assign node3936 = (inp[15]) ? 4'b0001 : 4'b0101;
															assign node3939 = (inp[15]) ? node3943 : node3940;
																assign node3940 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node3943 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node3946 = (inp[1]) ? node3954 : node3947;
														assign node3947 = (inp[7]) ? node3951 : node3948;
															assign node3948 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3951 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node3954 = (inp[15]) ? node3958 : node3955;
															assign node3955 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node3958 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node3961 = (inp[7]) ? node3981 : node3962;
													assign node3962 = (inp[1]) ? node3972 : node3963;
														assign node3963 = (inp[15]) ? node3967 : node3964;
															assign node3964 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node3967 = (inp[4]) ? 4'b1000 : node3968;
																assign node3968 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node3972 = (inp[15]) ? node3978 : node3973;
															assign node3973 = (inp[4]) ? node3975 : 4'b1000;
																assign node3975 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node3978 = (inp[4]) ? 4'b1000 : 4'b0100;
													assign node3981 = (inp[15]) ? node3991 : node3982;
														assign node3982 = (inp[4]) ? 4'b1000 : node3983;
															assign node3983 = (inp[1]) ? node3987 : node3984;
																assign node3984 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node3987 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node3991 = (inp[4]) ? node3999 : node3992;
															assign node3992 = (inp[14]) ? node3996 : node3993;
																assign node3993 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node3996 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node3999 = (inp[1]) ? node4003 : node4000;
																assign node4000 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node4003 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node4006 = (inp[10]) ? node4048 : node4007;
												assign node4007 = (inp[1]) ? node4027 : node4008;
													assign node4008 = (inp[14]) ? node4018 : node4009;
														assign node4009 = (inp[15]) ? node4013 : node4010;
															assign node4010 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node4013 = (inp[4]) ? node4015 : 4'b1000;
																assign node4015 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node4018 = (inp[4]) ? node4022 : node4019;
															assign node4019 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node4022 = (inp[15]) ? node4024 : 4'b1000;
																assign node4024 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4027 = (inp[15]) ? node4037 : node4028;
														assign node4028 = (inp[7]) ? node4032 : node4029;
															assign node4029 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node4032 = (inp[4]) ? 4'b0000 : node4033;
																assign node4033 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node4037 = (inp[14]) ? node4043 : node4038;
															assign node4038 = (inp[4]) ? node4040 : 4'b1001;
																assign node4040 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node4043 = (inp[7]) ? 4'b1000 : node4044;
																assign node4044 = (inp[4]) ? 4'b0000 : 4'b1000;
												assign node4048 = (inp[7]) ? node4066 : node4049;
													assign node4049 = (inp[1]) ? node4057 : node4050;
														assign node4050 = (inp[4]) ? node4054 : node4051;
															assign node4051 = (inp[15]) ? 4'b0100 : 4'b0000;
															assign node4054 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node4057 = (inp[15]) ? node4061 : node4058;
															assign node4058 = (inp[4]) ? 4'b0000 : 4'b1000;
															assign node4061 = (inp[4]) ? 4'b1000 : node4062;
																assign node4062 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node4066 = (inp[14]) ? node4082 : node4067;
														assign node4067 = (inp[1]) ? node4075 : node4068;
															assign node4068 = (inp[15]) ? node4072 : node4069;
																assign node4069 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node4072 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node4075 = (inp[15]) ? node4079 : node4076;
																assign node4076 = (inp[4]) ? 4'b1000 : 4'b0101;
																assign node4079 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node4082 = (inp[1]) ? node4088 : node4083;
															assign node4083 = (inp[15]) ? 4'b1001 : node4084;
																assign node4084 = (inp[4]) ? 4'b0000 : 4'b1101;
															assign node4088 = (inp[4]) ? node4092 : node4089;
																assign node4089 = (inp[15]) ? 4'b0000 : 4'b0100;
																assign node4092 = (inp[15]) ? 4'b0100 : 4'b1000;
										assign node4095 = (inp[10]) ? node4159 : node4096;
											assign node4096 = (inp[7]) ? node4132 : node4097;
												assign node4097 = (inp[4]) ? node4117 : node4098;
													assign node4098 = (inp[15]) ? node4104 : node4099;
														assign node4099 = (inp[1]) ? 4'b0000 : node4100;
															assign node4100 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4104 = (inp[12]) ? node4112 : node4105;
															assign node4105 = (inp[14]) ? node4109 : node4106;
																assign node4106 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node4109 = (inp[1]) ? 4'b1100 : 4'b0101;
															assign node4112 = (inp[1]) ? 4'b0101 : node4113;
																assign node4113 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node4117 = (inp[15]) ? node4127 : node4118;
														assign node4118 = (inp[14]) ? node4124 : node4119;
															assign node4119 = (inp[1]) ? 4'b0000 : node4120;
																assign node4120 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node4124 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node4127 = (inp[1]) ? 4'b0000 : node4128;
															assign node4128 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node4132 = (inp[4]) ? node4148 : node4133;
													assign node4133 = (inp[15]) ? node4139 : node4134;
														assign node4134 = (inp[1]) ? 4'b0000 : node4135;
															assign node4135 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node4139 = (inp[1]) ? node4141 : 4'b0001;
															assign node4141 = (inp[12]) ? node4145 : node4142;
																assign node4142 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node4145 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4148 = (inp[1]) ? node4154 : node4149;
														assign node4149 = (inp[12]) ? node4151 : 4'b0100;
															assign node4151 = (inp[15]) ? 4'b0100 : 4'b1000;
														assign node4154 = (inp[15]) ? 4'b0000 : node4155;
															assign node4155 = (inp[14]) ? 4'b0100 : 4'b0000;
											assign node4159 = (inp[1]) ? node4179 : node4160;
												assign node4160 = (inp[4]) ? node4172 : node4161;
													assign node4161 = (inp[15]) ? node4165 : node4162;
														assign node4162 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4165 = (inp[7]) ? node4169 : node4166;
															assign node4166 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node4169 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node4172 = (inp[15]) ? node4176 : node4173;
														assign node4173 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node4176 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4179 = (inp[15]) ? node4187 : node4180;
													assign node4180 = (inp[4]) ? node4182 : 4'b1000;
														assign node4182 = (inp[14]) ? node4184 : 4'b1000;
															assign node4184 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4187 = (inp[4]) ? 4'b1000 : node4188;
														assign node4188 = (inp[14]) ? node4192 : node4189;
															assign node4189 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4192 = (inp[7]) ? 4'b1000 : 4'b1100;
								assign node4196 = (inp[1]) ? node4384 : node4197;
									assign node4197 = (inp[4]) ? node4285 : node4198;
										assign node4198 = (inp[15]) ? node4244 : node4199;
											assign node4199 = (inp[7]) ? node4223 : node4200;
												assign node4200 = (inp[0]) ? node4208 : node4201;
													assign node4201 = (inp[10]) ? node4205 : node4202;
														assign node4202 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node4205 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node4208 = (inp[13]) ? node4216 : node4209;
														assign node4209 = (inp[12]) ? node4213 : node4210;
															assign node4210 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4213 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node4216 = (inp[12]) ? node4220 : node4217;
															assign node4217 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4220 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node4223 = (inp[13]) ? node4233 : node4224;
													assign node4224 = (inp[10]) ? node4230 : node4225;
														assign node4225 = (inp[0]) ? node4227 : 4'b0100;
															assign node4227 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node4230 = (inp[0]) ? 4'b0100 : 4'b0001;
													assign node4233 = (inp[10]) ? node4239 : node4234;
														assign node4234 = (inp[12]) ? node4236 : 4'b0001;
															assign node4236 = (inp[0]) ? 4'b0100 : 4'b0001;
														assign node4239 = (inp[0]) ? node4241 : 4'b0101;
															assign node4241 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node4244 = (inp[7]) ? node4264 : node4245;
												assign node4245 = (inp[0]) ? node4253 : node4246;
													assign node4246 = (inp[13]) ? 4'b0001 : node4247;
														assign node4247 = (inp[12]) ? node4249 : 4'b0100;
															assign node4249 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node4253 = (inp[13]) ? node4259 : node4254;
														assign node4254 = (inp[12]) ? node4256 : 4'b0100;
															assign node4256 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node4259 = (inp[12]) ? node4261 : 4'b1100;
															assign node4261 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node4264 = (inp[0]) ? node4274 : node4265;
													assign node4265 = (inp[10]) ? node4269 : node4266;
														assign node4266 = (inp[13]) ? 4'b1100 : 4'b0000;
														assign node4269 = (inp[13]) ? 4'b0001 : node4270;
															assign node4270 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node4274 = (inp[13]) ? node4280 : node4275;
														assign node4275 = (inp[12]) ? node4277 : 4'b0000;
															assign node4277 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node4280 = (inp[12]) ? node4282 : 4'b1000;
															assign node4282 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node4285 = (inp[15]) ? node4335 : node4286;
											assign node4286 = (inp[10]) ? node4306 : node4287;
												assign node4287 = (inp[13]) ? node4297 : node4288;
													assign node4288 = (inp[0]) ? node4292 : node4289;
														assign node4289 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4292 = (inp[12]) ? 4'b1001 : node4293;
															assign node4293 = (inp[14]) ? 4'b0101 : 4'b0001;
													assign node4297 = (inp[0]) ? node4301 : node4298;
														assign node4298 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4301 = (inp[7]) ? node4303 : 4'b1000;
															assign node4303 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node4306 = (inp[13]) ? node4320 : node4307;
													assign node4307 = (inp[7]) ? node4315 : node4308;
														assign node4308 = (inp[12]) ? node4312 : node4309;
															assign node4309 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4312 = (inp[0]) ? 4'b0101 : 4'b1100;
														assign node4315 = (inp[0]) ? node4317 : 4'b1000;
															assign node4317 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4320 = (inp[7]) ? node4328 : node4321;
														assign node4321 = (inp[0]) ? node4325 : node4322;
															assign node4322 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node4325 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4328 = (inp[12]) ? node4332 : node4329;
															assign node4329 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node4332 = (inp[0]) ? 4'b0000 : 4'b1001;
											assign node4335 = (inp[7]) ? node4359 : node4336;
												assign node4336 = (inp[10]) ? node4350 : node4337;
													assign node4337 = (inp[12]) ? node4343 : node4338;
														assign node4338 = (inp[0]) ? 4'b0001 : node4339;
															assign node4339 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node4343 = (inp[13]) ? node4347 : node4344;
															assign node4344 = (inp[0]) ? 4'b1100 : 4'b0101;
															assign node4347 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node4350 = (inp[0]) ? node4356 : node4351;
														assign node4351 = (inp[13]) ? node4353 : 4'b1000;
															assign node4353 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node4356 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node4359 = (inp[10]) ? node4373 : node4360;
													assign node4360 = (inp[0]) ? node4366 : node4361;
														assign node4361 = (inp[13]) ? node4363 : 4'b0001;
															assign node4363 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4366 = (inp[12]) ? node4370 : node4367;
															assign node4367 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node4370 = (inp[13]) ? 4'b0100 : 4'b1000;
													assign node4373 = (inp[13]) ? node4377 : node4374;
														assign node4374 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node4377 = (inp[0]) ? node4381 : node4378;
															assign node4378 = (inp[12]) ? 4'b0100 : 4'b0001;
															assign node4381 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node4384 = (inp[13]) ? node4498 : node4385;
										assign node4385 = (inp[0]) ? node4423 : node4386;
											assign node4386 = (inp[15]) ? node4406 : node4387;
												assign node4387 = (inp[7]) ? node4395 : node4388;
													assign node4388 = (inp[4]) ? node4390 : 4'b1001;
														assign node4390 = (inp[10]) ? 4'b1001 : node4391;
															assign node4391 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node4395 = (inp[4]) ? node4401 : node4396;
														assign node4396 = (inp[10]) ? 4'b1001 : node4397;
															assign node4397 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node4401 = (inp[10]) ? 4'b0101 : node4402;
															assign node4402 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node4406 = (inp[10]) ? node4420 : node4407;
													assign node4407 = (inp[7]) ? node4415 : node4408;
														assign node4408 = (inp[4]) ? node4412 : node4409;
															assign node4409 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node4412 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node4415 = (inp[4]) ? 4'b1001 : node4416;
															assign node4416 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node4420 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node4423 = (inp[12]) ? node4469 : node4424;
												assign node4424 = (inp[10]) ? node4454 : node4425;
													assign node4425 = (inp[15]) ? node4439 : node4426;
														assign node4426 = (inp[14]) ? node4432 : node4427;
															assign node4427 = (inp[7]) ? 4'b0001 : node4428;
																assign node4428 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node4432 = (inp[4]) ? node4436 : node4433;
																assign node4433 = (inp[7]) ? 4'b0101 : 4'b0001;
																assign node4436 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node4439 = (inp[14]) ? node4447 : node4440;
															assign node4440 = (inp[7]) ? node4444 : node4441;
																assign node4441 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node4444 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node4447 = (inp[7]) ? node4451 : node4448;
																assign node4448 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node4451 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4454 = (inp[15]) ? node4462 : node4455;
														assign node4455 = (inp[7]) ? node4459 : node4456;
															assign node4456 = (inp[4]) ? 4'b0001 : 4'b1001;
															assign node4459 = (inp[4]) ? 4'b1001 : 4'b0101;
														assign node4462 = (inp[4]) ? node4466 : node4463;
															assign node4463 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node4466 = (inp[7]) ? 4'b0101 : 4'b1001;
												assign node4469 = (inp[15]) ? node4485 : node4470;
													assign node4470 = (inp[7]) ? node4478 : node4471;
														assign node4471 = (inp[10]) ? node4475 : node4472;
															assign node4472 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node4475 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node4478 = (inp[4]) ? node4482 : node4479;
															assign node4479 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node4482 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4485 = (inp[10]) ? node4491 : node4486;
														assign node4486 = (inp[7]) ? 4'b1001 : node4487;
															assign node4487 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node4491 = (inp[4]) ? node4495 : node4492;
															assign node4492 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node4495 = (inp[7]) ? 4'b0101 : 4'b1001;
										assign node4498 = (inp[10]) ? node4542 : node4499;
											assign node4499 = (inp[4]) ? node4525 : node4500;
												assign node4500 = (inp[0]) ? node4516 : node4501;
													assign node4501 = (inp[12]) ? node4509 : node4502;
														assign node4502 = (inp[15]) ? node4506 : node4503;
															assign node4503 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4506 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node4509 = (inp[15]) ? node4513 : node4510;
															assign node4510 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4513 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node4516 = (inp[15]) ? node4518 : 4'b0001;
														assign node4518 = (inp[12]) ? node4522 : node4519;
															assign node4519 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node4522 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4525 = (inp[15]) ? node4535 : node4526;
													assign node4526 = (inp[12]) ? node4528 : 4'b0001;
														assign node4528 = (inp[14]) ? 4'b0101 : node4529;
															assign node4529 = (inp[7]) ? 4'b0101 : node4530;
																assign node4530 = (inp[0]) ? 4'b1001 : 4'b0101;
													assign node4535 = (inp[12]) ? 4'b0001 : node4536;
														assign node4536 = (inp[7]) ? node4538 : 4'b0001;
															assign node4538 = (inp[0]) ? 4'b0001 : 4'b1001;
											assign node4542 = (inp[4]) ? 4'b1001 : node4543;
												assign node4543 = (inp[14]) ? node4555 : node4544;
													assign node4544 = (inp[0]) ? node4550 : node4545;
														assign node4545 = (inp[15]) ? 4'b1001 : node4546;
															assign node4546 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node4550 = (inp[15]) ? node4552 : 4'b1001;
															assign node4552 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4555 = (inp[0]) ? node4561 : node4556;
														assign node4556 = (inp[7]) ? node4558 : 4'b1001;
															assign node4558 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node4561 = (inp[7]) ? 4'b1001 : node4562;
															assign node4562 = (inp[15]) ? 4'b1101 : 4'b1001;
							assign node4567 = (inp[0]) ? node5009 : node4568;
								assign node4568 = (inp[4]) ? node4810 : node4569;
									assign node4569 = (inp[11]) ? node4709 : node4570;
										assign node4570 = (inp[15]) ? node4656 : node4571;
											assign node4571 = (inp[13]) ? node4609 : node4572;
												assign node4572 = (inp[7]) ? node4596 : node4573;
													assign node4573 = (inp[1]) ? node4585 : node4574;
														assign node4574 = (inp[14]) ? node4580 : node4575;
															assign node4575 = (inp[10]) ? 4'b1001 : node4576;
																assign node4576 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node4580 = (inp[10]) ? 4'b1000 : node4581;
																assign node4581 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node4585 = (inp[14]) ? node4591 : node4586;
															assign node4586 = (inp[12]) ? 4'b0000 : node4587;
																assign node4587 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node4591 = (inp[12]) ? node4593 : 4'b0001;
																assign node4593 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node4596 = (inp[1]) ? node4604 : node4597;
														assign node4597 = (inp[10]) ? node4601 : node4598;
															assign node4598 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node4601 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node4604 = (inp[10]) ? node4606 : 4'b0100;
															assign node4606 = (inp[14]) ? 4'b1100 : 4'b0000;
												assign node4609 = (inp[7]) ? node4633 : node4610;
													assign node4610 = (inp[10]) ? node4624 : node4611;
														assign node4611 = (inp[14]) ? node4619 : node4612;
															assign node4612 = (inp[1]) ? node4616 : node4613;
																assign node4613 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node4616 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node4619 = (inp[1]) ? 4'b1001 : node4620;
																assign node4620 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4624 = (inp[1]) ? node4628 : node4625;
															assign node4625 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node4628 = (inp[14]) ? node4630 : 4'b1100;
																assign node4630 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node4633 = (inp[1]) ? node4645 : node4634;
														assign node4634 = (inp[14]) ? node4640 : node4635;
															assign node4635 = (inp[12]) ? 4'b0001 : node4636;
																assign node4636 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node4640 = (inp[10]) ? 4'b0000 : node4641;
																assign node4641 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node4645 = (inp[14]) ? node4651 : node4646;
															assign node4646 = (inp[10]) ? 4'b1000 : node4647;
																assign node4647 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node4651 = (inp[10]) ? node4653 : 4'b1001;
																assign node4653 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node4656 = (inp[10]) ? node4678 : node4657;
												assign node4657 = (inp[1]) ? node4669 : node4658;
													assign node4658 = (inp[12]) ? node4664 : node4659;
														assign node4659 = (inp[13]) ? 4'b0100 : node4660;
															assign node4660 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4664 = (inp[7]) ? 4'b1000 : node4665;
															assign node4665 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node4669 = (inp[13]) ? node4673 : node4670;
														assign node4670 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4673 = (inp[14]) ? 4'b0100 : node4674;
															assign node4674 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node4678 = (inp[1]) ? node4698 : node4679;
													assign node4679 = (inp[12]) ? node4689 : node4680;
														assign node4680 = (inp[7]) ? node4686 : node4681;
															assign node4681 = (inp[13]) ? node4683 : 4'b1100;
																assign node4683 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4686 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node4689 = (inp[7]) ? node4695 : node4690;
															assign node4690 = (inp[13]) ? node4692 : 4'b0100;
																assign node4692 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node4695 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node4698 = (inp[13]) ? node4702 : node4699;
														assign node4699 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node4702 = (inp[7]) ? 4'b1100 : node4703;
															assign node4703 = (inp[14]) ? node4705 : 4'b1000;
																assign node4705 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node4709 = (inp[1]) ? node4763 : node4710;
											assign node4710 = (inp[15]) ? node4734 : node4711;
												assign node4711 = (inp[13]) ? node4725 : node4712;
													assign node4712 = (inp[7]) ? node4718 : node4713;
														assign node4713 = (inp[10]) ? node4715 : 4'b0000;
															assign node4715 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node4718 = (inp[10]) ? node4722 : node4719;
															assign node4719 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node4722 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node4725 = (inp[10]) ? node4727 : 4'b1000;
														assign node4727 = (inp[7]) ? node4731 : node4728;
															assign node4728 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node4731 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node4734 = (inp[7]) ? node4748 : node4735;
													assign node4735 = (inp[10]) ? node4741 : node4736;
														assign node4736 = (inp[12]) ? node4738 : 4'b0101;
															assign node4738 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node4741 = (inp[13]) ? node4745 : node4742;
															assign node4742 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node4745 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node4748 = (inp[13]) ? node4756 : node4749;
														assign node4749 = (inp[12]) ? node4753 : node4750;
															assign node4750 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node4753 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node4756 = (inp[10]) ? node4760 : node4757;
															assign node4757 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node4760 = (inp[12]) ? 4'b0101 : 4'b1101;
											assign node4763 = (inp[10]) ? node4797 : node4764;
												assign node4764 = (inp[15]) ? node4778 : node4765;
													assign node4765 = (inp[7]) ? node4773 : node4766;
														assign node4766 = (inp[13]) ? node4770 : node4767;
															assign node4767 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node4770 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node4773 = (inp[13]) ? node4775 : 4'b0101;
															assign node4775 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node4778 = (inp[12]) ? node4792 : node4779;
														assign node4779 = (inp[14]) ? node4785 : node4780;
															assign node4780 = (inp[13]) ? node4782 : 4'b0001;
																assign node4782 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node4785 = (inp[13]) ? node4789 : node4786;
																assign node4786 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node4789 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node4792 = (inp[7]) ? node4794 : 4'b0101;
															assign node4794 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node4797 = (inp[15]) ? node4803 : node4798;
													assign node4798 = (inp[13]) ? node4800 : 4'b0001;
														assign node4800 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node4803 = (inp[13]) ? node4807 : node4804;
														assign node4804 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node4807 = (inp[7]) ? 4'b1101 : 4'b1001;
									assign node4810 = (inp[1]) ? node4914 : node4811;
										assign node4811 = (inp[11]) ? node4887 : node4812;
											assign node4812 = (inp[12]) ? node4846 : node4813;
												assign node4813 = (inp[15]) ? node4829 : node4814;
													assign node4814 = (inp[10]) ? node4826 : node4815;
														assign node4815 = (inp[14]) ? node4823 : node4816;
															assign node4816 = (inp[7]) ? node4820 : node4817;
																assign node4817 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node4820 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node4823 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node4826 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node4829 = (inp[14]) ? node4837 : node4830;
														assign node4830 = (inp[7]) ? node4832 : 4'b0001;
															assign node4832 = (inp[13]) ? node4834 : 4'b1001;
																assign node4834 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node4837 = (inp[13]) ? node4841 : node4838;
															assign node4838 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node4841 = (inp[10]) ? 4'b0001 : node4842;
																assign node4842 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node4846 = (inp[14]) ? node4866 : node4847;
													assign node4847 = (inp[13]) ? node4859 : node4848;
														assign node4848 = (inp[10]) ? node4854 : node4849;
															assign node4849 = (inp[7]) ? 4'b1100 : node4850;
																assign node4850 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node4854 = (inp[7]) ? node4856 : 4'b1001;
																assign node4856 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node4859 = (inp[15]) ? node4861 : 4'b1001;
															assign node4861 = (inp[7]) ? node4863 : 4'b1001;
																assign node4863 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node4866 = (inp[15]) ? node4876 : node4867;
														assign node4867 = (inp[13]) ? 4'b1001 : node4868;
															assign node4868 = (inp[7]) ? node4872 : node4869;
																assign node4869 = (inp[10]) ? 4'b1001 : 4'b1100;
																assign node4872 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node4876 = (inp[13]) ? node4880 : node4877;
															assign node4877 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node4880 = (inp[10]) ? node4884 : node4881;
																assign node4881 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node4884 = (inp[7]) ? 4'b0100 : 4'b1001;
											assign node4887 = (inp[15]) ? node4903 : node4888;
												assign node4888 = (inp[13]) ? node4894 : node4889;
													assign node4889 = (inp[7]) ? node4891 : 4'b0001;
														assign node4891 = (inp[10]) ? 4'b0001 : 4'b0100;
													assign node4894 = (inp[10]) ? 4'b0000 : node4895;
														assign node4895 = (inp[12]) ? node4899 : node4896;
															assign node4896 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node4899 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4903 = (inp[13]) ? node4909 : node4904;
													assign node4904 = (inp[10]) ? node4906 : 4'b0000;
														assign node4906 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node4909 = (inp[7]) ? node4911 : 4'b0001;
														assign node4911 = (inp[10]) ? 4'b0001 : 4'b1000;
										assign node4914 = (inp[11]) ? node4980 : node4915;
											assign node4915 = (inp[12]) ? node4949 : node4916;
												assign node4916 = (inp[13]) ? node4940 : node4917;
													assign node4917 = (inp[14]) ? node4929 : node4918;
														assign node4918 = (inp[15]) ? node4924 : node4919;
															assign node4919 = (inp[7]) ? node4921 : 4'b1001;
																assign node4921 = (inp[10]) ? 4'b1001 : 4'b1100;
															assign node4924 = (inp[10]) ? node4926 : 4'b1000;
																assign node4926 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node4929 = (inp[15]) ? node4935 : node4930;
															assign node4930 = (inp[7]) ? node4932 : 4'b1001;
																assign node4932 = (inp[10]) ? 4'b1001 : 4'b0101;
															assign node4935 = (inp[7]) ? 4'b0001 : node4936;
																assign node4936 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node4940 = (inp[15]) ? 4'b1001 : node4941;
														assign node4941 = (inp[14]) ? node4943 : 4'b1001;
															assign node4943 = (inp[7]) ? node4945 : 4'b0000;
																assign node4945 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node4949 = (inp[15]) ? node4961 : node4950;
													assign node4950 = (inp[13]) ? node4958 : node4951;
														assign node4951 = (inp[7]) ? node4953 : 4'b0001;
															assign node4953 = (inp[10]) ? 4'b0001 : node4954;
																assign node4954 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node4958 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node4961 = (inp[14]) ? node4971 : node4962;
														assign node4962 = (inp[13]) ? node4966 : node4963;
															assign node4963 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node4966 = (inp[10]) ? 4'b0001 : node4967;
																assign node4967 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node4971 = (inp[10]) ? node4977 : node4972;
															assign node4972 = (inp[13]) ? node4974 : 4'b0001;
																assign node4974 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node4977 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node4980 = (inp[13]) ? node4996 : node4981;
												assign node4981 = (inp[15]) ? node4989 : node4982;
													assign node4982 = (inp[7]) ? node4984 : 4'b1001;
														assign node4984 = (inp[10]) ? 4'b1001 : node4985;
															assign node4985 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node4989 = (inp[10]) ? node4993 : node4990;
														assign node4990 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node4993 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node4996 = (inp[10]) ? 4'b1001 : node4997;
													assign node4997 = (inp[12]) ? node5003 : node4998;
														assign node4998 = (inp[15]) ? node5000 : 4'b1001;
															assign node5000 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node5003 = (inp[7]) ? 4'b1001 : node5004;
															assign node5004 = (inp[15]) ? 4'b1001 : 4'b0001;
								assign node5009 = (inp[15]) ? 4'b1001 : node5010;
									assign node5010 = (inp[4]) ? node5070 : node5011;
										assign node5011 = (inp[7]) ? 4'b1101 : node5012;
											assign node5012 = (inp[13]) ? node5038 : node5013;
												assign node5013 = (inp[10]) ? node5025 : node5014;
													assign node5014 = (inp[12]) ? 4'b1101 : node5015;
														assign node5015 = (inp[1]) ? node5019 : node5016;
															assign node5016 = (inp[11]) ? 4'b0000 : 4'b1101;
															assign node5019 = (inp[11]) ? 4'b0001 : node5020;
																assign node5020 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5025 = (inp[1]) ? node5033 : node5026;
														assign node5026 = (inp[14]) ? node5028 : 4'b0000;
															assign node5028 = (inp[11]) ? 4'b0000 : node5029;
																assign node5029 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node5033 = (inp[14]) ? node5035 : 4'b0001;
															assign node5035 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node5038 = (inp[10]) ? node5056 : node5039;
													assign node5039 = (inp[12]) ? node5045 : node5040;
														assign node5040 = (inp[11]) ? node5042 : 4'b1000;
															assign node5042 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node5045 = (inp[1]) ? node5051 : node5046;
															assign node5046 = (inp[14]) ? node5048 : 4'b0000;
																assign node5048 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node5051 = (inp[11]) ? 4'b0001 : node5052;
																assign node5052 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5056 = (inp[1]) ? node5064 : node5057;
														assign node5057 = (inp[14]) ? node5059 : 4'b1000;
															assign node5059 = (inp[11]) ? 4'b1000 : node5060;
																assign node5060 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5064 = (inp[11]) ? 4'b1001 : node5065;
															assign node5065 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node5070 = (inp[1]) ? node5112 : node5071;
											assign node5071 = (inp[11]) ? node5099 : node5072;
												assign node5072 = (inp[14]) ? node5086 : node5073;
													assign node5073 = (inp[13]) ? node5081 : node5074;
														assign node5074 = (inp[10]) ? 4'b0000 : node5075;
															assign node5075 = (inp[12]) ? node5077 : 4'b0000;
																assign node5077 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node5081 = (inp[10]) ? 4'b1000 : node5082;
															assign node5082 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node5086 = (inp[13]) ? node5094 : node5087;
														assign node5087 = (inp[7]) ? 4'b1101 : node5088;
															assign node5088 = (inp[12]) ? 4'b1001 : node5089;
																assign node5089 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node5094 = (inp[10]) ? node5096 : 4'b0001;
															assign node5096 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node5099 = (inp[13]) ? node5107 : node5100;
													assign node5100 = (inp[12]) ? node5102 : 4'b0000;
														assign node5102 = (inp[10]) ? 4'b0000 : node5103;
															assign node5103 = (inp[7]) ? 4'b1101 : 4'b1000;
													assign node5107 = (inp[10]) ? 4'b1000 : node5108;
														assign node5108 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node5112 = (inp[14]) ? node5126 : node5113;
												assign node5113 = (inp[13]) ? node5121 : node5114;
													assign node5114 = (inp[12]) ? node5116 : 4'b0001;
														assign node5116 = (inp[10]) ? 4'b0001 : node5117;
															assign node5117 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node5121 = (inp[10]) ? 4'b1001 : node5122;
														assign node5122 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node5126 = (inp[11]) ? node5140 : node5127;
													assign node5127 = (inp[13]) ? node5135 : node5128;
														assign node5128 = (inp[12]) ? node5130 : 4'b0000;
															assign node5130 = (inp[10]) ? 4'b0000 : node5131;
																assign node5131 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node5135 = (inp[12]) ? node5137 : 4'b1000;
															assign node5137 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node5140 = (inp[12]) ? node5144 : node5141;
														assign node5141 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node5144 = (inp[7]) ? node5150 : node5145;
															assign node5145 = (inp[13]) ? 4'b0001 : node5146;
																assign node5146 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node5150 = (inp[10]) ? node5154 : node5151;
																assign node5151 = (inp[13]) ? 4'b0001 : 4'b1101;
																assign node5154 = (inp[13]) ? 4'b1001 : 4'b0001;
						assign node5158 = (inp[4]) ? node6028 : node5159;
							assign node5159 = (inp[1]) ? node5631 : node5160;
								assign node5160 = (inp[2]) ? node5400 : node5161;
									assign node5161 = (inp[11]) ? node5295 : node5162;
										assign node5162 = (inp[0]) ? node5230 : node5163;
											assign node5163 = (inp[13]) ? node5189 : node5164;
												assign node5164 = (inp[10]) ? node5172 : node5165;
													assign node5165 = (inp[7]) ? node5167 : 4'b0001;
														assign node5167 = (inp[14]) ? 4'b0000 : node5168;
															assign node5168 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node5172 = (inp[7]) ? node5180 : node5173;
														assign node5173 = (inp[15]) ? 4'b0001 : node5174;
															assign node5174 = (inp[14]) ? node5176 : 4'b1000;
																assign node5176 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5180 = (inp[15]) ? node5182 : 4'b0001;
															assign node5182 = (inp[14]) ? node5186 : node5183;
																assign node5183 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node5186 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node5189 = (inp[10]) ? node5211 : node5190;
													assign node5190 = (inp[15]) ? node5200 : node5191;
														assign node5191 = (inp[7]) ? node5197 : node5192;
															assign node5192 = (inp[14]) ? 4'b0000 : node5193;
																assign node5193 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node5197 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5200 = (inp[14]) ? node5208 : node5201;
															assign node5201 = (inp[7]) ? node5205 : node5202;
																assign node5202 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node5205 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node5208 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node5211 = (inp[15]) ? node5223 : node5212;
														assign node5212 = (inp[12]) ? node5218 : node5213;
															assign node5213 = (inp[7]) ? 4'b1001 : node5214;
																assign node5214 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node5218 = (inp[14]) ? 4'b0001 : node5219;
																assign node5219 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node5223 = (inp[7]) ? node5227 : node5224;
															assign node5224 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5227 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node5230 = (inp[12]) ? node5264 : node5231;
												assign node5231 = (inp[15]) ? node5243 : node5232;
													assign node5232 = (inp[13]) ? node5234 : 4'b0001;
														assign node5234 = (inp[7]) ? node5240 : node5235;
															assign node5235 = (inp[14]) ? node5237 : 4'b1000;
																assign node5237 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node5240 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node5243 = (inp[13]) ? node5255 : node5244;
														assign node5244 = (inp[10]) ? node5250 : node5245;
															assign node5245 = (inp[14]) ? 4'b0000 : node5246;
																assign node5246 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node5250 = (inp[14]) ? 4'b1000 : node5251;
																assign node5251 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node5255 = (inp[10]) ? node5261 : node5256;
															assign node5256 = (inp[7]) ? node5258 : 4'b0001;
																assign node5258 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5261 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node5264 = (inp[15]) ? node5284 : node5265;
													assign node5265 = (inp[10]) ? node5273 : node5266;
														assign node5266 = (inp[13]) ? node5270 : node5267;
															assign node5267 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5270 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node5273 = (inp[13]) ? node5279 : node5274;
															assign node5274 = (inp[7]) ? node5276 : 4'b1001;
																assign node5276 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node5279 = (inp[14]) ? node5281 : 4'b1000;
																assign node5281 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node5284 = (inp[13]) ? node5288 : node5285;
														assign node5285 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node5288 = (inp[14]) ? node5290 : 4'b0001;
															assign node5290 = (inp[10]) ? node5292 : 4'b0000;
																assign node5292 = (inp[7]) ? 4'b0000 : 4'b1001;
										assign node5295 = (inp[10]) ? node5347 : node5296;
											assign node5296 = (inp[0]) ? node5324 : node5297;
												assign node5297 = (inp[13]) ? node5313 : node5298;
													assign node5298 = (inp[12]) ? node5306 : node5299;
														assign node5299 = (inp[7]) ? node5303 : node5300;
															assign node5300 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node5303 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node5306 = (inp[15]) ? node5310 : node5307;
															assign node5307 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node5310 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node5313 = (inp[15]) ? node5319 : node5314;
														assign node5314 = (inp[7]) ? node5316 : 4'b1000;
															assign node5316 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5319 = (inp[12]) ? 4'b0000 : node5320;
															assign node5320 = (inp[7]) ? 4'b1000 : 4'b0001;
												assign node5324 = (inp[13]) ? node5334 : node5325;
													assign node5325 = (inp[7]) ? node5329 : node5326;
														assign node5326 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node5329 = (inp[15]) ? node5331 : 4'b0000;
															assign node5331 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node5334 = (inp[12]) ? node5340 : node5335;
														assign node5335 = (inp[15]) ? node5337 : 4'b0000;
															assign node5337 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node5340 = (inp[15]) ? node5344 : node5341;
															assign node5341 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node5344 = (inp[7]) ? 4'b1000 : 4'b0001;
											assign node5347 = (inp[0]) ? node5363 : node5348;
												assign node5348 = (inp[15]) ? node5356 : node5349;
													assign node5349 = (inp[12]) ? 4'b0000 : node5350;
														assign node5350 = (inp[7]) ? 4'b0000 : node5351;
															assign node5351 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node5356 = (inp[7]) ? node5360 : node5357;
														assign node5357 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node5360 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5363 = (inp[7]) ? node5377 : node5364;
													assign node5364 = (inp[15]) ? node5372 : node5365;
														assign node5365 = (inp[12]) ? node5369 : node5366;
															assign node5366 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node5369 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node5372 = (inp[12]) ? node5374 : 4'b0000;
															assign node5374 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node5377 = (inp[14]) ? node5389 : node5378;
														assign node5378 = (inp[13]) ? node5384 : node5379;
															assign node5379 = (inp[15]) ? node5381 : 4'b0001;
																assign node5381 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node5384 = (inp[15]) ? 4'b0001 : node5385;
																assign node5385 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node5389 = (inp[12]) ? node5395 : node5390;
															assign node5390 = (inp[13]) ? 4'b0001 : node5391;
																assign node5391 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node5395 = (inp[13]) ? node5397 : 4'b0001;
																assign node5397 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node5400 = (inp[15]) ? node5542 : node5401;
										assign node5401 = (inp[11]) ? node5481 : node5402;
											assign node5402 = (inp[14]) ? node5438 : node5403;
												assign node5403 = (inp[13]) ? node5421 : node5404;
													assign node5404 = (inp[12]) ? node5414 : node5405;
														assign node5405 = (inp[10]) ? node5407 : 4'b0000;
															assign node5407 = (inp[7]) ? node5411 : node5408;
																assign node5408 = (inp[0]) ? 4'b1000 : 4'b0001;
																assign node5411 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node5414 = (inp[10]) ? node5418 : node5415;
															assign node5415 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node5418 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node5421 = (inp[10]) ? node5431 : node5422;
														assign node5422 = (inp[0]) ? node5426 : node5423;
															assign node5423 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node5426 = (inp[12]) ? node5428 : 4'b0000;
																assign node5428 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node5431 = (inp[0]) ? node5433 : 4'b0000;
															assign node5433 = (inp[7]) ? node5435 : 4'b0001;
																assign node5435 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5438 = (inp[7]) ? node5458 : node5439;
													assign node5439 = (inp[12]) ? node5447 : node5440;
														assign node5440 = (inp[0]) ? node5442 : 4'b0000;
															assign node5442 = (inp[10]) ? node5444 : 4'b0000;
																assign node5444 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node5447 = (inp[0]) ? node5453 : node5448;
															assign node5448 = (inp[10]) ? 4'b1001 : node5449;
																assign node5449 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node5453 = (inp[10]) ? 4'b0000 : node5454;
																assign node5454 = (inp[13]) ? 4'b1000 : 4'b1001;
													assign node5458 = (inp[13]) ? node5468 : node5459;
														assign node5459 = (inp[10]) ? node5465 : node5460;
															assign node5460 = (inp[12]) ? 4'b1001 : node5461;
																assign node5461 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node5465 = (inp[0]) ? 4'b0001 : 4'b1000;
														assign node5468 = (inp[12]) ? node5476 : node5469;
															assign node5469 = (inp[0]) ? node5473 : node5470;
																assign node5470 = (inp[10]) ? 4'b0001 : 4'b1000;
																assign node5473 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node5476 = (inp[10]) ? 4'b0001 : node5477;
																assign node5477 = (inp[0]) ? 4'b0001 : 4'b1000;
											assign node5481 = (inp[7]) ? node5517 : node5482;
												assign node5482 = (inp[10]) ? node5494 : node5483;
													assign node5483 = (inp[0]) ? node5489 : node5484;
														assign node5484 = (inp[13]) ? 4'b1001 : node5485;
															assign node5485 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5489 = (inp[12]) ? node5491 : 4'b0001;
															assign node5491 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node5494 = (inp[12]) ? node5510 : node5495;
														assign node5495 = (inp[14]) ? node5503 : node5496;
															assign node5496 = (inp[0]) ? node5500 : node5497;
																assign node5497 = (inp[13]) ? 4'b1001 : 4'b1000;
																assign node5500 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node5503 = (inp[13]) ? node5507 : node5504;
																assign node5504 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node5507 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5510 = (inp[13]) ? node5514 : node5511;
															assign node5511 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node5514 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node5517 = (inp[10]) ? node5531 : node5518;
													assign node5518 = (inp[13]) ? node5526 : node5519;
														assign node5519 = (inp[12]) ? node5523 : node5520;
															assign node5520 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node5523 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node5526 = (inp[0]) ? node5528 : 4'b0000;
															assign node5528 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node5531 = (inp[13]) ? node5537 : node5532;
														assign node5532 = (inp[0]) ? 4'b0000 : node5533;
															assign node5533 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5537 = (inp[0]) ? node5539 : 4'b1000;
															assign node5539 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node5542 = (inp[0]) ? node5596 : node5543;
											assign node5543 = (inp[11]) ? node5573 : node5544;
												assign node5544 = (inp[13]) ? node5562 : node5545;
													assign node5545 = (inp[14]) ? node5557 : node5546;
														assign node5546 = (inp[7]) ? node5552 : node5547;
															assign node5547 = (inp[10]) ? node5549 : 4'b0000;
																assign node5549 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node5552 = (inp[10]) ? 4'b1000 : node5553;
																assign node5553 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5557 = (inp[12]) ? node5559 : 4'b0001;
															assign node5559 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node5562 = (inp[10]) ? node5564 : 4'b0000;
														assign node5564 = (inp[7]) ? node5566 : 4'b0001;
															assign node5566 = (inp[14]) ? node5570 : node5567;
																assign node5567 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node5570 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node5573 = (inp[10]) ? node5583 : node5574;
													assign node5574 = (inp[7]) ? node5580 : node5575;
														assign node5575 = (inp[12]) ? 4'b0000 : node5576;
															assign node5576 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node5580 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5583 = (inp[7]) ? node5591 : node5584;
														assign node5584 = (inp[12]) ? node5588 : node5585;
															assign node5585 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node5588 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node5591 = (inp[12]) ? 4'b1000 : node5592;
															assign node5592 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node5596 = (inp[7]) ? 4'b1001 : node5597;
												assign node5597 = (inp[14]) ? node5609 : node5598;
													assign node5598 = (inp[13]) ? node5604 : node5599;
														assign node5599 = (inp[12]) ? node5601 : 4'b0000;
															assign node5601 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node5604 = (inp[12]) ? node5606 : 4'b1000;
															assign node5606 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node5609 = (inp[11]) ? node5621 : node5610;
														assign node5610 = (inp[13]) ? node5616 : node5611;
															assign node5611 = (inp[10]) ? node5613 : 4'b1001;
																assign node5613 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5616 = (inp[12]) ? 4'b0001 : node5617;
																assign node5617 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node5621 = (inp[13]) ? node5625 : node5622;
															assign node5622 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node5625 = (inp[12]) ? node5627 : 4'b1000;
																assign node5627 = (inp[10]) ? 4'b1000 : 4'b0000;
								assign node5631 = (inp[11]) ? node5885 : node5632;
									assign node5632 = (inp[15]) ? node5754 : node5633;
										assign node5633 = (inp[2]) ? node5697 : node5634;
											assign node5634 = (inp[13]) ? node5664 : node5635;
												assign node5635 = (inp[7]) ? node5649 : node5636;
													assign node5636 = (inp[10]) ? node5642 : node5637;
														assign node5637 = (inp[12]) ? 4'b0001 : node5638;
															assign node5638 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node5642 = (inp[0]) ? node5644 : 4'b0000;
															assign node5644 = (inp[12]) ? 4'b0001 : node5645;
																assign node5645 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5649 = (inp[10]) ? node5657 : node5650;
														assign node5650 = (inp[14]) ? 4'b0001 : node5651;
															assign node5651 = (inp[0]) ? node5653 : 4'b0001;
																assign node5653 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5657 = (inp[14]) ? node5659 : 4'b1001;
															assign node5659 = (inp[0]) ? node5661 : 4'b1000;
																assign node5661 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node5664 = (inp[10]) ? node5682 : node5665;
													assign node5665 = (inp[0]) ? node5675 : node5666;
														assign node5666 = (inp[14]) ? 4'b0001 : node5667;
															assign node5667 = (inp[7]) ? node5671 : node5668;
																assign node5668 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node5671 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5675 = (inp[14]) ? 4'b0000 : node5676;
															assign node5676 = (inp[12]) ? 4'b0001 : node5677;
																assign node5677 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node5682 = (inp[0]) ? node5690 : node5683;
														assign node5683 = (inp[12]) ? node5685 : 4'b0000;
															assign node5685 = (inp[14]) ? 4'b1000 : node5686;
																assign node5686 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node5690 = (inp[14]) ? node5694 : node5691;
															assign node5691 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node5694 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node5697 = (inp[0]) ? node5729 : node5698;
												assign node5698 = (inp[13]) ? node5714 : node5699;
													assign node5699 = (inp[12]) ? node5705 : node5700;
														assign node5700 = (inp[10]) ? node5702 : 4'b0000;
															assign node5702 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node5705 = (inp[10]) ? node5711 : node5706;
															assign node5706 = (inp[14]) ? 4'b1000 : node5707;
																assign node5707 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node5711 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node5714 = (inp[10]) ? node5722 : node5715;
														assign node5715 = (inp[12]) ? 4'b0001 : node5716;
															assign node5716 = (inp[7]) ? 4'b0001 : node5717;
																assign node5717 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5722 = (inp[7]) ? 4'b0000 : node5723;
															assign node5723 = (inp[14]) ? node5725 : 4'b0000;
																assign node5725 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node5729 = (inp[10]) ? node5741 : node5730;
													assign node5730 = (inp[7]) ? node5732 : 4'b0000;
														assign node5732 = (inp[13]) ? 4'b0000 : node5733;
															assign node5733 = (inp[14]) ? node5737 : node5734;
																assign node5734 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node5737 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node5741 = (inp[13]) ? node5747 : node5742;
														assign node5742 = (inp[7]) ? node5744 : 4'b1000;
															assign node5744 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node5747 = (inp[7]) ? 4'b1000 : node5748;
															assign node5748 = (inp[14]) ? node5750 : 4'b1000;
																assign node5750 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node5754 = (inp[10]) ? node5838 : node5755;
											assign node5755 = (inp[2]) ? node5795 : node5756;
												assign node5756 = (inp[13]) ? node5776 : node5757;
													assign node5757 = (inp[14]) ? node5765 : node5758;
														assign node5758 = (inp[0]) ? node5760 : 4'b0000;
															assign node5760 = (inp[7]) ? 4'b0000 : node5761;
																assign node5761 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node5765 = (inp[12]) ? node5771 : node5766;
															assign node5766 = (inp[7]) ? node5768 : 4'b0001;
																assign node5768 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node5771 = (inp[7]) ? node5773 : 4'b1001;
																assign node5773 = (inp[0]) ? 4'b0000 : 4'b1000;
													assign node5776 = (inp[0]) ? node5786 : node5777;
														assign node5777 = (inp[7]) ? node5779 : 4'b1000;
															assign node5779 = (inp[12]) ? node5783 : node5780;
																assign node5780 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node5783 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node5786 = (inp[14]) ? 4'b1001 : node5787;
															assign node5787 = (inp[7]) ? node5791 : node5788;
																assign node5788 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node5791 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node5795 = (inp[13]) ? node5815 : node5796;
													assign node5796 = (inp[14]) ? node5808 : node5797;
														assign node5797 = (inp[7]) ? node5803 : node5798;
															assign node5798 = (inp[0]) ? node5800 : 4'b1001;
																assign node5800 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node5803 = (inp[0]) ? 4'b1001 : node5804;
																assign node5804 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node5808 = (inp[7]) ? node5812 : node5809;
															assign node5809 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node5812 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5815 = (inp[0]) ? node5829 : node5816;
														assign node5816 = (inp[14]) ? node5822 : node5817;
															assign node5817 = (inp[12]) ? 4'b1000 : node5818;
																assign node5818 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node5822 = (inp[7]) ? node5826 : node5823;
																assign node5823 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node5826 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node5829 = (inp[7]) ? 4'b1001 : node5830;
															assign node5830 = (inp[14]) ? node5834 : node5831;
																assign node5831 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node5834 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node5838 = (inp[0]) ? node5864 : node5839;
												assign node5839 = (inp[2]) ? node5849 : node5840;
													assign node5840 = (inp[13]) ? node5842 : 4'b0001;
														assign node5842 = (inp[12]) ? node5844 : 4'b0001;
															assign node5844 = (inp[14]) ? 4'b1001 : node5845;
																assign node5845 = (inp[7]) ? 4'b0000 : 4'b1001;
													assign node5849 = (inp[13]) ? node5859 : node5850;
														assign node5850 = (inp[7]) ? node5854 : node5851;
															assign node5851 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node5854 = (inp[14]) ? 4'b0000 : node5855;
																assign node5855 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5859 = (inp[14]) ? node5861 : 4'b0001;
															assign node5861 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node5864 = (inp[2]) ? node5876 : node5865;
													assign node5865 = (inp[13]) ? node5873 : node5866;
														assign node5866 = (inp[14]) ? node5868 : 4'b0000;
															assign node5868 = (inp[12]) ? node5870 : 4'b0001;
																assign node5870 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node5873 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node5876 = (inp[7]) ? 4'b1001 : node5877;
														assign node5877 = (inp[13]) ? node5881 : node5878;
															assign node5878 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node5881 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node5885 = (inp[13]) ? node5991 : node5886;
										assign node5886 = (inp[10]) ? node5922 : node5887;
											assign node5887 = (inp[2]) ? node5907 : node5888;
												assign node5888 = (inp[15]) ? node5900 : node5889;
													assign node5889 = (inp[0]) ? node5895 : node5890;
														assign node5890 = (inp[12]) ? 4'b1001 : node5891;
															assign node5891 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node5895 = (inp[12]) ? node5897 : 4'b1001;
															assign node5897 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node5900 = (inp[12]) ? 4'b0001 : node5901;
														assign node5901 = (inp[7]) ? node5903 : 4'b1001;
															assign node5903 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node5907 = (inp[12]) ? node5915 : node5908;
													assign node5908 = (inp[7]) ? node5910 : 4'b0001;
														assign node5910 = (inp[15]) ? node5912 : 4'b0001;
															assign node5912 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node5915 = (inp[15]) ? 4'b1001 : node5916;
														assign node5916 = (inp[0]) ? node5918 : 4'b0001;
															assign node5918 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node5922 = (inp[14]) ? node5964 : node5923;
												assign node5923 = (inp[2]) ? node5943 : node5924;
													assign node5924 = (inp[7]) ? node5930 : node5925;
														assign node5925 = (inp[0]) ? 4'b0001 : node5926;
															assign node5926 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node5930 = (inp[12]) ? node5938 : node5931;
															assign node5931 = (inp[0]) ? node5935 : node5932;
																assign node5932 = (inp[15]) ? 4'b1001 : 4'b0001;
																assign node5935 = (inp[15]) ? 4'b0001 : 4'b1001;
															assign node5938 = (inp[15]) ? 4'b0001 : node5939;
																assign node5939 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node5943 = (inp[7]) ? node5959 : node5944;
														assign node5944 = (inp[12]) ? node5952 : node5945;
															assign node5945 = (inp[0]) ? node5949 : node5946;
																assign node5946 = (inp[15]) ? 4'b1001 : 4'b0001;
																assign node5949 = (inp[15]) ? 4'b0001 : 4'b1001;
															assign node5952 = (inp[0]) ? node5956 : node5953;
																assign node5953 = (inp[15]) ? 4'b1001 : 4'b0001;
																assign node5956 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node5959 = (inp[0]) ? node5961 : 4'b0001;
															assign node5961 = (inp[15]) ? 4'b1001 : 4'b0001;
												assign node5964 = (inp[7]) ? node5978 : node5965;
													assign node5965 = (inp[15]) ? node5973 : node5966;
														assign node5966 = (inp[2]) ? node5970 : node5967;
															assign node5967 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node5970 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node5973 = (inp[0]) ? 4'b0001 : node5974;
															assign node5974 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node5978 = (inp[15]) ? node5984 : node5979;
														assign node5979 = (inp[0]) ? node5981 : 4'b0001;
															assign node5981 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node5984 = (inp[2]) ? node5988 : node5985;
															assign node5985 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node5988 = (inp[0]) ? 4'b1001 : 4'b0001;
										assign node5991 = (inp[10]) ? 4'b1001 : node5992;
											assign node5992 = (inp[15]) ? node6008 : node5993;
												assign node5993 = (inp[0]) ? node6001 : node5994;
													assign node5994 = (inp[7]) ? 4'b1001 : node5995;
														assign node5995 = (inp[2]) ? node5997 : 4'b1001;
															assign node5997 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node6001 = (inp[12]) ? 4'b0001 : node6002;
														assign node6002 = (inp[2]) ? 4'b0001 : node6003;
															assign node6003 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node6008 = (inp[0]) ? node6016 : node6009;
													assign node6009 = (inp[2]) ? node6011 : 4'b0001;
														assign node6011 = (inp[12]) ? node6013 : 4'b0001;
															assign node6013 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node6016 = (inp[7]) ? node6022 : node6017;
														assign node6017 = (inp[2]) ? node6019 : 4'b1001;
															assign node6019 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6022 = (inp[2]) ? 4'b1001 : node6023;
															assign node6023 = (inp[12]) ? 4'b1001 : 4'b0001;
							assign node6028 = (inp[13]) ? node6504 : node6029;
								assign node6029 = (inp[1]) ? node6293 : node6030;
									assign node6030 = (inp[10]) ? node6168 : node6031;
										assign node6031 = (inp[0]) ? node6097 : node6032;
											assign node6032 = (inp[2]) ? node6062 : node6033;
												assign node6033 = (inp[7]) ? node6045 : node6034;
													assign node6034 = (inp[15]) ? 4'b1000 : node6035;
														assign node6035 = (inp[12]) ? node6041 : node6036;
															assign node6036 = (inp[11]) ? 4'b0001 : node6037;
																assign node6037 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node6041 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node6045 = (inp[11]) ? node6055 : node6046;
														assign node6046 = (inp[14]) ? node6050 : node6047;
															assign node6047 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node6050 = (inp[15]) ? node6052 : 4'b1000;
																assign node6052 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6055 = (inp[12]) ? node6059 : node6056;
															assign node6056 = (inp[15]) ? 4'b1001 : 4'b0000;
															assign node6059 = (inp[15]) ? 4'b0001 : 4'b1001;
												assign node6062 = (inp[12]) ? node6078 : node6063;
													assign node6063 = (inp[7]) ? node6071 : node6064;
														assign node6064 = (inp[11]) ? node6068 : node6065;
															assign node6065 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node6068 = (inp[15]) ? 4'b0000 : 4'b1000;
														assign node6071 = (inp[11]) ? 4'b0001 : node6072;
															assign node6072 = (inp[15]) ? node6074 : 4'b1000;
																assign node6074 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node6078 = (inp[15]) ? node6088 : node6079;
														assign node6079 = (inp[14]) ? node6081 : 4'b0001;
															assign node6081 = (inp[7]) ? node6085 : node6082;
																assign node6082 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node6085 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node6088 = (inp[11]) ? node6094 : node6089;
															assign node6089 = (inp[14]) ? node6091 : 4'b0000;
																assign node6091 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6094 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node6097 = (inp[7]) ? node6133 : node6098;
												assign node6098 = (inp[15]) ? node6118 : node6099;
													assign node6099 = (inp[12]) ? node6105 : node6100;
														assign node6100 = (inp[11]) ? node6102 : 4'b0001;
															assign node6102 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node6105 = (inp[14]) ? node6113 : node6106;
															assign node6106 = (inp[2]) ? node6110 : node6107;
																assign node6107 = (inp[11]) ? 4'b1001 : 4'b0001;
																assign node6110 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node6113 = (inp[11]) ? 4'b0001 : node6114;
																assign node6114 = (inp[2]) ? 4'b1000 : 4'b0001;
													assign node6118 = (inp[11]) ? node6126 : node6119;
														assign node6119 = (inp[12]) ? node6121 : 4'b0000;
															assign node6121 = (inp[2]) ? node6123 : 4'b0000;
																assign node6123 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6126 = (inp[2]) ? node6130 : node6127;
															assign node6127 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node6130 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node6133 = (inp[11]) ? node6157 : node6134;
													assign node6134 = (inp[2]) ? node6150 : node6135;
														assign node6135 = (inp[12]) ? node6143 : node6136;
															assign node6136 = (inp[15]) ? node6140 : node6137;
																assign node6137 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node6140 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6143 = (inp[14]) ? node6147 : node6144;
																assign node6144 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node6147 = (inp[15]) ? 4'b1001 : 4'b0000;
														assign node6150 = (inp[15]) ? node6152 : 4'b1000;
															assign node6152 = (inp[12]) ? 4'b1001 : node6153;
																assign node6153 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node6157 = (inp[2]) ? node6163 : node6158;
														assign node6158 = (inp[15]) ? node6160 : 4'b1000;
															assign node6160 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node6163 = (inp[15]) ? node6165 : 4'b0000;
															assign node6165 = (inp[12]) ? 4'b1001 : 4'b0000;
										assign node6168 = (inp[11]) ? node6244 : node6169;
											assign node6169 = (inp[12]) ? node6201 : node6170;
												assign node6170 = (inp[7]) ? node6182 : node6171;
													assign node6171 = (inp[2]) ? node6177 : node6172;
														assign node6172 = (inp[14]) ? node6174 : 4'b0001;
															assign node6174 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node6177 = (inp[0]) ? 4'b1000 : node6178;
															assign node6178 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node6182 = (inp[0]) ? node6194 : node6183;
														assign node6183 = (inp[2]) ? node6189 : node6184;
															assign node6184 = (inp[14]) ? node6186 : 4'b1000;
																assign node6186 = (inp[15]) ? 4'b1000 : 4'b0001;
															assign node6189 = (inp[15]) ? 4'b1001 : node6190;
																assign node6190 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6194 = (inp[2]) ? 4'b0001 : node6195;
															assign node6195 = (inp[14]) ? 4'b0000 : node6196;
																assign node6196 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node6201 = (inp[2]) ? node6225 : node6202;
													assign node6202 = (inp[0]) ? node6214 : node6203;
														assign node6203 = (inp[7]) ? node6209 : node6204;
															assign node6204 = (inp[14]) ? 4'b1000 : node6205;
																assign node6205 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node6209 = (inp[14]) ? node6211 : 4'b0000;
																assign node6211 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node6214 = (inp[7]) ? node6220 : node6215;
															assign node6215 = (inp[15]) ? 4'b0001 : node6216;
																assign node6216 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node6220 = (inp[14]) ? node6222 : 4'b1000;
																assign node6222 = (inp[15]) ? 4'b1000 : 4'b0001;
													assign node6225 = (inp[15]) ? node6239 : node6226;
														assign node6226 = (inp[0]) ? node6234 : node6227;
															assign node6227 = (inp[14]) ? node6231 : node6228;
																assign node6228 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node6231 = (inp[7]) ? 4'b0000 : 4'b1001;
															assign node6234 = (inp[7]) ? node6236 : 4'b0000;
																assign node6236 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6239 = (inp[7]) ? node6241 : 4'b0000;
															assign node6241 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node6244 = (inp[0]) ? node6270 : node6245;
												assign node6245 = (inp[15]) ? node6257 : node6246;
													assign node6246 = (inp[7]) ? node6252 : node6247;
														assign node6247 = (inp[2]) ? node6249 : 4'b0000;
															assign node6249 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node6252 = (inp[2]) ? 4'b0000 : node6253;
															assign node6253 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node6257 = (inp[2]) ? node6263 : node6258;
														assign node6258 = (inp[12]) ? node6260 : 4'b0001;
															assign node6260 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node6263 = (inp[12]) ? node6267 : node6264;
															assign node6264 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node6267 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node6270 = (inp[15]) ? node6282 : node6271;
													assign node6271 = (inp[12]) ? node6277 : node6272;
														assign node6272 = (inp[2]) ? 4'b0001 : node6273;
															assign node6273 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6277 = (inp[2]) ? node6279 : 4'b0001;
															assign node6279 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node6282 = (inp[12]) ? node6288 : node6283;
														assign node6283 = (inp[7]) ? node6285 : 4'b0000;
															assign node6285 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node6288 = (inp[2]) ? node6290 : 4'b0000;
															assign node6290 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node6293 = (inp[11]) ? node6443 : node6294;
										assign node6294 = (inp[10]) ? node6370 : node6295;
											assign node6295 = (inp[15]) ? node6329 : node6296;
												assign node6296 = (inp[0]) ? node6310 : node6297;
													assign node6297 = (inp[12]) ? 4'b0000 : node6298;
														assign node6298 = (inp[7]) ? node6304 : node6299;
															assign node6299 = (inp[14]) ? node6301 : 4'b1000;
																assign node6301 = (inp[2]) ? 4'b1000 : 4'b0001;
															assign node6304 = (inp[2]) ? node6306 : 4'b0000;
																assign node6306 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6310 = (inp[12]) ? node6320 : node6311;
														assign node6311 = (inp[7]) ? node6315 : node6312;
															assign node6312 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node6315 = (inp[2]) ? node6317 : 4'b0001;
																assign node6317 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node6320 = (inp[7]) ? node6324 : node6321;
															assign node6321 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node6324 = (inp[14]) ? 4'b0001 : node6325;
																assign node6325 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node6329 = (inp[12]) ? node6351 : node6330;
													assign node6330 = (inp[7]) ? node6340 : node6331;
														assign node6331 = (inp[0]) ? node6337 : node6332;
															assign node6332 = (inp[14]) ? node6334 : 4'b0001;
																assign node6334 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node6337 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node6340 = (inp[14]) ? node6346 : node6341;
															assign node6341 = (inp[2]) ? node6343 : 4'b0000;
																assign node6343 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node6346 = (inp[0]) ? 4'b0000 : node6347;
																assign node6347 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node6351 = (inp[7]) ? node6363 : node6352;
														assign node6352 = (inp[0]) ? node6358 : node6353;
															assign node6353 = (inp[14]) ? 4'b1001 : node6354;
																assign node6354 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6358 = (inp[2]) ? 4'b0000 : node6359;
																assign node6359 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node6363 = (inp[0]) ? node6365 : 4'b1000;
															assign node6365 = (inp[2]) ? 4'b1001 : node6366;
																assign node6366 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node6370 = (inp[12]) ? node6398 : node6371;
												assign node6371 = (inp[14]) ? node6379 : node6372;
													assign node6372 = (inp[7]) ? node6376 : node6373;
														assign node6373 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node6376 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node6379 = (inp[2]) ? node6389 : node6380;
														assign node6380 = (inp[0]) ? node6386 : node6381;
															assign node6381 = (inp[7]) ? node6383 : 4'b0001;
																assign node6383 = (inp[15]) ? 4'b1000 : 4'b0000;
															assign node6386 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6389 = (inp[0]) ? node6393 : node6390;
															assign node6390 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6393 = (inp[7]) ? 4'b0000 : node6394;
																assign node6394 = (inp[15]) ? 4'b0001 : 4'b1000;
												assign node6398 = (inp[15]) ? node6420 : node6399;
													assign node6399 = (inp[7]) ? node6411 : node6400;
														assign node6400 = (inp[0]) ? node6406 : node6401;
															assign node6401 = (inp[2]) ? 4'b0001 : node6402;
																assign node6402 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node6406 = (inp[2]) ? 4'b0000 : node6407;
																assign node6407 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node6411 = (inp[0]) ? node6417 : node6412;
															assign node6412 = (inp[14]) ? node6414 : 4'b0000;
																assign node6414 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node6417 = (inp[2]) ? 4'b0001 : 4'b1000;
													assign node6420 = (inp[2]) ? node6428 : node6421;
														assign node6421 = (inp[7]) ? node6425 : node6422;
															assign node6422 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6425 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node6428 = (inp[0]) ? node6436 : node6429;
															assign node6429 = (inp[7]) ? node6433 : node6430;
																assign node6430 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node6433 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6436 = (inp[7]) ? node6440 : node6437;
																assign node6437 = (inp[14]) ? 4'b1000 : 4'b0000;
																assign node6440 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node6443 = (inp[10]) ? 4'b0001 : node6444;
											assign node6444 = (inp[12]) ? node6476 : node6445;
												assign node6445 = (inp[7]) ? node6463 : node6446;
													assign node6446 = (inp[14]) ? node6454 : node6447;
														assign node6447 = (inp[2]) ? 4'b0001 : node6448;
															assign node6448 = (inp[15]) ? node6450 : 4'b0001;
																assign node6450 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node6454 = (inp[2]) ? node6458 : node6455;
															assign node6455 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node6458 = (inp[0]) ? 4'b0001 : node6459;
																assign node6459 = (inp[15]) ? 4'b0001 : 4'b1001;
													assign node6463 = (inp[15]) ? node6471 : node6464;
														assign node6464 = (inp[0]) ? node6468 : node6465;
															assign node6465 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node6468 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node6471 = (inp[2]) ? node6473 : 4'b0001;
															assign node6473 = (inp[0]) ? 4'b0001 : 4'b1001;
												assign node6476 = (inp[0]) ? node6490 : node6477;
													assign node6477 = (inp[15]) ? node6483 : node6478;
														assign node6478 = (inp[7]) ? 4'b0001 : node6479;
															assign node6479 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node6483 = (inp[7]) ? node6487 : node6484;
															assign node6484 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node6487 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node6490 = (inp[7]) ? node6496 : node6491;
														assign node6491 = (inp[2]) ? node6493 : 4'b0001;
															assign node6493 = (inp[15]) ? 4'b0001 : 4'b1001;
														assign node6496 = (inp[15]) ? node6500 : node6497;
															assign node6497 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node6500 = (inp[2]) ? 4'b1001 : 4'b0001;
								assign node6504 = (inp[10]) ? node6728 : node6505;
									assign node6505 = (inp[1]) ? node6657 : node6506;
										assign node6506 = (inp[11]) ? node6590 : node6507;
											assign node6507 = (inp[14]) ? node6545 : node6508;
												assign node6508 = (inp[0]) ? node6522 : node6509;
													assign node6509 = (inp[7]) ? node6515 : node6510;
														assign node6510 = (inp[2]) ? node6512 : 4'b0001;
															assign node6512 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node6515 = (inp[2]) ? node6517 : 4'b0000;
															assign node6517 = (inp[12]) ? 4'b0001 : node6518;
																assign node6518 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node6522 = (inp[15]) ? node6532 : node6523;
														assign node6523 = (inp[2]) ? node6527 : node6524;
															assign node6524 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node6527 = (inp[12]) ? node6529 : 4'b0000;
																assign node6529 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6532 = (inp[12]) ? node6540 : node6533;
															assign node6533 = (inp[2]) ? node6537 : node6534;
																assign node6534 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node6537 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node6540 = (inp[7]) ? 4'b0000 : node6541;
																assign node6541 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node6545 = (inp[15]) ? node6569 : node6546;
													assign node6546 = (inp[2]) ? node6554 : node6547;
														assign node6547 = (inp[7]) ? 4'b0000 : node6548;
															assign node6548 = (inp[12]) ? node6550 : 4'b0000;
																assign node6550 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node6554 = (inp[12]) ? node6562 : node6555;
															assign node6555 = (inp[7]) ? node6559 : node6556;
																assign node6556 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node6559 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6562 = (inp[7]) ? node6566 : node6563;
																assign node6563 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node6566 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node6569 = (inp[2]) ? node6577 : node6570;
														assign node6570 = (inp[7]) ? node6574 : node6571;
															assign node6571 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node6574 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node6577 = (inp[12]) ? node6585 : node6578;
															assign node6578 = (inp[7]) ? node6582 : node6579;
																assign node6579 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node6582 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6585 = (inp[7]) ? node6587 : 4'b0000;
																assign node6587 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node6590 = (inp[15]) ? node6624 : node6591;
												assign node6591 = (inp[0]) ? node6603 : node6592;
													assign node6592 = (inp[12]) ? node6598 : node6593;
														assign node6593 = (inp[2]) ? 4'b0000 : node6594;
															assign node6594 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6598 = (inp[2]) ? node6600 : 4'b0000;
															assign node6600 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node6603 = (inp[7]) ? node6619 : node6604;
														assign node6604 = (inp[14]) ? node6612 : node6605;
															assign node6605 = (inp[12]) ? node6609 : node6606;
																assign node6606 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node6609 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node6612 = (inp[2]) ? node6616 : node6613;
																assign node6613 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node6616 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node6619 = (inp[12]) ? 4'b0000 : node6620;
															assign node6620 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node6624 = (inp[2]) ? node6644 : node6625;
													assign node6625 = (inp[0]) ? node6639 : node6626;
														assign node6626 = (inp[14]) ? node6634 : node6627;
															assign node6627 = (inp[7]) ? node6631 : node6628;
																assign node6628 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node6631 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node6634 = (inp[12]) ? 4'b0001 : node6635;
																assign node6635 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6639 = (inp[12]) ? node6641 : 4'b0000;
															assign node6641 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node6644 = (inp[12]) ? node6652 : node6645;
														assign node6645 = (inp[0]) ? node6649 : node6646;
															assign node6646 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node6649 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6652 = (inp[7]) ? 4'b0000 : node6653;
															assign node6653 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node6657 = (inp[11]) ? 4'b0001 : node6658;
											assign node6658 = (inp[15]) ? node6694 : node6659;
												assign node6659 = (inp[0]) ? node6675 : node6660;
													assign node6660 = (inp[2]) ? node6668 : node6661;
														assign node6661 = (inp[12]) ? 4'b0000 : node6662;
															assign node6662 = (inp[14]) ? node6664 : 4'b0000;
																assign node6664 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6668 = (inp[14]) ? 4'b0000 : node6669;
															assign node6669 = (inp[12]) ? node6671 : 4'b0000;
																assign node6671 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6675 = (inp[14]) ? node6687 : node6676;
														assign node6676 = (inp[7]) ? node6682 : node6677;
															assign node6677 = (inp[2]) ? node6679 : 4'b0001;
																assign node6679 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node6682 = (inp[12]) ? 4'b0001 : node6683;
																assign node6683 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node6687 = (inp[12]) ? node6689 : 4'b0000;
															assign node6689 = (inp[7]) ? node6691 : 4'b0001;
																assign node6691 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node6694 = (inp[0]) ? node6712 : node6695;
													assign node6695 = (inp[2]) ? node6701 : node6696;
														assign node6696 = (inp[12]) ? 4'b0001 : node6697;
															assign node6697 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node6701 = (inp[14]) ? node6707 : node6702;
															assign node6702 = (inp[7]) ? node6704 : 4'b0000;
																assign node6704 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node6707 = (inp[7]) ? 4'b0001 : node6708;
																assign node6708 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node6712 = (inp[12]) ? node6720 : node6713;
														assign node6713 = (inp[14]) ? node6715 : 4'b0000;
															assign node6715 = (inp[2]) ? 4'b0000 : node6716;
																assign node6716 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6720 = (inp[7]) ? 4'b0000 : node6721;
															assign node6721 = (inp[2]) ? node6723 : 4'b0000;
																assign node6723 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node6728 = (inp[11]) ? 4'b0000 : node6729;
										assign node6729 = (inp[1]) ? 4'b0000 : node6730;
											assign node6730 = (inp[14]) ? node6774 : node6731;
												assign node6731 = (inp[0]) ? node6759 : node6732;
													assign node6732 = (inp[7]) ? node6746 : node6733;
														assign node6733 = (inp[15]) ? node6741 : node6734;
															assign node6734 = (inp[2]) ? node6738 : node6735;
																assign node6735 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node6738 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node6741 = (inp[12]) ? node6743 : 4'b0000;
																assign node6743 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node6746 = (inp[12]) ? node6754 : node6747;
															assign node6747 = (inp[15]) ? node6751 : node6748;
																assign node6748 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node6751 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node6754 = (inp[15]) ? node6756 : 4'b0000;
																assign node6756 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node6759 = (inp[7]) ? node6761 : 4'b0000;
														assign node6761 = (inp[15]) ? node6769 : node6762;
															assign node6762 = (inp[2]) ? node6766 : node6763;
																assign node6763 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node6766 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node6769 = (inp[12]) ? node6771 : 4'b0000;
																assign node6771 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node6774 = (inp[2]) ? node6790 : node6775;
													assign node6775 = (inp[15]) ? node6779 : node6776;
														assign node6776 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node6779 = (inp[7]) ? node6785 : node6780;
															assign node6780 = (inp[12]) ? node6782 : 4'b0000;
																assign node6782 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6785 = (inp[0]) ? 4'b0001 : node6786;
																assign node6786 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node6790 = (inp[12]) ? node6804 : node6791;
														assign node6791 = (inp[7]) ? node6799 : node6792;
															assign node6792 = (inp[15]) ? node6796 : node6793;
																assign node6793 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node6796 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node6799 = (inp[15]) ? node6801 : 4'b0000;
																assign node6801 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node6804 = (inp[15]) ? node6806 : 4'b0000;
															assign node6806 = (inp[0]) ? node6808 : 4'b0000;
																assign node6808 = (inp[7]) ? 4'b0000 : 4'b0001;
			assign node6813 = (inp[15]) ? node10681 : node6814;
				assign node6814 = (inp[6]) ? node7756 : node6815;
					assign node6815 = (inp[0]) ? 4'b0101 : node6816;
						assign node6816 = (inp[5]) ? node7186 : node6817;
							assign node6817 = (inp[2]) ? 4'b0111 : node6818;
								assign node6818 = (inp[3]) ? node6942 : node6819;
									assign node6819 = (inp[4]) ? node6849 : node6820;
										assign node6820 = (inp[7]) ? 4'b0111 : node6821;
											assign node6821 = (inp[13]) ? node6823 : 4'b0111;
												assign node6823 = (inp[10]) ? node6835 : node6824;
													assign node6824 = (inp[12]) ? 4'b0111 : node6825;
														assign node6825 = (inp[1]) ? node6829 : node6826;
															assign node6826 = (inp[14]) ? 4'b0111 : 4'b0000;
															assign node6829 = (inp[14]) ? node6831 : 4'b0001;
																assign node6831 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node6835 = (inp[1]) ? node6843 : node6836;
														assign node6836 = (inp[11]) ? 4'b0000 : node6837;
															assign node6837 = (inp[14]) ? node6839 : 4'b0000;
																assign node6839 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node6843 = (inp[11]) ? 4'b0001 : node6844;
															assign node6844 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node6849 = (inp[7]) ? node6915 : node6850;
											assign node6850 = (inp[13]) ? node6880 : node6851;
												assign node6851 = (inp[10]) ? node6867 : node6852;
													assign node6852 = (inp[12]) ? node6858 : node6853;
														assign node6853 = (inp[1]) ? node6855 : 4'b0001;
															assign node6855 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6858 = (inp[1]) ? node6862 : node6859;
															assign node6859 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node6862 = (inp[11]) ? 4'b0001 : node6863;
																assign node6863 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6867 = (inp[1]) ? node6875 : node6868;
														assign node6868 = (inp[14]) ? node6870 : 4'b1000;
															assign node6870 = (inp[11]) ? 4'b1000 : node6871;
																assign node6871 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6875 = (inp[11]) ? 4'b1001 : node6876;
															assign node6876 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6880 = (inp[1]) ? node6898 : node6881;
													assign node6881 = (inp[11]) ? node6893 : node6882;
														assign node6882 = (inp[14]) ? node6888 : node6883;
															assign node6883 = (inp[10]) ? 4'b0000 : node6884;
																assign node6884 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node6888 = (inp[10]) ? node6890 : 4'b1001;
																assign node6890 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node6893 = (inp[10]) ? 4'b0000 : node6894;
															assign node6894 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node6898 = (inp[11]) ? node6910 : node6899;
														assign node6899 = (inp[14]) ? node6905 : node6900;
															assign node6900 = (inp[12]) ? node6902 : 4'b0001;
																assign node6902 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node6905 = (inp[12]) ? node6907 : 4'b0000;
																assign node6907 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node6910 = (inp[12]) ? node6912 : 4'b0001;
															assign node6912 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node6915 = (inp[13]) ? node6917 : 4'b0111;
												assign node6917 = (inp[10]) ? node6929 : node6918;
													assign node6918 = (inp[12]) ? 4'b0111 : node6919;
														assign node6919 = (inp[11]) ? 4'b0000 : node6920;
															assign node6920 = (inp[14]) ? node6924 : node6921;
																assign node6921 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node6924 = (inp[1]) ? 4'b0000 : 4'b0111;
													assign node6929 = (inp[1]) ? node6937 : node6930;
														assign node6930 = (inp[11]) ? 4'b0000 : node6931;
															assign node6931 = (inp[14]) ? node6933 : 4'b0000;
																assign node6933 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node6937 = (inp[14]) ? node6939 : 4'b0001;
															assign node6939 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node6942 = (inp[7]) ? node7074 : node6943;
										assign node6943 = (inp[4]) ? node7015 : node6944;
											assign node6944 = (inp[13]) ? node6980 : node6945;
												assign node6945 = (inp[10]) ? node6967 : node6946;
													assign node6946 = (inp[12]) ? node6956 : node6947;
														assign node6947 = (inp[1]) ? node6951 : node6948;
															assign node6948 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node6951 = (inp[11]) ? 4'b1001 : node6952;
																assign node6952 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6956 = (inp[1]) ? node6962 : node6957;
															assign node6957 = (inp[11]) ? 4'b0000 : node6958;
																assign node6958 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node6962 = (inp[11]) ? 4'b0001 : node6963;
																assign node6963 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6967 = (inp[1]) ? node6975 : node6968;
														assign node6968 = (inp[14]) ? node6970 : 4'b1000;
															assign node6970 = (inp[11]) ? 4'b1000 : node6971;
																assign node6971 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node6975 = (inp[11]) ? 4'b1001 : node6976;
															assign node6976 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6980 = (inp[10]) ? node7002 : node6981;
													assign node6981 = (inp[12]) ? node6991 : node6982;
														assign node6982 = (inp[1]) ? node6988 : node6983;
															assign node6983 = (inp[14]) ? node6985 : 4'b0100;
																assign node6985 = (inp[11]) ? 4'b0100 : 4'b1001;
															assign node6988 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node6991 = (inp[1]) ? node6997 : node6992;
															assign node6992 = (inp[11]) ? 4'b1000 : node6993;
																assign node6993 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node6997 = (inp[11]) ? 4'b1001 : node6998;
																assign node6998 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7002 = (inp[1]) ? node7010 : node7003;
														assign node7003 = (inp[14]) ? node7005 : 4'b0100;
															assign node7005 = (inp[11]) ? 4'b0100 : node7006;
																assign node7006 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node7010 = (inp[14]) ? node7012 : 4'b0101;
															assign node7012 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node7015 = (inp[1]) ? node7045 : node7016;
												assign node7016 = (inp[14]) ? node7028 : node7017;
													assign node7017 = (inp[13]) ? node7023 : node7018;
														assign node7018 = (inp[10]) ? 4'b1100 : node7019;
															assign node7019 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7023 = (inp[12]) ? node7025 : 4'b0100;
															assign node7025 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node7028 = (inp[11]) ? node7036 : node7029;
														assign node7029 = (inp[13]) ? 4'b1101 : node7030;
															assign node7030 = (inp[10]) ? node7032 : 4'b0101;
																assign node7032 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7036 = (inp[12]) ? node7040 : node7037;
															assign node7037 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node7040 = (inp[10]) ? 4'b1100 : node7041;
																assign node7041 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node7045 = (inp[11]) ? node7063 : node7046;
													assign node7046 = (inp[14]) ? node7052 : node7047;
														assign node7047 = (inp[13]) ? node7049 : 4'b1101;
															assign node7049 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node7052 = (inp[13]) ? node7058 : node7053;
															assign node7053 = (inp[10]) ? 4'b1100 : node7054;
																assign node7054 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node7058 = (inp[12]) ? node7060 : 4'b0100;
																assign node7060 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node7063 = (inp[13]) ? node7069 : node7064;
														assign node7064 = (inp[10]) ? 4'b1101 : node7065;
															assign node7065 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7069 = (inp[10]) ? 4'b0101 : node7070;
															assign node7070 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node7074 = (inp[13]) ? node7112 : node7075;
											assign node7075 = (inp[10]) ? node7099 : node7076;
												assign node7076 = (inp[12]) ? node7088 : node7077;
													assign node7077 = (inp[1]) ? node7083 : node7078;
														assign node7078 = (inp[11]) ? 4'b1000 : node7079;
															assign node7079 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node7083 = (inp[11]) ? 4'b1001 : node7084;
															assign node7084 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7088 = (inp[1]) ? node7094 : node7089;
														assign node7089 = (inp[11]) ? 4'b0000 : node7090;
															assign node7090 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node7094 = (inp[11]) ? 4'b0001 : node7095;
															assign node7095 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node7099 = (inp[1]) ? node7107 : node7100;
													assign node7100 = (inp[14]) ? node7102 : 4'b1000;
														assign node7102 = (inp[11]) ? 4'b1000 : node7103;
															assign node7103 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7107 = (inp[14]) ? node7109 : 4'b1001;
														assign node7109 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node7112 = (inp[4]) ? node7148 : node7113;
												assign node7113 = (inp[10]) ? node7135 : node7114;
													assign node7114 = (inp[12]) ? node7124 : node7115;
														assign node7115 = (inp[1]) ? node7119 : node7116;
															assign node7116 = (inp[11]) ? 4'b0000 : 4'b1001;
															assign node7119 = (inp[11]) ? 4'b0001 : node7120;
																assign node7120 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node7124 = (inp[1]) ? node7130 : node7125;
															assign node7125 = (inp[11]) ? 4'b1000 : node7126;
																assign node7126 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node7130 = (inp[14]) ? node7132 : 4'b1001;
																assign node7132 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node7135 = (inp[1]) ? node7143 : node7136;
														assign node7136 = (inp[14]) ? node7138 : 4'b0000;
															assign node7138 = (inp[11]) ? 4'b0000 : node7139;
																assign node7139 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node7143 = (inp[14]) ? node7145 : 4'b0001;
															assign node7145 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node7148 = (inp[12]) ? node7162 : node7149;
													assign node7149 = (inp[1]) ? node7157 : node7150;
														assign node7150 = (inp[14]) ? node7152 : 4'b0100;
															assign node7152 = (inp[11]) ? 4'b0100 : node7153;
																assign node7153 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node7157 = (inp[11]) ? 4'b0101 : node7158;
															assign node7158 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node7162 = (inp[10]) ? node7174 : node7163;
														assign node7163 = (inp[1]) ? node7169 : node7164;
															assign node7164 = (inp[14]) ? node7166 : 4'b1000;
																assign node7166 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node7169 = (inp[11]) ? 4'b1001 : node7170;
																assign node7170 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node7174 = (inp[1]) ? node7180 : node7175;
															assign node7175 = (inp[14]) ? node7177 : 4'b0100;
																assign node7177 = (inp[11]) ? 4'b0100 : 4'b1001;
															assign node7180 = (inp[14]) ? node7182 : 4'b0101;
																assign node7182 = (inp[11]) ? 4'b0101 : 4'b0100;
							assign node7186 = (inp[1]) ? node7478 : node7187;
								assign node7187 = (inp[11]) ? node7387 : node7188;
									assign node7188 = (inp[14]) ? node7288 : node7189;
										assign node7189 = (inp[3]) ? node7253 : node7190;
											assign node7190 = (inp[2]) ? node7226 : node7191;
												assign node7191 = (inp[13]) ? node7209 : node7192;
													assign node7192 = (inp[4]) ? node7198 : node7193;
														assign node7193 = (inp[10]) ? 4'b1100 : node7194;
															assign node7194 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node7198 = (inp[7]) ? node7204 : node7199;
															assign node7199 = (inp[10]) ? 4'b1000 : node7200;
																assign node7200 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node7204 = (inp[12]) ? node7206 : 4'b1100;
																assign node7206 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node7209 = (inp[7]) ? node7215 : node7210;
														assign node7210 = (inp[12]) ? node7212 : 4'b0000;
															assign node7212 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node7215 = (inp[4]) ? node7221 : node7216;
															assign node7216 = (inp[10]) ? 4'b0100 : node7217;
																assign node7217 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node7221 = (inp[10]) ? 4'b0000 : node7222;
																assign node7222 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node7226 = (inp[4]) ? node7234 : node7227;
													assign node7227 = (inp[7]) ? 4'b0111 : node7228;
														assign node7228 = (inp[13]) ? node7230 : 4'b0111;
															assign node7230 = (inp[10]) ? 4'b0000 : 4'b0111;
													assign node7234 = (inp[7]) ? node7246 : node7235;
														assign node7235 = (inp[13]) ? node7241 : node7236;
															assign node7236 = (inp[10]) ? 4'b1000 : node7237;
																assign node7237 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node7241 = (inp[12]) ? node7243 : 4'b0000;
																assign node7243 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node7246 = (inp[13]) ? node7248 : 4'b0111;
															assign node7248 = (inp[12]) ? node7250 : 4'b0000;
																assign node7250 = (inp[10]) ? 4'b0000 : 4'b0111;
											assign node7253 = (inp[13]) ? node7271 : node7254;
												assign node7254 = (inp[4]) ? node7260 : node7255;
													assign node7255 = (inp[10]) ? 4'b1000 : node7256;
														assign node7256 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node7260 = (inp[7]) ? node7266 : node7261;
														assign node7261 = (inp[12]) ? node7263 : 4'b1100;
															assign node7263 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node7266 = (inp[10]) ? 4'b1000 : node7267;
															assign node7267 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node7271 = (inp[12]) ? node7277 : node7272;
													assign node7272 = (inp[7]) ? node7274 : 4'b0100;
														assign node7274 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node7277 = (inp[10]) ? node7283 : node7278;
														assign node7278 = (inp[7]) ? 4'b1000 : node7279;
															assign node7279 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node7283 = (inp[7]) ? node7285 : 4'b0100;
															assign node7285 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node7288 = (inp[3]) ? node7352 : node7289;
											assign node7289 = (inp[2]) ? node7325 : node7290;
												assign node7290 = (inp[7]) ? node7312 : node7291;
													assign node7291 = (inp[4]) ? node7301 : node7292;
														assign node7292 = (inp[13]) ? node7298 : node7293;
															assign node7293 = (inp[10]) ? node7295 : 4'b0101;
																assign node7295 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7298 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node7301 = (inp[13]) ? node7307 : node7302;
															assign node7302 = (inp[10]) ? node7304 : 4'b0001;
																assign node7304 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7307 = (inp[12]) ? 4'b1001 : node7308;
																assign node7308 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node7312 = (inp[13]) ? node7318 : node7313;
														assign node7313 = (inp[10]) ? node7315 : 4'b0101;
															assign node7315 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7318 = (inp[12]) ? 4'b1101 : node7319;
															assign node7319 = (inp[10]) ? node7321 : 4'b1101;
																assign node7321 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node7325 = (inp[4]) ? node7335 : node7326;
													assign node7326 = (inp[7]) ? 4'b0111 : node7327;
														assign node7327 = (inp[10]) ? node7329 : 4'b0111;
															assign node7329 = (inp[13]) ? node7331 : 4'b0111;
																assign node7331 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node7335 = (inp[7]) ? node7345 : node7336;
														assign node7336 = (inp[13]) ? node7342 : node7337;
															assign node7337 = (inp[10]) ? node7339 : 4'b0001;
																assign node7339 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node7342 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node7345 = (inp[10]) ? node7347 : 4'b0111;
															assign node7347 = (inp[12]) ? 4'b0111 : node7348;
																assign node7348 = (inp[13]) ? 4'b0001 : 4'b0111;
											assign node7352 = (inp[13]) ? node7370 : node7353;
												assign node7353 = (inp[12]) ? node7365 : node7354;
													assign node7354 = (inp[10]) ? node7360 : node7355;
														assign node7355 = (inp[7]) ? 4'b0001 : node7356;
															assign node7356 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node7360 = (inp[4]) ? node7362 : 4'b1001;
															assign node7362 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7365 = (inp[7]) ? 4'b0001 : node7366;
														assign node7366 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node7370 = (inp[10]) ? node7376 : node7371;
													assign node7371 = (inp[4]) ? node7373 : 4'b1001;
														assign node7373 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node7376 = (inp[12]) ? node7382 : node7377;
														assign node7377 = (inp[7]) ? node7379 : 4'b0101;
															assign node7379 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node7382 = (inp[4]) ? node7384 : 4'b1001;
															assign node7384 = (inp[7]) ? 4'b1001 : 4'b1101;
									assign node7387 = (inp[13]) ? node7433 : node7388;
										assign node7388 = (inp[3]) ? node7416 : node7389;
											assign node7389 = (inp[2]) ? node7407 : node7390;
												assign node7390 = (inp[12]) ? node7396 : node7391;
													assign node7391 = (inp[7]) ? 4'b1100 : node7392;
														assign node7392 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node7396 = (inp[10]) ? node7402 : node7397;
														assign node7397 = (inp[7]) ? 4'b0100 : node7398;
															assign node7398 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7402 = (inp[4]) ? node7404 : 4'b1100;
															assign node7404 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node7407 = (inp[4]) ? node7409 : 4'b0111;
													assign node7409 = (inp[7]) ? 4'b0111 : node7410;
														assign node7410 = (inp[12]) ? node7412 : 4'b1000;
															assign node7412 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node7416 = (inp[12]) ? node7422 : node7417;
												assign node7417 = (inp[7]) ? 4'b1000 : node7418;
													assign node7418 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node7422 = (inp[10]) ? node7428 : node7423;
													assign node7423 = (inp[7]) ? 4'b0000 : node7424;
														assign node7424 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node7428 = (inp[7]) ? 4'b1000 : node7429;
														assign node7429 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node7433 = (inp[10]) ? node7465 : node7434;
											assign node7434 = (inp[12]) ? node7448 : node7435;
												assign node7435 = (inp[3]) ? node7443 : node7436;
													assign node7436 = (inp[7]) ? node7438 : 4'b0000;
														assign node7438 = (inp[2]) ? 4'b0111 : node7439;
															assign node7439 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node7443 = (inp[4]) ? 4'b0100 : node7444;
														assign node7444 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node7448 = (inp[3]) ? node7460 : node7449;
													assign node7449 = (inp[2]) ? node7455 : node7450;
														assign node7450 = (inp[7]) ? 4'b1100 : node7451;
															assign node7451 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node7455 = (inp[4]) ? node7457 : 4'b0111;
															assign node7457 = (inp[7]) ? 4'b0111 : 4'b1000;
													assign node7460 = (inp[7]) ? 4'b1000 : node7461;
														assign node7461 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node7465 = (inp[3]) ? node7473 : node7466;
												assign node7466 = (inp[7]) ? node7468 : 4'b0000;
													assign node7468 = (inp[4]) ? 4'b0000 : node7469;
														assign node7469 = (inp[2]) ? 4'b0111 : 4'b0100;
												assign node7473 = (inp[4]) ? 4'b0100 : node7474;
													assign node7474 = (inp[7]) ? 4'b0000 : 4'b0100;
								assign node7478 = (inp[11]) ? node7664 : node7479;
									assign node7479 = (inp[14]) ? node7575 : node7480;
										assign node7480 = (inp[3]) ? node7536 : node7481;
											assign node7481 = (inp[2]) ? node7515 : node7482;
												assign node7482 = (inp[7]) ? node7502 : node7483;
													assign node7483 = (inp[13]) ? node7495 : node7484;
														assign node7484 = (inp[4]) ? node7490 : node7485;
															assign node7485 = (inp[10]) ? 4'b1101 : node7486;
																assign node7486 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node7490 = (inp[10]) ? 4'b1001 : node7491;
																assign node7491 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node7495 = (inp[12]) ? node7497 : 4'b0001;
															assign node7497 = (inp[10]) ? 4'b0001 : node7498;
																assign node7498 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node7502 = (inp[13]) ? node7508 : node7503;
														assign node7503 = (inp[12]) ? node7505 : 4'b1101;
															assign node7505 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node7508 = (inp[12]) ? node7512 : node7509;
															assign node7509 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node7512 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node7515 = (inp[7]) ? node7527 : node7516;
													assign node7516 = (inp[4]) ? node7520 : node7517;
														assign node7517 = (inp[13]) ? 4'b0001 : 4'b0111;
														assign node7520 = (inp[13]) ? 4'b0001 : node7521;
															assign node7521 = (inp[10]) ? 4'b1001 : node7522;
																assign node7522 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7527 = (inp[4]) ? node7529 : 4'b0111;
														assign node7529 = (inp[13]) ? node7531 : 4'b0111;
															assign node7531 = (inp[12]) ? node7533 : 4'b0001;
																assign node7533 = (inp[10]) ? 4'b0001 : 4'b0111;
											assign node7536 = (inp[4]) ? node7552 : node7537;
												assign node7537 = (inp[13]) ? node7543 : node7538;
													assign node7538 = (inp[12]) ? node7540 : 4'b1001;
														assign node7540 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node7543 = (inp[10]) ? node7549 : node7544;
														assign node7544 = (inp[12]) ? 4'b1001 : node7545;
															assign node7545 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node7549 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7552 = (inp[7]) ? node7564 : node7553;
													assign node7553 = (inp[13]) ? node7559 : node7554;
														assign node7554 = (inp[10]) ? 4'b1101 : node7555;
															assign node7555 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node7559 = (inp[12]) ? node7561 : 4'b0101;
															assign node7561 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node7564 = (inp[13]) ? node7570 : node7565;
														assign node7565 = (inp[12]) ? node7567 : 4'b1001;
															assign node7567 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node7570 = (inp[12]) ? node7572 : 4'b0101;
															assign node7572 = (inp[10]) ? 4'b0101 : 4'b1001;
										assign node7575 = (inp[3]) ? node7629 : node7576;
											assign node7576 = (inp[2]) ? node7610 : node7577;
												assign node7577 = (inp[13]) ? node7595 : node7578;
													assign node7578 = (inp[10]) ? node7590 : node7579;
														assign node7579 = (inp[12]) ? node7585 : node7580;
															assign node7580 = (inp[4]) ? node7582 : 4'b1100;
																assign node7582 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node7585 = (inp[7]) ? 4'b0100 : node7586;
																assign node7586 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7590 = (inp[7]) ? 4'b1100 : node7591;
															assign node7591 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node7595 = (inp[10]) ? node7605 : node7596;
														assign node7596 = (inp[12]) ? node7600 : node7597;
															assign node7597 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node7600 = (inp[7]) ? 4'b1100 : node7601;
																assign node7601 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node7605 = (inp[7]) ? node7607 : 4'b0000;
															assign node7607 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node7610 = (inp[7]) ? node7620 : node7611;
													assign node7611 = (inp[4]) ? node7615 : node7612;
														assign node7612 = (inp[13]) ? 4'b0000 : 4'b0111;
														assign node7615 = (inp[13]) ? node7617 : 4'b1000;
															assign node7617 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node7620 = (inp[4]) ? node7622 : 4'b0111;
														assign node7622 = (inp[13]) ? node7624 : 4'b0111;
															assign node7624 = (inp[12]) ? node7626 : 4'b0000;
																assign node7626 = (inp[10]) ? 4'b0000 : 4'b0111;
											assign node7629 = (inp[13]) ? node7647 : node7630;
												assign node7630 = (inp[12]) ? node7636 : node7631;
													assign node7631 = (inp[4]) ? node7633 : 4'b1000;
														assign node7633 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node7636 = (inp[10]) ? node7642 : node7637;
														assign node7637 = (inp[4]) ? node7639 : 4'b0000;
															assign node7639 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7642 = (inp[4]) ? node7644 : 4'b1000;
															assign node7644 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node7647 = (inp[10]) ? node7659 : node7648;
													assign node7648 = (inp[12]) ? node7654 : node7649;
														assign node7649 = (inp[7]) ? node7651 : 4'b0100;
															assign node7651 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node7654 = (inp[4]) ? node7656 : 4'b1000;
															assign node7656 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node7659 = (inp[4]) ? 4'b0100 : node7660;
														assign node7660 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node7664 = (inp[13]) ? node7710 : node7665;
										assign node7665 = (inp[3]) ? node7693 : node7666;
											assign node7666 = (inp[2]) ? node7684 : node7667;
												assign node7667 = (inp[10]) ? node7679 : node7668;
													assign node7668 = (inp[12]) ? node7674 : node7669;
														assign node7669 = (inp[4]) ? node7671 : 4'b1101;
															assign node7671 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node7674 = (inp[7]) ? 4'b0101 : node7675;
															assign node7675 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node7679 = (inp[4]) ? node7681 : 4'b1101;
														assign node7681 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node7684 = (inp[7]) ? 4'b0111 : node7685;
													assign node7685 = (inp[4]) ? node7687 : 4'b0111;
														assign node7687 = (inp[12]) ? node7689 : 4'b1001;
															assign node7689 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node7693 = (inp[7]) ? node7705 : node7694;
												assign node7694 = (inp[4]) ? node7700 : node7695;
													assign node7695 = (inp[10]) ? 4'b1001 : node7696;
														assign node7696 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node7700 = (inp[10]) ? 4'b1101 : node7701;
														assign node7701 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node7705 = (inp[10]) ? 4'b1001 : node7706;
													assign node7706 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node7710 = (inp[10]) ? node7742 : node7711;
											assign node7711 = (inp[12]) ? node7725 : node7712;
												assign node7712 = (inp[3]) ? node7720 : node7713;
													assign node7713 = (inp[4]) ? 4'b0001 : node7714;
														assign node7714 = (inp[7]) ? node7716 : 4'b0001;
															assign node7716 = (inp[2]) ? 4'b0111 : 4'b0101;
													assign node7720 = (inp[4]) ? 4'b0101 : node7721;
														assign node7721 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node7725 = (inp[3]) ? node7737 : node7726;
													assign node7726 = (inp[2]) ? node7732 : node7727;
														assign node7727 = (inp[7]) ? 4'b1101 : node7728;
															assign node7728 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node7732 = (inp[7]) ? 4'b0111 : node7733;
															assign node7733 = (inp[4]) ? 4'b1001 : 4'b0111;
													assign node7737 = (inp[7]) ? 4'b1001 : node7738;
														assign node7738 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node7742 = (inp[3]) ? node7750 : node7743;
												assign node7743 = (inp[7]) ? node7745 : 4'b0001;
													assign node7745 = (inp[4]) ? 4'b0001 : node7746;
														assign node7746 = (inp[2]) ? 4'b0111 : 4'b0101;
												assign node7750 = (inp[7]) ? node7752 : 4'b0101;
													assign node7752 = (inp[4]) ? 4'b0101 : 4'b0001;
					assign node7756 = (inp[5]) ? node8946 : node7757;
						assign node7757 = (inp[0]) ? node8615 : node7758;
							assign node7758 = (inp[11]) ? node8272 : node7759;
								assign node7759 = (inp[3]) ? node8049 : node7760;
									assign node7760 = (inp[2]) ? node7858 : node7761;
										assign node7761 = (inp[10]) ? node7815 : node7762;
											assign node7762 = (inp[4]) ? node7798 : node7763;
												assign node7763 = (inp[13]) ? node7781 : node7764;
													assign node7764 = (inp[12]) ? node7774 : node7765;
														assign node7765 = (inp[7]) ? node7767 : 4'b0101;
															assign node7767 = (inp[14]) ? node7771 : node7768;
																assign node7768 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node7771 = (inp[1]) ? 4'b1100 : 4'b0101;
														assign node7774 = (inp[14]) ? node7778 : node7775;
															assign node7775 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node7778 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node7781 = (inp[7]) ? node7787 : node7782;
														assign node7782 = (inp[1]) ? 4'b1000 : node7783;
															assign node7783 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node7787 = (inp[12]) ? node7793 : node7788;
															assign node7788 = (inp[1]) ? node7790 : 4'b0100;
																assign node7790 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node7793 = (inp[14]) ? node7795 : 4'b1100;
																assign node7795 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node7798 = (inp[12]) ? node7804 : node7799;
													assign node7799 = (inp[7]) ? 4'b1000 : node7800;
														assign node7800 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node7804 = (inp[1]) ? node7810 : node7805;
														assign node7805 = (inp[7]) ? 4'b0000 : node7806;
															assign node7806 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node7810 = (inp[7]) ? 4'b1000 : node7811;
															assign node7811 = (inp[14]) ? 4'b1000 : 4'b1100;
											assign node7815 = (inp[4]) ? node7841 : node7816;
												assign node7816 = (inp[7]) ? node7826 : node7817;
													assign node7817 = (inp[12]) ? node7819 : 4'b0000;
														assign node7819 = (inp[1]) ? 4'b0000 : node7820;
															assign node7820 = (inp[13]) ? 4'b1000 : node7821;
																assign node7821 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node7826 = (inp[13]) ? node7834 : node7827;
														assign node7827 = (inp[14]) ? node7831 : node7828;
															assign node7828 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7831 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node7834 = (inp[1]) ? 4'b0000 : node7835;
															assign node7835 = (inp[12]) ? node7837 : 4'b0000;
																assign node7837 = (inp[14]) ? 4'b1101 : 4'b0100;
												assign node7841 = (inp[1]) ? node7853 : node7842;
													assign node7842 = (inp[12]) ? node7848 : node7843;
														assign node7843 = (inp[13]) ? 4'b0100 : node7844;
															assign node7844 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node7848 = (inp[13]) ? node7850 : 4'b1000;
															assign node7850 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node7853 = (inp[13]) ? 4'b0100 : node7854;
														assign node7854 = (inp[7]) ? 4'b0000 : 4'b0100;
										assign node7858 = (inp[7]) ? node7964 : node7859;
											assign node7859 = (inp[4]) ? node7909 : node7860;
												assign node7860 = (inp[13]) ? node7884 : node7861;
													assign node7861 = (inp[12]) ? node7871 : node7862;
														assign node7862 = (inp[14]) ? node7866 : node7863;
															assign node7863 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7866 = (inp[1]) ? 4'b1100 : node7867;
																assign node7867 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node7871 = (inp[10]) ? node7879 : node7872;
															assign node7872 = (inp[1]) ? node7876 : node7873;
																assign node7873 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node7876 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node7879 = (inp[1]) ? node7881 : 4'b0101;
																assign node7881 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7884 = (inp[12]) ? node7894 : node7885;
														assign node7885 = (inp[14]) ? node7889 : node7886;
															assign node7886 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node7889 = (inp[1]) ? 4'b0000 : node7890;
																assign node7890 = (inp[10]) ? 4'b0001 : 4'b1101;
														assign node7894 = (inp[10]) ? node7902 : node7895;
															assign node7895 = (inp[14]) ? node7899 : node7896;
																assign node7896 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node7899 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node7902 = (inp[1]) ? node7906 : node7903;
																assign node7903 = (inp[14]) ? 4'b1101 : 4'b0000;
																assign node7906 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node7909 = (inp[13]) ? node7941 : node7910;
													assign node7910 = (inp[12]) ? node7926 : node7911;
														assign node7911 = (inp[10]) ? node7919 : node7912;
															assign node7912 = (inp[1]) ? node7916 : node7913;
																assign node7913 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node7916 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node7919 = (inp[14]) ? node7923 : node7920;
																assign node7920 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node7923 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7926 = (inp[10]) ? node7934 : node7927;
															assign node7927 = (inp[14]) ? node7931 : node7928;
																assign node7928 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node7931 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node7934 = (inp[1]) ? node7938 : node7935;
																assign node7935 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node7938 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node7941 = (inp[12]) ? node7951 : node7942;
														assign node7942 = (inp[1]) ? node7948 : node7943;
															assign node7943 = (inp[14]) ? node7945 : 4'b0000;
																assign node7945 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node7948 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node7951 = (inp[10]) ? node7959 : node7952;
															assign node7952 = (inp[14]) ? node7956 : node7953;
																assign node7953 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node7956 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node7959 = (inp[14]) ? node7961 : 4'b0000;
																assign node7961 = (inp[1]) ? 4'b0000 : 4'b1001;
											assign node7964 = (inp[13]) ? node7990 : node7965;
												assign node7965 = (inp[12]) ? node7975 : node7966;
													assign node7966 = (inp[1]) ? node7972 : node7967;
														assign node7967 = (inp[14]) ? node7969 : 4'b1100;
															assign node7969 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node7972 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node7975 = (inp[10]) ? node7983 : node7976;
														assign node7976 = (inp[14]) ? node7980 : node7977;
															assign node7977 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node7980 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node7983 = (inp[14]) ? node7987 : node7984;
															assign node7984 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7987 = (inp[1]) ? 4'b1100 : 4'b0101;
												assign node7990 = (inp[4]) ? node8022 : node7991;
													assign node7991 = (inp[10]) ? node8007 : node7992;
														assign node7992 = (inp[12]) ? node8000 : node7993;
															assign node7993 = (inp[1]) ? node7997 : node7994;
																assign node7994 = (inp[14]) ? 4'b1101 : 4'b0100;
																assign node7997 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8000 = (inp[1]) ? node8004 : node8001;
																assign node8001 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node8004 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node8007 = (inp[12]) ? node8015 : node8008;
															assign node8008 = (inp[1]) ? node8012 : node8009;
																assign node8009 = (inp[14]) ? 4'b0101 : 4'b0100;
																assign node8012 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8015 = (inp[1]) ? node8019 : node8016;
																assign node8016 = (inp[14]) ? 4'b1101 : 4'b0100;
																assign node8019 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node8022 = (inp[10]) ? node8034 : node8023;
														assign node8023 = (inp[12]) ? node8029 : node8024;
															assign node8024 = (inp[14]) ? node8026 : 4'b0000;
																assign node8026 = (inp[1]) ? 4'b0000 : 4'b1101;
															assign node8029 = (inp[14]) ? node8031 : 4'b1100;
																assign node8031 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node8034 = (inp[12]) ? node8042 : node8035;
															assign node8035 = (inp[1]) ? node8039 : node8036;
																assign node8036 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node8039 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8042 = (inp[1]) ? node8046 : node8043;
																assign node8043 = (inp[14]) ? 4'b1101 : 4'b0000;
																assign node8046 = (inp[14]) ? 4'b0000 : 4'b0001;
									assign node8049 = (inp[10]) ? node8175 : node8050;
										assign node8050 = (inp[1]) ? node8116 : node8051;
											assign node8051 = (inp[12]) ? node8087 : node8052;
												assign node8052 = (inp[2]) ? node8070 : node8053;
													assign node8053 = (inp[4]) ? node8059 : node8054;
														assign node8054 = (inp[7]) ? 4'b1100 : node8055;
															assign node8055 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node8059 = (inp[13]) ? node8063 : node8060;
															assign node8060 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node8063 = (inp[7]) ? node8067 : node8064;
																assign node8064 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node8067 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node8070 = (inp[4]) ? node8082 : node8071;
														assign node8071 = (inp[14]) ? node8077 : node8072;
															assign node8072 = (inp[13]) ? node8074 : 4'b1000;
																assign node8074 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node8077 = (inp[13]) ? node8079 : 4'b0001;
																assign node8079 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node8082 = (inp[7]) ? 4'b1000 : node8083;
															assign node8083 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node8087 = (inp[13]) ? node8099 : node8088;
													assign node8088 = (inp[4]) ? node8092 : node8089;
														assign node8089 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node8092 = (inp[14]) ? 4'b0000 : node8093;
															assign node8093 = (inp[2]) ? 4'b0000 : node8094;
																assign node8094 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node8099 = (inp[4]) ? node8109 : node8100;
														assign node8100 = (inp[2]) ? node8104 : node8101;
															assign node8101 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node8104 = (inp[7]) ? node8106 : 4'b0000;
																assign node8106 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node8109 = (inp[2]) ? node8113 : node8110;
															assign node8110 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node8113 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node8116 = (inp[2]) ? node8146 : node8117;
												assign node8117 = (inp[4]) ? node8123 : node8118;
													assign node8118 = (inp[7]) ? 4'b1100 : node8119;
														assign node8119 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node8123 = (inp[14]) ? node8139 : node8124;
														assign node8124 = (inp[7]) ? node8132 : node8125;
															assign node8125 = (inp[13]) ? node8129 : node8126;
																assign node8126 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node8129 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node8132 = (inp[12]) ? node8136 : node8133;
																assign node8133 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node8136 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node8139 = (inp[13]) ? node8143 : node8140;
															assign node8140 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node8143 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node8146 = (inp[4]) ? node8170 : node8147;
													assign node8147 = (inp[14]) ? node8161 : node8148;
														assign node8148 = (inp[7]) ? node8154 : node8149;
															assign node8149 = (inp[13]) ? 4'b1000 : node8150;
																assign node8150 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8154 = (inp[12]) ? node8158 : node8155;
																assign node8155 = (inp[13]) ? 4'b0001 : 4'b1001;
																assign node8158 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node8161 = (inp[12]) ? node8167 : node8162;
															assign node8162 = (inp[7]) ? node8164 : 4'b1000;
																assign node8164 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node8167 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node8170 = (inp[13]) ? node8172 : 4'b1000;
														assign node8172 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node8175 = (inp[1]) ? node8239 : node8176;
											assign node8176 = (inp[12]) ? node8206 : node8177;
												assign node8177 = (inp[4]) ? node8191 : node8178;
													assign node8178 = (inp[2]) ? node8184 : node8179;
														assign node8179 = (inp[7]) ? node8181 : 4'b0000;
															assign node8181 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node8184 = (inp[13]) ? 4'b0000 : node8185;
															assign node8185 = (inp[7]) ? node8187 : 4'b0000;
																assign node8187 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node8191 = (inp[2]) ? node8201 : node8192;
														assign node8192 = (inp[13]) ? node8196 : node8193;
															assign node8193 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8196 = (inp[7]) ? node8198 : 4'b1101;
																assign node8198 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8201 = (inp[13]) ? 4'b0100 : node8202;
															assign node8202 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node8206 = (inp[2]) ? node8222 : node8207;
													assign node8207 = (inp[4]) ? node8213 : node8208;
														assign node8208 = (inp[7]) ? 4'b1100 : node8209;
															assign node8209 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node8213 = (inp[13]) ? node8217 : node8214;
															assign node8214 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node8217 = (inp[7]) ? 4'b1000 : node8218;
																assign node8218 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node8222 = (inp[4]) ? node8234 : node8223;
														assign node8223 = (inp[14]) ? node8229 : node8224;
															assign node8224 = (inp[7]) ? node8226 : 4'b1000;
																assign node8226 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node8229 = (inp[13]) ? node8231 : 4'b0001;
																assign node8231 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node8234 = (inp[13]) ? node8236 : 4'b1000;
															assign node8236 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node8239 = (inp[4]) ? node8253 : node8240;
												assign node8240 = (inp[7]) ? node8248 : node8241;
													assign node8241 = (inp[14]) ? node8243 : 4'b0000;
														assign node8243 = (inp[12]) ? 4'b0000 : node8244;
															assign node8244 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node8248 = (inp[13]) ? 4'b0000 : node8249;
														assign node8249 = (inp[2]) ? 4'b1001 : 4'b0100;
												assign node8253 = (inp[13]) ? node8263 : node8254;
													assign node8254 = (inp[2]) ? node8260 : node8255;
														assign node8255 = (inp[14]) ? node8257 : 4'b1000;
															assign node8257 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8260 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node8263 = (inp[14]) ? node8265 : 4'b0100;
														assign node8265 = (inp[2]) ? 4'b0100 : node8266;
															assign node8266 = (inp[12]) ? node8268 : 4'b0101;
																assign node8268 = (inp[7]) ? 4'b1001 : 4'b1101;
								assign node8272 = (inp[1]) ? node8486 : node8273;
									assign node8273 = (inp[3]) ? node8359 : node8274;
										assign node8274 = (inp[2]) ? node8328 : node8275;
											assign node8275 = (inp[4]) ? node8305 : node8276;
												assign node8276 = (inp[13]) ? node8290 : node8277;
													assign node8277 = (inp[7]) ? node8285 : node8278;
														assign node8278 = (inp[12]) ? node8282 : node8279;
															assign node8279 = (inp[10]) ? 4'b0001 : 4'b1100;
															assign node8282 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node8285 = (inp[10]) ? 4'b1100 : node8286;
															assign node8286 = (inp[14]) ? 4'b1100 : 4'b0100;
													assign node8290 = (inp[7]) ? node8298 : node8291;
														assign node8291 = (inp[14]) ? node8293 : 4'b1001;
															assign node8293 = (inp[10]) ? node8295 : 4'b1001;
																assign node8295 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8298 = (inp[10]) ? node8302 : node8299;
															assign node8299 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node8302 = (inp[12]) ? 4'b0100 : 4'b0001;
												assign node8305 = (inp[13]) ? node8313 : node8306;
													assign node8306 = (inp[12]) ? node8310 : node8307;
														assign node8307 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8310 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8313 = (inp[7]) ? node8321 : node8314;
														assign node8314 = (inp[10]) ? node8318 : node8315;
															assign node8315 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node8318 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node8321 = (inp[12]) ? node8325 : node8322;
															assign node8322 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node8325 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node8328 = (inp[13]) ? node8342 : node8329;
												assign node8329 = (inp[7]) ? node8337 : node8330;
													assign node8330 = (inp[4]) ? node8332 : 4'b1100;
														assign node8332 = (inp[10]) ? 4'b1000 : node8333;
															assign node8333 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8337 = (inp[12]) ? node8339 : 4'b1100;
														assign node8339 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node8342 = (inp[10]) ? node8354 : node8343;
													assign node8343 = (inp[12]) ? node8349 : node8344;
														assign node8344 = (inp[7]) ? node8346 : 4'b0000;
															assign node8346 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node8349 = (inp[7]) ? 4'b1100 : node8350;
															assign node8350 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node8354 = (inp[4]) ? 4'b0000 : node8355;
														assign node8355 = (inp[7]) ? 4'b0100 : 4'b0000;
										assign node8359 = (inp[2]) ? node8419 : node8360;
											assign node8360 = (inp[4]) ? node8394 : node8361;
												assign node8361 = (inp[13]) ? node8379 : node8362;
													assign node8362 = (inp[7]) ? node8370 : node8363;
														assign node8363 = (inp[10]) ? node8367 : node8364;
															assign node8364 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node8367 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node8370 = (inp[14]) ? 4'b1101 : node8371;
															assign node8371 = (inp[12]) ? node8375 : node8372;
																assign node8372 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node8375 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node8379 = (inp[7]) ? node8387 : node8380;
														assign node8380 = (inp[10]) ? node8384 : node8381;
															assign node8381 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8384 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node8387 = (inp[12]) ? node8391 : node8388;
															assign node8388 = (inp[10]) ? 4'b0001 : 4'b1101;
															assign node8391 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node8394 = (inp[13]) ? node8408 : node8395;
													assign node8395 = (inp[12]) ? node8401 : node8396;
														assign node8396 = (inp[10]) ? 4'b1000 : node8397;
															assign node8397 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node8401 = (inp[7]) ? node8405 : node8402;
															assign node8402 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8405 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node8408 = (inp[7]) ? node8414 : node8409;
														assign node8409 = (inp[10]) ? node8411 : 4'b0100;
															assign node8411 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node8414 = (inp[10]) ? node8416 : 4'b0000;
															assign node8416 = (inp[12]) ? 4'b1000 : 4'b0100;
											assign node8419 = (inp[4]) ? node8445 : node8420;
												assign node8420 = (inp[13]) ? node8430 : node8421;
													assign node8421 = (inp[12]) ? node8427 : node8422;
														assign node8422 = (inp[7]) ? 4'b1000 : node8423;
															assign node8423 = (inp[10]) ? 4'b0001 : 4'b1000;
														assign node8427 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node8430 = (inp[7]) ? node8438 : node8431;
														assign node8431 = (inp[12]) ? node8435 : node8432;
															assign node8432 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8435 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node8438 = (inp[12]) ? node8442 : node8439;
															assign node8439 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node8442 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node8445 = (inp[13]) ? node8465 : node8446;
													assign node8446 = (inp[7]) ? node8454 : node8447;
														assign node8447 = (inp[12]) ? node8451 : node8448;
															assign node8448 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node8451 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node8454 = (inp[14]) ? node8460 : node8455;
															assign node8455 = (inp[12]) ? 4'b1001 : node8456;
																assign node8456 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node8460 = (inp[10]) ? 4'b1001 : node8461;
																assign node8461 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node8465 = (inp[7]) ? node8479 : node8466;
														assign node8466 = (inp[14]) ? node8474 : node8467;
															assign node8467 = (inp[12]) ? node8471 : node8468;
																assign node8468 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node8471 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node8474 = (inp[12]) ? 4'b0101 : node8475;
																assign node8475 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node8479 = (inp[10]) ? node8483 : node8480;
															assign node8480 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8483 = (inp[12]) ? 4'b1001 : 4'b0101;
									assign node8486 = (inp[10]) ? node8576 : node8487;
										assign node8487 = (inp[4]) ? node8521 : node8488;
											assign node8488 = (inp[3]) ? node8506 : node8489;
												assign node8489 = (inp[7]) ? node8499 : node8490;
													assign node8490 = (inp[13]) ? node8494 : node8491;
														assign node8491 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node8494 = (inp[2]) ? node8496 : 4'b1001;
															assign node8496 = (inp[12]) ? 4'b1101 : 4'b0001;
													assign node8499 = (inp[12]) ? node8503 : node8500;
														assign node8500 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node8503 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node8506 = (inp[2]) ? node8512 : node8507;
													assign node8507 = (inp[13]) ? node8509 : 4'b1101;
														assign node8509 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node8512 = (inp[13]) ? node8516 : node8513;
														assign node8513 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8516 = (inp[12]) ? 4'b1001 : node8517;
															assign node8517 = (inp[7]) ? 4'b0001 : 4'b1001;
											assign node8521 = (inp[13]) ? node8553 : node8522;
												assign node8522 = (inp[7]) ? node8542 : node8523;
													assign node8523 = (inp[14]) ? node8535 : node8524;
														assign node8524 = (inp[3]) ? node8530 : node8525;
															assign node8525 = (inp[12]) ? node8527 : 4'b1001;
																assign node8527 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node8530 = (inp[2]) ? 4'b1001 : node8531;
																assign node8531 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8535 = (inp[3]) ? node8539 : node8536;
															assign node8536 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node8539 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node8542 = (inp[3]) ? node8548 : node8543;
														assign node8543 = (inp[2]) ? node8545 : 4'b1001;
															assign node8545 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node8548 = (inp[2]) ? 4'b1001 : node8549;
															assign node8549 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node8553 = (inp[7]) ? node8565 : node8554;
													assign node8554 = (inp[3]) ? node8560 : node8555;
														assign node8555 = (inp[2]) ? node8557 : 4'b1101;
															assign node8557 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8560 = (inp[2]) ? 4'b1101 : node8561;
															assign node8561 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node8565 = (inp[3]) ? node8571 : node8566;
														assign node8566 = (inp[2]) ? node8568 : 4'b1001;
															assign node8568 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node8571 = (inp[2]) ? 4'b1001 : node8572;
															assign node8572 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node8576 = (inp[13]) ? node8602 : node8577;
											assign node8577 = (inp[3]) ? node8591 : node8578;
												assign node8578 = (inp[2]) ? node8586 : node8579;
													assign node8579 = (inp[4]) ? node8583 : node8580;
														assign node8580 = (inp[7]) ? 4'b1101 : 4'b0001;
														assign node8583 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node8586 = (inp[7]) ? 4'b1101 : node8587;
														assign node8587 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node8591 = (inp[4]) ? node8597 : node8592;
													assign node8592 = (inp[7]) ? node8594 : 4'b0001;
														assign node8594 = (inp[2]) ? 4'b1001 : 4'b0101;
													assign node8597 = (inp[2]) ? node8599 : 4'b1001;
														assign node8599 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node8602 = (inp[4]) ? node8610 : node8603;
												assign node8603 = (inp[2]) ? node8605 : 4'b0001;
													assign node8605 = (inp[7]) ? node8607 : 4'b0001;
														assign node8607 = (inp[3]) ? 4'b0001 : 4'b0101;
												assign node8610 = (inp[3]) ? 4'b0101 : node8611;
													assign node8611 = (inp[2]) ? 4'b0001 : 4'b0101;
							assign node8615 = (inp[2]) ? 4'b0101 : node8616;
								assign node8616 = (inp[3]) ? node8734 : node8617;
									assign node8617 = (inp[4]) ? node8647 : node8618;
										assign node8618 = (inp[13]) ? node8620 : 4'b0101;
											assign node8620 = (inp[7]) ? 4'b0101 : node8621;
												assign node8621 = (inp[12]) ? node8633 : node8622;
													assign node8622 = (inp[1]) ? node8628 : node8623;
														assign node8623 = (inp[11]) ? 4'b0000 : node8624;
															assign node8624 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node8628 = (inp[14]) ? node8630 : 4'b0001;
															assign node8630 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node8633 = (inp[10]) ? node8635 : 4'b0101;
														assign node8635 = (inp[1]) ? node8641 : node8636;
															assign node8636 = (inp[11]) ? 4'b0000 : node8637;
																assign node8637 = (inp[14]) ? 4'b0101 : 4'b0000;
															assign node8641 = (inp[11]) ? 4'b0001 : node8642;
																assign node8642 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node8647 = (inp[7]) ? node8707 : node8648;
											assign node8648 = (inp[1]) ? node8678 : node8649;
												assign node8649 = (inp[14]) ? node8661 : node8650;
													assign node8650 = (inp[13]) ? node8656 : node8651;
														assign node8651 = (inp[12]) ? node8653 : 4'b1000;
															assign node8653 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node8656 = (inp[10]) ? 4'b0000 : node8657;
															assign node8657 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node8661 = (inp[11]) ? node8669 : node8662;
														assign node8662 = (inp[13]) ? node8664 : 4'b0001;
															assign node8664 = (inp[10]) ? node8666 : 4'b1001;
																assign node8666 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node8669 = (inp[13]) ? node8673 : node8670;
															assign node8670 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node8673 = (inp[10]) ? 4'b0000 : node8674;
																assign node8674 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node8678 = (inp[13]) ? node8690 : node8679;
													assign node8679 = (inp[12]) ? node8685 : node8680;
														assign node8680 = (inp[11]) ? 4'b1001 : node8681;
															assign node8681 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8685 = (inp[10]) ? 4'b1001 : node8686;
															assign node8686 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node8690 = (inp[14]) ? node8696 : node8691;
														assign node8691 = (inp[12]) ? node8693 : 4'b0001;
															assign node8693 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node8696 = (inp[11]) ? node8702 : node8697;
															assign node8697 = (inp[12]) ? node8699 : 4'b0000;
																assign node8699 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node8702 = (inp[12]) ? node8704 : 4'b0001;
																assign node8704 = (inp[10]) ? 4'b0001 : 4'b1001;
											assign node8707 = (inp[13]) ? node8709 : 4'b0101;
												assign node8709 = (inp[12]) ? node8721 : node8710;
													assign node8710 = (inp[1]) ? node8716 : node8711;
														assign node8711 = (inp[14]) ? node8713 : 4'b0000;
															assign node8713 = (inp[11]) ? 4'b0000 : 4'b0101;
														assign node8716 = (inp[14]) ? node8718 : 4'b0001;
															assign node8718 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node8721 = (inp[10]) ? node8723 : 4'b0101;
														assign node8723 = (inp[1]) ? node8729 : node8724;
															assign node8724 = (inp[14]) ? node8726 : 4'b0000;
																assign node8726 = (inp[11]) ? 4'b0000 : 4'b0101;
															assign node8729 = (inp[14]) ? node8731 : 4'b0001;
																assign node8731 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node8734 = (inp[4]) ? node8824 : node8735;
										assign node8735 = (inp[1]) ? node8779 : node8736;
											assign node8736 = (inp[11]) ? node8764 : node8737;
												assign node8737 = (inp[14]) ? node8751 : node8738;
													assign node8738 = (inp[13]) ? node8744 : node8739;
														assign node8739 = (inp[10]) ? 4'b1000 : node8740;
															assign node8740 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8744 = (inp[7]) ? node8746 : 4'b0100;
															assign node8746 = (inp[12]) ? node8748 : 4'b0000;
																assign node8748 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node8751 = (inp[13]) ? node8757 : node8752;
														assign node8752 = (inp[10]) ? node8754 : 4'b0001;
															assign node8754 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8757 = (inp[10]) ? node8759 : 4'b1001;
															assign node8759 = (inp[7]) ? node8761 : 4'b0101;
																assign node8761 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node8764 = (inp[13]) ? node8770 : node8765;
													assign node8765 = (inp[10]) ? 4'b1000 : node8766;
														assign node8766 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node8770 = (inp[10]) ? node8776 : node8771;
														assign node8771 = (inp[12]) ? 4'b1000 : node8772;
															assign node8772 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node8776 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node8779 = (inp[13]) ? node8797 : node8780;
												assign node8780 = (inp[12]) ? node8786 : node8781;
													assign node8781 = (inp[14]) ? node8783 : 4'b1001;
														assign node8783 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node8786 = (inp[10]) ? node8792 : node8787;
														assign node8787 = (inp[11]) ? 4'b0001 : node8788;
															assign node8788 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8792 = (inp[11]) ? 4'b1001 : node8793;
															assign node8793 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node8797 = (inp[7]) ? node8811 : node8798;
													assign node8798 = (inp[10]) ? node8806 : node8799;
														assign node8799 = (inp[12]) ? node8803 : node8800;
															assign node8800 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8803 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node8806 = (inp[11]) ? 4'b0101 : node8807;
															assign node8807 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node8811 = (inp[12]) ? node8817 : node8812;
														assign node8812 = (inp[11]) ? 4'b0001 : node8813;
															assign node8813 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node8817 = (inp[10]) ? 4'b0001 : node8818;
															assign node8818 = (inp[11]) ? 4'b1001 : node8819;
																assign node8819 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node8824 = (inp[7]) ? node8880 : node8825;
											assign node8825 = (inp[1]) ? node8853 : node8826;
												assign node8826 = (inp[11]) ? node8842 : node8827;
													assign node8827 = (inp[14]) ? node8835 : node8828;
														assign node8828 = (inp[13]) ? 4'b0100 : node8829;
															assign node8829 = (inp[12]) ? node8831 : 4'b1100;
																assign node8831 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node8835 = (inp[13]) ? node8837 : 4'b0101;
															assign node8837 = (inp[10]) ? node8839 : 4'b1101;
																assign node8839 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node8842 = (inp[13]) ? node8848 : node8843;
														assign node8843 = (inp[12]) ? node8845 : 4'b1100;
															assign node8845 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node8848 = (inp[12]) ? node8850 : 4'b0100;
															assign node8850 = (inp[10]) ? 4'b0100 : 4'b1100;
												assign node8853 = (inp[13]) ? node8869 : node8854;
													assign node8854 = (inp[11]) ? node8864 : node8855;
														assign node8855 = (inp[14]) ? node8859 : node8856;
															assign node8856 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node8859 = (inp[12]) ? node8861 : 4'b1100;
																assign node8861 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node8864 = (inp[12]) ? node8866 : 4'b1101;
															assign node8866 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node8869 = (inp[14]) ? node8875 : node8870;
														assign node8870 = (inp[12]) ? node8872 : 4'b0101;
															assign node8872 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node8875 = (inp[11]) ? 4'b0101 : node8876;
															assign node8876 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node8880 = (inp[13]) ? node8910 : node8881;
												assign node8881 = (inp[1]) ? node8895 : node8882;
													assign node8882 = (inp[14]) ? node8888 : node8883;
														assign node8883 = (inp[10]) ? 4'b1000 : node8884;
															assign node8884 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node8888 = (inp[11]) ? 4'b1000 : node8889;
															assign node8889 = (inp[12]) ? 4'b0001 : node8890;
																assign node8890 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node8895 = (inp[14]) ? node8901 : node8896;
														assign node8896 = (inp[10]) ? 4'b1001 : node8897;
															assign node8897 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8901 = (inp[11]) ? node8907 : node8902;
															assign node8902 = (inp[12]) ? node8904 : 4'b1000;
																assign node8904 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node8907 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node8910 = (inp[12]) ? node8924 : node8911;
													assign node8911 = (inp[1]) ? node8919 : node8912;
														assign node8912 = (inp[14]) ? node8914 : 4'b0100;
															assign node8914 = (inp[11]) ? 4'b0100 : node8915;
																assign node8915 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node8919 = (inp[14]) ? node8921 : 4'b0101;
															assign node8921 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node8924 = (inp[10]) ? node8936 : node8925;
														assign node8925 = (inp[1]) ? node8931 : node8926;
															assign node8926 = (inp[14]) ? node8928 : 4'b1000;
																assign node8928 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node8931 = (inp[14]) ? node8933 : 4'b1001;
																assign node8933 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node8936 = (inp[1]) ? node8940 : node8937;
															assign node8937 = (inp[11]) ? 4'b0100 : 4'b1001;
															assign node8940 = (inp[14]) ? node8942 : 4'b0101;
																assign node8942 = (inp[11]) ? 4'b0101 : 4'b0100;
						assign node8946 = (inp[3]) ? node9774 : node8947;
							assign node8947 = (inp[4]) ? node9353 : node8948;
								assign node8948 = (inp[13]) ? node9148 : node8949;
									assign node8949 = (inp[7]) ? node9053 : node8950;
										assign node8950 = (inp[0]) ? node9016 : node8951;
											assign node8951 = (inp[10]) ? node8989 : node8952;
												assign node8952 = (inp[1]) ? node8972 : node8953;
													assign node8953 = (inp[12]) ? node8963 : node8954;
														assign node8954 = (inp[14]) ? 4'b1100 : node8955;
															assign node8955 = (inp[11]) ? node8959 : node8956;
																assign node8956 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node8959 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node8963 = (inp[2]) ? node8969 : node8964;
															assign node8964 = (inp[11]) ? 4'b1100 : node8965;
																assign node8965 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node8969 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node8972 = (inp[11]) ? node8984 : node8973;
														assign node8973 = (inp[12]) ? node8979 : node8974;
															assign node8974 = (inp[2]) ? node8976 : 4'b0001;
																assign node8976 = (inp[14]) ? 4'b1100 : 4'b0000;
															assign node8979 = (inp[2]) ? 4'b1100 : node8980;
																assign node8980 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node8984 = (inp[12]) ? node8986 : 4'b0001;
															assign node8986 = (inp[2]) ? 4'b1101 : 4'b0001;
												assign node8989 = (inp[2]) ? node9001 : node8990;
													assign node8990 = (inp[1]) ? node8996 : node8991;
														assign node8991 = (inp[11]) ? 4'b1001 : node8992;
															assign node8992 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node8996 = (inp[12]) ? node8998 : 4'b0001;
															assign node8998 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node9001 = (inp[1]) ? node9011 : node9002;
														assign node9002 = (inp[14]) ? node9006 : node9003;
															assign node9003 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node9006 = (inp[12]) ? 4'b0000 : node9007;
																assign node9007 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node9011 = (inp[11]) ? 4'b1001 : node9012;
															assign node9012 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node9016 = (inp[2]) ? 4'b0101 : node9017;
												assign node9017 = (inp[10]) ? node9039 : node9018;
													assign node9018 = (inp[12]) ? node9028 : node9019;
														assign node9019 = (inp[1]) ? node9023 : node9020;
															assign node9020 = (inp[11]) ? 4'b1100 : 4'b0101;
															assign node9023 = (inp[11]) ? 4'b1101 : node9024;
																assign node9024 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node9028 = (inp[1]) ? node9034 : node9029;
															assign node9029 = (inp[14]) ? node9031 : 4'b0100;
																assign node9031 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node9034 = (inp[14]) ? node9036 : 4'b0101;
																assign node9036 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node9039 = (inp[1]) ? node9049 : node9040;
														assign node9040 = (inp[12]) ? node9044 : node9041;
															assign node9041 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node9044 = (inp[14]) ? node9046 : 4'b1100;
																assign node9046 = (inp[11]) ? 4'b1100 : 4'b0101;
														assign node9049 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node9053 = (inp[2]) ? node9127 : node9054;
											assign node9054 = (inp[1]) ? node9094 : node9055;
												assign node9055 = (inp[11]) ? node9085 : node9056;
													assign node9056 = (inp[12]) ? node9072 : node9057;
														assign node9057 = (inp[10]) ? node9065 : node9058;
															assign node9058 = (inp[0]) ? node9062 : node9059;
																assign node9059 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node9062 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node9065 = (inp[0]) ? node9069 : node9066;
																assign node9066 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node9069 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node9072 = (inp[10]) ? node9078 : node9073;
															assign node9073 = (inp[14]) ? 4'b0101 : node9074;
																assign node9074 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node9078 = (inp[0]) ? node9082 : node9079;
																assign node9079 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node9082 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node9085 = (inp[12]) ? node9087 : 4'b1100;
														assign node9087 = (inp[10]) ? node9091 : node9088;
															assign node9088 = (inp[0]) ? 4'b0100 : 4'b1100;
															assign node9091 = (inp[0]) ? 4'b1100 : 4'b0100;
												assign node9094 = (inp[11]) ? node9116 : node9095;
													assign node9095 = (inp[0]) ? node9105 : node9096;
														assign node9096 = (inp[14]) ? node9100 : node9097;
															assign node9097 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node9100 = (inp[10]) ? node9102 : 4'b1101;
																assign node9102 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node9105 = (inp[14]) ? node9111 : node9106;
															assign node9106 = (inp[12]) ? node9108 : 4'b1101;
																assign node9108 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node9111 = (inp[10]) ? 4'b1100 : node9112;
																assign node9112 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node9116 = (inp[10]) ? node9124 : node9117;
														assign node9117 = (inp[0]) ? node9121 : node9118;
															assign node9118 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node9121 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node9124 = (inp[0]) ? 4'b1101 : 4'b0001;
											assign node9127 = (inp[0]) ? 4'b0101 : node9128;
												assign node9128 = (inp[11]) ? node9140 : node9129;
													assign node9129 = (inp[10]) ? node9135 : node9130;
														assign node9130 = (inp[1]) ? 4'b1100 : node9131;
															assign node9131 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node9135 = (inp[1]) ? 4'b0100 : node9136;
															assign node9136 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node9140 = (inp[10]) ? 4'b0101 : node9141;
														assign node9141 = (inp[12]) ? node9143 : 4'b1101;
															assign node9143 = (inp[1]) ? 4'b1101 : 4'b0101;
									assign node9148 = (inp[0]) ? node9268 : node9149;
										assign node9149 = (inp[2]) ? node9209 : node9150;
											assign node9150 = (inp[1]) ? node9168 : node9151;
												assign node9151 = (inp[7]) ? node9163 : node9152;
													assign node9152 = (inp[10]) ? node9158 : node9153;
														assign node9153 = (inp[12]) ? node9155 : 4'b1001;
															assign node9155 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node9158 = (inp[12]) ? node9160 : 4'b1101;
															assign node9160 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node9163 = (inp[11]) ? 4'b1001 : node9164;
														assign node9164 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9168 = (inp[12]) ? node9194 : node9169;
													assign node9169 = (inp[14]) ? node9185 : node9170;
														assign node9170 = (inp[11]) ? node9178 : node9171;
															assign node9171 = (inp[7]) ? node9175 : node9172;
																assign node9172 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node9175 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node9178 = (inp[10]) ? node9182 : node9179;
																assign node9179 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node9182 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node9185 = (inp[10]) ? node9189 : node9186;
															assign node9186 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node9189 = (inp[7]) ? 4'b0101 : node9190;
																assign node9190 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node9194 = (inp[11]) ? node9200 : node9195;
														assign node9195 = (inp[10]) ? node9197 : 4'b1001;
															assign node9197 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node9200 = (inp[14]) ? node9204 : node9201;
															assign node9201 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node9204 = (inp[10]) ? node9206 : 4'b0101;
																assign node9206 = (inp[7]) ? 4'b0101 : 4'b0001;
											assign node9209 = (inp[1]) ? node9229 : node9210;
												assign node9210 = (inp[10]) ? node9220 : node9211;
													assign node9211 = (inp[11]) ? 4'b0000 : node9212;
														assign node9212 = (inp[12]) ? node9216 : node9213;
															assign node9213 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9216 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node9220 = (inp[11]) ? node9224 : node9221;
														assign node9221 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9224 = (inp[12]) ? 4'b1000 : node9225;
															assign node9225 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9229 = (inp[7]) ? node9247 : node9230;
													assign node9230 = (inp[10]) ? node9240 : node9231;
														assign node9231 = (inp[12]) ? node9235 : node9232;
															assign node9232 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node9235 = (inp[14]) ? 4'b0001 : node9236;
																assign node9236 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node9240 = (inp[11]) ? 4'b0101 : node9241;
															assign node9241 = (inp[14]) ? node9243 : 4'b0100;
																assign node9243 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node9247 = (inp[14]) ? node9257 : node9248;
														assign node9248 = (inp[11]) ? node9252 : node9249;
															assign node9249 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node9252 = (inp[10]) ? 4'b0001 : node9253;
																assign node9253 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9257 = (inp[11]) ? node9263 : node9258;
															assign node9258 = (inp[12]) ? node9260 : 4'b0001;
																assign node9260 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node9263 = (inp[12]) ? 4'b0001 : node9264;
																assign node9264 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node9268 = (inp[7]) ? node9318 : node9269;
											assign node9269 = (inp[2]) ? node9293 : node9270;
												assign node9270 = (inp[11]) ? node9282 : node9271;
													assign node9271 = (inp[10]) ? node9277 : node9272;
														assign node9272 = (inp[12]) ? node9274 : 4'b1000;
															assign node9274 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node9277 = (inp[12]) ? node9279 : 4'b0000;
															assign node9279 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node9282 = (inp[10]) ? node9288 : node9283;
														assign node9283 = (inp[1]) ? 4'b1001 : node9284;
															assign node9284 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9288 = (inp[12]) ? node9290 : 4'b0001;
															assign node9290 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node9293 = (inp[12]) ? node9307 : node9294;
													assign node9294 = (inp[1]) ? node9302 : node9295;
														assign node9295 = (inp[11]) ? 4'b0000 : node9296;
															assign node9296 = (inp[14]) ? node9298 : 4'b0000;
																assign node9298 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node9302 = (inp[11]) ? 4'b0001 : node9303;
															assign node9303 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node9307 = (inp[10]) ? node9309 : 4'b0101;
														assign node9309 = (inp[1]) ? node9313 : node9310;
															assign node9310 = (inp[11]) ? 4'b0000 : 4'b0101;
															assign node9313 = (inp[11]) ? 4'b0001 : node9314;
																assign node9314 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node9318 = (inp[2]) ? 4'b0101 : node9319;
												assign node9319 = (inp[10]) ? node9339 : node9320;
													assign node9320 = (inp[12]) ? node9330 : node9321;
														assign node9321 = (inp[14]) ? node9325 : node9322;
															assign node9322 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node9325 = (inp[11]) ? 4'b0100 : node9326;
																assign node9326 = (inp[1]) ? 4'b0100 : 4'b1101;
														assign node9330 = (inp[1]) ? node9336 : node9331;
															assign node9331 = (inp[11]) ? 4'b1100 : node9332;
																assign node9332 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node9336 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9339 = (inp[11]) ? node9347 : node9340;
														assign node9340 = (inp[12]) ? node9342 : 4'b0000;
															assign node9342 = (inp[1]) ? 4'b0000 : node9343;
																assign node9343 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node9347 = (inp[1]) ? 4'b0001 : node9348;
															assign node9348 = (inp[12]) ? 4'b0100 : 4'b0001;
								assign node9353 = (inp[1]) ? node9583 : node9354;
									assign node9354 = (inp[7]) ? node9498 : node9355;
										assign node9355 = (inp[0]) ? node9427 : node9356;
											assign node9356 = (inp[2]) ? node9396 : node9357;
												assign node9357 = (inp[10]) ? node9377 : node9358;
													assign node9358 = (inp[12]) ? node9368 : node9359;
														assign node9359 = (inp[11]) ? node9365 : node9360;
															assign node9360 = (inp[14]) ? node9362 : 4'b1000;
																assign node9362 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node9365 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node9368 = (inp[13]) ? node9374 : node9369;
															assign node9369 = (inp[14]) ? node9371 : 4'b1000;
																assign node9371 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node9374 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node9377 = (inp[13]) ? node9385 : node9378;
														assign node9378 = (inp[11]) ? 4'b0100 : node9379;
															assign node9379 = (inp[14]) ? 4'b1001 : node9380;
																assign node9380 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node9385 = (inp[14]) ? node9389 : node9386;
															assign node9386 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node9389 = (inp[12]) ? node9393 : node9390;
																assign node9390 = (inp[11]) ? 4'b1000 : 4'b0000;
																assign node9393 = (inp[11]) ? 4'b0000 : 4'b0100;
												assign node9396 = (inp[11]) ? node9420 : node9397;
													assign node9397 = (inp[12]) ? node9409 : node9398;
														assign node9398 = (inp[10]) ? node9402 : node9399;
															assign node9399 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node9402 = (inp[14]) ? node9406 : node9403;
																assign node9403 = (inp[13]) ? 4'b1000 : 4'b1001;
																assign node9406 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node9409 = (inp[13]) ? node9415 : node9410;
															assign node9410 = (inp[10]) ? 4'b0001 : node9411;
																assign node9411 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node9415 = (inp[14]) ? 4'b0001 : node9416;
																assign node9416 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node9420 = (inp[13]) ? node9424 : node9421;
														assign node9421 = (inp[10]) ? 4'b1001 : 4'b1100;
														assign node9424 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node9427 = (inp[13]) ? node9469 : node9428;
												assign node9428 = (inp[14]) ? node9442 : node9429;
													assign node9429 = (inp[2]) ? node9437 : node9430;
														assign node9430 = (inp[11]) ? 4'b1001 : node9431;
															assign node9431 = (inp[10]) ? 4'b0100 : node9432;
																assign node9432 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9437 = (inp[10]) ? 4'b1000 : node9438;
															assign node9438 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node9442 = (inp[12]) ? node9454 : node9443;
														assign node9443 = (inp[2]) ? node9449 : node9444;
															assign node9444 = (inp[10]) ? 4'b0101 : node9445;
																assign node9445 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node9449 = (inp[11]) ? 4'b1000 : node9450;
																assign node9450 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9454 = (inp[10]) ? node9462 : node9455;
															assign node9455 = (inp[11]) ? node9459 : node9456;
																assign node9456 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node9459 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node9462 = (inp[11]) ? node9466 : node9463;
																assign node9463 = (inp[2]) ? 4'b0001 : 4'b1000;
																assign node9466 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node9469 = (inp[11]) ? node9489 : node9470;
													assign node9470 = (inp[10]) ? node9482 : node9471;
														assign node9471 = (inp[2]) ? node9477 : node9472;
															assign node9472 = (inp[12]) ? 4'b0100 : node9473;
																assign node9473 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9477 = (inp[14]) ? 4'b1001 : node9478;
																assign node9478 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node9482 = (inp[2]) ? node9486 : node9483;
															assign node9483 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9486 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node9489 = (inp[12]) ? node9491 : 4'b0000;
														assign node9491 = (inp[10]) ? node9495 : node9492;
															assign node9492 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node9495 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node9498 = (inp[2]) ? node9546 : node9499;
											assign node9499 = (inp[11]) ? node9523 : node9500;
												assign node9500 = (inp[0]) ? node9514 : node9501;
													assign node9501 = (inp[10]) ? node9509 : node9502;
														assign node9502 = (inp[13]) ? node9506 : node9503;
															assign node9503 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node9506 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node9509 = (inp[13]) ? 4'b0000 : node9510;
															assign node9510 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node9514 = (inp[10]) ? node9518 : node9515;
														assign node9515 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9518 = (inp[12]) ? 4'b1000 : node9519;
															assign node9519 = (inp[14]) ? 4'b0000 : 4'b0100;
												assign node9523 = (inp[0]) ? node9537 : node9524;
													assign node9524 = (inp[12]) ? node9530 : node9525;
														assign node9525 = (inp[13]) ? node9527 : 4'b0000;
															assign node9527 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9530 = (inp[10]) ? node9534 : node9531;
															assign node9531 = (inp[13]) ? 4'b0100 : 4'b1101;
															assign node9534 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node9537 = (inp[10]) ? node9541 : node9538;
														assign node9538 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node9541 = (inp[12]) ? 4'b1001 : node9542;
															assign node9542 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node9546 = (inp[0]) ? node9568 : node9547;
												assign node9547 = (inp[13]) ? node9563 : node9548;
													assign node9548 = (inp[10]) ? node9556 : node9549;
														assign node9549 = (inp[11]) ? 4'b1000 : node9550;
															assign node9550 = (inp[12]) ? node9552 : 4'b1001;
																assign node9552 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9556 = (inp[11]) ? node9560 : node9557;
															assign node9557 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node9560 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node9563 = (inp[11]) ? 4'b1001 : node9564;
														assign node9564 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9568 = (inp[13]) ? node9570 : 4'b0101;
													assign node9570 = (inp[10]) ? node9578 : node9571;
														assign node9571 = (inp[12]) ? 4'b0101 : node9572;
															assign node9572 = (inp[14]) ? node9574 : 4'b0000;
																assign node9574 = (inp[11]) ? 4'b0000 : 4'b0101;
														assign node9578 = (inp[11]) ? 4'b0000 : node9579;
															assign node9579 = (inp[14]) ? 4'b0101 : 4'b0000;
									assign node9583 = (inp[11]) ? node9707 : node9584;
										assign node9584 = (inp[2]) ? node9642 : node9585;
											assign node9585 = (inp[10]) ? node9603 : node9586;
												assign node9586 = (inp[0]) ? node9594 : node9587;
													assign node9587 = (inp[13]) ? node9591 : node9588;
														assign node9588 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node9591 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node9594 = (inp[13]) ? node9596 : 4'b1000;
														assign node9596 = (inp[7]) ? 4'b1000 : node9597;
															assign node9597 = (inp[14]) ? 4'b0001 : node9598;
																assign node9598 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node9603 = (inp[0]) ? node9629 : node9604;
													assign node9604 = (inp[13]) ? node9620 : node9605;
														assign node9605 = (inp[14]) ? node9613 : node9606;
															assign node9606 = (inp[12]) ? node9610 : node9607;
																assign node9607 = (inp[7]) ? 4'b1001 : 4'b0000;
																assign node9610 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node9613 = (inp[7]) ? node9617 : node9614;
																assign node9614 = (inp[12]) ? 4'b0100 : 4'b0000;
																assign node9617 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node9620 = (inp[12]) ? node9626 : node9621;
															assign node9621 = (inp[14]) ? node9623 : 4'b0000;
																assign node9623 = (inp[7]) ? 4'b0100 : 4'b1001;
															assign node9626 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node9629 = (inp[13]) ? node9633 : node9630;
														assign node9630 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9633 = (inp[14]) ? node9635 : 4'b0000;
															assign node9635 = (inp[7]) ? node9639 : node9636;
																assign node9636 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node9639 = (inp[12]) ? 4'b0100 : 4'b0001;
											assign node9642 = (inp[12]) ? node9674 : node9643;
												assign node9643 = (inp[14]) ? node9659 : node9644;
													assign node9644 = (inp[10]) ? 4'b0001 : node9645;
														assign node9645 = (inp[7]) ? node9653 : node9646;
															assign node9646 = (inp[13]) ? node9650 : node9647;
																assign node9647 = (inp[0]) ? 4'b1001 : 4'b0001;
																assign node9650 = (inp[0]) ? 4'b0001 : 4'b0101;
															assign node9653 = (inp[13]) ? 4'b0001 : node9654;
																assign node9654 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node9659 = (inp[13]) ? node9667 : node9660;
														assign node9660 = (inp[0]) ? node9664 : node9661;
															assign node9661 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node9664 = (inp[7]) ? 4'b0101 : 4'b1000;
														assign node9667 = (inp[0]) ? 4'b0000 : node9668;
															assign node9668 = (inp[10]) ? 4'b0000 : node9669;
																assign node9669 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node9674 = (inp[0]) ? node9686 : node9675;
													assign node9675 = (inp[13]) ? 4'b1001 : node9676;
														assign node9676 = (inp[7]) ? node9682 : node9677;
															assign node9677 = (inp[10]) ? 4'b1001 : node9678;
																assign node9678 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node9682 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node9686 = (inp[7]) ? node9700 : node9687;
														assign node9687 = (inp[14]) ? node9693 : node9688;
															assign node9688 = (inp[10]) ? node9690 : 4'b0001;
																assign node9690 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node9693 = (inp[13]) ? node9697 : node9694;
																assign node9694 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node9697 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node9700 = (inp[10]) ? node9702 : 4'b0101;
															assign node9702 = (inp[13]) ? node9704 : 4'b0101;
																assign node9704 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node9707 = (inp[10]) ? node9759 : node9708;
											assign node9708 = (inp[2]) ? node9732 : node9709;
												assign node9709 = (inp[12]) ? node9711 : 4'b1001;
													assign node9711 = (inp[7]) ? node9727 : node9712;
														assign node9712 = (inp[14]) ? node9720 : node9713;
															assign node9713 = (inp[0]) ? node9717 : node9714;
																assign node9714 = (inp[13]) ? 4'b1001 : 4'b0001;
																assign node9717 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node9720 = (inp[13]) ? node9724 : node9721;
																assign node9721 = (inp[0]) ? 4'b1001 : 4'b0001;
																assign node9724 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node9727 = (inp[0]) ? 4'b1001 : node9728;
															assign node9728 = (inp[13]) ? 4'b1001 : 4'b0001;
												assign node9732 = (inp[7]) ? node9746 : node9733;
													assign node9733 = (inp[0]) ? node9739 : node9734;
														assign node9734 = (inp[12]) ? node9736 : 4'b0001;
															assign node9736 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node9739 = (inp[13]) ? node9743 : node9740;
															assign node9740 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node9743 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node9746 = (inp[0]) ? node9754 : node9747;
														assign node9747 = (inp[12]) ? node9751 : node9748;
															assign node9748 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node9751 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node9754 = (inp[13]) ? node9756 : 4'b0101;
															assign node9756 = (inp[12]) ? 4'b0101 : 4'b0001;
											assign node9759 = (inp[13]) ? 4'b0001 : node9760;
												assign node9760 = (inp[0]) ? node9766 : node9761;
													assign node9761 = (inp[2]) ? 4'b0001 : node9762;
														assign node9762 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node9766 = (inp[2]) ? node9770 : node9767;
														assign node9767 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node9770 = (inp[7]) ? 4'b0101 : 4'b1001;
							assign node9774 = (inp[4]) ? node10242 : node9775;
								assign node9775 = (inp[1]) ? node10041 : node9776;
									assign node9776 = (inp[11]) ? node9950 : node9777;
										assign node9777 = (inp[12]) ? node9863 : node9778;
											assign node9778 = (inp[13]) ? node9822 : node9779;
												assign node9779 = (inp[10]) ? node9801 : node9780;
													assign node9780 = (inp[0]) ? node9794 : node9781;
														assign node9781 = (inp[7]) ? node9789 : node9782;
															assign node9782 = (inp[14]) ? node9786 : node9783;
																assign node9783 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node9786 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node9789 = (inp[14]) ? node9791 : 4'b1000;
																assign node9791 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node9794 = (inp[2]) ? node9798 : node9795;
															assign node9795 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9798 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node9801 = (inp[2]) ? node9817 : node9802;
														assign node9802 = (inp[14]) ? node9810 : node9803;
															assign node9803 = (inp[0]) ? node9807 : node9804;
																assign node9804 = (inp[7]) ? 4'b1001 : 4'b0000;
																assign node9807 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node9810 = (inp[7]) ? node9814 : node9811;
																assign node9811 = (inp[0]) ? 4'b1001 : 4'b0001;
																assign node9814 = (inp[0]) ? 4'b0000 : 4'b1001;
														assign node9817 = (inp[7]) ? node9819 : 4'b0000;
															assign node9819 = (inp[0]) ? 4'b1001 : 4'b0000;
												assign node9822 = (inp[7]) ? node9844 : node9823;
													assign node9823 = (inp[2]) ? node9833 : node9824;
														assign node9824 = (inp[14]) ? node9826 : 4'b0000;
															assign node9826 = (inp[10]) ? node9830 : node9827;
																assign node9827 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node9830 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node9833 = (inp[0]) ? node9841 : node9834;
															assign node9834 = (inp[10]) ? node9838 : node9835;
																assign node9835 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node9838 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node9841 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node9844 = (inp[10]) ? node9854 : node9845;
														assign node9845 = (inp[0]) ? node9851 : node9846;
															assign node9846 = (inp[14]) ? 4'b0000 : node9847;
																assign node9847 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node9851 = (inp[2]) ? 4'b0000 : 4'b1001;
														assign node9854 = (inp[0]) ? node9858 : node9855;
															assign node9855 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node9858 = (inp[14]) ? 4'b0001 : node9859;
																assign node9859 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node9863 = (inp[0]) ? node9905 : node9864;
												assign node9864 = (inp[2]) ? node9886 : node9865;
													assign node9865 = (inp[7]) ? node9875 : node9866;
														assign node9866 = (inp[10]) ? node9872 : node9867;
															assign node9867 = (inp[13]) ? 4'b1000 : node9868;
																assign node9868 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9872 = (inp[13]) ? 4'b1001 : 4'b0000;
														assign node9875 = (inp[13]) ? node9879 : node9876;
															assign node9876 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node9879 = (inp[14]) ? node9883 : node9880;
																assign node9880 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node9883 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node9886 = (inp[14]) ? node9894 : node9887;
														assign node9887 = (inp[13]) ? node9891 : node9888;
															assign node9888 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node9891 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node9894 = (inp[7]) ? node9900 : node9895;
															assign node9895 = (inp[13]) ? node9897 : 4'b0001;
																assign node9897 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node9900 = (inp[10]) ? 4'b0000 : node9901;
																assign node9901 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node9905 = (inp[2]) ? node9931 : node9906;
													assign node9906 = (inp[7]) ? node9918 : node9907;
														assign node9907 = (inp[13]) ? node9913 : node9908;
															assign node9908 = (inp[14]) ? node9910 : 4'b0001;
																assign node9910 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node9913 = (inp[10]) ? 4'b0000 : node9914;
																assign node9914 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node9918 = (inp[10]) ? node9924 : node9919;
															assign node9919 = (inp[13]) ? 4'b0001 : node9920;
																assign node9920 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node9924 = (inp[13]) ? node9928 : node9925;
																assign node9925 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node9928 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node9931 = (inp[14]) ? node9943 : node9932;
														assign node9932 = (inp[10]) ? node9938 : node9933;
															assign node9933 = (inp[13]) ? node9935 : 4'b0000;
																assign node9935 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node9938 = (inp[7]) ? node9940 : 4'b1000;
																assign node9940 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node9943 = (inp[13]) ? node9945 : 4'b0001;
															assign node9945 = (inp[7]) ? 4'b1001 : node9946;
																assign node9946 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node9950 = (inp[0]) ? node9994 : node9951;
											assign node9951 = (inp[10]) ? node9977 : node9952;
												assign node9952 = (inp[7]) ? node9966 : node9953;
													assign node9953 = (inp[12]) ? node9959 : node9954;
														assign node9954 = (inp[2]) ? 4'b0001 : node9955;
															assign node9955 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node9959 = (inp[2]) ? node9963 : node9960;
															assign node9960 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node9963 = (inp[13]) ? 4'b0001 : 4'b1000;
													assign node9966 = (inp[13]) ? node9972 : node9967;
														assign node9967 = (inp[12]) ? node9969 : 4'b0000;
															assign node9969 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node9972 = (inp[2]) ? 4'b1000 : node9973;
															assign node9973 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node9977 = (inp[2]) ? node9983 : node9978;
													assign node9978 = (inp[7]) ? node9980 : 4'b1000;
														assign node9980 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node9983 = (inp[13]) ? node9989 : node9984;
														assign node9984 = (inp[12]) ? 4'b0001 : node9985;
															assign node9985 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node9989 = (inp[7]) ? 4'b0000 : node9990;
															assign node9990 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node9994 = (inp[13]) ? node10012 : node9995;
												assign node9995 = (inp[10]) ? node10001 : node9996;
													assign node9996 = (inp[2]) ? node9998 : 4'b1000;
														assign node9998 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node10001 = (inp[7]) ? node10007 : node10002;
														assign node10002 = (inp[2]) ? node10004 : 4'b1001;
															assign node10004 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node10007 = (inp[12]) ? node10009 : 4'b1000;
															assign node10009 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node10012 = (inp[2]) ? node10028 : node10013;
													assign node10013 = (inp[12]) ? node10021 : node10014;
														assign node10014 = (inp[10]) ? node10018 : node10015;
															assign node10015 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node10018 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node10021 = (inp[7]) ? node10025 : node10022;
															assign node10022 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node10025 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node10028 = (inp[12]) ? node10034 : node10029;
														assign node10029 = (inp[10]) ? node10031 : 4'b0000;
															assign node10031 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10034 = (inp[7]) ? node10038 : node10035;
															assign node10035 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node10038 = (inp[10]) ? 4'b0000 : 4'b1000;
									assign node10041 = (inp[11]) ? node10175 : node10042;
										assign node10042 = (inp[13]) ? node10108 : node10043;
											assign node10043 = (inp[2]) ? node10077 : node10044;
												assign node10044 = (inp[10]) ? node10066 : node10045;
													assign node10045 = (inp[14]) ? node10055 : node10046;
														assign node10046 = (inp[7]) ? node10050 : node10047;
															assign node10047 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node10050 = (inp[12]) ? 4'b1000 : node10051;
																assign node10051 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node10055 = (inp[7]) ? node10061 : node10056;
															assign node10056 = (inp[0]) ? node10058 : 4'b1001;
																assign node10058 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node10061 = (inp[0]) ? 4'b1001 : node10062;
																assign node10062 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node10066 = (inp[0]) ? node10070 : node10067;
														assign node10067 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10070 = (inp[12]) ? node10072 : 4'b0001;
															assign node10072 = (inp[7]) ? node10074 : 4'b1001;
																assign node10074 = (inp[14]) ? 4'b0001 : 4'b1000;
												assign node10077 = (inp[14]) ? node10093 : node10078;
													assign node10078 = (inp[7]) ? node10084 : node10079;
														assign node10079 = (inp[12]) ? 4'b0000 : node10080;
															assign node10080 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node10084 = (inp[10]) ? node10090 : node10085;
															assign node10085 = (inp[12]) ? 4'b0001 : node10086;
																assign node10086 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node10090 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node10093 = (inp[12]) ? node10105 : node10094;
														assign node10094 = (inp[0]) ? node10100 : node10095;
															assign node10095 = (inp[10]) ? 4'b0001 : node10096;
																assign node10096 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node10100 = (inp[10]) ? node10102 : 4'b1000;
																assign node10102 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node10105 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node10108 = (inp[10]) ? node10142 : node10109;
												assign node10109 = (inp[7]) ? node10121 : node10110;
													assign node10110 = (inp[0]) ? node10118 : node10111;
														assign node10111 = (inp[2]) ? 4'b1001 : node10112;
															assign node10112 = (inp[14]) ? 4'b1001 : node10113;
																assign node10113 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node10118 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10121 = (inp[12]) ? node10131 : node10122;
														assign node10122 = (inp[14]) ? node10124 : 4'b0001;
															assign node10124 = (inp[0]) ? node10128 : node10125;
																assign node10125 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node10128 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node10131 = (inp[0]) ? node10137 : node10132;
															assign node10132 = (inp[2]) ? node10134 : 4'b0000;
																assign node10134 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node10137 = (inp[2]) ? node10139 : 4'b1001;
																assign node10139 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node10142 = (inp[0]) ? node10160 : node10143;
													assign node10143 = (inp[7]) ? node10149 : node10144;
														assign node10144 = (inp[2]) ? 4'b1000 : node10145;
															assign node10145 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node10149 = (inp[14]) ? node10155 : node10150;
															assign node10150 = (inp[12]) ? node10152 : 4'b1001;
																assign node10152 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node10155 = (inp[12]) ? node10157 : 4'b1000;
																assign node10157 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node10160 = (inp[2]) ? node10168 : node10161;
														assign node10161 = (inp[12]) ? node10163 : 4'b0000;
															assign node10163 = (inp[7]) ? node10165 : 4'b1000;
																assign node10165 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10168 = (inp[7]) ? 4'b0000 : node10169;
															assign node10169 = (inp[14]) ? node10171 : 4'b0000;
																assign node10171 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node10175 = (inp[13]) ? node10219 : node10176;
											assign node10176 = (inp[2]) ? node10188 : node10177;
												assign node10177 = (inp[7]) ? node10179 : 4'b0001;
													assign node10179 = (inp[0]) ? node10183 : node10180;
														assign node10180 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node10183 = (inp[12]) ? node10185 : 4'b0001;
															assign node10185 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node10188 = (inp[12]) ? node10198 : node10189;
													assign node10189 = (inp[10]) ? node10191 : 4'b1001;
														assign node10191 = (inp[7]) ? node10195 : node10192;
															assign node10192 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node10195 = (inp[0]) ? 4'b1001 : 4'b0001;
													assign node10198 = (inp[10]) ? node10204 : node10199;
														assign node10199 = (inp[7]) ? 4'b0001 : node10200;
															assign node10200 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node10204 = (inp[14]) ? node10212 : node10205;
															assign node10205 = (inp[7]) ? node10209 : node10206;
																assign node10206 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node10209 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node10212 = (inp[7]) ? node10216 : node10213;
																assign node10213 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node10216 = (inp[0]) ? 4'b1001 : 4'b0001;
											assign node10219 = (inp[10]) ? 4'b0001 : node10220;
												assign node10220 = (inp[0]) ? node10228 : node10221;
													assign node10221 = (inp[12]) ? 4'b0001 : node10222;
														assign node10222 = (inp[7]) ? node10224 : 4'b0001;
															assign node10224 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node10228 = (inp[7]) ? node10236 : node10229;
														assign node10229 = (inp[14]) ? node10231 : 4'b1001;
															assign node10231 = (inp[2]) ? 4'b1001 : node10232;
																assign node10232 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node10236 = (inp[2]) ? node10238 : 4'b0001;
															assign node10238 = (inp[12]) ? 4'b1001 : 4'b0001;
								assign node10242 = (inp[13]) ? node10522 : node10243;
									assign node10243 = (inp[1]) ? node10385 : node10244;
										assign node10244 = (inp[0]) ? node10320 : node10245;
											assign node10245 = (inp[2]) ? node10289 : node10246;
												assign node10246 = (inp[14]) ? node10264 : node10247;
													assign node10247 = (inp[10]) ? node10253 : node10248;
														assign node10248 = (inp[7]) ? 4'b0001 : node10249;
															assign node10249 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node10253 = (inp[12]) ? node10259 : node10254;
															assign node10254 = (inp[11]) ? node10256 : 4'b0000;
																assign node10256 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node10259 = (inp[11]) ? 4'b0001 : node10260;
																assign node10260 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node10264 = (inp[12]) ? node10278 : node10265;
														assign node10265 = (inp[7]) ? node10271 : node10266;
															assign node10266 = (inp[11]) ? node10268 : 4'b0001;
																assign node10268 = (inp[10]) ? 4'b0001 : 4'b1000;
															assign node10271 = (inp[11]) ? node10275 : node10272;
																assign node10272 = (inp[10]) ? 4'b1001 : 4'b0000;
																assign node10275 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node10278 = (inp[10]) ? node10284 : node10279;
															assign node10279 = (inp[7]) ? 4'b0000 : node10280;
																assign node10280 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node10284 = (inp[11]) ? 4'b0001 : node10285;
																assign node10285 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node10289 = (inp[12]) ? node10307 : node10290;
													assign node10290 = (inp[10]) ? node10300 : node10291;
														assign node10291 = (inp[11]) ? node10297 : node10292;
															assign node10292 = (inp[7]) ? node10294 : 4'b0001;
																assign node10294 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10297 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node10300 = (inp[14]) ? node10302 : 4'b0001;
															assign node10302 = (inp[11]) ? 4'b0001 : node10303;
																assign node10303 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node10307 = (inp[10]) ? node10313 : node10308;
														assign node10308 = (inp[7]) ? 4'b1000 : node10309;
															assign node10309 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10313 = (inp[11]) ? node10317 : node10314;
															assign node10314 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node10317 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node10320 = (inp[12]) ? node10346 : node10321;
												assign node10321 = (inp[10]) ? node10335 : node10322;
													assign node10322 = (inp[11]) ? node10328 : node10323;
														assign node10323 = (inp[14]) ? 4'b1000 : node10324;
															assign node10324 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node10328 = (inp[2]) ? node10332 : node10329;
															assign node10329 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node10332 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node10335 = (inp[7]) ? node10339 : node10336;
														assign node10336 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node10339 = (inp[2]) ? node10341 : 4'b0001;
															assign node10341 = (inp[11]) ? 4'b1000 : node10342;
																assign node10342 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node10346 = (inp[2]) ? node10368 : node10347;
													assign node10347 = (inp[7]) ? node10355 : node10348;
														assign node10348 = (inp[10]) ? 4'b0000 : node10349;
															assign node10349 = (inp[11]) ? 4'b0001 : node10350;
																assign node10350 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node10355 = (inp[14]) ? node10363 : node10356;
															assign node10356 = (inp[11]) ? node10360 : node10357;
																assign node10357 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node10360 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node10363 = (inp[11]) ? node10365 : 4'b1000;
																assign node10365 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node10368 = (inp[11]) ? node10380 : node10369;
														assign node10369 = (inp[14]) ? node10375 : node10370;
															assign node10370 = (inp[10]) ? 4'b0001 : node10371;
																assign node10371 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node10375 = (inp[10]) ? node10377 : 4'b0000;
																assign node10377 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node10380 = (inp[10]) ? 4'b0000 : node10381;
															assign node10381 = (inp[7]) ? 4'b0001 : 4'b1000;
										assign node10385 = (inp[11]) ? node10489 : node10386;
											assign node10386 = (inp[10]) ? node10434 : node10387;
												assign node10387 = (inp[12]) ? node10413 : node10388;
													assign node10388 = (inp[7]) ? node10400 : node10389;
														assign node10389 = (inp[0]) ? node10395 : node10390;
															assign node10390 = (inp[14]) ? node10392 : 4'b0000;
																assign node10392 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node10395 = (inp[14]) ? node10397 : 4'b0001;
																assign node10397 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node10400 = (inp[0]) ? node10406 : node10401;
															assign node10401 = (inp[14]) ? node10403 : 4'b1001;
																assign node10403 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node10406 = (inp[14]) ? node10410 : node10407;
																assign node10407 = (inp[2]) ? 4'b0000 : 4'b1000;
																assign node10410 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node10413 = (inp[7]) ? node10425 : node10414;
														assign node10414 = (inp[0]) ? node10420 : node10415;
															assign node10415 = (inp[14]) ? 4'b1000 : node10416;
																assign node10416 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node10420 = (inp[14]) ? 4'b1001 : node10421;
																assign node10421 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node10425 = (inp[2]) ? node10431 : node10426;
															assign node10426 = (inp[0]) ? 4'b0001 : node10427;
																assign node10427 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10431 = (inp[0]) ? 4'b1000 : 4'b0001;
												assign node10434 = (inp[12]) ? node10466 : node10435;
													assign node10435 = (inp[14]) ? node10451 : node10436;
														assign node10436 = (inp[0]) ? node10444 : node10437;
															assign node10437 = (inp[7]) ? node10441 : node10438;
																assign node10438 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node10441 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node10444 = (inp[2]) ? node10448 : node10445;
																assign node10445 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node10448 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10451 = (inp[2]) ? node10459 : node10452;
															assign node10452 = (inp[7]) ? node10456 : node10453;
																assign node10453 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node10456 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node10459 = (inp[0]) ? node10463 : node10460;
																assign node10460 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node10463 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node10466 = (inp[7]) ? node10478 : node10467;
														assign node10467 = (inp[0]) ? node10473 : node10468;
															assign node10468 = (inp[2]) ? node10470 : 4'b1000;
																assign node10470 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node10473 = (inp[2]) ? node10475 : 4'b0001;
																assign node10475 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10478 = (inp[0]) ? node10482 : node10479;
															assign node10479 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node10482 = (inp[2]) ? node10486 : node10483;
																assign node10483 = (inp[14]) ? 4'b1000 : 4'b0000;
																assign node10486 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node10489 = (inp[10]) ? 4'b0001 : node10490;
												assign node10490 = (inp[12]) ? node10502 : node10491;
													assign node10491 = (inp[2]) ? node10497 : node10492;
														assign node10492 = (inp[0]) ? node10494 : 4'b0001;
															assign node10494 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node10497 = (inp[0]) ? 4'b0001 : node10498;
															assign node10498 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node10502 = (inp[2]) ? node10508 : node10503;
														assign node10503 = (inp[0]) ? 4'b0001 : node10504;
															assign node10504 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node10508 = (inp[14]) ? node10516 : node10509;
															assign node10509 = (inp[7]) ? node10513 : node10510;
																assign node10510 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node10513 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node10516 = (inp[7]) ? node10518 : 4'b1001;
																assign node10518 = (inp[0]) ? 4'b1001 : 4'b0001;
									assign node10522 = (inp[10]) ? node10648 : node10523;
										assign node10523 = (inp[1]) ? node10607 : node10524;
											assign node10524 = (inp[11]) ? node10566 : node10525;
												assign node10525 = (inp[12]) ? node10543 : node10526;
													assign node10526 = (inp[2]) ? node10532 : node10527;
														assign node10527 = (inp[14]) ? node10529 : 4'b0000;
															assign node10529 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node10532 = (inp[0]) ? node10538 : node10533;
															assign node10533 = (inp[7]) ? node10535 : 4'b0000;
																assign node10535 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10538 = (inp[7]) ? node10540 : 4'b0001;
																assign node10540 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10543 = (inp[7]) ? node10555 : node10544;
														assign node10544 = (inp[0]) ? node10550 : node10545;
															assign node10545 = (inp[14]) ? node10547 : 4'b0000;
																assign node10547 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node10550 = (inp[14]) ? node10552 : 4'b0001;
																assign node10552 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node10555 = (inp[0]) ? node10561 : node10556;
															assign node10556 = (inp[14]) ? node10558 : 4'b0001;
																assign node10558 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node10561 = (inp[2]) ? node10563 : 4'b0000;
																assign node10563 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node10566 = (inp[14]) ? node10586 : node10567;
													assign node10567 = (inp[7]) ? node10577 : node10568;
														assign node10568 = (inp[12]) ? node10570 : 4'b0000;
															assign node10570 = (inp[0]) ? node10574 : node10571;
																assign node10571 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node10574 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node10577 = (inp[12]) ? 4'b0000 : node10578;
															assign node10578 = (inp[0]) ? node10582 : node10579;
																assign node10579 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node10582 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node10586 = (inp[0]) ? node10596 : node10587;
														assign node10587 = (inp[12]) ? 4'b0000 : node10588;
															assign node10588 = (inp[2]) ? node10592 : node10589;
																assign node10589 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node10592 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node10596 = (inp[12]) ? node10602 : node10597;
															assign node10597 = (inp[2]) ? node10599 : 4'b0000;
																assign node10599 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node10602 = (inp[2]) ? node10604 : 4'b0001;
																assign node10604 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node10607 = (inp[11]) ? 4'b0001 : node10608;
												assign node10608 = (inp[0]) ? node10628 : node10609;
													assign node10609 = (inp[2]) ? node10617 : node10610;
														assign node10610 = (inp[7]) ? 4'b0000 : node10611;
															assign node10611 = (inp[12]) ? 4'b0001 : node10612;
																assign node10612 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10617 = (inp[12]) ? node10623 : node10618;
															assign node10618 = (inp[7]) ? node10620 : 4'b0001;
																assign node10620 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10623 = (inp[7]) ? 4'b0001 : node10624;
																assign node10624 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node10628 = (inp[7]) ? node10636 : node10629;
														assign node10629 = (inp[2]) ? 4'b0000 : node10630;
															assign node10630 = (inp[12]) ? 4'b0000 : node10631;
																assign node10631 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node10636 = (inp[2]) ? node10642 : node10637;
															assign node10637 = (inp[12]) ? node10639 : 4'b0001;
																assign node10639 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node10642 = (inp[14]) ? node10644 : 4'b0000;
																assign node10644 = (inp[12]) ? 4'b0000 : 4'b0001;
										assign node10648 = (inp[1]) ? 4'b0000 : node10649;
											assign node10649 = (inp[11]) ? 4'b0000 : node10650;
												assign node10650 = (inp[0]) ? node10668 : node10651;
													assign node10651 = (inp[12]) ? node10659 : node10652;
														assign node10652 = (inp[2]) ? node10654 : 4'b0000;
															assign node10654 = (inp[14]) ? 4'b0001 : node10655;
																assign node10655 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10659 = (inp[2]) ? 4'b0000 : node10660;
															assign node10660 = (inp[14]) ? node10664 : node10661;
																assign node10661 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node10664 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node10668 = (inp[12]) ? node10670 : 4'b0000;
														assign node10670 = (inp[7]) ? node10672 : 4'b0000;
															assign node10672 = (inp[2]) ? node10676 : node10673;
																assign node10673 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node10676 = (inp[14]) ? 4'b0000 : 4'b0001;
				assign node10681 = (inp[0]) ? node13069 : node10682;
					assign node10682 = (inp[6]) ? node11304 : node10683;
						assign node10683 = (inp[2]) ? node11187 : node10684;
							assign node10684 = (inp[5]) ? node10798 : node10685;
								assign node10685 = (inp[3]) ? node10687 : 4'b0011;
									assign node10687 = (inp[4]) ? node10709 : node10688;
										assign node10688 = (inp[13]) ? node10690 : 4'b0011;
											assign node10690 = (inp[7]) ? 4'b0011 : node10691;
												assign node10691 = (inp[12]) ? node10699 : node10692;
													assign node10692 = (inp[1]) ? node10694 : 4'b0000;
														assign node10694 = (inp[14]) ? node10696 : 4'b0001;
															assign node10696 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node10699 = (inp[10]) ? node10701 : 4'b0011;
														assign node10701 = (inp[1]) ? 4'b0001 : node10702;
															assign node10702 = (inp[11]) ? 4'b0000 : node10703;
																assign node10703 = (inp[14]) ? 4'b0011 : 4'b0000;
										assign node10709 = (inp[7]) ? node10775 : node10710;
											assign node10710 = (inp[1]) ? node10742 : node10711;
												assign node10711 = (inp[11]) ? node10731 : node10712;
													assign node10712 = (inp[14]) ? node10720 : node10713;
														assign node10713 = (inp[13]) ? 4'b0000 : node10714;
															assign node10714 = (inp[12]) ? node10716 : 4'b1000;
																assign node10716 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10720 = (inp[13]) ? node10726 : node10721;
															assign node10721 = (inp[12]) ? 4'b0001 : node10722;
																assign node10722 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node10726 = (inp[10]) ? node10728 : 4'b1001;
																assign node10728 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node10731 = (inp[13]) ? node10737 : node10732;
														assign node10732 = (inp[12]) ? node10734 : 4'b1000;
															assign node10734 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node10737 = (inp[12]) ? node10739 : 4'b0000;
															assign node10739 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node10742 = (inp[11]) ? node10764 : node10743;
													assign node10743 = (inp[14]) ? node10753 : node10744;
														assign node10744 = (inp[10]) ? node10750 : node10745;
															assign node10745 = (inp[13]) ? 4'b1001 : node10746;
																assign node10746 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node10750 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node10753 = (inp[13]) ? node10759 : node10754;
															assign node10754 = (inp[12]) ? node10756 : 4'b1000;
																assign node10756 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node10759 = (inp[12]) ? node10761 : 4'b0000;
																assign node10761 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node10764 = (inp[13]) ? node10770 : node10765;
														assign node10765 = (inp[10]) ? 4'b1001 : node10766;
															assign node10766 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node10770 = (inp[10]) ? 4'b0001 : node10771;
															assign node10771 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node10775 = (inp[13]) ? node10777 : 4'b0011;
												assign node10777 = (inp[10]) ? node10787 : node10778;
													assign node10778 = (inp[12]) ? 4'b0011 : node10779;
														assign node10779 = (inp[1]) ? node10783 : node10780;
															assign node10780 = (inp[14]) ? 4'b0011 : 4'b0000;
															assign node10783 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node10787 = (inp[1]) ? node10793 : node10788;
														assign node10788 = (inp[14]) ? node10790 : 4'b0000;
															assign node10790 = (inp[11]) ? 4'b0000 : 4'b0011;
														assign node10793 = (inp[11]) ? 4'b0001 : node10794;
															assign node10794 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node10798 = (inp[1]) ? node10998 : node10799;
									assign node10799 = (inp[11]) ? node10927 : node10800;
										assign node10800 = (inp[14]) ? node10858 : node10801;
											assign node10801 = (inp[13]) ? node10827 : node10802;
												assign node10802 = (inp[3]) ? node10814 : node10803;
													assign node10803 = (inp[12]) ? node10805 : 4'b1000;
														assign node10805 = (inp[10]) ? node10811 : node10806;
															assign node10806 = (inp[7]) ? 4'b0000 : node10807;
																assign node10807 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node10811 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node10814 = (inp[4]) ? node10820 : node10815;
														assign node10815 = (inp[12]) ? node10817 : 4'b1100;
															assign node10817 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node10820 = (inp[7]) ? 4'b1100 : node10821;
															assign node10821 = (inp[10]) ? 4'b1000 : node10822;
																assign node10822 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node10827 = (inp[10]) ? node10847 : node10828;
													assign node10828 = (inp[12]) ? node10836 : node10829;
														assign node10829 = (inp[3]) ? node10831 : 4'b0100;
															assign node10831 = (inp[4]) ? 4'b0000 : node10832;
																assign node10832 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node10836 = (inp[3]) ? node10842 : node10837;
															assign node10837 = (inp[7]) ? 4'b1000 : node10838;
																assign node10838 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node10842 = (inp[4]) ? node10844 : 4'b1100;
																assign node10844 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node10847 = (inp[3]) ? node10853 : node10848;
														assign node10848 = (inp[7]) ? node10850 : 4'b0100;
															assign node10850 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10853 = (inp[7]) ? node10855 : 4'b0000;
															assign node10855 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node10858 = (inp[13]) ? node10892 : node10859;
												assign node10859 = (inp[10]) ? node10871 : node10860;
													assign node10860 = (inp[3]) ? node10866 : node10861;
														assign node10861 = (inp[4]) ? node10863 : 4'b0001;
															assign node10863 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node10866 = (inp[7]) ? 4'b0101 : node10867;
															assign node10867 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node10871 = (inp[12]) ? node10883 : node10872;
														assign node10872 = (inp[3]) ? node10878 : node10873;
															assign node10873 = (inp[4]) ? node10875 : 4'b1001;
																assign node10875 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node10878 = (inp[4]) ? node10880 : 4'b1101;
																assign node10880 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node10883 = (inp[7]) ? node10889 : node10884;
															assign node10884 = (inp[3]) ? node10886 : 4'b0101;
																assign node10886 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node10889 = (inp[3]) ? 4'b0101 : 4'b0001;
												assign node10892 = (inp[12]) ? node10916 : node10893;
													assign node10893 = (inp[10]) ? node10905 : node10894;
														assign node10894 = (inp[3]) ? node10900 : node10895;
															assign node10895 = (inp[4]) ? node10897 : 4'b1001;
																assign node10897 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node10900 = (inp[4]) ? node10902 : 4'b1101;
																assign node10902 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node10905 = (inp[3]) ? node10911 : node10906;
															assign node10906 = (inp[7]) ? node10908 : 4'b0101;
																assign node10908 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node10911 = (inp[7]) ? node10913 : 4'b0001;
																assign node10913 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node10916 = (inp[3]) ? node10922 : node10917;
														assign node10917 = (inp[7]) ? 4'b1001 : node10918;
															assign node10918 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node10922 = (inp[7]) ? 4'b1101 : node10923;
															assign node10923 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node10927 = (inp[13]) ? node10963 : node10928;
											assign node10928 = (inp[10]) ? node10952 : node10929;
												assign node10929 = (inp[12]) ? node10941 : node10930;
													assign node10930 = (inp[3]) ? node10936 : node10931;
														assign node10931 = (inp[7]) ? 4'b1000 : node10932;
															assign node10932 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node10936 = (inp[4]) ? node10938 : 4'b1100;
															assign node10938 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node10941 = (inp[3]) ? node10947 : node10942;
														assign node10942 = (inp[7]) ? 4'b0000 : node10943;
															assign node10943 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10947 = (inp[4]) ? node10949 : 4'b0100;
															assign node10949 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node10952 = (inp[3]) ? node10958 : node10953;
													assign node10953 = (inp[7]) ? 4'b1000 : node10954;
														assign node10954 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node10958 = (inp[4]) ? node10960 : 4'b1100;
														assign node10960 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node10963 = (inp[12]) ? node10975 : node10964;
												assign node10964 = (inp[3]) ? node10970 : node10965;
													assign node10965 = (inp[4]) ? 4'b0100 : node10966;
														assign node10966 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node10970 = (inp[7]) ? node10972 : 4'b0000;
														assign node10972 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node10975 = (inp[10]) ? node10987 : node10976;
													assign node10976 = (inp[3]) ? node10982 : node10977;
														assign node10977 = (inp[7]) ? 4'b1000 : node10978;
															assign node10978 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node10982 = (inp[7]) ? 4'b1100 : node10983;
															assign node10983 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node10987 = (inp[3]) ? node10993 : node10988;
														assign node10988 = (inp[7]) ? node10990 : 4'b0100;
															assign node10990 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10993 = (inp[7]) ? node10995 : 4'b0000;
															assign node10995 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node10998 = (inp[13]) ? node11090 : node10999;
										assign node10999 = (inp[3]) ? node11047 : node11000;
											assign node11000 = (inp[7]) ? node11030 : node11001;
												assign node11001 = (inp[4]) ? node11013 : node11002;
													assign node11002 = (inp[10]) ? node11008 : node11003;
														assign node11003 = (inp[12]) ? 4'b0001 : node11004;
															assign node11004 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11008 = (inp[14]) ? node11010 : 4'b1001;
															assign node11010 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11013 = (inp[12]) ? node11019 : node11014;
														assign node11014 = (inp[11]) ? 4'b1101 : node11015;
															assign node11015 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node11019 = (inp[10]) ? node11025 : node11020;
															assign node11020 = (inp[11]) ? 4'b0101 : node11021;
																assign node11021 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node11025 = (inp[11]) ? 4'b1101 : node11026;
																assign node11026 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node11030 = (inp[10]) ? node11042 : node11031;
													assign node11031 = (inp[12]) ? node11037 : node11032;
														assign node11032 = (inp[14]) ? node11034 : 4'b1001;
															assign node11034 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11037 = (inp[11]) ? 4'b0001 : node11038;
															assign node11038 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11042 = (inp[11]) ? 4'b1001 : node11043;
														assign node11043 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node11047 = (inp[14]) ? node11061 : node11048;
												assign node11048 = (inp[7]) ? node11056 : node11049;
													assign node11049 = (inp[4]) ? 4'b1001 : node11050;
														assign node11050 = (inp[10]) ? 4'b1101 : node11051;
															assign node11051 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node11056 = (inp[10]) ? 4'b1101 : node11057;
														assign node11057 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node11061 = (inp[11]) ? node11077 : node11062;
													assign node11062 = (inp[7]) ? node11072 : node11063;
														assign node11063 = (inp[4]) ? node11067 : node11064;
															assign node11064 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node11067 = (inp[12]) ? node11069 : 4'b1000;
																assign node11069 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node11072 = (inp[10]) ? 4'b1100 : node11073;
															assign node11073 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node11077 = (inp[12]) ? node11083 : node11078;
														assign node11078 = (inp[7]) ? 4'b1101 : node11079;
															assign node11079 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node11083 = (inp[10]) ? 4'b1101 : node11084;
															assign node11084 = (inp[4]) ? node11086 : 4'b0101;
																assign node11086 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node11090 = (inp[11]) ? node11152 : node11091;
											assign node11091 = (inp[14]) ? node11119 : node11092;
												assign node11092 = (inp[12]) ? node11104 : node11093;
													assign node11093 = (inp[3]) ? node11099 : node11094;
														assign node11094 = (inp[4]) ? 4'b0101 : node11095;
															assign node11095 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11099 = (inp[4]) ? 4'b0001 : node11100;
															assign node11100 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node11104 = (inp[10]) ? node11110 : node11105;
														assign node11105 = (inp[4]) ? 4'b1101 : node11106;
															assign node11106 = (inp[3]) ? 4'b1101 : 4'b1001;
														assign node11110 = (inp[3]) ? node11116 : node11111;
															assign node11111 = (inp[7]) ? node11113 : 4'b0101;
																assign node11113 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node11116 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node11119 = (inp[10]) ? node11141 : node11120;
													assign node11120 = (inp[12]) ? node11132 : node11121;
														assign node11121 = (inp[3]) ? node11127 : node11122;
															assign node11122 = (inp[4]) ? 4'b0100 : node11123;
																assign node11123 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node11127 = (inp[4]) ? 4'b0000 : node11128;
																assign node11128 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node11132 = (inp[3]) ? node11138 : node11133;
															assign node11133 = (inp[7]) ? 4'b1000 : node11134;
																assign node11134 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node11138 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node11141 = (inp[3]) ? node11147 : node11142;
														assign node11142 = (inp[4]) ? 4'b0100 : node11143;
															assign node11143 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11147 = (inp[7]) ? node11149 : 4'b0000;
															assign node11149 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node11152 = (inp[12]) ? node11164 : node11153;
												assign node11153 = (inp[3]) ? node11159 : node11154;
													assign node11154 = (inp[4]) ? 4'b0101 : node11155;
														assign node11155 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node11159 = (inp[7]) ? node11161 : 4'b0001;
														assign node11161 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node11164 = (inp[10]) ? node11176 : node11165;
													assign node11165 = (inp[3]) ? node11171 : node11166;
														assign node11166 = (inp[4]) ? node11168 : 4'b1001;
															assign node11168 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node11171 = (inp[7]) ? 4'b1101 : node11172;
															assign node11172 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node11176 = (inp[3]) ? node11182 : node11177;
														assign node11177 = (inp[7]) ? node11179 : 4'b0101;
															assign node11179 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node11182 = (inp[7]) ? node11184 : 4'b0001;
															assign node11184 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node11187 = (inp[5]) ? node11189 : 4'b0011;
								assign node11189 = (inp[3]) ? node11191 : 4'b0011;
									assign node11191 = (inp[7]) ? node11273 : node11192;
										assign node11192 = (inp[4]) ? node11216 : node11193;
											assign node11193 = (inp[13]) ? node11195 : 4'b0011;
												assign node11195 = (inp[12]) ? node11209 : node11196;
													assign node11196 = (inp[1]) ? node11204 : node11197;
														assign node11197 = (inp[14]) ? node11199 : 4'b0000;
															assign node11199 = (inp[11]) ? 4'b0000 : node11200;
																assign node11200 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node11204 = (inp[11]) ? 4'b0001 : node11205;
															assign node11205 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11209 = (inp[10]) ? node11211 : 4'b0011;
														assign node11211 = (inp[1]) ? 4'b0001 : node11212;
															assign node11212 = (inp[11]) ? 4'b0000 : 4'b0011;
											assign node11216 = (inp[1]) ? node11246 : node11217;
												assign node11217 = (inp[14]) ? node11229 : node11218;
													assign node11218 = (inp[13]) ? node11224 : node11219;
														assign node11219 = (inp[10]) ? 4'b1000 : node11220;
															assign node11220 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node11224 = (inp[12]) ? node11226 : 4'b0000;
															assign node11226 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node11229 = (inp[11]) ? node11241 : node11230;
														assign node11230 = (inp[13]) ? node11236 : node11231;
															assign node11231 = (inp[10]) ? node11233 : 4'b0001;
																assign node11233 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11236 = (inp[10]) ? node11238 : 4'b1001;
																assign node11238 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node11241 = (inp[13]) ? 4'b0000 : node11242;
															assign node11242 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node11246 = (inp[11]) ? node11262 : node11247;
													assign node11247 = (inp[14]) ? node11255 : node11248;
														assign node11248 = (inp[12]) ? node11252 : node11249;
															assign node11249 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node11252 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node11255 = (inp[13]) ? 4'b0000 : node11256;
															assign node11256 = (inp[12]) ? node11258 : 4'b1000;
																assign node11258 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node11262 = (inp[13]) ? node11268 : node11263;
														assign node11263 = (inp[10]) ? 4'b1001 : node11264;
															assign node11264 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node11268 = (inp[10]) ? 4'b0001 : node11269;
															assign node11269 = (inp[14]) ? 4'b1001 : 4'b0001;
										assign node11273 = (inp[13]) ? node11275 : 4'b0011;
											assign node11275 = (inp[4]) ? node11277 : 4'b0011;
												assign node11277 = (inp[12]) ? node11291 : node11278;
													assign node11278 = (inp[1]) ? node11286 : node11279;
														assign node11279 = (inp[11]) ? 4'b0000 : node11280;
															assign node11280 = (inp[14]) ? node11282 : 4'b0000;
																assign node11282 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node11286 = (inp[11]) ? 4'b0001 : node11287;
															assign node11287 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node11291 = (inp[10]) ? node11293 : 4'b0011;
														assign node11293 = (inp[1]) ? node11299 : node11294;
															assign node11294 = (inp[11]) ? 4'b0000 : node11295;
																assign node11295 = (inp[14]) ? 4'b0011 : 4'b0000;
															assign node11299 = (inp[14]) ? node11301 : 4'b0001;
																assign node11301 = (inp[11]) ? 4'b0001 : 4'b0000;
						assign node11304 = (inp[1]) ? node12290 : node11305;
							assign node11305 = (inp[5]) ? node11819 : node11306;
								assign node11306 = (inp[14]) ? node11546 : node11307;
									assign node11307 = (inp[13]) ? node11393 : node11308;
										assign node11308 = (inp[3]) ? node11330 : node11309;
											assign node11309 = (inp[7]) ? node11325 : node11310;
												assign node11310 = (inp[4]) ? node11316 : node11311;
													assign node11311 = (inp[12]) ? node11313 : 4'b1000;
														assign node11313 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node11316 = (inp[12]) ? node11322 : node11317;
														assign node11317 = (inp[2]) ? 4'b1100 : node11318;
															assign node11318 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node11322 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node11325 = (inp[12]) ? node11327 : 4'b1000;
													assign node11327 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node11330 = (inp[2]) ? node11372 : node11331;
												assign node11331 = (inp[11]) ? node11353 : node11332;
													assign node11332 = (inp[4]) ? node11344 : node11333;
														assign node11333 = (inp[7]) ? node11339 : node11334;
															assign node11334 = (inp[10]) ? 4'b0100 : node11335;
																assign node11335 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11339 = (inp[10]) ? node11341 : 4'b0000;
																assign node11341 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node11344 = (inp[10]) ? node11348 : node11345;
															assign node11345 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node11348 = (inp[12]) ? 4'b1100 : node11349;
																assign node11349 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node11353 = (inp[4]) ? node11363 : node11354;
														assign node11354 = (inp[12]) ? node11360 : node11355;
															assign node11355 = (inp[10]) ? node11357 : 4'b1001;
																assign node11357 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node11360 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node11363 = (inp[10]) ? node11367 : node11364;
															assign node11364 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node11367 = (inp[12]) ? 4'b1101 : node11368;
																assign node11368 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node11372 = (inp[7]) ? node11388 : node11373;
													assign node11373 = (inp[4]) ? node11379 : node11374;
														assign node11374 = (inp[12]) ? node11376 : 4'b1100;
															assign node11376 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node11379 = (inp[10]) ? node11383 : node11380;
															assign node11380 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11383 = (inp[12]) ? 4'b1000 : node11384;
																assign node11384 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node11388 = (inp[12]) ? node11390 : 4'b1100;
														assign node11390 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node11393 = (inp[12]) ? node11453 : node11394;
											assign node11394 = (inp[3]) ? node11414 : node11395;
												assign node11395 = (inp[2]) ? node11409 : node11396;
													assign node11396 = (inp[4]) ? node11400 : node11397;
														assign node11397 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11400 = (inp[7]) ? 4'b0100 : node11401;
															assign node11401 = (inp[11]) ? node11405 : node11402;
																assign node11402 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node11405 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node11409 = (inp[4]) ? 4'b0100 : node11410;
														assign node11410 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node11414 = (inp[4]) ? node11430 : node11415;
													assign node11415 = (inp[2]) ? node11427 : node11416;
														assign node11416 = (inp[10]) ? node11424 : node11417;
															assign node11417 = (inp[11]) ? node11421 : node11418;
																assign node11418 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node11421 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node11424 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node11427 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node11430 = (inp[7]) ? node11444 : node11431;
														assign node11431 = (inp[11]) ? node11439 : node11432;
															assign node11432 = (inp[2]) ? node11436 : node11433;
																assign node11433 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node11436 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node11439 = (inp[2]) ? node11441 : 4'b0000;
																assign node11441 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node11444 = (inp[10]) ? node11448 : node11445;
															assign node11445 = (inp[2]) ? 4'b0000 : 4'b1100;
															assign node11448 = (inp[2]) ? node11450 : 4'b0000;
																assign node11450 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node11453 = (inp[11]) ? node11503 : node11454;
												assign node11454 = (inp[10]) ? node11478 : node11455;
													assign node11455 = (inp[3]) ? node11465 : node11456;
														assign node11456 = (inp[7]) ? 4'b1000 : node11457;
															assign node11457 = (inp[2]) ? node11461 : node11458;
																assign node11458 = (inp[4]) ? 4'b0000 : 4'b1000;
																assign node11461 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node11465 = (inp[2]) ? node11473 : node11466;
															assign node11466 = (inp[7]) ? node11470 : node11467;
																assign node11467 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node11470 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node11473 = (inp[4]) ? node11475 : 4'b1100;
																assign node11475 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node11478 = (inp[3]) ? node11488 : node11479;
														assign node11479 = (inp[7]) ? node11485 : node11480;
															assign node11480 = (inp[4]) ? node11482 : 4'b0100;
																assign node11482 = (inp[2]) ? 4'b0100 : 4'b1000;
															assign node11485 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node11488 = (inp[2]) ? node11496 : node11489;
															assign node11489 = (inp[4]) ? node11493 : node11490;
																assign node11490 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node11493 = (inp[7]) ? 4'b1100 : 4'b1001;
															assign node11496 = (inp[7]) ? node11500 : node11497;
																assign node11497 = (inp[4]) ? 4'b1000 : 4'b0000;
																assign node11500 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node11503 = (inp[3]) ? node11519 : node11504;
													assign node11504 = (inp[10]) ? node11512 : node11505;
														assign node11505 = (inp[4]) ? node11507 : 4'b1000;
															assign node11507 = (inp[7]) ? 4'b1000 : node11508;
																assign node11508 = (inp[2]) ? 4'b1100 : 4'b0001;
														assign node11512 = (inp[7]) ? node11516 : node11513;
															assign node11513 = (inp[4]) ? 4'b1001 : 4'b0100;
															assign node11516 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node11519 = (inp[2]) ? node11535 : node11520;
														assign node11520 = (inp[10]) ? node11528 : node11521;
															assign node11521 = (inp[7]) ? node11525 : node11522;
																assign node11522 = (inp[4]) ? 4'b0000 : 4'b0101;
																assign node11525 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node11528 = (inp[4]) ? node11532 : node11529;
																assign node11529 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node11532 = (inp[7]) ? 4'b1101 : 4'b1000;
														assign node11535 = (inp[7]) ? node11541 : node11536;
															assign node11536 = (inp[4]) ? node11538 : 4'b0000;
																assign node11538 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node11541 = (inp[10]) ? node11543 : 4'b1100;
																assign node11543 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node11546 = (inp[11]) ? node11684 : node11547;
										assign node11547 = (inp[3]) ? node11599 : node11548;
											assign node11548 = (inp[13]) ? node11564 : node11549;
												assign node11549 = (inp[12]) ? node11559 : node11550;
													assign node11550 = (inp[10]) ? node11552 : 4'b0001;
														assign node11552 = (inp[7]) ? 4'b1001 : node11553;
															assign node11553 = (inp[2]) ? node11555 : 4'b0000;
																assign node11555 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node11559 = (inp[7]) ? 4'b0001 : node11560;
														assign node11560 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node11564 = (inp[2]) ? node11584 : node11565;
													assign node11565 = (inp[4]) ? node11571 : node11566;
														assign node11566 = (inp[10]) ? node11568 : 4'b1001;
															assign node11568 = (inp[7]) ? 4'b1001 : 4'b0101;
														assign node11571 = (inp[7]) ? node11579 : node11572;
															assign node11572 = (inp[10]) ? node11576 : node11573;
																assign node11573 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node11576 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node11579 = (inp[10]) ? node11581 : 4'b1001;
																assign node11581 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node11584 = (inp[12]) ? node11594 : node11585;
														assign node11585 = (inp[10]) ? node11589 : node11586;
															assign node11586 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node11589 = (inp[4]) ? 4'b0101 : node11590;
																assign node11590 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node11594 = (inp[7]) ? 4'b1001 : node11595;
															assign node11595 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node11599 = (inp[2]) ? node11645 : node11600;
												assign node11600 = (inp[4]) ? node11626 : node11601;
													assign node11601 = (inp[7]) ? node11617 : node11602;
														assign node11602 = (inp[13]) ? node11610 : node11603;
															assign node11603 = (inp[10]) ? node11607 : node11604;
																assign node11604 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node11607 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node11610 = (inp[10]) ? node11614 : node11611;
																assign node11611 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node11614 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node11617 = (inp[10]) ? node11621 : node11618;
															assign node11618 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11621 = (inp[12]) ? 4'b1000 : node11622;
																assign node11622 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node11626 = (inp[7]) ? node11638 : node11627;
														assign node11627 = (inp[13]) ? node11635 : node11628;
															assign node11628 = (inp[12]) ? node11632 : node11629;
																assign node11629 = (inp[10]) ? 4'b0000 : 4'b1100;
																assign node11632 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node11635 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node11638 = (inp[10]) ? node11642 : node11639;
															assign node11639 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node11642 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node11645 = (inp[4]) ? node11659 : node11646;
													assign node11646 = (inp[13]) ? node11652 : node11647;
														assign node11647 = (inp[12]) ? 4'b0101 : node11648;
															assign node11648 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node11652 = (inp[10]) ? node11654 : 4'b1101;
															assign node11654 = (inp[12]) ? 4'b1101 : node11655;
																assign node11655 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node11659 = (inp[7]) ? node11673 : node11660;
														assign node11660 = (inp[13]) ? node11666 : node11661;
															assign node11661 = (inp[10]) ? node11663 : 4'b0001;
																assign node11663 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node11666 = (inp[12]) ? node11670 : node11667;
																assign node11667 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node11670 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node11673 = (inp[13]) ? node11679 : node11674;
															assign node11674 = (inp[12]) ? 4'b0101 : node11675;
																assign node11675 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node11679 = (inp[12]) ? 4'b1101 : node11680;
																assign node11680 = (inp[10]) ? 4'b0000 : 4'b1101;
										assign node11684 = (inp[3]) ? node11738 : node11685;
											assign node11685 = (inp[13]) ? node11707 : node11686;
												assign node11686 = (inp[12]) ? node11696 : node11687;
													assign node11687 = (inp[4]) ? node11689 : 4'b1000;
														assign node11689 = (inp[7]) ? 4'b1000 : node11690;
															assign node11690 = (inp[2]) ? 4'b1100 : node11691;
																assign node11691 = (inp[10]) ? 4'b0001 : 4'b1100;
													assign node11696 = (inp[10]) ? node11702 : node11697;
														assign node11697 = (inp[4]) ? node11699 : 4'b0000;
															assign node11699 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11702 = (inp[4]) ? node11704 : 4'b1000;
															assign node11704 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node11707 = (inp[2]) ? node11727 : node11708;
													assign node11708 = (inp[4]) ? node11716 : node11709;
														assign node11709 = (inp[7]) ? node11711 : 4'b0100;
															assign node11711 = (inp[10]) ? 4'b0000 : node11712;
																assign node11712 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node11716 = (inp[7]) ? node11724 : node11717;
															assign node11717 = (inp[12]) ? node11721 : node11718;
																assign node11718 = (inp[10]) ? 4'b0001 : 4'b1001;
																assign node11721 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node11724 = (inp[10]) ? 4'b0100 : 4'b1000;
													assign node11727 = (inp[12]) ? node11733 : node11728;
														assign node11728 = (inp[7]) ? node11730 : 4'b0100;
															assign node11730 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node11733 = (inp[10]) ? 4'b0100 : node11734;
															assign node11734 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node11738 = (inp[2]) ? node11784 : node11739;
												assign node11739 = (inp[4]) ? node11761 : node11740;
													assign node11740 = (inp[7]) ? node11752 : node11741;
														assign node11741 = (inp[13]) ? node11745 : node11742;
															assign node11742 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node11745 = (inp[12]) ? node11749 : node11746;
																assign node11746 = (inp[10]) ? 4'b0101 : 4'b1101;
																assign node11749 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node11752 = (inp[10]) ? node11756 : node11753;
															assign node11753 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11756 = (inp[12]) ? 4'b1001 : node11757;
																assign node11757 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node11761 = (inp[13]) ? node11771 : node11762;
														assign node11762 = (inp[12]) ? node11768 : node11763;
															assign node11763 = (inp[7]) ? node11765 : 4'b0001;
																assign node11765 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node11768 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node11771 = (inp[7]) ? node11777 : node11772;
															assign node11772 = (inp[10]) ? node11774 : 4'b0000;
																assign node11774 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node11777 = (inp[12]) ? node11781 : node11778;
																assign node11778 = (inp[10]) ? 4'b0000 : 4'b1101;
																assign node11781 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node11784 = (inp[13]) ? node11798 : node11785;
													assign node11785 = (inp[7]) ? node11793 : node11786;
														assign node11786 = (inp[4]) ? node11790 : node11787;
															assign node11787 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node11790 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node11793 = (inp[10]) ? 4'b1100 : node11794;
															assign node11794 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node11798 = (inp[4]) ? node11806 : node11799;
														assign node11799 = (inp[12]) ? node11801 : 4'b0000;
															assign node11801 = (inp[10]) ? node11803 : 4'b1100;
																assign node11803 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node11806 = (inp[7]) ? node11812 : node11807;
															assign node11807 = (inp[10]) ? 4'b1001 : node11808;
																assign node11808 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node11812 = (inp[10]) ? node11816 : node11813;
																assign node11813 = (inp[12]) ? 4'b1100 : 4'b0000;
																assign node11816 = (inp[12]) ? 4'b0000 : 4'b0001;
								assign node11819 = (inp[3]) ? node12037 : node11820;
									assign node11820 = (inp[4]) ? node11930 : node11821;
										assign node11821 = (inp[13]) ? node11875 : node11822;
											assign node11822 = (inp[10]) ? node11842 : node11823;
												assign node11823 = (inp[12]) ? node11833 : node11824;
													assign node11824 = (inp[11]) ? node11830 : node11825;
														assign node11825 = (inp[14]) ? 4'b1000 : node11826;
															assign node11826 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node11830 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node11833 = (inp[2]) ? node11839 : node11834;
														assign node11834 = (inp[11]) ? 4'b1000 : node11835;
															assign node11835 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11839 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node11842 = (inp[7]) ? node11858 : node11843;
													assign node11843 = (inp[2]) ? node11851 : node11844;
														assign node11844 = (inp[11]) ? node11848 : node11845;
															assign node11845 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node11848 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node11851 = (inp[12]) ? node11855 : node11852;
															assign node11852 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node11855 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node11858 = (inp[11]) ? node11868 : node11859;
														assign node11859 = (inp[12]) ? node11865 : node11860;
															assign node11860 = (inp[2]) ? 4'b0000 : node11861;
																assign node11861 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11865 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node11868 = (inp[2]) ? node11872 : node11869;
															assign node11869 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node11872 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node11875 = (inp[10]) ? node11901 : node11876;
												assign node11876 = (inp[2]) ? node11886 : node11877;
													assign node11877 = (inp[11]) ? 4'b0100 : node11878;
														assign node11878 = (inp[12]) ? node11882 : node11879;
															assign node11879 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node11882 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node11886 = (inp[11]) ? node11894 : node11887;
														assign node11887 = (inp[12]) ? node11891 : node11888;
															assign node11888 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node11891 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node11894 = (inp[7]) ? node11898 : node11895;
															assign node11895 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node11898 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node11901 = (inp[12]) ? node11913 : node11902;
													assign node11902 = (inp[2]) ? node11908 : node11903;
														assign node11903 = (inp[7]) ? node11905 : 4'b1001;
															assign node11905 = (inp[11]) ? 4'b0100 : 4'b1101;
														assign node11908 = (inp[11]) ? node11910 : 4'b0100;
															assign node11910 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node11913 = (inp[7]) ? node11921 : node11914;
														assign node11914 = (inp[2]) ? node11918 : node11915;
															assign node11915 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node11918 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node11921 = (inp[2]) ? node11927 : node11922;
															assign node11922 = (inp[14]) ? 4'b1100 : node11923;
																assign node11923 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node11927 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node11930 = (inp[2]) ? node11984 : node11931;
											assign node11931 = (inp[13]) ? node11953 : node11932;
												assign node11932 = (inp[11]) ? node11948 : node11933;
													assign node11933 = (inp[12]) ? node11943 : node11934;
														assign node11934 = (inp[14]) ? node11940 : node11935;
															assign node11935 = (inp[7]) ? 4'b1001 : node11936;
																assign node11936 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node11940 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node11943 = (inp[7]) ? 4'b0001 : node11944;
															assign node11944 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node11948 = (inp[7]) ? 4'b1001 : node11949;
														assign node11949 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node11953 = (inp[11]) ? node11971 : node11954;
													assign node11954 = (inp[14]) ? node11962 : node11955;
														assign node11955 = (inp[12]) ? 4'b0000 : node11956;
															assign node11956 = (inp[10]) ? node11958 : 4'b0000;
																assign node11958 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node11962 = (inp[7]) ? node11966 : node11963;
															assign node11963 = (inp[10]) ? 4'b0000 : 4'b1001;
															assign node11966 = (inp[10]) ? 4'b0001 : node11967;
																assign node11967 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node11971 = (inp[12]) ? node11977 : node11972;
														assign node11972 = (inp[10]) ? node11974 : 4'b1000;
															assign node11974 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node11977 = (inp[7]) ? node11981 : node11978;
															assign node11978 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node11981 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node11984 = (inp[10]) ? node12018 : node11985;
												assign node11985 = (inp[13]) ? node12001 : node11986;
													assign node11986 = (inp[7]) ? node11994 : node11987;
														assign node11987 = (inp[11]) ? 4'b1000 : node11988;
															assign node11988 = (inp[12]) ? 4'b0000 : node11989;
																assign node11989 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11994 = (inp[12]) ? node11998 : node11995;
															assign node11995 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node11998 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node12001 = (inp[7]) ? node12009 : node12002;
														assign node12002 = (inp[12]) ? node12006 : node12003;
															assign node12003 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node12006 = (inp[11]) ? 4'b0100 : 4'b1001;
														assign node12009 = (inp[11]) ? 4'b0000 : node12010;
															assign node12010 = (inp[14]) ? node12014 : node12011;
																assign node12011 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node12014 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node12018 = (inp[13]) ? node12024 : node12019;
													assign node12019 = (inp[12]) ? 4'b0000 : node12020;
														assign node12020 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node12024 = (inp[7]) ? node12030 : node12025;
														assign node12025 = (inp[12]) ? node12027 : 4'b1001;
															assign node12027 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node12030 = (inp[11]) ? node12034 : node12031;
															assign node12031 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node12034 = (inp[12]) ? 4'b1000 : 4'b0100;
									assign node12037 = (inp[4]) ? node12171 : node12038;
										assign node12038 = (inp[10]) ? node12104 : node12039;
											assign node12039 = (inp[11]) ? node12077 : node12040;
												assign node12040 = (inp[12]) ? node12060 : node12041;
													assign node12041 = (inp[7]) ? node12055 : node12042;
														assign node12042 = (inp[14]) ? node12048 : node12043;
															assign node12043 = (inp[2]) ? node12045 : 4'b1000;
																assign node12045 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node12048 = (inp[2]) ? node12052 : node12049;
																assign node12049 = (inp[13]) ? 4'b0001 : 4'b1000;
																assign node12052 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node12055 = (inp[2]) ? 4'b1001 : node12056;
															assign node12056 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node12060 = (inp[2]) ? node12068 : node12061;
														assign node12061 = (inp[13]) ? node12063 : 4'b1000;
															assign node12063 = (inp[7]) ? 4'b1001 : node12064;
																assign node12064 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node12068 = (inp[13]) ? node12070 : 4'b0001;
															assign node12070 = (inp[14]) ? node12074 : node12071;
																assign node12071 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node12074 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node12077 = (inp[12]) ? node12091 : node12078;
													assign node12078 = (inp[7]) ? node12084 : node12079;
														assign node12079 = (inp[13]) ? node12081 : 4'b0000;
															assign node12081 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node12084 = (inp[13]) ? node12088 : node12085;
															assign node12085 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node12088 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node12091 = (inp[2]) ? node12099 : node12092;
														assign node12092 = (inp[7]) ? node12096 : node12093;
															assign node12093 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node12096 = (inp[13]) ? 4'b0001 : 4'b1001;
														assign node12099 = (inp[7]) ? node12101 : 4'b1001;
															assign node12101 = (inp[14]) ? 4'b0000 : 4'b1001;
											assign node12104 = (inp[7]) ? node12138 : node12105;
												assign node12105 = (inp[11]) ? node12129 : node12106;
													assign node12106 = (inp[14]) ? node12118 : node12107;
														assign node12107 = (inp[13]) ? node12113 : node12108;
															assign node12108 = (inp[2]) ? node12110 : 4'b1001;
																assign node12110 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node12113 = (inp[12]) ? node12115 : 4'b0001;
																assign node12115 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node12118 = (inp[13]) ? node12124 : node12119;
															assign node12119 = (inp[2]) ? 4'b1001 : node12120;
																assign node12120 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node12124 = (inp[2]) ? node12126 : 4'b0000;
																assign node12126 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node12129 = (inp[2]) ? node12135 : node12130;
														assign node12130 = (inp[13]) ? node12132 : 4'b0001;
															assign node12132 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node12135 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node12138 = (inp[12]) ? node12156 : node12139;
													assign node12139 = (inp[11]) ? node12151 : node12140;
														assign node12140 = (inp[2]) ? node12144 : node12141;
															assign node12141 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node12144 = (inp[14]) ? node12148 : node12145;
																assign node12145 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node12148 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node12151 = (inp[2]) ? node12153 : 4'b0000;
															assign node12153 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node12156 = (inp[2]) ? node12166 : node12157;
														assign node12157 = (inp[11]) ? node12163 : node12158;
															assign node12158 = (inp[14]) ? 4'b0000 : node12159;
																assign node12159 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node12163 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node12166 = (inp[13]) ? 4'b0000 : node12167;
															assign node12167 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node12171 = (inp[13]) ? node12231 : node12172;
											assign node12172 = (inp[2]) ? node12196 : node12173;
												assign node12173 = (inp[7]) ? node12181 : node12174;
													assign node12174 = (inp[10]) ? node12176 : 4'b0000;
														assign node12176 = (inp[14]) ? 4'b0000 : node12177;
															assign node12177 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node12181 = (inp[12]) ? node12185 : node12182;
														assign node12182 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node12185 = (inp[10]) ? node12193 : node12186;
															assign node12186 = (inp[14]) ? node12190 : node12187;
																assign node12187 = (inp[11]) ? 4'b1000 : 4'b0000;
																assign node12190 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node12193 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node12196 = (inp[7]) ? node12216 : node12197;
													assign node12197 = (inp[11]) ? node12211 : node12198;
														assign node12198 = (inp[14]) ? node12206 : node12199;
															assign node12199 = (inp[12]) ? node12203 : node12200;
																assign node12200 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node12203 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node12206 = (inp[12]) ? 4'b1001 : node12207;
																assign node12207 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node12211 = (inp[12]) ? 4'b0001 : node12212;
															assign node12212 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node12216 = (inp[11]) ? node12226 : node12217;
														assign node12217 = (inp[12]) ? node12223 : node12218;
															assign node12218 = (inp[10]) ? 4'b0001 : node12219;
																assign node12219 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node12223 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12226 = (inp[10]) ? 4'b0000 : node12227;
															assign node12227 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node12231 = (inp[10]) ? node12265 : node12232;
												assign node12232 = (inp[7]) ? node12246 : node12233;
													assign node12233 = (inp[2]) ? node12235 : 4'b0000;
														assign node12235 = (inp[12]) ? node12241 : node12236;
															assign node12236 = (inp[14]) ? node12238 : 4'b0000;
																assign node12238 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node12241 = (inp[11]) ? 4'b0001 : node12242;
																assign node12242 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node12246 = (inp[14]) ? node12252 : node12247;
														assign node12247 = (inp[2]) ? node12249 : 4'b0001;
															assign node12249 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node12252 = (inp[11]) ? node12258 : node12253;
															assign node12253 = (inp[2]) ? 4'b0000 : node12254;
																assign node12254 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node12258 = (inp[12]) ? node12262 : node12259;
																assign node12259 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node12262 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node12265 = (inp[11]) ? 4'b0000 : node12266;
													assign node12266 = (inp[14]) ? node12278 : node12267;
														assign node12267 = (inp[12]) ? node12273 : node12268;
															assign node12268 = (inp[7]) ? 4'b0000 : node12269;
																assign node12269 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node12273 = (inp[7]) ? node12275 : 4'b0000;
																assign node12275 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node12278 = (inp[2]) ? node12284 : node12279;
															assign node12279 = (inp[12]) ? node12281 : 4'b0000;
																assign node12281 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node12284 = (inp[7]) ? node12286 : 4'b0001;
																assign node12286 = (inp[12]) ? 4'b0000 : 4'b0001;
							assign node12290 = (inp[11]) ? node12778 : node12291;
								assign node12291 = (inp[5]) ? node12537 : node12292;
									assign node12292 = (inp[14]) ? node12416 : node12293;
										assign node12293 = (inp[2]) ? node12351 : node12294;
											assign node12294 = (inp[3]) ? node12326 : node12295;
												assign node12295 = (inp[4]) ? node12311 : node12296;
													assign node12296 = (inp[13]) ? node12302 : node12297;
														assign node12297 = (inp[10]) ? 4'b1001 : node12298;
															assign node12298 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12302 = (inp[7]) ? node12308 : node12303;
															assign node12303 = (inp[10]) ? 4'b0101 : node12304;
																assign node12304 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node12308 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12311 = (inp[10]) ? node12321 : node12312;
														assign node12312 = (inp[7]) ? node12316 : node12313;
															assign node12313 = (inp[13]) ? 4'b1000 : 4'b1101;
															assign node12316 = (inp[13]) ? 4'b0101 : node12317;
																assign node12317 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12321 = (inp[13]) ? 4'b0000 : node12322;
															assign node12322 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node12326 = (inp[10]) ? node12340 : node12327;
													assign node12327 = (inp[4]) ? node12333 : node12328;
														assign node12328 = (inp[7]) ? 4'b1000 : node12329;
															assign node12329 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node12333 = (inp[7]) ? 4'b1100 : node12334;
															assign node12334 = (inp[13]) ? node12336 : 4'b1100;
																assign node12336 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12340 = (inp[4]) ? node12346 : node12341;
														assign node12341 = (inp[7]) ? node12343 : 4'b0100;
															assign node12343 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node12346 = (inp[13]) ? 4'b0000 : node12347;
															assign node12347 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node12351 = (inp[13]) ? node12383 : node12352;
												assign node12352 = (inp[12]) ? node12364 : node12353;
													assign node12353 = (inp[3]) ? node12359 : node12354;
														assign node12354 = (inp[4]) ? node12356 : 4'b1001;
															assign node12356 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node12359 = (inp[4]) ? node12361 : 4'b1101;
															assign node12361 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node12364 = (inp[10]) ? node12374 : node12365;
														assign node12365 = (inp[3]) ? node12369 : node12366;
															assign node12366 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12369 = (inp[4]) ? node12371 : 4'b0101;
																assign node12371 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12374 = (inp[4]) ? node12376 : 4'b1101;
															assign node12376 = (inp[3]) ? node12380 : node12377;
																assign node12377 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node12380 = (inp[7]) ? 4'b1101 : 4'b0000;
												assign node12383 = (inp[10]) ? node12405 : node12384;
													assign node12384 = (inp[12]) ? node12396 : node12385;
														assign node12385 = (inp[3]) ? node12391 : node12386;
															assign node12386 = (inp[4]) ? 4'b0101 : node12387;
																assign node12387 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12391 = (inp[4]) ? 4'b1000 : node12392;
																assign node12392 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12396 = (inp[3]) ? node12400 : node12397;
															assign node12397 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node12400 = (inp[7]) ? 4'b1101 : node12401;
																assign node12401 = (inp[4]) ? 4'b1000 : 4'b1101;
													assign node12405 = (inp[4]) ? node12413 : node12406;
														assign node12406 = (inp[3]) ? node12410 : node12407;
															assign node12407 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12410 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12413 = (inp[3]) ? 4'b0000 : 4'b0101;
										assign node12416 = (inp[13]) ? node12472 : node12417;
											assign node12417 = (inp[3]) ? node12441 : node12418;
												assign node12418 = (inp[12]) ? node12428 : node12419;
													assign node12419 = (inp[4]) ? node12421 : 4'b1000;
														assign node12421 = (inp[7]) ? 4'b1000 : node12422;
															assign node12422 = (inp[2]) ? 4'b1100 : node12423;
																assign node12423 = (inp[10]) ? 4'b0000 : 4'b1100;
													assign node12428 = (inp[10]) ? node12434 : node12429;
														assign node12429 = (inp[7]) ? 4'b0000 : node12430;
															assign node12430 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node12434 = (inp[4]) ? node12436 : 4'b1000;
															assign node12436 = (inp[2]) ? 4'b1100 : node12437;
																assign node12437 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node12441 = (inp[7]) ? node12457 : node12442;
													assign node12442 = (inp[4]) ? node12450 : node12443;
														assign node12443 = (inp[10]) ? node12447 : node12444;
															assign node12444 = (inp[2]) ? 4'b0100 : 4'b1000;
															assign node12447 = (inp[2]) ? 4'b1100 : 4'b0100;
														assign node12450 = (inp[10]) ? 4'b0000 : node12451;
															assign node12451 = (inp[2]) ? node12453 : 4'b1100;
																assign node12453 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12457 = (inp[12]) ? node12465 : node12458;
														assign node12458 = (inp[2]) ? 4'b1100 : node12459;
															assign node12459 = (inp[4]) ? node12461 : 4'b1000;
																assign node12461 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node12465 = (inp[10]) ? node12469 : node12466;
															assign node12466 = (inp[2]) ? 4'b0100 : 4'b1100;
															assign node12469 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node12472 = (inp[10]) ? node12518 : node12473;
												assign node12473 = (inp[12]) ? node12499 : node12474;
													assign node12474 = (inp[3]) ? node12484 : node12475;
														assign node12475 = (inp[4]) ? node12479 : node12476;
															assign node12476 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node12479 = (inp[2]) ? 4'b0100 : node12480;
																assign node12480 = (inp[7]) ? 4'b0100 : 4'b1000;
														assign node12484 = (inp[2]) ? node12492 : node12485;
															assign node12485 = (inp[7]) ? node12489 : node12486;
																assign node12486 = (inp[4]) ? 4'b0001 : 4'b1100;
																assign node12489 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node12492 = (inp[4]) ? node12496 : node12493;
																assign node12493 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node12496 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node12499 = (inp[3]) ? node12507 : node12500;
														assign node12500 = (inp[7]) ? 4'b1000 : node12501;
															assign node12501 = (inp[2]) ? node12503 : 4'b1000;
																assign node12503 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node12507 = (inp[7]) ? node12513 : node12508;
															assign node12508 = (inp[4]) ? node12510 : 4'b1100;
																assign node12510 = (inp[2]) ? 4'b1000 : 4'b0001;
															assign node12513 = (inp[2]) ? 4'b1100 : node12514;
																assign node12514 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node12518 = (inp[4]) ? node12528 : node12519;
													assign node12519 = (inp[3]) ? node12523 : node12520;
														assign node12520 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node12523 = (inp[7]) ? 4'b0100 : node12524;
															assign node12524 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node12528 = (inp[2]) ? node12534 : node12529;
														assign node12529 = (inp[3]) ? node12531 : 4'b0000;
															assign node12531 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node12534 = (inp[3]) ? 4'b0000 : 4'b0100;
									assign node12537 = (inp[3]) ? node12659 : node12538;
										assign node12538 = (inp[2]) ? node12606 : node12539;
											assign node12539 = (inp[12]) ? node12573 : node12540;
												assign node12540 = (inp[13]) ? node12562 : node12541;
													assign node12541 = (inp[4]) ? node12555 : node12542;
														assign node12542 = (inp[14]) ? node12550 : node12543;
															assign node12543 = (inp[10]) ? node12547 : node12544;
																assign node12544 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node12547 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node12550 = (inp[7]) ? 4'b1001 : node12551;
																assign node12551 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node12555 = (inp[10]) ? node12559 : node12556;
															assign node12556 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12559 = (inp[7]) ? 4'b0101 : 4'b1000;
													assign node12562 = (inp[4]) ? node12568 : node12563;
														assign node12563 = (inp[10]) ? 4'b0001 : node12564;
															assign node12564 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node12568 = (inp[10]) ? 4'b0000 : node12569;
															assign node12569 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node12573 = (inp[4]) ? node12597 : node12574;
													assign node12574 = (inp[14]) ? node12586 : node12575;
														assign node12575 = (inp[13]) ? node12581 : node12576;
															assign node12576 = (inp[7]) ? 4'b1000 : node12577;
																assign node12577 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node12581 = (inp[7]) ? 4'b0100 : node12582;
																assign node12582 = (inp[10]) ? 4'b1001 : 4'b0100;
														assign node12586 = (inp[13]) ? node12592 : node12587;
															assign node12587 = (inp[10]) ? node12589 : 4'b1001;
																assign node12589 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12592 = (inp[10]) ? node12594 : 4'b0101;
																assign node12594 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node12597 = (inp[13]) ? node12603 : node12598;
														assign node12598 = (inp[10]) ? node12600 : 4'b1001;
															assign node12600 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node12603 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node12606 = (inp[4]) ? node12622 : node12607;
												assign node12607 = (inp[10]) ? node12613 : node12608;
													assign node12608 = (inp[7]) ? 4'b1000 : node12609;
														assign node12609 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node12613 = (inp[7]) ? node12619 : node12614;
														assign node12614 = (inp[13]) ? node12616 : 4'b0100;
															assign node12616 = (inp[14]) ? 4'b0100 : 4'b0000;
														assign node12619 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node12622 = (inp[13]) ? node12640 : node12623;
													assign node12623 = (inp[14]) ? node12633 : node12624;
														assign node12624 = (inp[12]) ? node12628 : node12625;
															assign node12625 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node12628 = (inp[10]) ? 4'b1000 : node12629;
																assign node12629 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node12633 = (inp[10]) ? node12637 : node12634;
															assign node12634 = (inp[7]) ? 4'b1100 : 4'b1001;
															assign node12637 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node12640 = (inp[14]) ? node12654 : node12641;
														assign node12641 = (inp[12]) ? node12647 : node12642;
															assign node12642 = (inp[10]) ? 4'b0001 : node12643;
																assign node12643 = (inp[7]) ? 4'b1000 : 4'b0001;
															assign node12647 = (inp[7]) ? node12651 : node12648;
																assign node12648 = (inp[10]) ? 4'b1001 : 4'b0100;
																assign node12651 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node12654 = (inp[12]) ? node12656 : 4'b0001;
															assign node12656 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node12659 = (inp[4]) ? node12727 : node12660;
											assign node12660 = (inp[10]) ? node12694 : node12661;
												assign node12661 = (inp[13]) ? node12679 : node12662;
													assign node12662 = (inp[2]) ? node12672 : node12663;
														assign node12663 = (inp[14]) ? node12665 : 4'b1000;
															assign node12665 = (inp[12]) ? node12669 : node12666;
																assign node12666 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node12669 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node12672 = (inp[7]) ? node12676 : node12673;
															assign node12673 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node12676 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12679 = (inp[12]) ? node12689 : node12680;
														assign node12680 = (inp[7]) ? node12686 : node12681;
															assign node12681 = (inp[2]) ? node12683 : 4'b0000;
																assign node12683 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node12686 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12689 = (inp[2]) ? 4'b0000 : node12690;
															assign node12690 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node12694 = (inp[13]) ? node12710 : node12695;
													assign node12695 = (inp[2]) ? node12703 : node12696;
														assign node12696 = (inp[7]) ? node12698 : 4'b1001;
															assign node12698 = (inp[14]) ? 4'b0001 : node12699;
																assign node12699 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node12703 = (inp[14]) ? node12705 : 4'b0001;
															assign node12705 = (inp[7]) ? node12707 : 4'b0000;
																assign node12707 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node12710 = (inp[14]) ? node12722 : node12711;
														assign node12711 = (inp[7]) ? node12717 : node12712;
															assign node12712 = (inp[2]) ? 4'b1001 : node12713;
																assign node12713 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node12717 = (inp[12]) ? 4'b1000 : node12718;
																assign node12718 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node12722 = (inp[2]) ? 4'b1001 : node12723;
															assign node12723 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node12727 = (inp[13]) ? node12761 : node12728;
												assign node12728 = (inp[7]) ? node12740 : node12729;
													assign node12729 = (inp[14]) ? 4'b0001 : node12730;
														assign node12730 = (inp[2]) ? node12736 : node12731;
															assign node12731 = (inp[10]) ? node12733 : 4'b0001;
																assign node12733 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node12736 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node12740 = (inp[2]) ? node12754 : node12741;
														assign node12741 = (inp[14]) ? node12747 : node12742;
															assign node12742 = (inp[10]) ? node12744 : 4'b0000;
																assign node12744 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node12747 = (inp[12]) ? node12751 : node12748;
																assign node12748 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node12751 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node12754 = (inp[10]) ? node12756 : 4'b0000;
															assign node12756 = (inp[12]) ? 4'b0000 : node12757;
																assign node12757 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node12761 = (inp[10]) ? 4'b0000 : node12762;
													assign node12762 = (inp[2]) ? node12770 : node12763;
														assign node12763 = (inp[14]) ? node12765 : 4'b0000;
															assign node12765 = (inp[12]) ? 4'b0000 : node12766;
																assign node12766 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node12770 = (inp[7]) ? 4'b0000 : node12771;
															assign node12771 = (inp[14]) ? 4'b0000 : node12772;
																assign node12772 = (inp[12]) ? 4'b0001 : 4'b0000;
								assign node12778 = (inp[5]) ? node12940 : node12779;
									assign node12779 = (inp[10]) ? node12881 : node12780;
										assign node12780 = (inp[3]) ? node12830 : node12781;
											assign node12781 = (inp[7]) ? node12799 : node12782;
												assign node12782 = (inp[4]) ? node12790 : node12783;
													assign node12783 = (inp[13]) ? node12787 : node12784;
														assign node12784 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12787 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node12790 = (inp[13]) ? node12794 : node12791;
														assign node12791 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node12794 = (inp[2]) ? node12796 : 4'b1001;
															assign node12796 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node12799 = (inp[4]) ? node12823 : node12800;
													assign node12800 = (inp[2]) ? node12808 : node12801;
														assign node12801 = (inp[13]) ? node12805 : node12802;
															assign node12802 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node12805 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node12808 = (inp[14]) ? node12816 : node12809;
															assign node12809 = (inp[12]) ? node12813 : node12810;
																assign node12810 = (inp[13]) ? 4'b0001 : 4'b1001;
																assign node12813 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node12816 = (inp[13]) ? node12820 : node12817;
																assign node12817 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node12820 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node12823 = (inp[12]) ? node12827 : node12824;
														assign node12824 = (inp[13]) ? 4'b0101 : 4'b1001;
														assign node12827 = (inp[13]) ? 4'b1001 : 4'b0001;
											assign node12830 = (inp[2]) ? node12844 : node12831;
												assign node12831 = (inp[4]) ? node12837 : node12832;
													assign node12832 = (inp[13]) ? node12834 : 4'b1001;
														assign node12834 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node12837 = (inp[13]) ? node12839 : 4'b1101;
														assign node12839 = (inp[7]) ? 4'b1101 : node12840;
															assign node12840 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node12844 = (inp[4]) ? node12868 : node12845;
													assign node12845 = (inp[7]) ? node12853 : node12846;
														assign node12846 = (inp[13]) ? node12850 : node12847;
															assign node12847 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node12850 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node12853 = (inp[14]) ? node12861 : node12854;
															assign node12854 = (inp[12]) ? node12858 : node12855;
																assign node12855 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node12858 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node12861 = (inp[12]) ? node12865 : node12862;
																assign node12862 = (inp[13]) ? 4'b0101 : 4'b1101;
																assign node12865 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node12868 = (inp[7]) ? node12874 : node12869;
														assign node12869 = (inp[13]) ? 4'b1001 : node12870;
															assign node12870 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node12874 = (inp[12]) ? node12878 : node12875;
															assign node12875 = (inp[13]) ? 4'b0001 : 4'b1101;
															assign node12878 = (inp[13]) ? 4'b1101 : 4'b0101;
										assign node12881 = (inp[13]) ? node12925 : node12882;
											assign node12882 = (inp[3]) ? node12892 : node12883;
												assign node12883 = (inp[4]) ? node12885 : 4'b1001;
													assign node12885 = (inp[2]) ? node12889 : node12886;
														assign node12886 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node12889 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node12892 = (inp[2]) ? node12920 : node12893;
													assign node12893 = (inp[12]) ? node12907 : node12894;
														assign node12894 = (inp[14]) ? node12902 : node12895;
															assign node12895 = (inp[7]) ? node12899 : node12896;
																assign node12896 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node12899 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node12902 = (inp[7]) ? 4'b0001 : node12903;
																assign node12903 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node12907 = (inp[14]) ? node12913 : node12908;
															assign node12908 = (inp[4]) ? 4'b0101 : node12909;
																assign node12909 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12913 = (inp[7]) ? node12917 : node12914;
																assign node12914 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node12917 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node12920 = (inp[4]) ? node12922 : 4'b1101;
														assign node12922 = (inp[7]) ? 4'b1101 : 4'b0001;
											assign node12925 = (inp[4]) ? node12935 : node12926;
												assign node12926 = (inp[3]) ? node12930 : node12927;
													assign node12927 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node12930 = (inp[7]) ? 4'b0101 : node12931;
														assign node12931 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node12935 = (inp[3]) ? 4'b0001 : node12936;
													assign node12936 = (inp[2]) ? 4'b0101 : 4'b0001;
									assign node12940 = (inp[3]) ? node13022 : node12941;
										assign node12941 = (inp[13]) ? node12993 : node12942;
											assign node12942 = (inp[12]) ? node12970 : node12943;
												assign node12943 = (inp[7]) ? node12957 : node12944;
													assign node12944 = (inp[4]) ? node12952 : node12945;
														assign node12945 = (inp[2]) ? node12949 : node12946;
															assign node12946 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node12949 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node12952 = (inp[10]) ? 4'b1001 : node12953;
															assign node12953 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node12957 = (inp[10]) ? node12963 : node12958;
														assign node12958 = (inp[4]) ? 4'b0001 : node12959;
															assign node12959 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node12963 = (inp[2]) ? node12967 : node12964;
															assign node12964 = (inp[4]) ? 4'b0101 : 4'b1001;
															assign node12967 = (inp[4]) ? 4'b1001 : 4'b0001;
												assign node12970 = (inp[2]) ? node12984 : node12971;
													assign node12971 = (inp[4]) ? node12977 : node12972;
														assign node12972 = (inp[10]) ? node12974 : 4'b1001;
															assign node12974 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node12977 = (inp[10]) ? node12981 : node12978;
															assign node12978 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node12981 = (inp[7]) ? 4'b0101 : 4'b1001;
													assign node12984 = (inp[4]) ? node12988 : node12985;
														assign node12985 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node12988 = (inp[7]) ? node12990 : 4'b1001;
															assign node12990 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node12993 = (inp[10]) ? node13015 : node12994;
												assign node12994 = (inp[4]) ? node13004 : node12995;
													assign node12995 = (inp[2]) ? node13001 : node12996;
														assign node12996 = (inp[7]) ? node12998 : 4'b0001;
															assign node12998 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node13001 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node13004 = (inp[12]) ? node13012 : node13005;
														assign node13005 = (inp[2]) ? node13009 : node13006;
															assign node13006 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node13009 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node13012 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node13015 = (inp[7]) ? node13017 : 4'b0001;
													assign node13017 = (inp[4]) ? 4'b0001 : node13018;
														assign node13018 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node13022 = (inp[4]) ? node13052 : node13023;
											assign node13023 = (inp[10]) ? node13045 : node13024;
												assign node13024 = (inp[13]) ? node13034 : node13025;
													assign node13025 = (inp[2]) ? node13029 : node13026;
														assign node13026 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13029 = (inp[7]) ? 4'b0001 : node13030;
															assign node13030 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13034 = (inp[12]) ? node13040 : node13035;
														assign node13035 = (inp[7]) ? node13037 : 4'b1001;
															assign node13037 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node13040 = (inp[2]) ? node13042 : 4'b1001;
															assign node13042 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node13045 = (inp[2]) ? node13047 : 4'b0001;
													assign node13047 = (inp[13]) ? 4'b0001 : node13048;
														assign node13048 = (inp[7]) ? 4'b1001 : 4'b0001;
											assign node13052 = (inp[10]) ? node13066 : node13053;
												assign node13053 = (inp[13]) ? 4'b0001 : node13054;
													assign node13054 = (inp[12]) ? node13060 : node13055;
														assign node13055 = (inp[2]) ? 4'b0001 : node13056;
															assign node13056 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node13060 = (inp[7]) ? node13062 : 4'b0001;
															assign node13062 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node13066 = (inp[13]) ? 4'b0000 : 4'b0001;
					assign node13069 = (inp[6]) ? node13071 : 4'b0001;
						assign node13071 = (inp[2]) ? node13631 : node13072;
							assign node13072 = (inp[5]) ? node13182 : node13073;
								assign node13073 = (inp[3]) ? node13075 : 4'b0001;
									assign node13075 = (inp[7]) ? node13157 : node13076;
										assign node13076 = (inp[4]) ? node13100 : node13077;
											assign node13077 = (inp[13]) ? node13079 : 4'b0001;
												assign node13079 = (inp[1]) ? node13093 : node13080;
													assign node13080 = (inp[11]) ? node13088 : node13081;
														assign node13081 = (inp[14]) ? 4'b0001 : node13082;
															assign node13082 = (inp[12]) ? node13084 : 4'b0000;
																assign node13084 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node13088 = (inp[10]) ? 4'b0000 : node13089;
															assign node13089 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node13093 = (inp[14]) ? node13095 : 4'b0001;
														assign node13095 = (inp[11]) ? 4'b0001 : node13096;
															assign node13096 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node13100 = (inp[1]) ? node13128 : node13101;
												assign node13101 = (inp[14]) ? node13113 : node13102;
													assign node13102 = (inp[13]) ? node13108 : node13103;
														assign node13103 = (inp[12]) ? node13105 : 4'b1000;
															assign node13105 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node13108 = (inp[12]) ? node13110 : 4'b0000;
															assign node13110 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node13113 = (inp[11]) ? node13117 : node13114;
														assign node13114 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node13117 = (inp[13]) ? node13123 : node13118;
															assign node13118 = (inp[10]) ? 4'b1000 : node13119;
																assign node13119 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13123 = (inp[12]) ? node13125 : 4'b0000;
																assign node13125 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node13128 = (inp[14]) ? node13140 : node13129;
													assign node13129 = (inp[13]) ? node13135 : node13130;
														assign node13130 = (inp[12]) ? node13132 : 4'b1001;
															assign node13132 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13135 = (inp[10]) ? 4'b0001 : node13136;
															assign node13136 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node13140 = (inp[11]) ? node13148 : node13141;
														assign node13141 = (inp[13]) ? 4'b0000 : node13142;
															assign node13142 = (inp[10]) ? 4'b1000 : node13143;
																assign node13143 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13148 = (inp[12]) ? node13150 : 4'b1001;
															assign node13150 = (inp[13]) ? node13154 : node13151;
																assign node13151 = (inp[10]) ? 4'b1001 : 4'b0001;
																assign node13154 = (inp[10]) ? 4'b0001 : 4'b1001;
										assign node13157 = (inp[13]) ? node13159 : 4'b0001;
											assign node13159 = (inp[4]) ? node13161 : 4'b0001;
												assign node13161 = (inp[1]) ? node13175 : node13162;
													assign node13162 = (inp[12]) ? node13168 : node13163;
														assign node13163 = (inp[11]) ? 4'b0000 : node13164;
															assign node13164 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node13168 = (inp[10]) ? node13170 : 4'b0001;
															assign node13170 = (inp[11]) ? 4'b0000 : node13171;
																assign node13171 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node13175 = (inp[14]) ? node13177 : 4'b0001;
														assign node13177 = (inp[12]) ? 4'b0001 : node13178;
															assign node13178 = (inp[11]) ? 4'b0001 : 4'b0000;
								assign node13182 = (inp[1]) ? node13428 : node13183;
									assign node13183 = (inp[3]) ? node13309 : node13184;
										assign node13184 = (inp[14]) ? node13236 : node13185;
											assign node13185 = (inp[13]) ? node13205 : node13186;
												assign node13186 = (inp[10]) ? node13198 : node13187;
													assign node13187 = (inp[12]) ? node13193 : node13188;
														assign node13188 = (inp[4]) ? node13190 : 4'b1000;
															assign node13190 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node13193 = (inp[4]) ? node13195 : 4'b0000;
															assign node13195 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node13198 = (inp[7]) ? 4'b1000 : node13199;
														assign node13199 = (inp[4]) ? node13201 : 4'b1000;
															assign node13201 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node13205 = (inp[10]) ? node13223 : node13206;
													assign node13206 = (inp[12]) ? node13216 : node13207;
														assign node13207 = (inp[7]) ? node13213 : node13208;
															assign node13208 = (inp[4]) ? node13210 : 4'b0100;
																assign node13210 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13213 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node13216 = (inp[4]) ? node13218 : 4'b1000;
															assign node13218 = (inp[7]) ? 4'b1000 : node13219;
																assign node13219 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node13223 = (inp[4]) ? node13227 : node13224;
														assign node13224 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node13227 = (inp[12]) ? node13231 : node13228;
															assign node13228 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node13231 = (inp[7]) ? 4'b0100 : node13232;
																assign node13232 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node13236 = (inp[11]) ? node13270 : node13237;
												assign node13237 = (inp[13]) ? node13251 : node13238;
													assign node13238 = (inp[10]) ? node13244 : node13239;
														assign node13239 = (inp[4]) ? node13241 : 4'b0001;
															assign node13241 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node13244 = (inp[12]) ? 4'b0001 : node13245;
															assign node13245 = (inp[7]) ? 4'b1001 : node13246;
																assign node13246 = (inp[4]) ? 4'b0000 : 4'b1001;
													assign node13251 = (inp[4]) ? node13257 : node13252;
														assign node13252 = (inp[10]) ? node13254 : 4'b1001;
															assign node13254 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13257 = (inp[7]) ? node13265 : node13258;
															assign node13258 = (inp[10]) ? node13262 : node13259;
																assign node13259 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node13262 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node13265 = (inp[12]) ? 4'b1001 : node13266;
																assign node13266 = (inp[10]) ? 4'b0000 : 4'b1001;
												assign node13270 = (inp[13]) ? node13288 : node13271;
													assign node13271 = (inp[4]) ? node13277 : node13272;
														assign node13272 = (inp[10]) ? 4'b1000 : node13273;
															assign node13273 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13277 = (inp[7]) ? node13285 : node13278;
															assign node13278 = (inp[12]) ? node13282 : node13279;
																assign node13279 = (inp[10]) ? 4'b0001 : 4'b1100;
																assign node13282 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node13285 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node13288 = (inp[4]) ? node13296 : node13289;
														assign node13289 = (inp[7]) ? 4'b0000 : node13290;
															assign node13290 = (inp[12]) ? node13292 : 4'b0100;
																assign node13292 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node13296 = (inp[7]) ? node13302 : node13297;
															assign node13297 = (inp[12]) ? node13299 : 4'b0001;
																assign node13299 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node13302 = (inp[12]) ? node13306 : node13303;
																assign node13303 = (inp[10]) ? 4'b0001 : 4'b0100;
																assign node13306 = (inp[10]) ? 4'b0100 : 4'b1000;
										assign node13309 = (inp[4]) ? node13363 : node13310;
											assign node13310 = (inp[10]) ? node13332 : node13311;
												assign node13311 = (inp[13]) ? node13319 : node13312;
													assign node13312 = (inp[11]) ? node13316 : node13313;
														assign node13313 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13316 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13319 = (inp[11]) ? 4'b0000 : node13320;
														assign node13320 = (inp[14]) ? node13326 : node13321;
															assign node13321 = (inp[7]) ? node13323 : 4'b1001;
																assign node13323 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node13326 = (inp[12]) ? node13328 : 4'b0000;
																assign node13328 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node13332 = (inp[13]) ? node13350 : node13333;
													assign node13333 = (inp[11]) ? node13343 : node13334;
														assign node13334 = (inp[12]) ? node13340 : node13335;
															assign node13335 = (inp[7]) ? 4'b0000 : node13336;
																assign node13336 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node13340 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node13343 = (inp[7]) ? node13347 : node13344;
															assign node13344 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13347 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node13350 = (inp[7]) ? node13356 : node13351;
														assign node13351 = (inp[12]) ? node13353 : 4'b1001;
															assign node13353 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node13356 = (inp[11]) ? node13360 : node13357;
															assign node13357 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node13360 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node13363 = (inp[13]) ? node13397 : node13364;
												assign node13364 = (inp[10]) ? node13384 : node13365;
													assign node13365 = (inp[14]) ? node13377 : node13366;
														assign node13366 = (inp[7]) ? node13372 : node13367;
															assign node13367 = (inp[11]) ? node13369 : 4'b1000;
																assign node13369 = (inp[12]) ? 4'b1000 : 4'b0001;
															assign node13372 = (inp[11]) ? 4'b1001 : node13373;
																assign node13373 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node13377 = (inp[11]) ? node13381 : node13378;
															assign node13378 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node13381 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node13384 = (inp[7]) ? node13392 : node13385;
														assign node13385 = (inp[12]) ? node13389 : node13386;
															assign node13386 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node13389 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node13392 = (inp[12]) ? node13394 : 4'b0000;
															assign node13394 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node13397 = (inp[11]) ? node13421 : node13398;
													assign node13398 = (inp[12]) ? node13408 : node13399;
														assign node13399 = (inp[7]) ? node13405 : node13400;
															assign node13400 = (inp[10]) ? node13402 : 4'b0001;
																assign node13402 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node13405 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node13408 = (inp[10]) ? node13416 : node13409;
															assign node13409 = (inp[7]) ? node13413 : node13410;
																assign node13410 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node13413 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node13416 = (inp[7]) ? 4'b0000 : node13417;
																assign node13417 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node13421 = (inp[10]) ? 4'b0000 : node13422;
														assign node13422 = (inp[7]) ? 4'b0000 : node13423;
															assign node13423 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node13428 = (inp[11]) ? node13562 : node13429;
										assign node13429 = (inp[14]) ? node13497 : node13430;
											assign node13430 = (inp[3]) ? node13458 : node13431;
												assign node13431 = (inp[13]) ? node13443 : node13432;
													assign node13432 = (inp[4]) ? node13438 : node13433;
														assign node13433 = (inp[12]) ? node13435 : 4'b1001;
															assign node13435 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13438 = (inp[7]) ? 4'b1001 : node13439;
															assign node13439 = (inp[10]) ? 4'b0000 : 4'b1101;
													assign node13443 = (inp[4]) ? node13451 : node13444;
														assign node13444 = (inp[7]) ? 4'b0001 : node13445;
															assign node13445 = (inp[10]) ? 4'b0101 : node13446;
																assign node13446 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node13451 = (inp[10]) ? 4'b0000 : node13452;
															assign node13452 = (inp[12]) ? node13454 : 4'b0101;
																assign node13454 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node13458 = (inp[4]) ? node13476 : node13459;
													assign node13459 = (inp[13]) ? node13469 : node13460;
														assign node13460 = (inp[7]) ? node13466 : node13461;
															assign node13461 = (inp[12]) ? 4'b1000 : node13462;
																assign node13462 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node13466 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node13469 = (inp[12]) ? node13471 : 4'b0001;
															assign node13471 = (inp[7]) ? 4'b0000 : node13472;
																assign node13472 = (inp[10]) ? 4'b1001 : 4'b0000;
													assign node13476 = (inp[10]) ? node13488 : node13477;
														assign node13477 = (inp[12]) ? node13483 : node13478;
															assign node13478 = (inp[7]) ? node13480 : 4'b0001;
																assign node13480 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node13483 = (inp[13]) ? 4'b0001 : node13484;
																assign node13484 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node13488 = (inp[7]) ? node13492 : node13489;
															assign node13489 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node13492 = (inp[13]) ? 4'b0000 : node13493;
																assign node13493 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node13497 = (inp[3]) ? node13533 : node13498;
												assign node13498 = (inp[13]) ? node13518 : node13499;
													assign node13499 = (inp[12]) ? node13507 : node13500;
														assign node13500 = (inp[7]) ? 4'b1000 : node13501;
															assign node13501 = (inp[10]) ? node13503 : 4'b1100;
																assign node13503 = (inp[4]) ? 4'b0000 : 4'b1000;
														assign node13507 = (inp[10]) ? node13513 : node13508;
															assign node13508 = (inp[7]) ? 4'b0000 : node13509;
																assign node13509 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node13513 = (inp[4]) ? node13515 : 4'b1000;
																assign node13515 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node13518 = (inp[10]) ? node13528 : node13519;
														assign node13519 = (inp[12]) ? 4'b1000 : node13520;
															assign node13520 = (inp[4]) ? node13524 : node13521;
																assign node13521 = (inp[7]) ? 4'b0000 : 4'b0100;
																assign node13524 = (inp[7]) ? 4'b0100 : 4'b1000;
														assign node13528 = (inp[4]) ? 4'b0000 : node13529;
															assign node13529 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node13533 = (inp[4]) ? node13545 : node13534;
													assign node13534 = (inp[13]) ? node13540 : node13535;
														assign node13535 = (inp[10]) ? node13537 : 4'b1000;
															assign node13537 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node13540 = (inp[10]) ? node13542 : 4'b0001;
															assign node13542 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node13545 = (inp[7]) ? node13557 : node13546;
														assign node13546 = (inp[13]) ? node13552 : node13547;
															assign node13547 = (inp[10]) ? 4'b0000 : node13548;
																assign node13548 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node13552 = (inp[12]) ? node13554 : 4'b0000;
																assign node13554 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node13557 = (inp[10]) ? node13559 : 4'b0000;
															assign node13559 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node13562 = (inp[13]) ? node13604 : node13563;
											assign node13563 = (inp[4]) ? node13583 : node13564;
												assign node13564 = (inp[3]) ? node13570 : node13565;
													assign node13565 = (inp[12]) ? node13567 : 4'b1001;
														assign node13567 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node13570 = (inp[12]) ? node13578 : node13571;
														assign node13571 = (inp[10]) ? node13575 : node13572;
															assign node13572 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node13575 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node13578 = (inp[7]) ? node13580 : 4'b1001;
															assign node13580 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node13583 = (inp[7]) ? node13593 : node13584;
													assign node13584 = (inp[10]) ? 4'b0001 : node13585;
														assign node13585 = (inp[3]) ? node13589 : node13586;
															assign node13586 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node13589 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node13593 = (inp[3]) ? node13599 : node13594;
														assign node13594 = (inp[12]) ? node13596 : 4'b1001;
															assign node13596 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node13599 = (inp[10]) ? 4'b0001 : node13600;
															assign node13600 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node13604 = (inp[10]) ? node13622 : node13605;
												assign node13605 = (inp[3]) ? node13615 : node13606;
													assign node13606 = (inp[12]) ? 4'b1001 : node13607;
														assign node13607 = (inp[7]) ? node13611 : node13608;
															assign node13608 = (inp[4]) ? 4'b1001 : 4'b0101;
															assign node13611 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node13615 = (inp[7]) ? node13617 : 4'b0001;
														assign node13617 = (inp[12]) ? 4'b0001 : node13618;
															assign node13618 = (inp[4]) ? 4'b0001 : 4'b1001;
												assign node13622 = (inp[3]) ? node13628 : node13623;
													assign node13623 = (inp[4]) ? 4'b0001 : node13624;
														assign node13624 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node13628 = (inp[4]) ? 4'b0000 : 4'b0001;
							assign node13631 = (inp[5]) ? node13633 : 4'b0001;
								assign node13633 = (inp[3]) ? node13635 : 4'b0001;
									assign node13635 = (inp[4]) ? node13659 : node13636;
										assign node13636 = (inp[13]) ? node13638 : 4'b0001;
											assign node13638 = (inp[7]) ? 4'b0001 : node13639;
												assign node13639 = (inp[1]) ? node13651 : node13640;
													assign node13640 = (inp[12]) ? node13646 : node13641;
														assign node13641 = (inp[11]) ? 4'b0000 : node13642;
															assign node13642 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node13646 = (inp[10]) ? node13648 : 4'b0001;
															assign node13648 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node13651 = (inp[14]) ? node13653 : 4'b0001;
														assign node13653 = (inp[11]) ? 4'b0001 : node13654;
															assign node13654 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node13659 = (inp[13]) ? node13701 : node13660;
											assign node13660 = (inp[7]) ? 4'b0001 : node13661;
												assign node13661 = (inp[1]) ? node13685 : node13662;
													assign node13662 = (inp[14]) ? node13672 : node13663;
														assign node13663 = (inp[11]) ? 4'b1000 : node13664;
															assign node13664 = (inp[10]) ? node13668 : node13665;
																assign node13665 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node13668 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node13672 = (inp[11]) ? node13678 : node13673;
															assign node13673 = (inp[12]) ? 4'b0001 : node13674;
																assign node13674 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node13678 = (inp[12]) ? node13682 : node13679;
																assign node13679 = (inp[10]) ? 4'b0001 : 4'b1000;
																assign node13682 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node13685 = (inp[11]) ? node13695 : node13686;
														assign node13686 = (inp[14]) ? node13690 : node13687;
															assign node13687 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node13690 = (inp[12]) ? 4'b0000 : node13691;
																assign node13691 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node13695 = (inp[10]) ? 4'b0001 : node13696;
															assign node13696 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node13701 = (inp[10]) ? node13727 : node13702;
												assign node13702 = (inp[1]) ? node13714 : node13703;
													assign node13703 = (inp[7]) ? node13709 : node13704;
														assign node13704 = (inp[11]) ? 4'b0000 : node13705;
															assign node13705 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node13709 = (inp[12]) ? 4'b0001 : node13710;
															assign node13710 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node13714 = (inp[11]) ? 4'b0001 : node13715;
														assign node13715 = (inp[7]) ? node13721 : node13716;
															assign node13716 = (inp[12]) ? node13718 : 4'b0001;
																assign node13718 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node13721 = (inp[12]) ? 4'b0001 : node13722;
																assign node13722 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node13727 = (inp[1]) ? 4'b0000 : node13728;
													assign node13728 = (inp[11]) ? 4'b0000 : node13729;
														assign node13729 = (inp[14]) ? node13731 : 4'b0000;
															assign node13731 = (inp[7]) ? node13733 : 4'b0000;
																assign node13733 = (inp[12]) ? 4'b0001 : 4'b0000;
		assign node13738 = (inp[9]) ? node20740 : node13739;
			assign node13739 = (inp[15]) ? node17459 : node13740;
				assign node13740 = (inp[6]) ? node14636 : node13741;
					assign node13741 = (inp[0]) ? 4'b1100 : node13742;
						assign node13742 = (inp[2]) ? node14246 : node13743;
							assign node13743 = (inp[1]) ? node13997 : node13744;
								assign node13744 = (inp[13]) ? node13892 : node13745;
									assign node13745 = (inp[14]) ? node13801 : node13746;
										assign node13746 = (inp[3]) ? node13782 : node13747;
											assign node13747 = (inp[5]) ? node13765 : node13748;
												assign node13748 = (inp[4]) ? node13754 : node13749;
													assign node13749 = (inp[12]) ? 4'b1110 : node13750;
														assign node13750 = (inp[7]) ? 4'b1110 : 4'b0001;
													assign node13754 = (inp[7]) ? node13760 : node13755;
														assign node13755 = (inp[10]) ? node13757 : 4'b1001;
															assign node13757 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node13760 = (inp[12]) ? 4'b1110 : node13761;
															assign node13761 = (inp[10]) ? 4'b0001 : 4'b1110;
												assign node13765 = (inp[12]) ? node13777 : node13766;
													assign node13766 = (inp[10]) ? node13772 : node13767;
														assign node13767 = (inp[4]) ? node13769 : 4'b1101;
															assign node13769 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node13772 = (inp[4]) ? 4'b0001 : node13773;
															assign node13773 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node13777 = (inp[7]) ? 4'b1101 : node13778;
														assign node13778 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node13782 = (inp[7]) ? node13794 : node13783;
												assign node13783 = (inp[4]) ? node13789 : node13784;
													assign node13784 = (inp[10]) ? node13786 : 4'b1001;
														assign node13786 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node13789 = (inp[12]) ? 4'b1101 : node13790;
														assign node13790 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node13794 = (inp[12]) ? 4'b1001 : node13795;
													assign node13795 = (inp[10]) ? node13797 : 4'b1001;
														assign node13797 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node13801 = (inp[11]) ? node13851 : node13802;
											assign node13802 = (inp[12]) ? node13834 : node13803;
												assign node13803 = (inp[10]) ? node13821 : node13804;
													assign node13804 = (inp[3]) ? node13816 : node13805;
														assign node13805 = (inp[5]) ? node13811 : node13806;
															assign node13806 = (inp[7]) ? 4'b1110 : node13807;
																assign node13807 = (inp[4]) ? 4'b1000 : 4'b1110;
															assign node13811 = (inp[7]) ? 4'b1100 : node13812;
																assign node13812 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node13816 = (inp[4]) ? node13818 : 4'b1000;
															assign node13818 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node13821 = (inp[3]) ? node13829 : node13822;
														assign node13822 = (inp[7]) ? node13824 : 4'b0000;
															assign node13824 = (inp[4]) ? 4'b0000 : node13825;
																assign node13825 = (inp[5]) ? 4'b0100 : 4'b1110;
														assign node13829 = (inp[7]) ? node13831 : 4'b0100;
															assign node13831 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node13834 = (inp[3]) ? node13846 : node13835;
													assign node13835 = (inp[5]) ? node13841 : node13836;
														assign node13836 = (inp[4]) ? node13838 : 4'b1110;
															assign node13838 = (inp[7]) ? 4'b1110 : 4'b1000;
														assign node13841 = (inp[4]) ? node13843 : 4'b1100;
															assign node13843 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node13846 = (inp[7]) ? 4'b1000 : node13847;
														assign node13847 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node13851 = (inp[3]) ? node13875 : node13852;
												assign node13852 = (inp[5]) ? node13860 : node13853;
													assign node13853 = (inp[4]) ? node13855 : 4'b1110;
														assign node13855 = (inp[7]) ? 4'b1110 : node13856;
															assign node13856 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node13860 = (inp[4]) ? node13868 : node13861;
														assign node13861 = (inp[12]) ? 4'b1101 : node13862;
															assign node13862 = (inp[10]) ? node13864 : 4'b1101;
																assign node13864 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node13868 = (inp[7]) ? node13870 : 4'b1001;
															assign node13870 = (inp[10]) ? node13872 : 4'b1101;
																assign node13872 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node13875 = (inp[10]) ? node13881 : node13876;
													assign node13876 = (inp[4]) ? node13878 : 4'b1001;
														assign node13878 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node13881 = (inp[12]) ? node13887 : node13882;
														assign node13882 = (inp[4]) ? 4'b0101 : node13883;
															assign node13883 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node13887 = (inp[7]) ? 4'b1001 : node13888;
															assign node13888 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node13892 = (inp[3]) ? node13944 : node13893;
										assign node13893 = (inp[7]) ? node13911 : node13894;
											assign node13894 = (inp[14]) ? node13900 : node13895;
												assign node13895 = (inp[12]) ? 4'b0001 : node13896;
													assign node13896 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node13900 = (inp[11]) ? node13906 : node13901;
													assign node13901 = (inp[10]) ? node13903 : 4'b0000;
														assign node13903 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node13906 = (inp[10]) ? node13908 : 4'b0001;
														assign node13908 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node13911 = (inp[4]) ? node13927 : node13912;
												assign node13912 = (inp[5]) ? node13914 : 4'b1110;
													assign node13914 = (inp[12]) ? node13922 : node13915;
														assign node13915 = (inp[10]) ? node13917 : 4'b0101;
															assign node13917 = (inp[11]) ? 4'b1101 : node13918;
																assign node13918 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13922 = (inp[11]) ? 4'b0101 : node13923;
															assign node13923 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node13927 = (inp[14]) ? node13933 : node13928;
													assign node13928 = (inp[10]) ? node13930 : 4'b0001;
														assign node13930 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node13933 = (inp[11]) ? node13939 : node13934;
														assign node13934 = (inp[10]) ? node13936 : 4'b0000;
															assign node13936 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node13939 = (inp[10]) ? node13941 : 4'b0001;
															assign node13941 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node13944 = (inp[14]) ? node13962 : node13945;
											assign node13945 = (inp[4]) ? node13957 : node13946;
												assign node13946 = (inp[7]) ? node13952 : node13947;
													assign node13947 = (inp[10]) ? node13949 : 4'b0101;
														assign node13949 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node13952 = (inp[12]) ? 4'b0001 : node13953;
														assign node13953 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node13957 = (inp[12]) ? 4'b0101 : node13958;
													assign node13958 = (inp[10]) ? 4'b1101 : 4'b0101;
											assign node13962 = (inp[11]) ? node13980 : node13963;
												assign node13963 = (inp[12]) ? node13975 : node13964;
													assign node13964 = (inp[10]) ? node13970 : node13965;
														assign node13965 = (inp[7]) ? node13967 : 4'b0100;
															assign node13967 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node13970 = (inp[7]) ? node13972 : 4'b1100;
															assign node13972 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node13975 = (inp[7]) ? node13977 : 4'b0100;
														assign node13977 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node13980 = (inp[12]) ? node13992 : node13981;
													assign node13981 = (inp[10]) ? node13987 : node13982;
														assign node13982 = (inp[7]) ? node13984 : 4'b0101;
															assign node13984 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node13987 = (inp[4]) ? 4'b1101 : node13988;
															assign node13988 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node13992 = (inp[7]) ? node13994 : 4'b0101;
														assign node13994 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node13997 = (inp[11]) ? node14163 : node13998;
									assign node13998 = (inp[14]) ? node14078 : node13999;
										assign node13999 = (inp[13]) ? node14045 : node14000;
											assign node14000 = (inp[12]) ? node14014 : node14001;
												assign node14001 = (inp[3]) ? node14009 : node14002;
													assign node14002 = (inp[4]) ? 4'b0000 : node14003;
														assign node14003 = (inp[5]) ? node14005 : 4'b1110;
															assign node14005 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node14009 = (inp[7]) ? node14011 : 4'b0100;
														assign node14011 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node14014 = (inp[10]) ? node14032 : node14015;
													assign node14015 = (inp[3]) ? node14027 : node14016;
														assign node14016 = (inp[5]) ? node14022 : node14017;
															assign node14017 = (inp[4]) ? node14019 : 4'b1110;
																assign node14019 = (inp[7]) ? 4'b1110 : 4'b1000;
															assign node14022 = (inp[7]) ? 4'b1100 : node14023;
																assign node14023 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node14027 = (inp[4]) ? node14029 : 4'b1000;
															assign node14029 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node14032 = (inp[3]) ? node14040 : node14033;
														assign node14033 = (inp[4]) ? 4'b0000 : node14034;
															assign node14034 = (inp[5]) ? node14036 : 4'b1110;
																assign node14036 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node14040 = (inp[7]) ? node14042 : 4'b0100;
															assign node14042 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node14045 = (inp[3]) ? node14061 : node14046;
												assign node14046 = (inp[7]) ? node14052 : node14047;
													assign node14047 = (inp[10]) ? 4'b1000 : node14048;
														assign node14048 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14052 = (inp[4]) ? node14056 : node14053;
														assign node14053 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node14056 = (inp[12]) ? node14058 : 4'b1000;
															assign node14058 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14061 = (inp[4]) ? node14073 : node14062;
													assign node14062 = (inp[7]) ? node14068 : node14063;
														assign node14063 = (inp[10]) ? 4'b1100 : node14064;
															assign node14064 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node14068 = (inp[10]) ? 4'b1000 : node14069;
															assign node14069 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node14073 = (inp[12]) ? node14075 : 4'b1100;
														assign node14075 = (inp[10]) ? 4'b1100 : 4'b0100;
										assign node14078 = (inp[13]) ? node14130 : node14079;
											assign node14079 = (inp[3]) ? node14113 : node14080;
												assign node14080 = (inp[5]) ? node14100 : node14081;
													assign node14081 = (inp[7]) ? node14093 : node14082;
														assign node14082 = (inp[4]) ? node14088 : node14083;
															assign node14083 = (inp[12]) ? 4'b1110 : node14084;
																assign node14084 = (inp[10]) ? 4'b0001 : 4'b1110;
															assign node14088 = (inp[10]) ? node14090 : 4'b1001;
																assign node14090 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14093 = (inp[12]) ? 4'b1110 : node14094;
															assign node14094 = (inp[10]) ? node14096 : 4'b1110;
																assign node14096 = (inp[4]) ? 4'b0001 : 4'b1110;
													assign node14100 = (inp[7]) ? node14108 : node14101;
														assign node14101 = (inp[4]) ? node14103 : 4'b1101;
															assign node14103 = (inp[10]) ? node14105 : 4'b1001;
																assign node14105 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14108 = (inp[10]) ? node14110 : 4'b1101;
															assign node14110 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node14113 = (inp[10]) ? node14119 : node14114;
													assign node14114 = (inp[7]) ? 4'b1001 : node14115;
														assign node14115 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node14119 = (inp[12]) ? node14125 : node14120;
														assign node14120 = (inp[7]) ? node14122 : 4'b0101;
															assign node14122 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node14125 = (inp[7]) ? 4'b1001 : node14126;
															assign node14126 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node14130 = (inp[3]) ? node14146 : node14131;
												assign node14131 = (inp[7]) ? node14137 : node14132;
													assign node14132 = (inp[10]) ? node14134 : 4'b0001;
														assign node14134 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14137 = (inp[4]) ? node14141 : node14138;
														assign node14138 = (inp[5]) ? 4'b0101 : 4'b1110;
														assign node14141 = (inp[12]) ? 4'b0001 : node14142;
															assign node14142 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node14146 = (inp[7]) ? node14152 : node14147;
													assign node14147 = (inp[12]) ? 4'b0101 : node14148;
														assign node14148 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node14152 = (inp[4]) ? node14158 : node14153;
														assign node14153 = (inp[12]) ? 4'b0001 : node14154;
															assign node14154 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node14158 = (inp[12]) ? 4'b0101 : node14159;
															assign node14159 = (inp[10]) ? 4'b1101 : 4'b0101;
									assign node14163 = (inp[13]) ? node14209 : node14164;
										assign node14164 = (inp[12]) ? node14178 : node14165;
											assign node14165 = (inp[3]) ? node14173 : node14166;
												assign node14166 = (inp[4]) ? 4'b0000 : node14167;
													assign node14167 = (inp[7]) ? node14169 : 4'b0000;
														assign node14169 = (inp[5]) ? 4'b0100 : 4'b1110;
												assign node14173 = (inp[4]) ? 4'b0100 : node14174;
													assign node14174 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node14178 = (inp[10]) ? node14196 : node14179;
												assign node14179 = (inp[3]) ? node14191 : node14180;
													assign node14180 = (inp[5]) ? node14186 : node14181;
														assign node14181 = (inp[7]) ? 4'b1110 : node14182;
															assign node14182 = (inp[4]) ? 4'b1000 : 4'b1110;
														assign node14186 = (inp[7]) ? 4'b1100 : node14187;
															assign node14187 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node14191 = (inp[4]) ? node14193 : 4'b1000;
														assign node14193 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node14196 = (inp[3]) ? node14204 : node14197;
													assign node14197 = (inp[4]) ? 4'b0000 : node14198;
														assign node14198 = (inp[7]) ? node14200 : 4'b0000;
															assign node14200 = (inp[5]) ? 4'b0100 : 4'b1110;
													assign node14204 = (inp[7]) ? node14206 : 4'b0100;
														assign node14206 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node14209 = (inp[3]) ? node14229 : node14210;
											assign node14210 = (inp[7]) ? node14216 : node14211;
												assign node14211 = (inp[10]) ? 4'b1000 : node14212;
													assign node14212 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node14216 = (inp[4]) ? node14224 : node14217;
													assign node14217 = (inp[5]) ? node14219 : 4'b1110;
														assign node14219 = (inp[12]) ? node14221 : 4'b1100;
															assign node14221 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node14224 = (inp[10]) ? 4'b1000 : node14225;
														assign node14225 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node14229 = (inp[4]) ? node14241 : node14230;
												assign node14230 = (inp[7]) ? node14236 : node14231;
													assign node14231 = (inp[10]) ? 4'b1100 : node14232;
														assign node14232 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node14236 = (inp[12]) ? node14238 : 4'b1000;
														assign node14238 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node14241 = (inp[12]) ? node14243 : 4'b1100;
													assign node14243 = (inp[10]) ? 4'b1100 : 4'b0100;
							assign node14246 = (inp[5]) ? node14248 : 4'b1110;
								assign node14248 = (inp[3]) ? node14438 : node14249;
									assign node14249 = (inp[4]) ? node14313 : node14250;
										assign node14250 = (inp[7]) ? 4'b1110 : node14251;
											assign node14251 = (inp[13]) ? node14279 : node14252;
												assign node14252 = (inp[12]) ? node14272 : node14253;
													assign node14253 = (inp[10]) ? node14261 : node14254;
														assign node14254 = (inp[1]) ? node14256 : 4'b1110;
															assign node14256 = (inp[11]) ? 4'b0000 : node14257;
																assign node14257 = (inp[14]) ? 4'b1110 : 4'b0000;
														assign node14261 = (inp[1]) ? node14267 : node14262;
															assign node14262 = (inp[14]) ? node14264 : 4'b0001;
																assign node14264 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node14267 = (inp[14]) ? node14269 : 4'b0000;
																assign node14269 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node14272 = (inp[11]) ? node14274 : 4'b1110;
														assign node14274 = (inp[1]) ? node14276 : 4'b1110;
															assign node14276 = (inp[10]) ? 4'b0000 : 4'b1110;
												assign node14279 = (inp[1]) ? node14295 : node14280;
													assign node14280 = (inp[14]) ? node14286 : node14281;
														assign node14281 = (inp[12]) ? 4'b0001 : node14282;
															assign node14282 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node14286 = (inp[11]) ? node14292 : node14287;
															assign node14287 = (inp[10]) ? node14289 : 4'b0000;
																assign node14289 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14292 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14295 = (inp[11]) ? node14307 : node14296;
														assign node14296 = (inp[14]) ? node14302 : node14297;
															assign node14297 = (inp[10]) ? 4'b1000 : node14298;
																assign node14298 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14302 = (inp[10]) ? node14304 : 4'b0001;
																assign node14304 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node14307 = (inp[12]) ? node14309 : 4'b1000;
															assign node14309 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node14313 = (inp[7]) ? node14379 : node14314;
											assign node14314 = (inp[1]) ? node14346 : node14315;
												assign node14315 = (inp[14]) ? node14327 : node14316;
													assign node14316 = (inp[13]) ? node14322 : node14317;
														assign node14317 = (inp[10]) ? node14319 : 4'b1001;
															assign node14319 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node14322 = (inp[11]) ? node14324 : 4'b0001;
															assign node14324 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node14327 = (inp[11]) ? node14339 : node14328;
														assign node14328 = (inp[13]) ? node14334 : node14329;
															assign node14329 = (inp[12]) ? 4'b1000 : node14330;
																assign node14330 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node14334 = (inp[10]) ? node14336 : 4'b0000;
																assign node14336 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14339 = (inp[13]) ? node14343 : node14340;
															assign node14340 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node14343 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node14346 = (inp[11]) ? node14368 : node14347;
													assign node14347 = (inp[14]) ? node14357 : node14348;
														assign node14348 = (inp[13]) ? node14354 : node14349;
															assign node14349 = (inp[10]) ? 4'b0000 : node14350;
																assign node14350 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node14354 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14357 = (inp[13]) ? node14363 : node14358;
															assign node14358 = (inp[12]) ? 4'b1001 : node14359;
																assign node14359 = (inp[10]) ? 4'b0001 : 4'b1001;
															assign node14363 = (inp[10]) ? node14365 : 4'b0001;
																assign node14365 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14368 = (inp[13]) ? node14374 : node14369;
														assign node14369 = (inp[10]) ? 4'b0000 : node14370;
															assign node14370 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node14374 = (inp[12]) ? node14376 : 4'b1000;
															assign node14376 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node14379 = (inp[13]) ? node14409 : node14380;
												assign node14380 = (inp[10]) ? node14390 : node14381;
													assign node14381 = (inp[12]) ? 4'b1110 : node14382;
														assign node14382 = (inp[1]) ? node14384 : 4'b1110;
															assign node14384 = (inp[11]) ? 4'b0000 : node14385;
																assign node14385 = (inp[14]) ? 4'b1110 : 4'b0000;
													assign node14390 = (inp[12]) ? node14402 : node14391;
														assign node14391 = (inp[1]) ? node14397 : node14392;
															assign node14392 = (inp[11]) ? 4'b0001 : node14393;
																assign node14393 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14397 = (inp[11]) ? 4'b0000 : node14398;
																assign node14398 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node14402 = (inp[11]) ? 4'b0000 : node14403;
															assign node14403 = (inp[14]) ? 4'b1110 : node14404;
																assign node14404 = (inp[1]) ? 4'b0000 : 4'b1110;
												assign node14409 = (inp[1]) ? node14425 : node14410;
													assign node14410 = (inp[14]) ? node14416 : node14411;
														assign node14411 = (inp[12]) ? 4'b0001 : node14412;
															assign node14412 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node14416 = (inp[11]) ? node14422 : node14417;
															assign node14417 = (inp[10]) ? node14419 : 4'b0000;
																assign node14419 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14422 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node14425 = (inp[14]) ? node14431 : node14426;
														assign node14426 = (inp[10]) ? 4'b1000 : node14427;
															assign node14427 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node14431 = (inp[11]) ? 4'b1000 : node14432;
															assign node14432 = (inp[12]) ? 4'b0001 : node14433;
																assign node14433 = (inp[10]) ? 4'b1001 : 4'b0001;
									assign node14438 = (inp[1]) ? node14532 : node14439;
										assign node14439 = (inp[13]) ? node14485 : node14440;
											assign node14440 = (inp[12]) ? node14468 : node14441;
												assign node14441 = (inp[10]) ? node14455 : node14442;
													assign node14442 = (inp[11]) ? node14450 : node14443;
														assign node14443 = (inp[14]) ? node14445 : 4'b1001;
															assign node14445 = (inp[7]) ? 4'b1000 : node14446;
																assign node14446 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node14450 = (inp[4]) ? node14452 : 4'b1001;
															assign node14452 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node14455 = (inp[7]) ? node14461 : node14456;
														assign node14456 = (inp[11]) ? 4'b0101 : node14457;
															assign node14457 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node14461 = (inp[4]) ? 4'b0101 : node14462;
															assign node14462 = (inp[11]) ? 4'b0001 : node14463;
																assign node14463 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node14468 = (inp[4]) ? node14474 : node14469;
													assign node14469 = (inp[11]) ? 4'b1001 : node14470;
														assign node14470 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node14474 = (inp[7]) ? node14480 : node14475;
														assign node14475 = (inp[14]) ? node14477 : 4'b1101;
															assign node14477 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14480 = (inp[14]) ? node14482 : 4'b1001;
															assign node14482 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node14485 = (inp[12]) ? node14515 : node14486;
												assign node14486 = (inp[10]) ? node14502 : node14487;
													assign node14487 = (inp[7]) ? node14493 : node14488;
														assign node14488 = (inp[14]) ? node14490 : 4'b0101;
															assign node14490 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node14493 = (inp[4]) ? node14499 : node14494;
															assign node14494 = (inp[11]) ? 4'b0001 : node14495;
																assign node14495 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14499 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node14502 = (inp[4]) ? node14510 : node14503;
														assign node14503 = (inp[7]) ? node14505 : 4'b1101;
															assign node14505 = (inp[14]) ? node14507 : 4'b1001;
																assign node14507 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node14510 = (inp[11]) ? 4'b1101 : node14511;
															assign node14511 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node14515 = (inp[14]) ? node14521 : node14516;
													assign node14516 = (inp[4]) ? 4'b0101 : node14517;
														assign node14517 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node14521 = (inp[11]) ? node14527 : node14522;
														assign node14522 = (inp[7]) ? node14524 : 4'b0100;
															assign node14524 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node14527 = (inp[4]) ? 4'b0101 : node14528;
															assign node14528 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node14532 = (inp[11]) ? node14600 : node14533;
											assign node14533 = (inp[14]) ? node14569 : node14534;
												assign node14534 = (inp[13]) ? node14552 : node14535;
													assign node14535 = (inp[10]) ? node14547 : node14536;
														assign node14536 = (inp[12]) ? node14542 : node14537;
															assign node14537 = (inp[7]) ? node14539 : 4'b0100;
																assign node14539 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node14542 = (inp[7]) ? 4'b1000 : node14543;
																assign node14543 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node14547 = (inp[7]) ? node14549 : 4'b0100;
															assign node14549 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node14552 = (inp[7]) ? node14558 : node14553;
														assign node14553 = (inp[12]) ? node14555 : 4'b1100;
															assign node14555 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node14558 = (inp[4]) ? node14564 : node14559;
															assign node14559 = (inp[10]) ? 4'b1000 : node14560;
																assign node14560 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node14564 = (inp[12]) ? node14566 : 4'b1100;
																assign node14566 = (inp[10]) ? 4'b1100 : 4'b0100;
												assign node14569 = (inp[13]) ? node14587 : node14570;
													assign node14570 = (inp[12]) ? node14582 : node14571;
														assign node14571 = (inp[10]) ? node14577 : node14572;
															assign node14572 = (inp[4]) ? node14574 : 4'b1001;
																assign node14574 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node14577 = (inp[7]) ? node14579 : 4'b0101;
																assign node14579 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node14582 = (inp[7]) ? 4'b1001 : node14583;
															assign node14583 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node14587 = (inp[7]) ? node14593 : node14588;
														assign node14588 = (inp[12]) ? 4'b0101 : node14589;
															assign node14589 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node14593 = (inp[4]) ? 4'b0101 : node14594;
															assign node14594 = (inp[10]) ? node14596 : 4'b0001;
																assign node14596 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node14600 = (inp[13]) ? node14618 : node14601;
												assign node14601 = (inp[10]) ? node14613 : node14602;
													assign node14602 = (inp[12]) ? node14608 : node14603;
														assign node14603 = (inp[4]) ? 4'b0100 : node14604;
															assign node14604 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node14608 = (inp[4]) ? node14610 : 4'b1000;
															assign node14610 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node14613 = (inp[7]) ? node14615 : 4'b0100;
														assign node14615 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node14618 = (inp[10]) ? node14630 : node14619;
													assign node14619 = (inp[12]) ? node14625 : node14620;
														assign node14620 = (inp[4]) ? 4'b1100 : node14621;
															assign node14621 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node14625 = (inp[4]) ? 4'b0100 : node14626;
															assign node14626 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node14630 = (inp[4]) ? 4'b1100 : node14631;
														assign node14631 = (inp[7]) ? 4'b1000 : 4'b1100;
					assign node14636 = (inp[5]) ? node15800 : node14637;
						assign node14637 = (inp[0]) ? node15445 : node14638;
							assign node14638 = (inp[11]) ? node15130 : node14639;
								assign node14639 = (inp[10]) ? node14871 : node14640;
									assign node14640 = (inp[13]) ? node14744 : node14641;
										assign node14641 = (inp[4]) ? node14689 : node14642;
											assign node14642 = (inp[3]) ? node14662 : node14643;
												assign node14643 = (inp[1]) ? node14647 : node14644;
													assign node14644 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node14647 = (inp[14]) ? node14655 : node14648;
														assign node14648 = (inp[12]) ? 4'b1100 : node14649;
															assign node14649 = (inp[7]) ? 4'b0100 : node14650;
																assign node14650 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node14655 = (inp[2]) ? 4'b1101 : node14656;
															assign node14656 = (inp[7]) ? 4'b1101 : node14657;
																assign node14657 = (inp[12]) ? 4'b1101 : 4'b0001;
												assign node14662 = (inp[2]) ? node14670 : node14663;
													assign node14663 = (inp[12]) ? 4'b1101 : node14664;
														assign node14664 = (inp[1]) ? node14666 : 4'b1101;
															assign node14666 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node14670 = (inp[12]) ? node14682 : node14671;
														assign node14671 = (inp[1]) ? node14675 : node14672;
															assign node14672 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14675 = (inp[14]) ? node14679 : node14676;
																assign node14676 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node14679 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node14682 = (inp[14]) ? node14686 : node14683;
															assign node14683 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node14686 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node14689 = (inp[1]) ? node14707 : node14690;
												assign node14690 = (inp[2]) ? node14698 : node14691;
													assign node14691 = (inp[3]) ? node14693 : 4'b1001;
														assign node14693 = (inp[14]) ? 4'b1001 : node14694;
															assign node14694 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node14698 = (inp[3]) ? 4'b1001 : node14699;
														assign node14699 = (inp[7]) ? node14703 : node14700;
															assign node14700 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14703 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node14707 = (inp[12]) ? node14729 : node14708;
													assign node14708 = (inp[14]) ? node14720 : node14709;
														assign node14709 = (inp[3]) ? node14715 : node14710;
															assign node14710 = (inp[2]) ? 4'b0000 : node14711;
																assign node14711 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node14715 = (inp[2]) ? node14717 : 4'b0001;
																assign node14717 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node14720 = (inp[3]) ? node14726 : node14721;
															assign node14721 = (inp[2]) ? node14723 : 4'b0001;
																assign node14723 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node14726 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node14729 = (inp[2]) ? node14735 : node14730;
														assign node14730 = (inp[3]) ? node14732 : 4'b1001;
															assign node14732 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node14735 = (inp[3]) ? 4'b1001 : node14736;
															assign node14736 = (inp[14]) ? node14740 : node14737;
																assign node14737 = (inp[7]) ? 4'b1100 : 4'b1000;
																assign node14740 = (inp[7]) ? 4'b1101 : 4'b1001;
										assign node14744 = (inp[2]) ? node14808 : node14745;
											assign node14745 = (inp[12]) ? node14779 : node14746;
												assign node14746 = (inp[1]) ? node14774 : node14747;
													assign node14747 = (inp[14]) ? node14761 : node14748;
														assign node14748 = (inp[4]) ? node14754 : node14749;
															assign node14749 = (inp[7]) ? node14751 : 4'b1001;
																assign node14751 = (inp[3]) ? 4'b1101 : 4'b0101;
															assign node14754 = (inp[7]) ? node14758 : node14755;
																assign node14755 = (inp[3]) ? 4'b1100 : 4'b1101;
																assign node14758 = (inp[3]) ? 4'b1000 : 4'b1001;
														assign node14761 = (inp[4]) ? node14767 : node14762;
															assign node14762 = (inp[7]) ? node14764 : 4'b1001;
																assign node14764 = (inp[3]) ? 4'b1101 : 4'b0100;
															assign node14767 = (inp[7]) ? node14771 : node14768;
																assign node14768 = (inp[3]) ? 4'b0101 : 4'b1101;
																assign node14771 = (inp[3]) ? 4'b0001 : 4'b1001;
													assign node14774 = (inp[4]) ? node14776 : 4'b0001;
														assign node14776 = (inp[3]) ? 4'b1001 : 4'b0101;
												assign node14779 = (inp[7]) ? node14789 : node14780;
													assign node14780 = (inp[4]) ? node14782 : 4'b1001;
														assign node14782 = (inp[3]) ? node14784 : 4'b1101;
															assign node14784 = (inp[1]) ? node14786 : 4'b0100;
																assign node14786 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node14789 = (inp[4]) ? node14799 : node14790;
														assign node14790 = (inp[3]) ? 4'b1101 : node14791;
															assign node14791 = (inp[1]) ? node14795 : node14792;
																assign node14792 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node14795 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node14799 = (inp[3]) ? node14801 : 4'b1001;
															assign node14801 = (inp[1]) ? node14805 : node14802;
																assign node14802 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node14805 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node14808 = (inp[3]) ? node14848 : node14809;
												assign node14809 = (inp[4]) ? node14833 : node14810;
													assign node14810 = (inp[7]) ? node14824 : node14811;
														assign node14811 = (inp[12]) ? node14817 : node14812;
															assign node14812 = (inp[1]) ? 4'b1000 : node14813;
																assign node14813 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14817 = (inp[1]) ? node14821 : node14818;
																assign node14818 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node14821 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node14824 = (inp[1]) ? node14828 : node14825;
															assign node14825 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node14828 = (inp[14]) ? 4'b0101 : node14829;
																assign node14829 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node14833 = (inp[12]) ? node14841 : node14834;
														assign node14834 = (inp[1]) ? node14838 : node14835;
															assign node14835 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node14838 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node14841 = (inp[14]) ? node14845 : node14842;
															assign node14842 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node14845 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node14848 = (inp[4]) ? node14864 : node14849;
													assign node14849 = (inp[7]) ? node14855 : node14850;
														assign node14850 = (inp[12]) ? 4'b1001 : node14851;
															assign node14851 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node14855 = (inp[14]) ? node14861 : node14856;
															assign node14856 = (inp[1]) ? node14858 : 4'b0001;
																assign node14858 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node14861 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node14864 = (inp[7]) ? node14866 : 4'b1101;
														assign node14866 = (inp[1]) ? node14868 : 4'b1001;
															assign node14868 = (inp[12]) ? 4'b1001 : 4'b0101;
									assign node14871 = (inp[4]) ? node15003 : node14872;
										assign node14872 = (inp[7]) ? node14934 : node14873;
											assign node14873 = (inp[12]) ? node14907 : node14874;
												assign node14874 = (inp[1]) ? node14892 : node14875;
													assign node14875 = (inp[13]) ? node14881 : node14876;
														assign node14876 = (inp[2]) ? node14878 : 4'b0001;
															assign node14878 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node14881 = (inp[2]) ? node14887 : node14882;
															assign node14882 = (inp[3]) ? node14884 : 4'b0001;
																assign node14884 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node14887 = (inp[14]) ? 4'b1000 : node14888;
																assign node14888 = (inp[3]) ? 4'b0001 : 4'b1001;
													assign node14892 = (inp[2]) ? node14900 : node14893;
														assign node14893 = (inp[3]) ? node14895 : 4'b1001;
															assign node14895 = (inp[13]) ? node14897 : 4'b1001;
																assign node14897 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node14900 = (inp[3]) ? 4'b1001 : node14901;
															assign node14901 = (inp[14]) ? 4'b1001 : node14902;
																assign node14902 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node14907 = (inp[3]) ? node14923 : node14908;
													assign node14908 = (inp[2]) ? node14910 : 4'b0001;
														assign node14910 = (inp[13]) ? node14918 : node14911;
															assign node14911 = (inp[14]) ? node14915 : node14912;
																assign node14912 = (inp[1]) ? 4'b0000 : 4'b1101;
																assign node14915 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node14918 = (inp[1]) ? 4'b0001 : node14919;
																assign node14919 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node14923 = (inp[2]) ? 4'b0001 : node14924;
														assign node14924 = (inp[13]) ? node14926 : 4'b0001;
															assign node14926 = (inp[14]) ? node14930 : node14927;
																assign node14927 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node14930 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node14934 = (inp[13]) ? node14978 : node14935;
												assign node14935 = (inp[2]) ? node14955 : node14936;
													assign node14936 = (inp[3]) ? node14950 : node14937;
														assign node14937 = (inp[12]) ? node14945 : node14938;
															assign node14938 = (inp[1]) ? node14942 : node14939;
																assign node14939 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node14942 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node14945 = (inp[1]) ? 4'b0100 : node14946;
																assign node14946 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node14950 = (inp[12]) ? 4'b0101 : node14951;
															assign node14951 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node14955 = (inp[3]) ? node14963 : node14956;
														assign node14956 = (inp[12]) ? 4'b1101 : node14957;
															assign node14957 = (inp[14]) ? 4'b0101 : node14958;
																assign node14958 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node14963 = (inp[12]) ? node14971 : node14964;
															assign node14964 = (inp[14]) ? node14968 : node14965;
																assign node14965 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node14968 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node14971 = (inp[14]) ? node14975 : node14972;
																assign node14972 = (inp[1]) ? 4'b0000 : 4'b1001;
																assign node14975 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node14978 = (inp[2]) ? node14984 : node14979;
													assign node14979 = (inp[12]) ? 4'b0001 : node14980;
														assign node14980 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node14984 = (inp[3]) ? node14998 : node14985;
														assign node14985 = (inp[12]) ? node14991 : node14986;
															assign node14986 = (inp[14]) ? node14988 : 4'b1101;
																assign node14988 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node14991 = (inp[14]) ? node14995 : node14992;
																assign node14992 = (inp[1]) ? 4'b1100 : 4'b0101;
																assign node14995 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node14998 = (inp[1]) ? node15000 : 4'b0001;
															assign node15000 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node15003 = (inp[13]) ? node15085 : node15004;
											assign node15004 = (inp[7]) ? node15046 : node15005;
												assign node15005 = (inp[2]) ? node15025 : node15006;
													assign node15006 = (inp[3]) ? node15012 : node15007;
														assign node15007 = (inp[12]) ? 4'b0101 : node15008;
															assign node15008 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node15012 = (inp[12]) ? node15018 : node15013;
															assign node15013 = (inp[1]) ? node15015 : 4'b1001;
																assign node15015 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node15018 = (inp[1]) ? node15022 : node15019;
																assign node15019 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node15022 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node15025 = (inp[3]) ? node15041 : node15026;
														assign node15026 = (inp[12]) ? node15034 : node15027;
															assign node15027 = (inp[14]) ? node15031 : node15028;
																assign node15028 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node15031 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node15034 = (inp[1]) ? node15038 : node15035;
																assign node15035 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node15038 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node15041 = (inp[12]) ? 4'b0101 : node15042;
															assign node15042 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node15046 = (inp[3]) ? node15066 : node15047;
													assign node15047 = (inp[2]) ? node15053 : node15048;
														assign node15048 = (inp[12]) ? 4'b0001 : node15049;
															assign node15049 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node15053 = (inp[12]) ? node15059 : node15054;
															assign node15054 = (inp[1]) ? 4'b0000 : node15055;
																assign node15055 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node15059 = (inp[1]) ? node15063 : node15060;
																assign node15060 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node15063 = (inp[14]) ? 4'b1101 : 4'b0000;
													assign node15066 = (inp[2]) ? node15080 : node15067;
														assign node15067 = (inp[14]) ? node15073 : node15068;
															assign node15068 = (inp[1]) ? node15070 : 4'b1000;
																assign node15070 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node15073 = (inp[1]) ? node15077 : node15074;
																assign node15074 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node15077 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node15080 = (inp[1]) ? node15082 : 4'b0001;
															assign node15082 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node15085 = (inp[2]) ? node15109 : node15086;
												assign node15086 = (inp[3]) ? node15092 : node15087;
													assign node15087 = (inp[1]) ? node15089 : 4'b0101;
														assign node15089 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node15092 = (inp[12]) ? node15100 : node15093;
														assign node15093 = (inp[1]) ? node15097 : node15094;
															assign node15094 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node15097 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node15100 = (inp[1]) ? node15106 : node15101;
															assign node15101 = (inp[14]) ? node15103 : 4'b0100;
																assign node15103 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node15106 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node15109 = (inp[3]) ? node15125 : node15110;
													assign node15110 = (inp[12]) ? node15118 : node15111;
														assign node15111 = (inp[1]) ? node15115 : node15112;
															assign node15112 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node15115 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node15118 = (inp[14]) ? node15122 : node15119;
															assign node15119 = (inp[1]) ? 4'b1000 : 4'b0001;
															assign node15122 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node15125 = (inp[1]) ? node15127 : 4'b0101;
														assign node15127 = (inp[12]) ? 4'b0101 : 4'b1101;
								assign node15130 = (inp[1]) ? node15324 : node15131;
									assign node15131 = (inp[13]) ? node15237 : node15132;
										assign node15132 = (inp[3]) ? node15182 : node15133;
											assign node15133 = (inp[2]) ? node15165 : node15134;
												assign node15134 = (inp[4]) ? node15148 : node15135;
													assign node15135 = (inp[7]) ? node15143 : node15136;
														assign node15136 = (inp[12]) ? node15140 : node15137;
															assign node15137 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15140 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node15143 = (inp[12]) ? 4'b1101 : node15144;
															assign node15144 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node15148 = (inp[7]) ? node15156 : node15149;
														assign node15149 = (inp[10]) ? node15153 : node15150;
															assign node15150 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node15153 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node15156 = (inp[14]) ? node15158 : 4'b0000;
															assign node15158 = (inp[10]) ? node15162 : node15159;
																assign node15159 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node15162 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node15165 = (inp[7]) ? node15175 : node15166;
													assign node15166 = (inp[12]) ? node15172 : node15167;
														assign node15167 = (inp[10]) ? 4'b0001 : node15168;
															assign node15168 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node15172 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node15175 = (inp[12]) ? 4'b1101 : node15176;
														assign node15176 = (inp[10]) ? node15178 : 4'b1101;
															assign node15178 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node15182 = (inp[4]) ? node15212 : node15183;
												assign node15183 = (inp[2]) ? node15199 : node15184;
													assign node15184 = (inp[7]) ? node15192 : node15185;
														assign node15185 = (inp[10]) ? node15189 : node15186;
															assign node15186 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node15189 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15192 = (inp[10]) ? node15196 : node15193;
															assign node15193 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node15196 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node15199 = (inp[7]) ? node15207 : node15200;
														assign node15200 = (inp[12]) ? node15204 : node15201;
															assign node15201 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15204 = (inp[10]) ? 4'b0000 : 4'b1001;
														assign node15207 = (inp[10]) ? node15209 : 4'b1001;
															assign node15209 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node15212 = (inp[2]) ? node15220 : node15213;
													assign node15213 = (inp[10]) ? 4'b1001 : node15214;
														assign node15214 = (inp[12]) ? node15216 : 4'b0001;
															assign node15216 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node15220 = (inp[7]) ? node15228 : node15221;
														assign node15221 = (inp[12]) ? node15225 : node15222;
															assign node15222 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node15225 = (inp[14]) ? 4'b0100 : 4'b1000;
														assign node15228 = (inp[14]) ? node15230 : 4'b1000;
															assign node15230 = (inp[10]) ? node15234 : node15231;
																assign node15231 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node15234 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node15237 = (inp[4]) ? node15289 : node15238;
											assign node15238 = (inp[3]) ? node15272 : node15239;
												assign node15239 = (inp[2]) ? node15261 : node15240;
													assign node15240 = (inp[7]) ? node15254 : node15241;
														assign node15241 = (inp[14]) ? node15247 : node15242;
															assign node15242 = (inp[12]) ? 4'b1000 : node15243;
																assign node15243 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15247 = (inp[12]) ? node15251 : node15248;
																assign node15248 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node15251 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node15254 = (inp[12]) ? node15258 : node15255;
															assign node15255 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15258 = (inp[10]) ? 4'b0000 : 4'b0101;
													assign node15261 = (inp[7]) ? node15267 : node15262;
														assign node15262 = (inp[10]) ? node15264 : 4'b0001;
															assign node15264 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15267 = (inp[10]) ? node15269 : 4'b0101;
															assign node15269 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node15272 = (inp[10]) ? node15280 : node15273;
													assign node15273 = (inp[12]) ? node15275 : 4'b0000;
														assign node15275 = (inp[7]) ? node15277 : 4'b1000;
															assign node15277 = (inp[2]) ? 4'b0001 : 4'b1100;
													assign node15280 = (inp[7]) ? node15286 : node15281;
														assign node15281 = (inp[2]) ? node15283 : 4'b0001;
															assign node15283 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15286 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node15289 = (inp[3]) ? node15305 : node15290;
												assign node15290 = (inp[2]) ? node15300 : node15291;
													assign node15291 = (inp[10]) ? node15297 : node15292;
														assign node15292 = (inp[12]) ? node15294 : 4'b0100;
															assign node15294 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node15297 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node15300 = (inp[10]) ? node15302 : 4'b0001;
														assign node15302 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node15305 = (inp[2]) ? node15315 : node15306;
													assign node15306 = (inp[10]) ? 4'b0101 : node15307;
														assign node15307 = (inp[7]) ? node15311 : node15308;
															assign node15308 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node15311 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15315 = (inp[12]) ? node15319 : node15316;
														assign node15316 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node15319 = (inp[10]) ? 4'b0100 : node15320;
															assign node15320 = (inp[7]) ? 4'b1000 : 4'b1100;
									assign node15324 = (inp[10]) ? node15404 : node15325;
										assign node15325 = (inp[4]) ? node15357 : node15326;
											assign node15326 = (inp[3]) ? node15346 : node15327;
												assign node15327 = (inp[7]) ? node15337 : node15328;
													assign node15328 = (inp[2]) ? node15330 : 4'b0000;
														assign node15330 = (inp[12]) ? node15334 : node15331;
															assign node15331 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node15334 = (inp[13]) ? 4'b0000 : 4'b1100;
													assign node15337 = (inp[13]) ? node15341 : node15338;
														assign node15338 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node15341 = (inp[2]) ? node15343 : 4'b0000;
															assign node15343 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node15346 = (inp[13]) ? 4'b0000 : node15347;
													assign node15347 = (inp[2]) ? node15351 : node15348;
														assign node15348 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node15351 = (inp[12]) ? node15353 : 4'b0000;
															assign node15353 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node15357 = (inp[13]) ? node15391 : node15358;
												assign node15358 = (inp[7]) ? node15380 : node15359;
													assign node15359 = (inp[14]) ? node15369 : node15360;
														assign node15360 = (inp[12]) ? node15362 : 4'b0100;
															assign node15362 = (inp[2]) ? node15366 : node15363;
																assign node15363 = (inp[3]) ? 4'b0000 : 4'b0100;
																assign node15366 = (inp[3]) ? 4'b0100 : 4'b1000;
														assign node15369 = (inp[12]) ? node15373 : node15370;
															assign node15370 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node15373 = (inp[2]) ? node15377 : node15374;
																assign node15374 = (inp[3]) ? 4'b0000 : 4'b0100;
																assign node15377 = (inp[3]) ? 4'b0100 : 4'b1000;
													assign node15380 = (inp[3]) ? node15386 : node15381;
														assign node15381 = (inp[2]) ? node15383 : 4'b0000;
															assign node15383 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node15386 = (inp[12]) ? 4'b0000 : node15387;
															assign node15387 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node15391 = (inp[3]) ? node15397 : node15392;
													assign node15392 = (inp[2]) ? node15394 : 4'b0100;
														assign node15394 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node15397 = (inp[2]) ? 4'b0100 : node15398;
														assign node15398 = (inp[12]) ? node15400 : 4'b0100;
															assign node15400 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node15404 = (inp[13]) ? node15432 : node15405;
											assign node15405 = (inp[2]) ? node15419 : node15406;
												assign node15406 = (inp[7]) ? node15412 : node15407;
													assign node15407 = (inp[4]) ? node15409 : 4'b1000;
														assign node15409 = (inp[3]) ? 4'b0100 : 4'b1100;
													assign node15412 = (inp[4]) ? node15416 : node15413;
														assign node15413 = (inp[3]) ? 4'b1100 : 4'b0100;
														assign node15416 = (inp[3]) ? 4'b0000 : 4'b1000;
												assign node15419 = (inp[3]) ? node15425 : node15420;
													assign node15420 = (inp[7]) ? node15422 : 4'b0000;
														assign node15422 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node15425 = (inp[7]) ? node15429 : node15426;
														assign node15426 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node15429 = (inp[4]) ? 4'b1000 : 4'b0000;
											assign node15432 = (inp[4]) ? node15440 : node15433;
												assign node15433 = (inp[2]) ? node15435 : 4'b1000;
													assign node15435 = (inp[3]) ? 4'b1000 : node15436;
														assign node15436 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node15440 = (inp[2]) ? node15442 : 4'b1100;
													assign node15442 = (inp[3]) ? 4'b1100 : 4'b1000;
							assign node15445 = (inp[2]) ? 4'b1100 : node15446;
								assign node15446 = (inp[1]) ? node15612 : node15447;
									assign node15447 = (inp[13]) ? node15529 : node15448;
										assign node15448 = (inp[3]) ? node15488 : node15449;
											assign node15449 = (inp[7]) ? node15477 : node15450;
												assign node15450 = (inp[4]) ? node15460 : node15451;
													assign node15451 = (inp[10]) ? node15453 : 4'b1100;
														assign node15453 = (inp[12]) ? 4'b1100 : node15454;
															assign node15454 = (inp[11]) ? 4'b0001 : node15455;
																assign node15455 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node15460 = (inp[14]) ? node15466 : node15461;
														assign node15461 = (inp[10]) ? node15463 : 4'b1001;
															assign node15463 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node15466 = (inp[11]) ? node15472 : node15467;
															assign node15467 = (inp[10]) ? node15469 : 4'b1000;
																assign node15469 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node15472 = (inp[12]) ? 4'b1001 : node15473;
																assign node15473 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node15477 = (inp[12]) ? 4'b1100 : node15478;
													assign node15478 = (inp[10]) ? node15480 : 4'b1100;
														assign node15480 = (inp[4]) ? node15482 : 4'b1100;
															assign node15482 = (inp[14]) ? node15484 : 4'b0001;
																assign node15484 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node15488 = (inp[10]) ? node15506 : node15489;
												assign node15489 = (inp[14]) ? node15495 : node15490;
													assign node15490 = (inp[4]) ? node15492 : 4'b1001;
														assign node15492 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node15495 = (inp[11]) ? node15501 : node15496;
														assign node15496 = (inp[7]) ? 4'b1000 : node15497;
															assign node15497 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node15501 = (inp[4]) ? node15503 : 4'b1001;
															assign node15503 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node15506 = (inp[12]) ? node15518 : node15507;
													assign node15507 = (inp[4]) ? node15513 : node15508;
														assign node15508 = (inp[7]) ? node15510 : 4'b0101;
															assign node15510 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node15513 = (inp[14]) ? node15515 : 4'b0101;
															assign node15515 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node15518 = (inp[7]) ? node15524 : node15519;
														assign node15519 = (inp[4]) ? 4'b1101 : node15520;
															assign node15520 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15524 = (inp[11]) ? 4'b1001 : node15525;
															assign node15525 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node15529 = (inp[3]) ? node15561 : node15530;
											assign node15530 = (inp[7]) ? node15548 : node15531;
												assign node15531 = (inp[10]) ? node15537 : node15532;
													assign node15532 = (inp[14]) ? node15534 : 4'b0001;
														assign node15534 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node15537 = (inp[12]) ? node15543 : node15538;
														assign node15538 = (inp[14]) ? node15540 : 4'b1001;
															assign node15540 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15543 = (inp[14]) ? node15545 : 4'b0001;
															assign node15545 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node15548 = (inp[4]) ? node15550 : 4'b1100;
													assign node15550 = (inp[12]) ? node15556 : node15551;
														assign node15551 = (inp[10]) ? node15553 : 4'b0001;
															assign node15553 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15556 = (inp[11]) ? 4'b0001 : node15557;
															assign node15557 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node15561 = (inp[7]) ? node15579 : node15562;
												assign node15562 = (inp[12]) ? node15574 : node15563;
													assign node15563 = (inp[10]) ? node15569 : node15564;
														assign node15564 = (inp[14]) ? node15566 : 4'b0101;
															assign node15566 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node15569 = (inp[11]) ? 4'b1101 : node15570;
															assign node15570 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node15574 = (inp[14]) ? node15576 : 4'b0101;
														assign node15576 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node15579 = (inp[4]) ? node15597 : node15580;
													assign node15580 = (inp[11]) ? node15592 : node15581;
														assign node15581 = (inp[14]) ? node15587 : node15582;
															assign node15582 = (inp[10]) ? node15584 : 4'b0001;
																assign node15584 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node15587 = (inp[12]) ? 4'b0000 : node15588;
																assign node15588 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node15592 = (inp[10]) ? node15594 : 4'b0001;
															assign node15594 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15597 = (inp[14]) ? node15603 : node15598;
														assign node15598 = (inp[10]) ? node15600 : 4'b0101;
															assign node15600 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node15603 = (inp[11]) ? node15609 : node15604;
															assign node15604 = (inp[12]) ? 4'b0100 : node15605;
																assign node15605 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node15609 = (inp[12]) ? 4'b0101 : 4'b1101;
									assign node15612 = (inp[14]) ? node15680 : node15613;
										assign node15613 = (inp[13]) ? node15649 : node15614;
											assign node15614 = (inp[10]) ? node15638 : node15615;
												assign node15615 = (inp[12]) ? node15627 : node15616;
													assign node15616 = (inp[3]) ? node15622 : node15617;
														assign node15617 = (inp[7]) ? node15619 : 4'b0000;
															assign node15619 = (inp[4]) ? 4'b0000 : 4'b1100;
														assign node15622 = (inp[4]) ? 4'b0100 : node15623;
															assign node15623 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node15627 = (inp[3]) ? node15633 : node15628;
														assign node15628 = (inp[7]) ? 4'b1100 : node15629;
															assign node15629 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node15633 = (inp[7]) ? 4'b1000 : node15634;
															assign node15634 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node15638 = (inp[3]) ? node15644 : node15639;
													assign node15639 = (inp[4]) ? 4'b0000 : node15640;
														assign node15640 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node15644 = (inp[4]) ? 4'b0100 : node15645;
														assign node15645 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node15649 = (inp[3]) ? node15663 : node15650;
												assign node15650 = (inp[7]) ? node15656 : node15651;
													assign node15651 = (inp[12]) ? node15653 : 4'b1000;
														assign node15653 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node15656 = (inp[4]) ? node15658 : 4'b1100;
														assign node15658 = (inp[10]) ? 4'b1000 : node15659;
															assign node15659 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node15663 = (inp[12]) ? node15669 : node15664;
													assign node15664 = (inp[4]) ? 4'b1100 : node15665;
														assign node15665 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node15669 = (inp[10]) ? node15675 : node15670;
														assign node15670 = (inp[4]) ? 4'b0100 : node15671;
															assign node15671 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node15675 = (inp[4]) ? 4'b1100 : node15676;
															assign node15676 = (inp[7]) ? 4'b1000 : 4'b1100;
										assign node15680 = (inp[11]) ? node15742 : node15681;
											assign node15681 = (inp[13]) ? node15715 : node15682;
												assign node15682 = (inp[3]) ? node15702 : node15683;
													assign node15683 = (inp[7]) ? node15695 : node15684;
														assign node15684 = (inp[4]) ? node15690 : node15685;
															assign node15685 = (inp[10]) ? node15687 : 4'b1100;
																assign node15687 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node15690 = (inp[12]) ? 4'b1001 : node15691;
																assign node15691 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node15695 = (inp[4]) ? node15697 : 4'b1100;
															assign node15697 = (inp[12]) ? 4'b1100 : node15698;
																assign node15698 = (inp[10]) ? 4'b0001 : 4'b1100;
													assign node15702 = (inp[4]) ? node15708 : node15703;
														assign node15703 = (inp[10]) ? node15705 : 4'b1001;
															assign node15705 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node15708 = (inp[12]) ? node15712 : node15709;
															assign node15709 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node15712 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node15715 = (inp[3]) ? node15725 : node15716;
													assign node15716 = (inp[7]) ? node15722 : node15717;
														assign node15717 = (inp[10]) ? node15719 : 4'b0001;
															assign node15719 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15722 = (inp[4]) ? 4'b0001 : 4'b1100;
													assign node15725 = (inp[10]) ? node15731 : node15726;
														assign node15726 = (inp[7]) ? node15728 : 4'b0101;
															assign node15728 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node15731 = (inp[12]) ? node15737 : node15732;
															assign node15732 = (inp[7]) ? node15734 : 4'b1101;
																assign node15734 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node15737 = (inp[4]) ? 4'b0101 : node15738;
																assign node15738 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node15742 = (inp[13]) ? node15772 : node15743;
												assign node15743 = (inp[10]) ? node15761 : node15744;
													assign node15744 = (inp[12]) ? node15754 : node15745;
														assign node15745 = (inp[3]) ? node15749 : node15746;
															assign node15746 = (inp[7]) ? 4'b1100 : 4'b0000;
															assign node15749 = (inp[7]) ? node15751 : 4'b0100;
																assign node15751 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node15754 = (inp[3]) ? node15756 : 4'b1100;
															assign node15756 = (inp[4]) ? node15758 : 4'b1000;
																assign node15758 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node15761 = (inp[3]) ? node15767 : node15762;
														assign node15762 = (inp[4]) ? 4'b0000 : node15763;
															assign node15763 = (inp[7]) ? 4'b1100 : 4'b0000;
														assign node15767 = (inp[4]) ? 4'b0100 : node15768;
															assign node15768 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node15772 = (inp[3]) ? node15782 : node15773;
													assign node15773 = (inp[7]) ? node15779 : node15774;
														assign node15774 = (inp[12]) ? node15776 : 4'b1000;
															assign node15776 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node15779 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node15782 = (inp[7]) ? node15788 : node15783;
														assign node15783 = (inp[12]) ? node15785 : 4'b1100;
															assign node15785 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node15788 = (inp[4]) ? node15794 : node15789;
															assign node15789 = (inp[10]) ? 4'b1000 : node15790;
																assign node15790 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15794 = (inp[12]) ? node15796 : 4'b1100;
																assign node15796 = (inp[10]) ? 4'b1100 : 4'b0100;
						assign node15800 = (inp[3]) ? node16600 : node15801;
							assign node15801 = (inp[4]) ? node16177 : node15802;
								assign node15802 = (inp[7]) ? node16002 : node15803;
									assign node15803 = (inp[1]) ? node15903 : node15804;
										assign node15804 = (inp[2]) ? node15844 : node15805;
											assign node15805 = (inp[0]) ? node15827 : node15806;
												assign node15806 = (inp[13]) ? node15816 : node15807;
													assign node15807 = (inp[12]) ? node15809 : 4'b0000;
														assign node15809 = (inp[11]) ? 4'b0000 : node15810;
															assign node15810 = (inp[10]) ? 4'b1000 : node15811;
																assign node15811 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node15816 = (inp[12]) ? node15822 : node15817;
														assign node15817 = (inp[11]) ? node15819 : 4'b0100;
															assign node15819 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node15822 = (inp[11]) ? 4'b0100 : node15823;
															assign node15823 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node15827 = (inp[11]) ? node15835 : node15828;
													assign node15828 = (inp[10]) ? 4'b0001 : node15829;
														assign node15829 = (inp[13]) ? 4'b1001 : node15830;
															assign node15830 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node15835 = (inp[12]) ? node15839 : node15836;
														assign node15836 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node15839 = (inp[10]) ? 4'b0000 : node15840;
															assign node15840 = (inp[13]) ? 4'b1000 : 4'b1101;
											assign node15844 = (inp[13]) ? node15870 : node15845;
												assign node15845 = (inp[10]) ? node15855 : node15846;
													assign node15846 = (inp[0]) ? 4'b1100 : node15847;
														assign node15847 = (inp[14]) ? node15851 : node15848;
															assign node15848 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node15851 = (inp[11]) ? 4'b0001 : 4'b1101;
													assign node15855 = (inp[0]) ? node15863 : node15856;
														assign node15856 = (inp[11]) ? 4'b1001 : node15857;
															assign node15857 = (inp[14]) ? node15859 : 4'b1000;
																assign node15859 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15863 = (inp[12]) ? 4'b1100 : node15864;
															assign node15864 = (inp[11]) ? 4'b0001 : node15865;
																assign node15865 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node15870 = (inp[0]) ? node15890 : node15871;
													assign node15871 = (inp[10]) ? node15883 : node15872;
														assign node15872 = (inp[14]) ? node15878 : node15873;
															assign node15873 = (inp[12]) ? node15875 : 4'b1000;
																assign node15875 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node15878 = (inp[11]) ? node15880 : 4'b0001;
																assign node15880 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node15883 = (inp[11]) ? 4'b0101 : node15884;
															assign node15884 = (inp[14]) ? node15886 : 4'b0100;
																assign node15886 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node15890 = (inp[12]) ? node15898 : node15891;
														assign node15891 = (inp[10]) ? node15893 : 4'b0001;
															assign node15893 = (inp[11]) ? 4'b1001 : node15894;
																assign node15894 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15898 = (inp[11]) ? 4'b0001 : node15899;
															assign node15899 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node15903 = (inp[11]) ? node15971 : node15904;
											assign node15904 = (inp[0]) ? node15944 : node15905;
												assign node15905 = (inp[13]) ? node15921 : node15906;
													assign node15906 = (inp[2]) ? node15910 : node15907;
														assign node15907 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node15910 = (inp[14]) ? node15916 : node15911;
															assign node15911 = (inp[10]) ? node15913 : 4'b0001;
																assign node15913 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node15916 = (inp[10]) ? node15918 : 4'b0000;
																assign node15918 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node15921 = (inp[12]) ? node15933 : node15922;
														assign node15922 = (inp[10]) ? node15928 : node15923;
															assign node15923 = (inp[2]) ? node15925 : 4'b1100;
																assign node15925 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node15928 = (inp[2]) ? 4'b1101 : node15929;
																assign node15929 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node15933 = (inp[2]) ? node15939 : node15934;
															assign node15934 = (inp[10]) ? node15936 : 4'b0100;
																assign node15936 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node15939 = (inp[10]) ? 4'b0100 : node15940;
																assign node15940 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node15944 = (inp[2]) ? node15956 : node15945;
													assign node15945 = (inp[10]) ? node15953 : node15946;
														assign node15946 = (inp[12]) ? node15948 : 4'b0001;
															assign node15948 = (inp[13]) ? 4'b1001 : node15949;
																assign node15949 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node15953 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node15956 = (inp[13]) ? node15960 : node15957;
														assign node15957 = (inp[14]) ? 4'b1100 : 4'b0000;
														assign node15960 = (inp[14]) ? node15966 : node15961;
															assign node15961 = (inp[12]) ? node15963 : 4'b1000;
																assign node15963 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node15966 = (inp[12]) ? 4'b0001 : node15967;
																assign node15967 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node15971 = (inp[13]) ? node15987 : node15972;
												assign node15972 = (inp[2]) ? node15978 : node15973;
													assign node15973 = (inp[0]) ? node15975 : 4'b1000;
														assign node15975 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node15978 = (inp[10]) ? 4'b0000 : node15979;
														assign node15979 = (inp[0]) ? node15983 : node15980;
															assign node15980 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node15983 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node15987 = (inp[0]) ? node15997 : node15988;
													assign node15988 = (inp[10]) ? node15994 : node15989;
														assign node15989 = (inp[2]) ? node15991 : 4'b1100;
															assign node15991 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node15994 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node15997 = (inp[10]) ? 4'b1000 : node15998;
														assign node15998 = (inp[2]) ? 4'b1000 : 4'b0000;
									assign node16002 = (inp[0]) ? node16110 : node16003;
										assign node16003 = (inp[13]) ? node16055 : node16004;
											assign node16004 = (inp[10]) ? node16032 : node16005;
												assign node16005 = (inp[11]) ? node16021 : node16006;
													assign node16006 = (inp[2]) ? node16016 : node16007;
														assign node16007 = (inp[1]) ? node16013 : node16008;
															assign node16008 = (inp[14]) ? 4'b1101 : node16009;
																assign node16009 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node16013 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node16016 = (inp[1]) ? node16018 : 4'b1101;
															assign node16018 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node16021 = (inp[2]) ? node16029 : node16022;
														assign node16022 = (inp[1]) ? node16026 : node16023;
															assign node16023 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node16026 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node16029 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node16032 = (inp[2]) ? node16044 : node16033;
													assign node16033 = (inp[1]) ? node16039 : node16034;
														assign node16034 = (inp[12]) ? node16036 : 4'b0000;
															assign node16036 = (inp[11]) ? 4'b0000 : 4'b0101;
														assign node16039 = (inp[12]) ? node16041 : 4'b1000;
															assign node16041 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node16044 = (inp[11]) ? node16052 : node16045;
														assign node16045 = (inp[12]) ? 4'b0101 : node16046;
															assign node16046 = (inp[1]) ? node16048 : 4'b0101;
																assign node16048 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node16052 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node16055 = (inp[2]) ? node16079 : node16056;
												assign node16056 = (inp[10]) ? node16068 : node16057;
													assign node16057 = (inp[1]) ? node16063 : node16058;
														assign node16058 = (inp[11]) ? 4'b0000 : node16059;
															assign node16059 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16063 = (inp[11]) ? 4'b1000 : node16064;
															assign node16064 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16068 = (inp[1]) ? node16074 : node16069;
														assign node16069 = (inp[11]) ? 4'b0100 : node16070;
															assign node16070 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node16074 = (inp[11]) ? 4'b1100 : node16075;
															assign node16075 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node16079 = (inp[1]) ? node16097 : node16080;
													assign node16080 = (inp[11]) ? node16092 : node16081;
														assign node16081 = (inp[14]) ? node16087 : node16082;
															assign node16082 = (inp[12]) ? 4'b0000 : node16083;
																assign node16083 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node16087 = (inp[10]) ? node16089 : 4'b0001;
																assign node16089 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16092 = (inp[10]) ? 4'b0001 : node16093;
															assign node16093 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16097 = (inp[11]) ? node16105 : node16098;
														assign node16098 = (inp[14]) ? node16102 : node16099;
															assign node16099 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node16102 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16105 = (inp[12]) ? 4'b1000 : node16106;
															assign node16106 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node16110 = (inp[2]) ? 4'b1100 : node16111;
											assign node16111 = (inp[13]) ? node16145 : node16112;
												assign node16112 = (inp[1]) ? node16130 : node16113;
													assign node16113 = (inp[10]) ? node16119 : node16114;
														assign node16114 = (inp[11]) ? 4'b1101 : node16115;
															assign node16115 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node16119 = (inp[12]) ? node16125 : node16120;
															assign node16120 = (inp[14]) ? node16122 : 4'b0101;
																assign node16122 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node16125 = (inp[11]) ? 4'b1101 : node16126;
																assign node16126 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node16130 = (inp[14]) ? node16136 : node16131;
														assign node16131 = (inp[10]) ? 4'b0100 : node16132;
															assign node16132 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node16136 = (inp[11]) ? node16142 : node16137;
															assign node16137 = (inp[12]) ? 4'b1101 : node16138;
																assign node16138 = (inp[10]) ? 4'b0101 : 4'b1101;
															assign node16142 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node16145 = (inp[11]) ? node16165 : node16146;
													assign node16146 = (inp[10]) ? node16160 : node16147;
														assign node16147 = (inp[12]) ? node16153 : node16148;
															assign node16148 = (inp[1]) ? 4'b0001 : node16149;
																assign node16149 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node16153 = (inp[14]) ? node16157 : node16154;
																assign node16154 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node16157 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node16160 = (inp[12]) ? 4'b0001 : node16161;
															assign node16161 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node16165 = (inp[10]) ? node16171 : node16166;
														assign node16166 = (inp[12]) ? node16168 : 4'b0000;
															assign node16168 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node16171 = (inp[1]) ? 4'b1000 : node16172;
															assign node16172 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node16177 = (inp[1]) ? node16411 : node16178;
									assign node16178 = (inp[0]) ? node16310 : node16179;
										assign node16179 = (inp[2]) ? node16249 : node16180;
											assign node16180 = (inp[13]) ? node16216 : node16181;
												assign node16181 = (inp[11]) ? node16207 : node16182;
													assign node16182 = (inp[14]) ? node16194 : node16183;
														assign node16183 = (inp[12]) ? node16189 : node16184;
															assign node16184 = (inp[7]) ? 4'b0001 : node16185;
																assign node16185 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node16189 = (inp[10]) ? node16191 : 4'b1100;
																assign node16191 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16194 = (inp[12]) ? node16200 : node16195;
															assign node16195 = (inp[7]) ? 4'b0000 : node16196;
																assign node16196 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node16200 = (inp[10]) ? node16204 : node16201;
																assign node16201 = (inp[7]) ? 4'b1100 : 4'b1000;
																assign node16204 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node16207 = (inp[10]) ? node16209 : 4'b0001;
														assign node16209 = (inp[7]) ? node16213 : node16210;
															assign node16210 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node16213 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node16216 = (inp[11]) ? node16236 : node16217;
													assign node16217 = (inp[12]) ? node16225 : node16218;
														assign node16218 = (inp[10]) ? node16220 : 4'b0001;
															assign node16220 = (inp[7]) ? 4'b1001 : node16221;
																assign node16221 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node16225 = (inp[7]) ? node16231 : node16226;
															assign node16226 = (inp[10]) ? node16228 : 4'b1001;
																assign node16228 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node16231 = (inp[10]) ? 4'b0001 : node16232;
																assign node16232 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node16236 = (inp[7]) ? node16242 : node16237;
														assign node16237 = (inp[10]) ? 4'b1001 : node16238;
															assign node16238 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16242 = (inp[12]) ? node16246 : node16243;
															assign node16243 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node16246 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node16249 = (inp[11]) ? node16285 : node16250;
												assign node16250 = (inp[12]) ? node16266 : node16251;
													assign node16251 = (inp[13]) ? node16257 : node16252;
														assign node16252 = (inp[10]) ? 4'b0000 : node16253;
															assign node16253 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node16257 = (inp[7]) ? node16263 : node16258;
															assign node16258 = (inp[10]) ? node16260 : 4'b0100;
																assign node16260 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node16263 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node16266 = (inp[13]) ? node16280 : node16267;
														assign node16267 = (inp[14]) ? node16273 : node16268;
															assign node16268 = (inp[10]) ? 4'b1000 : node16269;
																assign node16269 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node16273 = (inp[10]) ? node16277 : node16274;
																assign node16274 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node16277 = (inp[7]) ? 4'b0101 : 4'b1000;
														assign node16280 = (inp[7]) ? 4'b1000 : node16281;
															assign node16281 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node16285 = (inp[12]) ? node16297 : node16286;
													assign node16286 = (inp[10]) ? node16294 : node16287;
														assign node16287 = (inp[7]) ? node16291 : node16288;
															assign node16288 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node16291 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node16294 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node16297 = (inp[13]) ? node16303 : node16298;
														assign node16298 = (inp[10]) ? 4'b0000 : node16299;
															assign node16299 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node16303 = (inp[7]) ? node16307 : node16304;
															assign node16304 = (inp[10]) ? 4'b1001 : 4'b0100;
															assign node16307 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node16310 = (inp[13]) ? node16356 : node16311;
											assign node16311 = (inp[10]) ? node16331 : node16312;
												assign node16312 = (inp[7]) ? node16324 : node16313;
													assign node16313 = (inp[2]) ? node16319 : node16314;
														assign node16314 = (inp[11]) ? node16316 : 4'b1001;
															assign node16316 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node16319 = (inp[11]) ? 4'b1001 : node16320;
															assign node16320 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node16324 = (inp[2]) ? 4'b1100 : node16325;
														assign node16325 = (inp[11]) ? node16327 : 4'b1001;
															assign node16327 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node16331 = (inp[2]) ? node16343 : node16332;
													assign node16332 = (inp[11]) ? node16336 : node16333;
														assign node16333 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node16336 = (inp[7]) ? node16340 : node16337;
															assign node16337 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node16340 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16343 = (inp[12]) ? node16349 : node16344;
														assign node16344 = (inp[14]) ? node16346 : 4'b0001;
															assign node16346 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node16349 = (inp[7]) ? 4'b1100 : node16350;
															assign node16350 = (inp[11]) ? 4'b1001 : node16351;
																assign node16351 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node16356 = (inp[11]) ? node16390 : node16357;
												assign node16357 = (inp[12]) ? node16373 : node16358;
													assign node16358 = (inp[14]) ? node16368 : node16359;
														assign node16359 = (inp[2]) ? node16365 : node16360;
															assign node16360 = (inp[10]) ? 4'b0000 : node16361;
																assign node16361 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node16365 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node16368 = (inp[2]) ? node16370 : 4'b0001;
															assign node16370 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node16373 = (inp[2]) ? node16387 : node16374;
														assign node16374 = (inp[14]) ? node16380 : node16375;
															assign node16375 = (inp[10]) ? 4'b0000 : node16376;
																assign node16376 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node16380 = (inp[10]) ? node16384 : node16381;
																assign node16381 = (inp[7]) ? 4'b1001 : 4'b0001;
																assign node16384 = (inp[7]) ? 4'b0101 : 4'b1001;
														assign node16387 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node16390 = (inp[7]) ? node16400 : node16391;
													assign node16391 = (inp[12]) ? 4'b0001 : node16392;
														assign node16392 = (inp[10]) ? node16396 : node16393;
															assign node16393 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node16396 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node16400 = (inp[10]) ? node16406 : node16401;
														assign node16401 = (inp[2]) ? 4'b0001 : node16402;
															assign node16402 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node16406 = (inp[2]) ? node16408 : 4'b0001;
															assign node16408 = (inp[12]) ? 4'b0001 : 4'b1001;
									assign node16411 = (inp[11]) ? node16539 : node16412;
										assign node16412 = (inp[2]) ? node16476 : node16413;
											assign node16413 = (inp[10]) ? node16441 : node16414;
												assign node16414 = (inp[0]) ? node16424 : node16415;
													assign node16415 = (inp[14]) ? node16419 : node16416;
														assign node16416 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node16419 = (inp[12]) ? node16421 : 4'b1001;
															assign node16421 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node16424 = (inp[12]) ? node16434 : node16425;
														assign node16425 = (inp[13]) ? node16429 : node16426;
															assign node16426 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node16429 = (inp[7]) ? 4'b0101 : node16430;
																assign node16430 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node16434 = (inp[13]) ? node16436 : 4'b1001;
															assign node16436 = (inp[14]) ? node16438 : 4'b1001;
																assign node16438 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node16441 = (inp[14]) ? node16463 : node16442;
													assign node16442 = (inp[7]) ? node16454 : node16443;
														assign node16443 = (inp[12]) ? node16449 : node16444;
															assign node16444 = (inp[0]) ? node16446 : 4'b0001;
																assign node16446 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node16449 = (inp[13]) ? 4'b0001 : node16450;
																assign node16450 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node16454 = (inp[0]) ? node16460 : node16455;
															assign node16455 = (inp[13]) ? 4'b0001 : node16456;
																assign node16456 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node16460 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16463 = (inp[13]) ? node16471 : node16464;
														assign node16464 = (inp[7]) ? node16468 : node16465;
															assign node16465 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node16468 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16471 = (inp[0]) ? node16473 : 4'b0000;
															assign node16473 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node16476 = (inp[14]) ? node16512 : node16477;
												assign node16477 = (inp[13]) ? node16499 : node16478;
													assign node16478 = (inp[7]) ? node16488 : node16479;
														assign node16479 = (inp[10]) ? 4'b0000 : node16480;
															assign node16480 = (inp[12]) ? node16484 : node16481;
																assign node16481 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node16484 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node16488 = (inp[10]) ? node16494 : node16489;
															assign node16489 = (inp[0]) ? node16491 : 4'b0101;
																assign node16491 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node16494 = (inp[0]) ? 4'b0000 : node16495;
																assign node16495 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16499 = (inp[12]) ? node16507 : node16500;
														assign node16500 = (inp[10]) ? 4'b1000 : node16501;
															assign node16501 = (inp[7]) ? 4'b1000 : node16502;
																assign node16502 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node16507 = (inp[10]) ? node16509 : 4'b0000;
															assign node16509 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node16512 = (inp[13]) ? node16524 : node16513;
													assign node16513 = (inp[0]) ? node16519 : node16514;
														assign node16514 = (inp[12]) ? 4'b0000 : node16515;
															assign node16515 = (inp[10]) ? 4'b1000 : 4'b0100;
														assign node16519 = (inp[7]) ? node16521 : 4'b1001;
															assign node16521 = (inp[10]) ? 4'b0001 : 4'b1100;
													assign node16524 = (inp[10]) ? node16534 : node16525;
														assign node16525 = (inp[0]) ? 4'b0001 : node16526;
															assign node16526 = (inp[7]) ? node16530 : node16527;
																assign node16527 = (inp[12]) ? 4'b0100 : 4'b0001;
																assign node16530 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16534 = (inp[0]) ? node16536 : 4'b0001;
															assign node16536 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node16539 = (inp[10]) ? node16587 : node16540;
											assign node16540 = (inp[2]) ? node16560 : node16541;
												assign node16541 = (inp[12]) ? node16547 : node16542;
													assign node16542 = (inp[13]) ? 4'b0000 : node16543;
														assign node16543 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node16547 = (inp[0]) ? node16553 : node16548;
														assign node16548 = (inp[13]) ? node16550 : 4'b1000;
															assign node16550 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node16553 = (inp[13]) ? node16557 : node16554;
															assign node16554 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node16557 = (inp[7]) ? 4'b0100 : 4'b1000;
												assign node16560 = (inp[7]) ? node16574 : node16561;
													assign node16561 = (inp[0]) ? node16567 : node16562;
														assign node16562 = (inp[13]) ? node16564 : 4'b1000;
															assign node16564 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16567 = (inp[13]) ? node16571 : node16568;
															assign node16568 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node16571 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16574 = (inp[13]) ? node16582 : node16575;
														assign node16575 = (inp[12]) ? node16579 : node16576;
															assign node16576 = (inp[0]) ? 4'b0000 : 4'b1100;
															assign node16579 = (inp[0]) ? 4'b1100 : 4'b0100;
														assign node16582 = (inp[0]) ? node16584 : 4'b1000;
															assign node16584 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node16587 = (inp[13]) ? 4'b1000 : node16588;
												assign node16588 = (inp[0]) ? node16594 : node16589;
													assign node16589 = (inp[7]) ? node16591 : 4'b1000;
														assign node16591 = (inp[2]) ? 4'b1000 : 4'b0100;
													assign node16594 = (inp[2]) ? 4'b0000 : node16595;
														assign node16595 = (inp[7]) ? 4'b1000 : 4'b0000;
							assign node16600 = (inp[4]) ? node17058 : node16601;
								assign node16601 = (inp[11]) ? node16885 : node16602;
									assign node16602 = (inp[2]) ? node16740 : node16603;
										assign node16603 = (inp[13]) ? node16679 : node16604;
											assign node16604 = (inp[14]) ? node16640 : node16605;
												assign node16605 = (inp[10]) ? node16619 : node16606;
													assign node16606 = (inp[0]) ? node16608 : 4'b0000;
														assign node16608 = (inp[12]) ? node16616 : node16609;
															assign node16609 = (inp[7]) ? node16613 : node16610;
																assign node16610 = (inp[1]) ? 4'b1000 : 4'b0000;
																assign node16613 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node16616 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node16619 = (inp[0]) ? node16627 : node16620;
														assign node16620 = (inp[1]) ? 4'b1000 : node16621;
															assign node16621 = (inp[7]) ? 4'b0000 : node16622;
																assign node16622 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16627 = (inp[7]) ? node16633 : node16628;
															assign node16628 = (inp[12]) ? node16630 : 4'b0000;
																assign node16630 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node16633 = (inp[12]) ? node16637 : node16634;
																assign node16634 = (inp[1]) ? 4'b1000 : 4'b0000;
																assign node16637 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node16640 = (inp[0]) ? node16658 : node16641;
													assign node16641 = (inp[10]) ? node16649 : node16642;
														assign node16642 = (inp[7]) ? node16644 : 4'b0000;
															assign node16644 = (inp[1]) ? 4'b0000 : node16645;
																assign node16645 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node16649 = (inp[1]) ? node16653 : node16650;
															assign node16650 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node16653 = (inp[7]) ? node16655 : 4'b0001;
																assign node16655 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node16658 = (inp[1]) ? node16672 : node16659;
														assign node16659 = (inp[10]) ? node16665 : node16660;
															assign node16660 = (inp[7]) ? 4'b1001 : node16661;
																assign node16661 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node16665 = (inp[7]) ? node16669 : node16666;
																assign node16666 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node16669 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node16672 = (inp[12]) ? 4'b0000 : node16673;
															assign node16673 = (inp[7]) ? node16675 : 4'b1000;
																assign node16675 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node16679 = (inp[10]) ? node16711 : node16680;
												assign node16680 = (inp[0]) ? node16696 : node16681;
													assign node16681 = (inp[1]) ? node16689 : node16682;
														assign node16682 = (inp[14]) ? 4'b0001 : node16683;
															assign node16683 = (inp[7]) ? 4'b0001 : node16684;
																assign node16684 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node16689 = (inp[14]) ? 4'b0000 : node16690;
															assign node16690 = (inp[12]) ? 4'b0001 : node16691;
																assign node16691 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node16696 = (inp[1]) ? node16706 : node16697;
														assign node16697 = (inp[7]) ? node16703 : node16698;
															assign node16698 = (inp[14]) ? 4'b1000 : node16699;
																assign node16699 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node16703 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16706 = (inp[12]) ? 4'b0000 : node16707;
															assign node16707 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node16711 = (inp[0]) ? node16727 : node16712;
													assign node16712 = (inp[1]) ? node16720 : node16713;
														assign node16713 = (inp[7]) ? node16717 : node16714;
															assign node16714 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16717 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16720 = (inp[7]) ? node16722 : 4'b1001;
															assign node16722 = (inp[14]) ? 4'b1001 : node16723;
																assign node16723 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node16727 = (inp[1]) ? node16737 : node16728;
														assign node16728 = (inp[12]) ? node16734 : node16729;
															assign node16729 = (inp[14]) ? node16731 : 4'b1001;
																assign node16731 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node16734 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node16737 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node16740 = (inp[13]) ? node16824 : node16741;
											assign node16741 = (inp[10]) ? node16779 : node16742;
												assign node16742 = (inp[12]) ? node16766 : node16743;
													assign node16743 = (inp[7]) ? node16753 : node16744;
														assign node16744 = (inp[1]) ? node16750 : node16745;
															assign node16745 = (inp[0]) ? node16747 : 4'b0001;
																assign node16747 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node16750 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node16753 = (inp[0]) ? node16759 : node16754;
															assign node16754 = (inp[1]) ? 4'b1000 : node16755;
																assign node16755 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16759 = (inp[14]) ? node16763 : node16760;
																assign node16760 = (inp[1]) ? 4'b0000 : 4'b1001;
																assign node16763 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node16766 = (inp[14]) ? node16772 : node16767;
														assign node16767 = (inp[1]) ? node16769 : 4'b1001;
															assign node16769 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node16772 = (inp[1]) ? node16774 : 4'b1000;
															assign node16774 = (inp[7]) ? node16776 : 4'b1001;
																assign node16776 = (inp[0]) ? 4'b1001 : 4'b0001;
												assign node16779 = (inp[14]) ? node16803 : node16780;
													assign node16780 = (inp[7]) ? node16792 : node16781;
														assign node16781 = (inp[1]) ? node16787 : node16782;
															assign node16782 = (inp[0]) ? 4'b0001 : node16783;
																assign node16783 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node16787 = (inp[12]) ? node16789 : 4'b1001;
																assign node16789 = (inp[0]) ? 4'b0001 : 4'b1001;
														assign node16792 = (inp[1]) ? node16800 : node16793;
															assign node16793 = (inp[12]) ? node16797 : node16794;
																assign node16794 = (inp[0]) ? 4'b0001 : 4'b1001;
																assign node16797 = (inp[0]) ? 4'b1001 : 4'b0001;
															assign node16800 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node16803 = (inp[1]) ? node16813 : node16804;
														assign node16804 = (inp[7]) ? node16806 : 4'b0001;
															assign node16806 = (inp[0]) ? node16810 : node16807;
																assign node16807 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node16810 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node16813 = (inp[0]) ? node16817 : node16814;
															assign node16814 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node16817 = (inp[7]) ? node16821 : node16818;
																assign node16818 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node16821 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node16824 = (inp[0]) ? node16850 : node16825;
												assign node16825 = (inp[10]) ? node16833 : node16826;
													assign node16826 = (inp[7]) ? node16828 : 4'b0000;
														assign node16828 = (inp[1]) ? 4'b0000 : node16829;
															assign node16829 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node16833 = (inp[12]) ? node16841 : node16834;
														assign node16834 = (inp[14]) ? node16836 : 4'b0001;
															assign node16836 = (inp[1]) ? node16838 : 4'b0000;
																assign node16838 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node16841 = (inp[7]) ? node16847 : node16842;
															assign node16842 = (inp[14]) ? node16844 : 4'b1001;
																assign node16844 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node16847 = (inp[14]) ? 4'b1001 : 4'b0000;
												assign node16850 = (inp[7]) ? node16868 : node16851;
													assign node16851 = (inp[10]) ? node16857 : node16852;
														assign node16852 = (inp[12]) ? 4'b1001 : node16853;
															assign node16853 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node16857 = (inp[1]) ? node16861 : node16858;
															assign node16858 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node16861 = (inp[14]) ? node16865 : node16862;
																assign node16862 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node16865 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16868 = (inp[10]) ? node16880 : node16869;
														assign node16869 = (inp[12]) ? node16875 : node16870;
															assign node16870 = (inp[1]) ? 4'b0001 : node16871;
																assign node16871 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node16875 = (inp[14]) ? node16877 : 4'b0000;
																assign node16877 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node16880 = (inp[12]) ? 4'b0001 : node16881;
															assign node16881 = (inp[1]) ? 4'b1001 : 4'b0001;
									assign node16885 = (inp[1]) ? node16991 : node16886;
										assign node16886 = (inp[7]) ? node16936 : node16887;
											assign node16887 = (inp[10]) ? node16911 : node16888;
												assign node16888 = (inp[13]) ? node16900 : node16889;
													assign node16889 = (inp[0]) ? node16895 : node16890;
														assign node16890 = (inp[2]) ? node16892 : 4'b1000;
															assign node16892 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node16895 = (inp[2]) ? node16897 : 4'b0000;
															assign node16897 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node16900 = (inp[2]) ? node16906 : node16901;
														assign node16901 = (inp[12]) ? node16903 : 4'b1001;
															assign node16903 = (inp[0]) ? 4'b1001 : 4'b0001;
														assign node16906 = (inp[12]) ? 4'b1000 : node16907;
															assign node16907 = (inp[0]) ? 4'b0000 : 4'b1000;
												assign node16911 = (inp[0]) ? node16925 : node16912;
													assign node16912 = (inp[13]) ? node16918 : node16913;
														assign node16913 = (inp[12]) ? node16915 : 4'b0001;
															assign node16915 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node16918 = (inp[2]) ? node16922 : node16919;
															assign node16919 = (inp[12]) ? 4'b1001 : 4'b0000;
															assign node16922 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node16925 = (inp[2]) ? node16931 : node16926;
														assign node16926 = (inp[12]) ? node16928 : 4'b0000;
															assign node16928 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node16931 = (inp[13]) ? 4'b0001 : node16932;
															assign node16932 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node16936 = (inp[13]) ? node16962 : node16937;
												assign node16937 = (inp[10]) ? node16949 : node16938;
													assign node16938 = (inp[0]) ? node16944 : node16939;
														assign node16939 = (inp[12]) ? 4'b0001 : node16940;
															assign node16940 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node16944 = (inp[2]) ? 4'b1001 : node16945;
															assign node16945 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node16949 = (inp[12]) ? node16957 : node16950;
														assign node16950 = (inp[0]) ? node16954 : node16951;
															assign node16951 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node16954 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node16957 = (inp[0]) ? node16959 : 4'b1000;
															assign node16959 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node16962 = (inp[2]) ? node16976 : node16963;
													assign node16963 = (inp[10]) ? node16969 : node16964;
														assign node16964 = (inp[12]) ? node16966 : 4'b0000;
															assign node16966 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node16969 = (inp[0]) ? node16973 : node16970;
															assign node16970 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node16973 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node16976 = (inp[0]) ? node16984 : node16977;
														assign node16977 = (inp[10]) ? node16981 : node16978;
															assign node16978 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node16981 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node16984 = (inp[10]) ? node16988 : node16985;
															assign node16985 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node16988 = (inp[12]) ? 4'b0000 : 4'b1000;
										assign node16991 = (inp[13]) ? node17037 : node16992;
											assign node16992 = (inp[2]) ? node17022 : node16993;
												assign node16993 = (inp[10]) ? node17005 : node16994;
													assign node16994 = (inp[0]) ? node17000 : node16995;
														assign node16995 = (inp[7]) ? 4'b1000 : node16996;
															assign node16996 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node17000 = (inp[7]) ? node17002 : 4'b1000;
															assign node17002 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17005 = (inp[12]) ? node17013 : node17006;
														assign node17006 = (inp[7]) ? node17010 : node17007;
															assign node17007 = (inp[0]) ? 4'b0000 : 4'b1000;
															assign node17010 = (inp[0]) ? 4'b1000 : 4'b0000;
														assign node17013 = (inp[14]) ? 4'b1000 : node17014;
															assign node17014 = (inp[0]) ? node17018 : node17015;
																assign node17015 = (inp[7]) ? 4'b0000 : 4'b1000;
																assign node17018 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node17022 = (inp[0]) ? node17024 : 4'b0000;
													assign node17024 = (inp[12]) ? node17030 : node17025;
														assign node17025 = (inp[7]) ? 4'b0000 : node17026;
															assign node17026 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node17030 = (inp[7]) ? node17034 : node17031;
															assign node17031 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node17034 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node17037 = (inp[10]) ? 4'b1000 : node17038;
												assign node17038 = (inp[0]) ? node17050 : node17039;
													assign node17039 = (inp[12]) ? node17045 : node17040;
														assign node17040 = (inp[7]) ? node17042 : 4'b1000;
															assign node17042 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node17045 = (inp[2]) ? node17047 : 4'b1000;
															assign node17047 = (inp[7]) ? 4'b1000 : 4'b0000;
													assign node17050 = (inp[7]) ? node17052 : 4'b0000;
														assign node17052 = (inp[2]) ? 4'b0000 : node17053;
															assign node17053 = (inp[12]) ? 4'b0000 : 4'b1000;
								assign node17058 = (inp[13]) ? node17312 : node17059;
									assign node17059 = (inp[1]) ? node17203 : node17060;
										assign node17060 = (inp[10]) ? node17124 : node17061;
											assign node17061 = (inp[2]) ? node17091 : node17062;
												assign node17062 = (inp[0]) ? node17078 : node17063;
													assign node17063 = (inp[12]) ? node17069 : node17064;
														assign node17064 = (inp[11]) ? node17066 : 4'b1000;
															assign node17066 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17069 = (inp[11]) ? node17075 : node17070;
															assign node17070 = (inp[14]) ? node17072 : 4'b1000;
																assign node17072 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node17075 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node17078 = (inp[11]) ? node17086 : node17079;
														assign node17079 = (inp[14]) ? node17081 : 4'b0000;
															assign node17081 = (inp[7]) ? node17083 : 4'b0000;
																assign node17083 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node17086 = (inp[7]) ? node17088 : 4'b1000;
															assign node17088 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node17091 = (inp[11]) ? node17113 : node17092;
													assign node17092 = (inp[7]) ? node17106 : node17093;
														assign node17093 = (inp[14]) ? node17101 : node17094;
															assign node17094 = (inp[12]) ? node17098 : node17095;
																assign node17095 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node17098 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node17101 = (inp[12]) ? node17103 : 4'b0000;
																assign node17103 = (inp[0]) ? 4'b1001 : 4'b0000;
														assign node17106 = (inp[0]) ? 4'b1001 : node17107;
															assign node17107 = (inp[14]) ? 4'b0001 : node17108;
																assign node17108 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17113 = (inp[0]) ? node17117 : node17114;
														assign node17114 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17117 = (inp[12]) ? node17121 : node17118;
															assign node17118 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17121 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node17124 = (inp[0]) ? node17160 : node17125;
												assign node17125 = (inp[2]) ? node17141 : node17126;
													assign node17126 = (inp[7]) ? node17136 : node17127;
														assign node17127 = (inp[12]) ? node17133 : node17128;
															assign node17128 = (inp[11]) ? 4'b0001 : node17129;
																assign node17129 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node17133 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node17136 = (inp[11]) ? 4'b0001 : node17137;
															assign node17137 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17141 = (inp[7]) ? node17151 : node17142;
														assign node17142 = (inp[12]) ? node17148 : node17143;
															assign node17143 = (inp[11]) ? 4'b1000 : node17144;
																assign node17144 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17148 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node17151 = (inp[14]) ? 4'b0001 : node17152;
															assign node17152 = (inp[11]) ? node17156 : node17153;
																assign node17153 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node17156 = (inp[12]) ? 4'b1000 : 4'b0001;
												assign node17160 = (inp[11]) ? node17190 : node17161;
													assign node17161 = (inp[7]) ? node17177 : node17162;
														assign node17162 = (inp[12]) ? node17170 : node17163;
															assign node17163 = (inp[2]) ? node17167 : node17164;
																assign node17164 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node17167 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17170 = (inp[14]) ? node17174 : node17171;
																assign node17171 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node17174 = (inp[2]) ? 4'b0000 : 4'b1001;
														assign node17177 = (inp[2]) ? node17185 : node17178;
															assign node17178 = (inp[12]) ? node17182 : node17179;
																assign node17179 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node17182 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node17185 = (inp[12]) ? node17187 : 4'b0000;
																assign node17187 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node17190 = (inp[2]) ? node17198 : node17191;
														assign node17191 = (inp[14]) ? 4'b0000 : node17192;
															assign node17192 = (inp[12]) ? 4'b0000 : node17193;
																assign node17193 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17198 = (inp[12]) ? node17200 : 4'b0000;
															assign node17200 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node17203 = (inp[11]) ? node17277 : node17204;
											assign node17204 = (inp[0]) ? node17240 : node17205;
												assign node17205 = (inp[7]) ? node17223 : node17206;
													assign node17206 = (inp[10]) ? node17212 : node17207;
														assign node17207 = (inp[14]) ? node17209 : 4'b0001;
															assign node17209 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node17212 = (inp[12]) ? node17218 : node17213;
															assign node17213 = (inp[14]) ? node17215 : 4'b0000;
																assign node17215 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node17218 = (inp[2]) ? 4'b0000 : node17219;
																assign node17219 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17223 = (inp[12]) ? node17233 : node17224;
														assign node17224 = (inp[2]) ? node17226 : 4'b0001;
															assign node17226 = (inp[10]) ? node17230 : node17227;
																assign node17227 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node17230 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17233 = (inp[14]) ? 4'b0001 : node17234;
															assign node17234 = (inp[2]) ? node17236 : 4'b1000;
																assign node17236 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node17240 = (inp[7]) ? node17260 : node17241;
													assign node17241 = (inp[10]) ? node17253 : node17242;
														assign node17242 = (inp[12]) ? node17248 : node17243;
															assign node17243 = (inp[2]) ? 4'b1000 : node17244;
																assign node17244 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node17248 = (inp[14]) ? node17250 : 4'b0000;
																assign node17250 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node17253 = (inp[14]) ? 4'b0001 : node17254;
															assign node17254 = (inp[2]) ? 4'b0001 : node17255;
																assign node17255 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node17260 = (inp[14]) ? node17270 : node17261;
														assign node17261 = (inp[10]) ? node17265 : node17262;
															assign node17262 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node17265 = (inp[12]) ? node17267 : 4'b0000;
																assign node17267 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node17270 = (inp[12]) ? 4'b0000 : node17271;
															assign node17271 = (inp[10]) ? node17273 : 4'b0000;
																assign node17273 = (inp[2]) ? 4'b1000 : 4'b0000;
											assign node17277 = (inp[10]) ? 4'b0000 : node17278;
												assign node17278 = (inp[2]) ? node17300 : node17279;
													assign node17279 = (inp[12]) ? node17285 : node17280;
														assign node17280 = (inp[0]) ? 4'b0000 : node17281;
															assign node17281 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node17285 = (inp[14]) ? node17293 : node17286;
															assign node17286 = (inp[7]) ? node17290 : node17287;
																assign node17287 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node17290 = (inp[0]) ? 4'b1000 : 4'b0000;
															assign node17293 = (inp[7]) ? node17297 : node17294;
																assign node17294 = (inp[0]) ? 4'b0000 : 4'b1000;
																assign node17297 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node17300 = (inp[12]) ? node17306 : node17301;
														assign node17301 = (inp[7]) ? 4'b1000 : node17302;
															assign node17302 = (inp[0]) ? 4'b0000 : 4'b1000;
														assign node17306 = (inp[7]) ? 4'b0000 : node17307;
															assign node17307 = (inp[0]) ? 4'b1000 : 4'b0000;
									assign node17312 = (inp[10]) ? node17408 : node17313;
										assign node17313 = (inp[1]) ? node17373 : node17314;
											assign node17314 = (inp[12]) ? node17340 : node17315;
												assign node17315 = (inp[7]) ? node17329 : node17316;
													assign node17316 = (inp[0]) ? node17324 : node17317;
														assign node17317 = (inp[2]) ? node17319 : 4'b0000;
															assign node17319 = (inp[14]) ? 4'b0001 : node17320;
																assign node17320 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17324 = (inp[2]) ? 4'b0000 : node17325;
															assign node17325 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node17329 = (inp[2]) ? node17337 : node17330;
														assign node17330 = (inp[0]) ? 4'b0000 : node17331;
															assign node17331 = (inp[14]) ? node17333 : 4'b0001;
																assign node17333 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17337 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node17340 = (inp[2]) ? node17360 : node17341;
													assign node17341 = (inp[7]) ? node17353 : node17342;
														assign node17342 = (inp[0]) ? node17348 : node17343;
															assign node17343 = (inp[14]) ? 4'b0001 : node17344;
																assign node17344 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node17348 = (inp[11]) ? 4'b0000 : node17349;
																assign node17349 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17353 = (inp[11]) ? 4'b0001 : node17354;
															assign node17354 = (inp[14]) ? 4'b0001 : node17355;
																assign node17355 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node17360 = (inp[7]) ? node17368 : node17361;
														assign node17361 = (inp[0]) ? node17365 : node17362;
															assign node17362 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node17365 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17368 = (inp[11]) ? 4'b0000 : node17369;
															assign node17369 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node17373 = (inp[11]) ? 4'b0000 : node17374;
												assign node17374 = (inp[0]) ? node17394 : node17375;
													assign node17375 = (inp[2]) ? node17383 : node17376;
														assign node17376 = (inp[14]) ? node17378 : 4'b0001;
															assign node17378 = (inp[7]) ? node17380 : 4'b0001;
																assign node17380 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node17383 = (inp[7]) ? node17389 : node17384;
															assign node17384 = (inp[12]) ? 4'b0000 : node17385;
																assign node17385 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node17389 = (inp[12]) ? node17391 : 4'b0001;
																assign node17391 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node17394 = (inp[14]) ? node17400 : node17395;
														assign node17395 = (inp[2]) ? node17397 : 4'b0000;
															assign node17397 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17400 = (inp[12]) ? 4'b0000 : node17401;
															assign node17401 = (inp[7]) ? node17403 : 4'b0000;
																assign node17403 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node17408 = (inp[11]) ? 4'b0000 : node17409;
											assign node17409 = (inp[1]) ? 4'b0000 : node17410;
												assign node17410 = (inp[2]) ? node17432 : node17411;
													assign node17411 = (inp[14]) ? node17419 : node17412;
														assign node17412 = (inp[12]) ? 4'b0000 : node17413;
															assign node17413 = (inp[0]) ? node17415 : 4'b0000;
																assign node17415 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17419 = (inp[7]) ? node17425 : node17420;
															assign node17420 = (inp[12]) ? node17422 : 4'b0000;
																assign node17422 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node17425 = (inp[12]) ? node17429 : node17426;
																assign node17426 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node17429 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node17432 = (inp[12]) ? node17446 : node17433;
														assign node17433 = (inp[7]) ? node17439 : node17434;
															assign node17434 = (inp[14]) ? node17436 : 4'b0000;
																assign node17436 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node17439 = (inp[0]) ? node17443 : node17440;
																assign node17440 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node17443 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node17446 = (inp[14]) ? node17452 : node17447;
															assign node17447 = (inp[7]) ? node17449 : 4'b0001;
																assign node17449 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node17452 = (inp[0]) ? node17454 : 4'b0000;
																assign node17454 = (inp[7]) ? 4'b0000 : 4'b0001;
				assign node17459 = (inp[0]) ? node19963 : node17460;
					assign node17460 = (inp[6]) ? node18148 : node17461;
						assign node17461 = (inp[5]) ? node17609 : node17462;
							assign node17462 = (inp[3]) ? node17464 : 4'b1010;
								assign node17464 = (inp[2]) ? 4'b1010 : node17465;
									assign node17465 = (inp[7]) ? node17553 : node17466;
										assign node17466 = (inp[1]) ? node17508 : node17467;
											assign node17467 = (inp[13]) ? node17491 : node17468;
												assign node17468 = (inp[4]) ? node17478 : node17469;
													assign node17469 = (inp[12]) ? 4'b1010 : node17470;
														assign node17470 = (inp[10]) ? node17472 : 4'b1010;
															assign node17472 = (inp[11]) ? 4'b0001 : node17473;
																assign node17473 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node17478 = (inp[12]) ? node17486 : node17479;
														assign node17479 = (inp[10]) ? node17481 : 4'b1001;
															assign node17481 = (inp[14]) ? node17483 : 4'b0001;
																assign node17483 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17486 = (inp[11]) ? 4'b1001 : node17487;
															assign node17487 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node17491 = (inp[12]) ? node17503 : node17492;
													assign node17492 = (inp[10]) ? node17498 : node17493;
														assign node17493 = (inp[11]) ? 4'b0001 : node17494;
															assign node17494 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17498 = (inp[14]) ? node17500 : 4'b1001;
															assign node17500 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node17503 = (inp[14]) ? node17505 : 4'b0001;
														assign node17505 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node17508 = (inp[11]) ? node17540 : node17509;
												assign node17509 = (inp[14]) ? node17523 : node17510;
													assign node17510 = (inp[13]) ? node17518 : node17511;
														assign node17511 = (inp[10]) ? 4'b0000 : node17512;
															assign node17512 = (inp[12]) ? node17514 : 4'b0000;
																assign node17514 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node17518 = (inp[12]) ? node17520 : 4'b1000;
															assign node17520 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node17523 = (inp[13]) ? node17535 : node17524;
														assign node17524 = (inp[4]) ? node17530 : node17525;
															assign node17525 = (inp[10]) ? node17527 : 4'b1010;
																assign node17527 = (inp[12]) ? 4'b1010 : 4'b0001;
															assign node17530 = (inp[10]) ? node17532 : 4'b1001;
																assign node17532 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node17535 = (inp[10]) ? node17537 : 4'b0001;
															assign node17537 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node17540 = (inp[13]) ? node17548 : node17541;
													assign node17541 = (inp[10]) ? 4'b0000 : node17542;
														assign node17542 = (inp[12]) ? node17544 : 4'b0000;
															assign node17544 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node17548 = (inp[12]) ? node17550 : 4'b1000;
														assign node17550 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node17553 = (inp[4]) ? node17555 : 4'b1010;
											assign node17555 = (inp[13]) ? node17583 : node17556;
												assign node17556 = (inp[10]) ? node17566 : node17557;
													assign node17557 = (inp[1]) ? node17559 : 4'b1010;
														assign node17559 = (inp[12]) ? 4'b1010 : node17560;
															assign node17560 = (inp[11]) ? 4'b0000 : node17561;
																assign node17561 = (inp[14]) ? 4'b1010 : 4'b0000;
													assign node17566 = (inp[12]) ? node17576 : node17567;
														assign node17567 = (inp[14]) ? node17571 : node17568;
															assign node17568 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node17571 = (inp[11]) ? 4'b0000 : node17572;
																assign node17572 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node17576 = (inp[1]) ? node17578 : 4'b1010;
															assign node17578 = (inp[14]) ? node17580 : 4'b0000;
																assign node17580 = (inp[11]) ? 4'b0000 : 4'b1010;
												assign node17583 = (inp[12]) ? node17597 : node17584;
													assign node17584 = (inp[1]) ? node17592 : node17585;
														assign node17585 = (inp[10]) ? node17587 : 4'b0001;
															assign node17587 = (inp[11]) ? 4'b1001 : node17588;
																assign node17588 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node17592 = (inp[14]) ? node17594 : 4'b1000;
															assign node17594 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node17597 = (inp[1]) ? node17603 : node17598;
														assign node17598 = (inp[11]) ? 4'b0001 : node17599;
															assign node17599 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node17603 = (inp[11]) ? node17605 : 4'b0001;
															assign node17605 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node17609 = (inp[2]) ? node18009 : node17610;
								assign node17610 = (inp[1]) ? node17806 : node17611;
									assign node17611 = (inp[11]) ? node17735 : node17612;
										assign node17612 = (inp[14]) ? node17674 : node17613;
											assign node17613 = (inp[13]) ? node17641 : node17614;
												assign node17614 = (inp[12]) ? node17634 : node17615;
													assign node17615 = (inp[10]) ? node17625 : node17616;
														assign node17616 = (inp[4]) ? node17618 : 4'b1101;
															assign node17618 = (inp[3]) ? node17622 : node17619;
																assign node17619 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node17622 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node17625 = (inp[3]) ? node17629 : node17626;
															assign node17626 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node17629 = (inp[4]) ? 4'b0001 : node17630;
																assign node17630 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node17634 = (inp[3]) ? node17636 : 4'b1001;
														assign node17636 = (inp[7]) ? 4'b1101 : node17637;
															assign node17637 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node17641 = (inp[10]) ? node17653 : node17642;
													assign node17642 = (inp[3]) ? node17648 : node17643;
														assign node17643 = (inp[4]) ? 4'b0101 : node17644;
															assign node17644 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17648 = (inp[4]) ? 4'b0001 : node17649;
															assign node17649 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node17653 = (inp[12]) ? node17665 : node17654;
														assign node17654 = (inp[3]) ? node17660 : node17655;
															assign node17655 = (inp[4]) ? 4'b1101 : node17656;
																assign node17656 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node17660 = (inp[7]) ? node17662 : 4'b1001;
																assign node17662 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17665 = (inp[7]) ? node17669 : node17666;
															assign node17666 = (inp[3]) ? 4'b0001 : 4'b0101;
															assign node17669 = (inp[3]) ? node17671 : 4'b0001;
																assign node17671 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node17674 = (inp[13]) ? node17704 : node17675;
												assign node17675 = (inp[10]) ? node17687 : node17676;
													assign node17676 = (inp[3]) ? node17682 : node17677;
														assign node17677 = (inp[7]) ? 4'b1000 : node17678;
															assign node17678 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node17682 = (inp[4]) ? node17684 : 4'b1100;
															assign node17684 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node17687 = (inp[12]) ? node17699 : node17688;
														assign node17688 = (inp[3]) ? node17694 : node17689;
															assign node17689 = (inp[4]) ? 4'b0100 : node17690;
																assign node17690 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node17694 = (inp[4]) ? 4'b0000 : node17695;
																assign node17695 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node17699 = (inp[3]) ? 4'b1100 : node17700;
															assign node17700 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node17704 = (inp[10]) ? node17716 : node17705;
													assign node17705 = (inp[3]) ? node17711 : node17706;
														assign node17706 = (inp[7]) ? node17708 : 4'b0100;
															assign node17708 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node17711 = (inp[4]) ? 4'b0000 : node17712;
															assign node17712 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node17716 = (inp[12]) ? node17726 : node17717;
														assign node17717 = (inp[3]) ? node17721 : node17718;
															assign node17718 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node17721 = (inp[7]) ? node17723 : 4'b1000;
																assign node17723 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node17726 = (inp[3]) ? node17730 : node17727;
															assign node17727 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node17730 = (inp[4]) ? 4'b0000 : node17731;
																assign node17731 = (inp[7]) ? 4'b0100 : 4'b0000;
										assign node17735 = (inp[13]) ? node17771 : node17736;
											assign node17736 = (inp[12]) ? node17760 : node17737;
												assign node17737 = (inp[10]) ? node17749 : node17738;
													assign node17738 = (inp[3]) ? node17744 : node17739;
														assign node17739 = (inp[4]) ? node17741 : 4'b1001;
															assign node17741 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node17744 = (inp[4]) ? node17746 : 4'b1101;
															assign node17746 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node17749 = (inp[3]) ? node17755 : node17750;
														assign node17750 = (inp[4]) ? 4'b0101 : node17751;
															assign node17751 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17755 = (inp[7]) ? node17757 : 4'b0001;
															assign node17757 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node17760 = (inp[3]) ? node17766 : node17761;
													assign node17761 = (inp[7]) ? 4'b1001 : node17762;
														assign node17762 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node17766 = (inp[4]) ? node17768 : 4'b1101;
														assign node17768 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node17771 = (inp[10]) ? node17783 : node17772;
												assign node17772 = (inp[3]) ? node17778 : node17773;
													assign node17773 = (inp[7]) ? node17775 : 4'b0101;
														assign node17775 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node17778 = (inp[4]) ? 4'b0001 : node17779;
														assign node17779 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node17783 = (inp[12]) ? node17795 : node17784;
													assign node17784 = (inp[3]) ? node17790 : node17785;
														assign node17785 = (inp[4]) ? 4'b1101 : node17786;
															assign node17786 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node17790 = (inp[4]) ? 4'b1001 : node17791;
															assign node17791 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node17795 = (inp[3]) ? node17801 : node17796;
														assign node17796 = (inp[7]) ? node17798 : 4'b0101;
															assign node17798 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node17801 = (inp[7]) ? node17803 : 4'b0001;
															assign node17803 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node17806 = (inp[14]) ? node17872 : node17807;
										assign node17807 = (inp[13]) ? node17841 : node17808;
											assign node17808 = (inp[10]) ? node17830 : node17809;
												assign node17809 = (inp[12]) ? node17821 : node17810;
													assign node17810 = (inp[3]) ? node17816 : node17811;
														assign node17811 = (inp[7]) ? node17813 : 4'b0100;
															assign node17813 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node17816 = (inp[4]) ? 4'b0000 : node17817;
															assign node17817 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node17821 = (inp[3]) ? node17825 : node17822;
														assign node17822 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node17825 = (inp[4]) ? node17827 : 4'b1100;
															assign node17827 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node17830 = (inp[3]) ? node17836 : node17831;
													assign node17831 = (inp[7]) ? node17833 : 4'b0100;
														assign node17833 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node17836 = (inp[7]) ? node17838 : 4'b0000;
														assign node17838 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node17841 = (inp[10]) ? node17861 : node17842;
												assign node17842 = (inp[12]) ? node17850 : node17843;
													assign node17843 = (inp[3]) ? 4'b1000 : node17844;
														assign node17844 = (inp[7]) ? node17846 : 4'b1100;
															assign node17846 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node17850 = (inp[3]) ? node17856 : node17851;
														assign node17851 = (inp[4]) ? 4'b0100 : node17852;
															assign node17852 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node17856 = (inp[4]) ? 4'b0000 : node17857;
															assign node17857 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node17861 = (inp[3]) ? node17867 : node17862;
													assign node17862 = (inp[4]) ? 4'b1100 : node17863;
														assign node17863 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node17867 = (inp[7]) ? node17869 : 4'b1000;
														assign node17869 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node17872 = (inp[11]) ? node17940 : node17873;
											assign node17873 = (inp[13]) ? node17909 : node17874;
												assign node17874 = (inp[10]) ? node17886 : node17875;
													assign node17875 = (inp[3]) ? node17881 : node17876;
														assign node17876 = (inp[7]) ? 4'b1001 : node17877;
															assign node17877 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node17881 = (inp[4]) ? node17883 : 4'b1101;
															assign node17883 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node17886 = (inp[12]) ? node17898 : node17887;
														assign node17887 = (inp[3]) ? node17893 : node17888;
															assign node17888 = (inp[4]) ? 4'b0101 : node17889;
																assign node17889 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node17893 = (inp[4]) ? 4'b0001 : node17894;
																assign node17894 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node17898 = (inp[3]) ? node17904 : node17899;
															assign node17899 = (inp[7]) ? 4'b1001 : node17900;
																assign node17900 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node17904 = (inp[4]) ? node17906 : 4'b1101;
																assign node17906 = (inp[7]) ? 4'b1101 : 4'b1001;
												assign node17909 = (inp[10]) ? node17921 : node17910;
													assign node17910 = (inp[3]) ? node17916 : node17911;
														assign node17911 = (inp[4]) ? 4'b0101 : node17912;
															assign node17912 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node17916 = (inp[7]) ? node17918 : 4'b0001;
															assign node17918 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node17921 = (inp[12]) ? node17933 : node17922;
														assign node17922 = (inp[3]) ? node17928 : node17923;
															assign node17923 = (inp[7]) ? node17925 : 4'b1101;
																assign node17925 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node17928 = (inp[4]) ? 4'b1001 : node17929;
																assign node17929 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node17933 = (inp[7]) ? node17935 : 4'b0001;
															assign node17935 = (inp[4]) ? node17937 : 4'b0101;
																assign node17937 = (inp[3]) ? 4'b0001 : 4'b0101;
											assign node17940 = (inp[13]) ? node17976 : node17941;
												assign node17941 = (inp[12]) ? node17953 : node17942;
													assign node17942 = (inp[3]) ? node17948 : node17943;
														assign node17943 = (inp[7]) ? node17945 : 4'b0100;
															assign node17945 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node17948 = (inp[4]) ? 4'b0000 : node17949;
															assign node17949 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node17953 = (inp[10]) ? node17965 : node17954;
														assign node17954 = (inp[3]) ? node17960 : node17955;
															assign node17955 = (inp[7]) ? 4'b1000 : node17956;
																assign node17956 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node17960 = (inp[7]) ? 4'b1100 : node17961;
																assign node17961 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node17965 = (inp[3]) ? node17971 : node17966;
															assign node17966 = (inp[7]) ? node17968 : 4'b0100;
																assign node17968 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node17971 = (inp[7]) ? node17973 : 4'b0000;
																assign node17973 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node17976 = (inp[10]) ? node17998 : node17977;
													assign node17977 = (inp[12]) ? node17987 : node17978;
														assign node17978 = (inp[3]) ? node17982 : node17979;
															assign node17979 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node17982 = (inp[4]) ? 4'b1000 : node17983;
																assign node17983 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node17987 = (inp[3]) ? node17993 : node17988;
															assign node17988 = (inp[4]) ? 4'b0100 : node17989;
																assign node17989 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node17993 = (inp[4]) ? 4'b0000 : node17994;
																assign node17994 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node17998 = (inp[3]) ? node18004 : node17999;
														assign node17999 = (inp[4]) ? 4'b1100 : node18000;
															assign node18000 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node18004 = (inp[7]) ? node18006 : 4'b1000;
															assign node18006 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node18009 = (inp[3]) ? node18011 : 4'b1010;
									assign node18011 = (inp[4]) ? node18073 : node18012;
										assign node18012 = (inp[7]) ? 4'b1010 : node18013;
											assign node18013 = (inp[13]) ? node18043 : node18014;
												assign node18014 = (inp[12]) ? node18034 : node18015;
													assign node18015 = (inp[10]) ? node18023 : node18016;
														assign node18016 = (inp[1]) ? node18018 : 4'b1010;
															assign node18018 = (inp[11]) ? 4'b0000 : node18019;
																assign node18019 = (inp[14]) ? 4'b1010 : 4'b0000;
														assign node18023 = (inp[1]) ? node18029 : node18024;
															assign node18024 = (inp[14]) ? node18026 : 4'b0001;
																assign node18026 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node18029 = (inp[14]) ? node18031 : 4'b0000;
																assign node18031 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node18034 = (inp[10]) ? node18036 : 4'b1010;
														assign node18036 = (inp[1]) ? node18038 : 4'b1010;
															assign node18038 = (inp[14]) ? node18040 : 4'b0000;
																assign node18040 = (inp[11]) ? 4'b0000 : 4'b1010;
												assign node18043 = (inp[10]) ? node18057 : node18044;
													assign node18044 = (inp[1]) ? node18050 : node18045;
														assign node18045 = (inp[14]) ? node18047 : 4'b0001;
															assign node18047 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node18050 = (inp[14]) ? node18054 : node18051;
															assign node18051 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node18054 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node18057 = (inp[1]) ? node18065 : node18058;
														assign node18058 = (inp[12]) ? 4'b0001 : node18059;
															assign node18059 = (inp[14]) ? node18061 : 4'b1001;
																assign node18061 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18065 = (inp[14]) ? node18067 : 4'b1000;
															assign node18067 = (inp[11]) ? 4'b1000 : node18068;
																assign node18068 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node18073 = (inp[1]) ? node18111 : node18074;
											assign node18074 = (inp[13]) ? node18098 : node18075;
												assign node18075 = (inp[7]) ? node18089 : node18076;
													assign node18076 = (inp[12]) ? node18084 : node18077;
														assign node18077 = (inp[10]) ? node18079 : 4'b1001;
															assign node18079 = (inp[11]) ? 4'b0001 : node18080;
																assign node18080 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18084 = (inp[11]) ? 4'b1001 : node18085;
															assign node18085 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18089 = (inp[12]) ? 4'b1010 : node18090;
														assign node18090 = (inp[10]) ? node18092 : 4'b1010;
															assign node18092 = (inp[11]) ? 4'b0001 : node18093;
																assign node18093 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18098 = (inp[12]) ? node18106 : node18099;
													assign node18099 = (inp[10]) ? node18101 : 4'b0001;
														assign node18101 = (inp[11]) ? 4'b1001 : node18102;
															assign node18102 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node18106 = (inp[11]) ? 4'b0001 : node18107;
														assign node18107 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node18111 = (inp[11]) ? node18135 : node18112;
												assign node18112 = (inp[14]) ? node18126 : node18113;
													assign node18113 = (inp[13]) ? node18121 : node18114;
														assign node18114 = (inp[12]) ? node18116 : 4'b0000;
															assign node18116 = (inp[10]) ? 4'b0000 : node18117;
																assign node18117 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node18121 = (inp[12]) ? node18123 : 4'b1000;
															assign node18123 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node18126 = (inp[13]) ? node18132 : node18127;
														assign node18127 = (inp[7]) ? node18129 : 4'b1001;
															assign node18129 = (inp[12]) ? 4'b1010 : 4'b0001;
														assign node18132 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node18135 = (inp[13]) ? node18143 : node18136;
													assign node18136 = (inp[10]) ? 4'b0000 : node18137;
														assign node18137 = (inp[12]) ? node18139 : 4'b0000;
															assign node18139 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node18143 = (inp[10]) ? 4'b1000 : node18144;
														assign node18144 = (inp[12]) ? 4'b0000 : 4'b1000;
						assign node18148 = (inp[5]) ? node19104 : node18149;
							assign node18149 = (inp[11]) ? node18721 : node18150;
								assign node18150 = (inp[2]) ? node18416 : node18151;
									assign node18151 = (inp[3]) ? node18329 : node18152;
										assign node18152 = (inp[4]) ? node18266 : node18153;
											assign node18153 = (inp[7]) ? node18207 : node18154;
												assign node18154 = (inp[13]) ? node18182 : node18155;
													assign node18155 = (inp[10]) ? node18167 : node18156;
														assign node18156 = (inp[12]) ? node18162 : node18157;
															assign node18157 = (inp[14]) ? node18159 : 4'b1001;
																assign node18159 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node18162 = (inp[14]) ? node18164 : 4'b1000;
																assign node18164 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node18167 = (inp[12]) ? node18175 : node18168;
															assign node18168 = (inp[1]) ? node18172 : node18169;
																assign node18169 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node18172 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node18175 = (inp[14]) ? node18179 : node18176;
																assign node18176 = (inp[1]) ? 4'b0100 : 4'b1001;
																assign node18179 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node18182 = (inp[12]) ? node18196 : node18183;
														assign node18183 = (inp[10]) ? node18189 : node18184;
															assign node18184 = (inp[14]) ? node18186 : 4'b1100;
																assign node18186 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node18189 = (inp[14]) ? node18193 : node18190;
																assign node18190 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node18193 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node18196 = (inp[10]) ? node18202 : node18197;
															assign node18197 = (inp[14]) ? 4'b0101 : node18198;
																assign node18198 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node18202 = (inp[1]) ? 4'b0101 : node18203;
																assign node18203 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node18207 = (inp[13]) ? node18237 : node18208;
													assign node18208 = (inp[10]) ? node18224 : node18209;
														assign node18209 = (inp[12]) ? node18217 : node18210;
															assign node18210 = (inp[1]) ? node18214 : node18211;
																assign node18211 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node18214 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node18217 = (inp[14]) ? node18221 : node18218;
																assign node18218 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node18221 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node18224 = (inp[12]) ? node18230 : node18225;
															assign node18225 = (inp[14]) ? node18227 : 4'b0000;
																assign node18227 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node18230 = (inp[1]) ? node18234 : node18231;
																assign node18231 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node18234 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node18237 = (inp[10]) ? node18253 : node18238;
														assign node18238 = (inp[12]) ? node18246 : node18239;
															assign node18239 = (inp[1]) ? node18243 : node18240;
																assign node18240 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18243 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node18246 = (inp[1]) ? node18250 : node18247;
																assign node18247 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18250 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18253 = (inp[12]) ? node18261 : node18254;
															assign node18254 = (inp[1]) ? node18258 : node18255;
																assign node18255 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node18258 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node18261 = (inp[14]) ? 4'b0001 : node18262;
																assign node18262 = (inp[1]) ? 4'b1000 : 4'b0001;
											assign node18266 = (inp[13]) ? node18304 : node18267;
												assign node18267 = (inp[10]) ? node18285 : node18268;
													assign node18268 = (inp[7]) ? node18276 : node18269;
														assign node18269 = (inp[1]) ? node18273 : node18270;
															assign node18270 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node18273 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node18276 = (inp[14]) ? node18282 : node18277;
															assign node18277 = (inp[1]) ? node18279 : 4'b1001;
																assign node18279 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node18282 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node18285 = (inp[7]) ? node18291 : node18286;
														assign node18286 = (inp[12]) ? 4'b0001 : node18287;
															assign node18287 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node18291 = (inp[12]) ? node18299 : node18292;
															assign node18292 = (inp[14]) ? node18296 : node18293;
																assign node18293 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node18296 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node18299 = (inp[1]) ? 4'b0100 : node18300;
																assign node18300 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node18304 = (inp[7]) ? node18316 : node18305;
													assign node18305 = (inp[10]) ? node18311 : node18306;
														assign node18306 = (inp[12]) ? 4'b1001 : node18307;
															assign node18307 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node18311 = (inp[12]) ? 4'b0001 : node18312;
															assign node18312 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node18316 = (inp[10]) ? node18324 : node18317;
														assign node18317 = (inp[1]) ? node18321 : node18318;
															assign node18318 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node18321 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node18324 = (inp[1]) ? node18326 : 4'b0001;
															assign node18326 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node18329 = (inp[10]) ? node18373 : node18330;
											assign node18330 = (inp[12]) ? node18358 : node18331;
												assign node18331 = (inp[1]) ? node18343 : node18332;
													assign node18332 = (inp[4]) ? node18338 : node18333;
														assign node18333 = (inp[7]) ? 4'b1001 : node18334;
															assign node18334 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node18338 = (inp[7]) ? 4'b1101 : node18339;
															assign node18339 = (inp[14]) ? 4'b1101 : 4'b1000;
													assign node18343 = (inp[4]) ? node18349 : node18344;
														assign node18344 = (inp[7]) ? node18346 : 4'b0101;
															assign node18346 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node18349 = (inp[7]) ? node18355 : node18350;
															assign node18350 = (inp[13]) ? node18352 : 4'b0001;
																assign node18352 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node18355 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node18358 = (inp[4]) ? node18364 : node18359;
													assign node18359 = (inp[7]) ? 4'b1001 : node18360;
														assign node18360 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node18364 = (inp[13]) ? node18366 : 4'b1101;
														assign node18366 = (inp[7]) ? 4'b1101 : node18367;
															assign node18367 = (inp[1]) ? 4'b1001 : node18368;
																assign node18368 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node18373 = (inp[4]) ? node18391 : node18374;
												assign node18374 = (inp[13]) ? node18386 : node18375;
													assign node18375 = (inp[7]) ? node18381 : node18376;
														assign node18376 = (inp[1]) ? node18378 : 4'b0101;
															assign node18378 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node18381 = (inp[1]) ? node18383 : 4'b0001;
															assign node18383 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node18386 = (inp[1]) ? node18388 : 4'b0101;
														assign node18388 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node18391 = (inp[13]) ? node18401 : node18392;
													assign node18392 = (inp[7]) ? node18398 : node18393;
														assign node18393 = (inp[1]) ? node18395 : 4'b0001;
															assign node18395 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18398 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node18401 = (inp[1]) ? node18409 : node18402;
														assign node18402 = (inp[14]) ? node18404 : 4'b0000;
															assign node18404 = (inp[7]) ? 4'b0001 : node18405;
																assign node18405 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node18409 = (inp[14]) ? node18413 : node18410;
															assign node18410 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node18413 = (inp[12]) ? 4'b0000 : 4'b1000;
									assign node18416 = (inp[13]) ? node18586 : node18417;
										assign node18417 = (inp[12]) ? node18517 : node18418;
											assign node18418 = (inp[10]) ? node18468 : node18419;
												assign node18419 = (inp[1]) ? node18443 : node18420;
													assign node18420 = (inp[14]) ? node18432 : node18421;
														assign node18421 = (inp[3]) ? node18427 : node18422;
															assign node18422 = (inp[7]) ? 4'b1001 : node18423;
																assign node18423 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node18427 = (inp[4]) ? node18429 : 4'b1101;
																assign node18429 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node18432 = (inp[3]) ? node18438 : node18433;
															assign node18433 = (inp[4]) ? node18435 : 4'b1000;
																assign node18435 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node18438 = (inp[7]) ? 4'b1100 : node18439;
																assign node18439 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node18443 = (inp[14]) ? node18457 : node18444;
														assign node18444 = (inp[3]) ? node18450 : node18445;
															assign node18445 = (inp[4]) ? 4'b0100 : node18446;
																assign node18446 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node18450 = (inp[4]) ? node18454 : node18451;
																assign node18451 = (inp[7]) ? 4'b0100 : 4'b0000;
																assign node18454 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node18457 = (inp[3]) ? node18463 : node18458;
															assign node18458 = (inp[7]) ? 4'b1001 : node18459;
																assign node18459 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node18463 = (inp[7]) ? 4'b1101 : node18464;
																assign node18464 = (inp[4]) ? 4'b0001 : 4'b1101;
												assign node18468 = (inp[3]) ? node18490 : node18469;
													assign node18469 = (inp[7]) ? node18477 : node18470;
														assign node18470 = (inp[14]) ? node18474 : node18471;
															assign node18471 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node18474 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node18477 = (inp[4]) ? node18485 : node18478;
															assign node18478 = (inp[1]) ? node18482 : node18479;
																assign node18479 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18482 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node18485 = (inp[14]) ? 4'b0101 : node18486;
																assign node18486 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node18490 = (inp[4]) ? node18506 : node18491;
														assign node18491 = (inp[7]) ? node18499 : node18492;
															assign node18492 = (inp[1]) ? node18496 : node18493;
																assign node18493 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18496 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node18499 = (inp[1]) ? node18503 : node18500;
																assign node18500 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node18503 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node18506 = (inp[7]) ? node18510 : node18507;
															assign node18507 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node18510 = (inp[1]) ? node18514 : node18511;
																assign node18511 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18514 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node18517 = (inp[3]) ? node18549 : node18518;
												assign node18518 = (inp[4]) ? node18528 : node18519;
													assign node18519 = (inp[1]) ? node18523 : node18520;
														assign node18520 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node18523 = (inp[14]) ? 4'b1001 : node18524;
															assign node18524 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node18528 = (inp[7]) ? node18538 : node18529;
														assign node18529 = (inp[1]) ? node18533 : node18530;
															assign node18530 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node18533 = (inp[14]) ? 4'b1101 : node18534;
																assign node18534 = (inp[10]) ? 4'b0100 : 4'b1100;
														assign node18538 = (inp[10]) ? node18544 : node18539;
															assign node18539 = (inp[1]) ? node18541 : 4'b1001;
																assign node18541 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node18544 = (inp[14]) ? node18546 : 4'b0100;
																assign node18546 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node18549 = (inp[4]) ? node18567 : node18550;
													assign node18550 = (inp[7]) ? node18558 : node18551;
														assign node18551 = (inp[14]) ? node18555 : node18552;
															assign node18552 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node18555 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node18558 = (inp[1]) ? node18562 : node18559;
															assign node18559 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node18562 = (inp[14]) ? 4'b1101 : node18563;
																assign node18563 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node18567 = (inp[7]) ? node18577 : node18568;
														assign node18568 = (inp[10]) ? 4'b0001 : node18569;
															assign node18569 = (inp[1]) ? node18573 : node18570;
																assign node18570 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node18573 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node18577 = (inp[14]) ? node18583 : node18578;
															assign node18578 = (inp[1]) ? node18580 : 4'b1101;
																assign node18580 = (inp[10]) ? 4'b0000 : 4'b1100;
															assign node18583 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node18586 = (inp[3]) ? node18652 : node18587;
											assign node18587 = (inp[7]) ? node18619 : node18588;
												assign node18588 = (inp[12]) ? node18604 : node18589;
													assign node18589 = (inp[10]) ? node18597 : node18590;
														assign node18590 = (inp[1]) ? node18594 : node18591;
															assign node18591 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node18594 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node18597 = (inp[14]) ? node18601 : node18598;
															assign node18598 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node18601 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node18604 = (inp[10]) ? node18612 : node18605;
														assign node18605 = (inp[14]) ? node18609 : node18606;
															assign node18606 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node18609 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node18612 = (inp[1]) ? node18616 : node18613;
															assign node18613 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node18616 = (inp[14]) ? 4'b0101 : 4'b1100;
												assign node18619 = (inp[4]) ? node18631 : node18620;
													assign node18620 = (inp[14]) ? node18628 : node18621;
														assign node18621 = (inp[1]) ? node18623 : 4'b0001;
															assign node18623 = (inp[12]) ? node18625 : 4'b1000;
																assign node18625 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18628 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node18631 = (inp[10]) ? node18639 : node18632;
														assign node18632 = (inp[12]) ? node18634 : 4'b0101;
															assign node18634 = (inp[14]) ? 4'b0100 : node18635;
																assign node18635 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node18639 = (inp[12]) ? node18645 : node18640;
															assign node18640 = (inp[14]) ? 4'b1100 : node18641;
																assign node18641 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node18645 = (inp[1]) ? node18649 : node18646;
																assign node18646 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node18649 = (inp[14]) ? 4'b0101 : 4'b1100;
											assign node18652 = (inp[4]) ? node18694 : node18653;
												assign node18653 = (inp[7]) ? node18675 : node18654;
													assign node18654 = (inp[12]) ? node18666 : node18655;
														assign node18655 = (inp[10]) ? node18661 : node18656;
															assign node18656 = (inp[1]) ? 4'b1000 : node18657;
																assign node18657 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18661 = (inp[1]) ? 4'b1001 : node18662;
																assign node18662 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node18666 = (inp[10]) ? node18668 : 4'b0001;
															assign node18668 = (inp[1]) ? node18672 : node18669;
																assign node18669 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node18672 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node18675 = (inp[10]) ? node18685 : node18676;
														assign node18676 = (inp[14]) ? node18682 : node18677;
															assign node18677 = (inp[1]) ? node18679 : 4'b0101;
																assign node18679 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node18682 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node18685 = (inp[1]) ? node18691 : node18686;
															assign node18686 = (inp[14]) ? 4'b1100 : node18687;
																assign node18687 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node18691 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node18694 = (inp[7]) ? node18706 : node18695;
													assign node18695 = (inp[10]) ? node18701 : node18696;
														assign node18696 = (inp[12]) ? 4'b1001 : node18697;
															assign node18697 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node18701 = (inp[12]) ? 4'b0001 : node18702;
															assign node18702 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node18706 = (inp[10]) ? node18716 : node18707;
														assign node18707 = (inp[1]) ? node18711 : node18708;
															assign node18708 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node18711 = (inp[12]) ? node18713 : 4'b0001;
																assign node18713 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18716 = (inp[12]) ? 4'b0001 : node18717;
															assign node18717 = (inp[1]) ? 4'b1001 : 4'b0001;
								assign node18721 = (inp[1]) ? node18907 : node18722;
									assign node18722 = (inp[2]) ? node18826 : node18723;
										assign node18723 = (inp[3]) ? node18765 : node18724;
											assign node18724 = (inp[4]) ? node18744 : node18725;
												assign node18725 = (inp[13]) ? node18733 : node18726;
													assign node18726 = (inp[12]) ? 4'b1001 : node18727;
														assign node18727 = (inp[10]) ? node18729 : 4'b1001;
															assign node18729 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node18733 = (inp[7]) ? node18739 : node18734;
														assign node18734 = (inp[12]) ? 4'b0101 : node18735;
															assign node18735 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node18739 = (inp[12]) ? 4'b0001 : node18740;
															assign node18740 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node18744 = (inp[13]) ? node18756 : node18745;
													assign node18745 = (inp[7]) ? node18751 : node18746;
														assign node18746 = (inp[14]) ? node18748 : 4'b0000;
															assign node18748 = (inp[10]) ? 4'b0000 : 4'b1101;
														assign node18751 = (inp[12]) ? 4'b1001 : node18752;
															assign node18752 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node18756 = (inp[10]) ? node18762 : node18757;
														assign node18757 = (inp[12]) ? node18759 : 4'b0000;
															assign node18759 = (inp[7]) ? 4'b0101 : 4'b1000;
														assign node18762 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node18765 = (inp[4]) ? node18801 : node18766;
												assign node18766 = (inp[7]) ? node18776 : node18767;
													assign node18767 = (inp[12]) ? node18771 : node18768;
														assign node18768 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node18771 = (inp[10]) ? 4'b0100 : node18772;
															assign node18772 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node18776 = (inp[13]) ? node18790 : node18777;
														assign node18777 = (inp[14]) ? node18785 : node18778;
															assign node18778 = (inp[10]) ? node18782 : node18779;
																assign node18779 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node18782 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node18785 = (inp[10]) ? 4'b1000 : node18786;
																assign node18786 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node18790 = (inp[14]) ? node18796 : node18791;
															assign node18791 = (inp[12]) ? 4'b0100 : node18792;
																assign node18792 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node18796 = (inp[10]) ? node18798 : 4'b1000;
																assign node18798 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node18801 = (inp[13]) ? node18817 : node18802;
													assign node18802 = (inp[7]) ? node18810 : node18803;
														assign node18803 = (inp[10]) ? node18807 : node18804;
															assign node18804 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node18807 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node18810 = (inp[12]) ? node18814 : node18811;
															assign node18811 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node18814 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node18817 = (inp[10]) ? 4'b0001 : node18818;
														assign node18818 = (inp[7]) ? node18822 : node18819;
															assign node18819 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node18822 = (inp[12]) ? 4'b1100 : 4'b0000;
										assign node18826 = (inp[13]) ? node18866 : node18827;
											assign node18827 = (inp[12]) ? node18853 : node18828;
												assign node18828 = (inp[10]) ? node18840 : node18829;
													assign node18829 = (inp[3]) ? node18835 : node18830;
														assign node18830 = (inp[4]) ? node18832 : 4'b1001;
															assign node18832 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node18835 = (inp[4]) ? node18837 : 4'b1101;
															assign node18837 = (inp[7]) ? 4'b1101 : 4'b0000;
													assign node18840 = (inp[3]) ? node18846 : node18841;
														assign node18841 = (inp[7]) ? node18843 : 4'b0101;
															assign node18843 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node18846 = (inp[4]) ? node18850 : node18847;
															assign node18847 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node18850 = (inp[7]) ? 4'b0001 : 4'b1000;
												assign node18853 = (inp[3]) ? node18859 : node18854;
													assign node18854 = (inp[7]) ? 4'b1001 : node18855;
														assign node18855 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node18859 = (inp[4]) ? node18861 : 4'b1101;
														assign node18861 = (inp[7]) ? 4'b1101 : node18862;
															assign node18862 = (inp[10]) ? 4'b0000 : 4'b1001;
											assign node18866 = (inp[3]) ? node18884 : node18867;
												assign node18867 = (inp[7]) ? node18873 : node18868;
													assign node18868 = (inp[10]) ? node18870 : 4'b0101;
														assign node18870 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node18873 = (inp[4]) ? node18879 : node18874;
														assign node18874 = (inp[12]) ? 4'b0001 : node18875;
															assign node18875 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node18879 = (inp[10]) ? node18881 : 4'b0101;
															assign node18881 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node18884 = (inp[4]) ? node18896 : node18885;
													assign node18885 = (inp[7]) ? node18891 : node18886;
														assign node18886 = (inp[10]) ? node18888 : 4'b0001;
															assign node18888 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node18891 = (inp[10]) ? node18893 : 4'b0101;
															assign node18893 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node18896 = (inp[12]) ? node18900 : node18897;
														assign node18897 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node18900 = (inp[7]) ? node18904 : node18901;
															assign node18901 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node18904 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node18907 = (inp[13]) ? node19031 : node18908;
										assign node18908 = (inp[12]) ? node18968 : node18909;
											assign node18909 = (inp[10]) ? node18943 : node18910;
												assign node18910 = (inp[3]) ? node18924 : node18911;
													assign node18911 = (inp[2]) ? node18919 : node18912;
														assign node18912 = (inp[4]) ? node18916 : node18913;
															assign node18913 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node18916 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node18919 = (inp[7]) ? node18921 : 4'b0100;
															assign node18921 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node18924 = (inp[2]) ? node18938 : node18925;
														assign node18925 = (inp[14]) ? node18931 : node18926;
															assign node18926 = (inp[7]) ? node18928 : 4'b0100;
																assign node18928 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node18931 = (inp[7]) ? node18935 : node18932;
																assign node18932 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node18935 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node18938 = (inp[4]) ? 4'b0000 : node18939;
															assign node18939 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node18943 = (inp[3]) ? node18953 : node18944;
													assign node18944 = (inp[4]) ? node18948 : node18945;
														assign node18945 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node18948 = (inp[2]) ? 4'b0100 : node18949;
															assign node18949 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node18953 = (inp[2]) ? node18961 : node18954;
														assign node18954 = (inp[4]) ? node18958 : node18955;
															assign node18955 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node18958 = (inp[7]) ? 4'b1100 : 4'b0000;
														assign node18961 = (inp[7]) ? node18965 : node18962;
															assign node18962 = (inp[4]) ? 4'b1000 : 4'b0000;
															assign node18965 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node18968 = (inp[10]) ? node19002 : node18969;
												assign node18969 = (inp[3]) ? node18981 : node18970;
													assign node18970 = (inp[2]) ? node18976 : node18971;
														assign node18971 = (inp[4]) ? node18973 : 4'b1000;
															assign node18973 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node18976 = (inp[7]) ? 4'b1000 : node18977;
															assign node18977 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node18981 = (inp[2]) ? node18997 : node18982;
														assign node18982 = (inp[14]) ? node18990 : node18983;
															assign node18983 = (inp[7]) ? node18987 : node18984;
																assign node18984 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node18987 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node18990 = (inp[7]) ? node18994 : node18991;
																assign node18991 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node18994 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node18997 = (inp[4]) ? node18999 : 4'b1100;
															assign node18999 = (inp[7]) ? 4'b1100 : 4'b0000;
												assign node19002 = (inp[2]) ? node19018 : node19003;
													assign node19003 = (inp[3]) ? node19011 : node19004;
														assign node19004 = (inp[4]) ? node19008 : node19005;
															assign node19005 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node19008 = (inp[7]) ? 4'b0100 : 4'b1000;
														assign node19011 = (inp[4]) ? node19015 : node19012;
															assign node19012 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node19015 = (inp[7]) ? 4'b1100 : 4'b0000;
													assign node19018 = (inp[3]) ? node19024 : node19019;
														assign node19019 = (inp[4]) ? 4'b0100 : node19020;
															assign node19020 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node19024 = (inp[4]) ? node19028 : node19025;
															assign node19025 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node19028 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node19031 = (inp[10]) ? node19071 : node19032;
											assign node19032 = (inp[12]) ? node19052 : node19033;
												assign node19033 = (inp[2]) ? node19041 : node19034;
													assign node19034 = (inp[4]) ? 4'b0000 : node19035;
														assign node19035 = (inp[3]) ? 4'b0100 : node19036;
															assign node19036 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node19041 = (inp[3]) ? node19047 : node19042;
														assign node19042 = (inp[7]) ? node19044 : 4'b1100;
															assign node19044 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node19047 = (inp[4]) ? 4'b0000 : node19048;
															assign node19048 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node19052 = (inp[4]) ? node19062 : node19053;
													assign node19053 = (inp[7]) ? node19059 : node19054;
														assign node19054 = (inp[3]) ? node19056 : 4'b0100;
															assign node19056 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node19059 = (inp[3]) ? 4'b0100 : 4'b0000;
													assign node19062 = (inp[2]) ? node19068 : node19063;
														assign node19063 = (inp[7]) ? 4'b0000 : node19064;
															assign node19064 = (inp[3]) ? 4'b1000 : 4'b0000;
														assign node19068 = (inp[3]) ? 4'b0000 : 4'b0100;
											assign node19071 = (inp[4]) ? node19099 : node19072;
												assign node19072 = (inp[2]) ? node19078 : node19073;
													assign node19073 = (inp[7]) ? node19075 : 4'b1100;
														assign node19075 = (inp[3]) ? 4'b1100 : 4'b1000;
													assign node19078 = (inp[12]) ? node19086 : node19079;
														assign node19079 = (inp[3]) ? node19083 : node19080;
															assign node19080 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node19083 = (inp[7]) ? 4'b1100 : 4'b1000;
														assign node19086 = (inp[14]) ? node19094 : node19087;
															assign node19087 = (inp[3]) ? node19091 : node19088;
																assign node19088 = (inp[7]) ? 4'b1000 : 4'b1100;
																assign node19091 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node19094 = (inp[7]) ? 4'b1000 : node19095;
																assign node19095 = (inp[3]) ? 4'b1000 : 4'b1100;
												assign node19099 = (inp[3]) ? 4'b1000 : node19100;
													assign node19100 = (inp[2]) ? 4'b1100 : 4'b1000;
							assign node19104 = (inp[3]) ? node19552 : node19105;
								assign node19105 = (inp[4]) ? node19339 : node19106;
									assign node19106 = (inp[11]) ? node19244 : node19107;
										assign node19107 = (inp[2]) ? node19185 : node19108;
											assign node19108 = (inp[13]) ? node19154 : node19109;
												assign node19109 = (inp[7]) ? node19129 : node19110;
													assign node19110 = (inp[10]) ? node19120 : node19111;
														assign node19111 = (inp[1]) ? node19117 : node19112;
															assign node19112 = (inp[14]) ? 4'b1001 : node19113;
																assign node19113 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node19117 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node19120 = (inp[14]) ? node19124 : node19121;
															assign node19121 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node19124 = (inp[1]) ? 4'b1100 : node19125;
																assign node19125 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node19129 = (inp[1]) ? node19141 : node19130;
														assign node19130 = (inp[14]) ? node19136 : node19131;
															assign node19131 = (inp[10]) ? 4'b1000 : node19132;
																assign node19132 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19136 = (inp[12]) ? node19138 : 4'b1001;
																assign node19138 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node19141 = (inp[14]) ? node19149 : node19142;
															assign node19142 = (inp[12]) ? node19146 : node19143;
																assign node19143 = (inp[10]) ? 4'b0101 : 4'b0001;
																assign node19146 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node19149 = (inp[10]) ? node19151 : 4'b0000;
																assign node19151 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node19154 = (inp[7]) ? node19166 : node19155;
													assign node19155 = (inp[12]) ? node19159 : node19156;
														assign node19156 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node19159 = (inp[1]) ? 4'b0000 : node19160;
															assign node19160 = (inp[10]) ? 4'b1000 : node19161;
																assign node19161 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node19166 = (inp[10]) ? node19176 : node19167;
														assign node19167 = (inp[1]) ? node19173 : node19168;
															assign node19168 = (inp[14]) ? 4'b0101 : node19169;
																assign node19169 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node19173 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node19176 = (inp[12]) ? node19180 : node19177;
															assign node19177 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node19180 = (inp[1]) ? 4'b0000 : node19181;
																assign node19181 = (inp[14]) ? 4'b1101 : 4'b0100;
											assign node19185 = (inp[10]) ? node19205 : node19186;
												assign node19186 = (inp[7]) ? node19198 : node19187;
													assign node19187 = (inp[13]) ? node19193 : node19188;
														assign node19188 = (inp[12]) ? 4'b1001 : node19189;
															assign node19189 = (inp[1]) ? 4'b0101 : 4'b1001;
														assign node19193 = (inp[1]) ? node19195 : 4'b1101;
															assign node19195 = (inp[12]) ? 4'b1101 : 4'b0101;
													assign node19198 = (inp[1]) ? node19200 : 4'b1001;
														assign node19200 = (inp[12]) ? 4'b1001 : node19201;
															assign node19201 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node19205 = (inp[1]) ? node19223 : node19206;
													assign node19206 = (inp[14]) ? node19214 : node19207;
														assign node19207 = (inp[7]) ? node19211 : node19208;
															assign node19208 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node19211 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node19214 = (inp[12]) ? 4'b0101 : node19215;
															assign node19215 = (inp[13]) ? node19219 : node19216;
																assign node19216 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node19219 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node19223 = (inp[12]) ? node19235 : node19224;
														assign node19224 = (inp[14]) ? node19232 : node19225;
															assign node19225 = (inp[13]) ? node19229 : node19226;
																assign node19226 = (inp[7]) ? 4'b1001 : 4'b1101;
																assign node19229 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node19232 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node19235 = (inp[7]) ? node19241 : node19236;
															assign node19236 = (inp[13]) ? node19238 : 4'b0101;
																assign node19238 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node19241 = (inp[13]) ? 4'b0101 : 4'b0001;
										assign node19244 = (inp[1]) ? node19304 : node19245;
											assign node19245 = (inp[2]) ? node19267 : node19246;
												assign node19246 = (inp[13]) ? node19260 : node19247;
													assign node19247 = (inp[7]) ? node19255 : node19248;
														assign node19248 = (inp[12]) ? node19252 : node19249;
															assign node19249 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node19252 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node19255 = (inp[10]) ? 4'b1001 : node19256;
															assign node19256 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node19260 = (inp[7]) ? node19262 : 4'b0000;
														assign node19262 = (inp[10]) ? 4'b0000 : node19263;
															assign node19263 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node19267 = (inp[7]) ? node19281 : node19268;
													assign node19268 = (inp[13]) ? node19276 : node19269;
														assign node19269 = (inp[10]) ? node19273 : node19270;
															assign node19270 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node19273 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19276 = (inp[10]) ? 4'b0001 : node19277;
															assign node19277 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node19281 = (inp[13]) ? node19297 : node19282;
														assign node19282 = (inp[14]) ? node19290 : node19283;
															assign node19283 = (inp[10]) ? node19287 : node19284;
																assign node19284 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node19287 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19290 = (inp[10]) ? node19294 : node19291;
																assign node19291 = (inp[12]) ? 4'b1000 : 4'b0000;
																assign node19294 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19297 = (inp[10]) ? node19301 : node19298;
															assign node19298 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node19301 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node19304 = (inp[10]) ? node19328 : node19305;
												assign node19305 = (inp[2]) ? node19319 : node19306;
													assign node19306 = (inp[7]) ? node19312 : node19307;
														assign node19307 = (inp[13]) ? 4'b1000 : node19308;
															assign node19308 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node19312 = (inp[13]) ? node19316 : node19313;
															assign node19313 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19316 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node19319 = (inp[7]) ? node19325 : node19320;
														assign node19320 = (inp[12]) ? 4'b0100 : node19321;
															assign node19321 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node19325 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node19328 = (inp[13]) ? node19334 : node19329;
													assign node19329 = (inp[2]) ? node19331 : 4'b0100;
														assign node19331 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node19334 = (inp[7]) ? node19336 : 4'b1000;
														assign node19336 = (inp[2]) ? 4'b1100 : 4'b1000;
									assign node19339 = (inp[1]) ? node19457 : node19340;
										assign node19340 = (inp[13]) ? node19392 : node19341;
											assign node19341 = (inp[2]) ? node19367 : node19342;
												assign node19342 = (inp[11]) ? node19358 : node19343;
													assign node19343 = (inp[12]) ? node19351 : node19344;
														assign node19344 = (inp[14]) ? 4'b0000 : node19345;
															assign node19345 = (inp[10]) ? node19347 : 4'b0100;
																assign node19347 = (inp[7]) ? 4'b0100 : 4'b0001;
														assign node19351 = (inp[7]) ? 4'b1000 : node19352;
															assign node19352 = (inp[14]) ? node19354 : 4'b0001;
																assign node19354 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node19358 = (inp[7]) ? node19364 : node19359;
														assign node19359 = (inp[10]) ? node19361 : 4'b0100;
															assign node19361 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node19364 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node19367 = (inp[10]) ? node19385 : node19368;
													assign node19368 = (inp[12]) ? node19378 : node19369;
														assign node19369 = (inp[14]) ? node19373 : node19370;
															assign node19370 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node19373 = (inp[11]) ? 4'b0001 : node19374;
																assign node19374 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node19378 = (inp[7]) ? node19382 : node19379;
															assign node19379 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node19382 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node19385 = (inp[11]) ? 4'b1001 : node19386;
														assign node19386 = (inp[14]) ? node19388 : 4'b1000;
															assign node19388 = (inp[12]) ? 4'b0001 : 4'b1001;
											assign node19392 = (inp[2]) ? node19424 : node19393;
												assign node19393 = (inp[14]) ? node19409 : node19394;
													assign node19394 = (inp[11]) ? node19402 : node19395;
														assign node19395 = (inp[12]) ? node19397 : 4'b1001;
															assign node19397 = (inp[10]) ? node19399 : 4'b0001;
																assign node19399 = (inp[7]) ? 4'b1001 : 4'b0001;
														assign node19402 = (inp[10]) ? node19404 : 4'b1001;
															assign node19404 = (inp[12]) ? node19406 : 4'b0000;
																assign node19406 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node19409 = (inp[11]) ? node19419 : node19410;
														assign node19410 = (inp[12]) ? node19416 : node19411;
															assign node19411 = (inp[10]) ? node19413 : 4'b1000;
																assign node19413 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node19416 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19419 = (inp[10]) ? node19421 : 4'b1001;
															assign node19421 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node19424 = (inp[7]) ? node19436 : node19425;
													assign node19425 = (inp[11]) ? 4'b0000 : node19426;
														assign node19426 = (inp[10]) ? node19432 : node19427;
															assign node19427 = (inp[12]) ? node19429 : 4'b0000;
																assign node19429 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node19432 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19436 = (inp[14]) ? node19448 : node19437;
														assign node19437 = (inp[11]) ? node19445 : node19438;
															assign node19438 = (inp[10]) ? node19442 : node19439;
																assign node19439 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node19442 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node19445 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node19448 = (inp[11]) ? 4'b1001 : node19449;
															assign node19449 = (inp[12]) ? node19453 : node19450;
																assign node19450 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node19453 = (inp[10]) ? 4'b1001 : 4'b0001;
										assign node19457 = (inp[11]) ? node19521 : node19458;
											assign node19458 = (inp[2]) ? node19492 : node19459;
												assign node19459 = (inp[13]) ? node19481 : node19460;
													assign node19460 = (inp[12]) ? node19474 : node19461;
														assign node19461 = (inp[14]) ? node19467 : node19462;
															assign node19462 = (inp[10]) ? 4'b0000 : node19463;
																assign node19463 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node19467 = (inp[7]) ? node19471 : node19468;
																assign node19468 = (inp[10]) ? 4'b1001 : 4'b1100;
																assign node19471 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node19474 = (inp[7]) ? node19478 : node19475;
															assign node19475 = (inp[10]) ? 4'b1000 : 4'b0100;
															assign node19478 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node19481 = (inp[10]) ? 4'b0001 : node19482;
														assign node19482 = (inp[14]) ? node19486 : node19483;
															assign node19483 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node19486 = (inp[12]) ? 4'b1001 : node19487;
																assign node19487 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node19492 = (inp[14]) ? node19504 : node19493;
													assign node19493 = (inp[13]) ? node19499 : node19494;
														assign node19494 = (inp[7]) ? node19496 : 4'b0101;
															assign node19496 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node19499 = (inp[12]) ? 4'b0000 : node19500;
															assign node19500 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node19504 = (inp[13]) ? node19514 : node19505;
														assign node19505 = (inp[12]) ? node19511 : node19506;
															assign node19506 = (inp[10]) ? node19508 : 4'b0000;
																assign node19508 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node19511 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node19514 = (inp[12]) ? node19516 : 4'b1000;
															assign node19516 = (inp[10]) ? 4'b0000 : node19517;
																assign node19517 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node19521 = (inp[13]) ? node19539 : node19522;
												assign node19522 = (inp[10]) ? node19534 : node19523;
													assign node19523 = (inp[12]) ? node19529 : node19524;
														assign node19524 = (inp[2]) ? 4'b1000 : node19525;
															assign node19525 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node19529 = (inp[2]) ? 4'b0000 : node19530;
															assign node19530 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node19534 = (inp[7]) ? 4'b0000 : node19535;
														assign node19535 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node19539 = (inp[10]) ? 4'b1000 : node19540;
													assign node19540 = (inp[2]) ? node19546 : node19541;
														assign node19541 = (inp[7]) ? node19543 : 4'b0000;
															assign node19543 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19546 = (inp[12]) ? 4'b1000 : node19547;
															assign node19547 = (inp[14]) ? 4'b0100 : 4'b1000;
								assign node19552 = (inp[1]) ? node19798 : node19553;
									assign node19553 = (inp[13]) ? node19681 : node19554;
										assign node19554 = (inp[7]) ? node19618 : node19555;
											assign node19555 = (inp[10]) ? node19593 : node19556;
												assign node19556 = (inp[2]) ? node19572 : node19557;
													assign node19557 = (inp[12]) ? node19565 : node19558;
														assign node19558 = (inp[4]) ? 4'b1001 : node19559;
															assign node19559 = (inp[11]) ? 4'b1001 : node19560;
																assign node19560 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19565 = (inp[4]) ? 4'b0001 : node19566;
															assign node19566 = (inp[14]) ? 4'b1001 : node19567;
																assign node19567 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node19572 = (inp[12]) ? node19580 : node19573;
														assign node19573 = (inp[14]) ? node19575 : 4'b0001;
															assign node19575 = (inp[4]) ? 4'b0001 : node19576;
																assign node19576 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node19580 = (inp[14]) ? node19588 : node19581;
															assign node19581 = (inp[11]) ? node19585 : node19582;
																assign node19582 = (inp[4]) ? 4'b0001 : 4'b1000;
																assign node19585 = (inp[4]) ? 4'b1000 : 4'b0001;
															assign node19588 = (inp[4]) ? node19590 : 4'b0001;
																assign node19590 = (inp[11]) ? 4'b1000 : 4'b0001;
												assign node19593 = (inp[2]) ? node19603 : node19594;
													assign node19594 = (inp[4]) ? node19598 : node19595;
														assign node19595 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node19598 = (inp[12]) ? node19600 : 4'b0000;
															assign node19600 = (inp[11]) ? 4'b0001 : 4'b1000;
													assign node19603 = (inp[12]) ? node19611 : node19604;
														assign node19604 = (inp[4]) ? 4'b0001 : node19605;
															assign node19605 = (inp[11]) ? 4'b0000 : node19606;
																assign node19606 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19611 = (inp[11]) ? 4'b0001 : node19612;
															assign node19612 = (inp[4]) ? node19614 : 4'b0001;
																assign node19614 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node19618 = (inp[10]) ? node19654 : node19619;
												assign node19619 = (inp[11]) ? node19641 : node19620;
													assign node19620 = (inp[2]) ? node19632 : node19621;
														assign node19621 = (inp[4]) ? node19625 : node19622;
															assign node19622 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node19625 = (inp[14]) ? node19629 : node19626;
																assign node19626 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node19629 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node19632 = (inp[12]) ? node19638 : node19633;
															assign node19633 = (inp[14]) ? 4'b0000 : node19634;
																assign node19634 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node19638 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node19641 = (inp[4]) ? node19647 : node19642;
														assign node19642 = (inp[12]) ? 4'b0000 : node19643;
															assign node19643 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node19647 = (inp[12]) ? node19651 : node19648;
															assign node19648 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node19651 = (inp[2]) ? 4'b1001 : 4'b0000;
												assign node19654 = (inp[4]) ? node19668 : node19655;
													assign node19655 = (inp[11]) ? node19663 : node19656;
														assign node19656 = (inp[2]) ? node19660 : node19657;
															assign node19657 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node19660 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node19663 = (inp[2]) ? node19665 : 4'b0001;
															assign node19665 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node19668 = (inp[12]) ? node19674 : node19669;
														assign node19669 = (inp[11]) ? 4'b0000 : node19670;
															assign node19670 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node19674 = (inp[2]) ? node19678 : node19675;
															assign node19675 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node19678 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node19681 = (inp[4]) ? node19747 : node19682;
											assign node19682 = (inp[7]) ? node19724 : node19683;
												assign node19683 = (inp[10]) ? node19707 : node19684;
													assign node19684 = (inp[11]) ? node19692 : node19685;
														assign node19685 = (inp[2]) ? node19689 : node19686;
															assign node19686 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node19689 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node19692 = (inp[14]) ? node19700 : node19693;
															assign node19693 = (inp[2]) ? node19697 : node19694;
																assign node19694 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node19697 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node19700 = (inp[12]) ? node19704 : node19701;
																assign node19701 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node19704 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node19707 = (inp[14]) ? node19715 : node19708;
														assign node19708 = (inp[11]) ? node19712 : node19709;
															assign node19709 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node19712 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node19715 = (inp[11]) ? node19721 : node19716;
															assign node19716 = (inp[2]) ? 4'b0000 : node19717;
																assign node19717 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node19721 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node19724 = (inp[10]) ? node19736 : node19725;
													assign node19725 = (inp[11]) ? node19731 : node19726;
														assign node19726 = (inp[2]) ? node19728 : 4'b0000;
															assign node19728 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node19731 = (inp[2]) ? node19733 : 4'b0001;
															assign node19733 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node19736 = (inp[2]) ? node19740 : node19737;
														assign node19737 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node19740 = (inp[11]) ? 4'b1001 : node19741;
															assign node19741 = (inp[14]) ? 4'b0001 : node19742;
																assign node19742 = (inp[12]) ? 4'b0000 : 4'b1000;
											assign node19747 = (inp[10]) ? node19777 : node19748;
												assign node19748 = (inp[2]) ? node19762 : node19749;
													assign node19749 = (inp[7]) ? node19755 : node19750;
														assign node19750 = (inp[11]) ? 4'b0000 : node19751;
															assign node19751 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19755 = (inp[14]) ? node19757 : 4'b0001;
															assign node19757 = (inp[11]) ? node19759 : 4'b0000;
																assign node19759 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node19762 = (inp[7]) ? node19770 : node19763;
														assign node19763 = (inp[12]) ? node19767 : node19764;
															assign node19764 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node19767 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node19770 = (inp[12]) ? node19774 : node19771;
															assign node19771 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node19774 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node19777 = (inp[11]) ? 4'b0000 : node19778;
													assign node19778 = (inp[12]) ? node19786 : node19779;
														assign node19779 = (inp[7]) ? node19781 : 4'b0000;
															assign node19781 = (inp[14]) ? node19783 : 4'b0000;
																assign node19783 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node19786 = (inp[2]) ? node19792 : node19787;
															assign node19787 = (inp[14]) ? node19789 : 4'b0000;
																assign node19789 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node19792 = (inp[14]) ? node19794 : 4'b0001;
																assign node19794 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node19798 = (inp[4]) ? node19896 : node19799;
										assign node19799 = (inp[11]) ? node19857 : node19800;
											assign node19800 = (inp[10]) ? node19842 : node19801;
												assign node19801 = (inp[13]) ? node19823 : node19802;
													assign node19802 = (inp[2]) ? node19812 : node19803;
														assign node19803 = (inp[12]) ? node19807 : node19804;
															assign node19804 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node19807 = (inp[14]) ? node19809 : 4'b1001;
																assign node19809 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19812 = (inp[14]) ? node19818 : node19813;
															assign node19813 = (inp[12]) ? node19815 : 4'b1000;
																assign node19815 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node19818 = (inp[12]) ? node19820 : 4'b1001;
																assign node19820 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node19823 = (inp[12]) ? node19835 : node19824;
														assign node19824 = (inp[2]) ? node19830 : node19825;
															assign node19825 = (inp[14]) ? 4'b1001 : node19826;
																assign node19826 = (inp[7]) ? 4'b0000 : 4'b1001;
															assign node19830 = (inp[7]) ? 4'b1001 : node19831;
																assign node19831 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node19835 = (inp[7]) ? 4'b1001 : node19836;
															assign node19836 = (inp[14]) ? node19838 : 4'b0001;
																assign node19838 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node19842 = (inp[2]) ? node19848 : node19843;
													assign node19843 = (inp[13]) ? node19845 : 4'b0000;
														assign node19845 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19848 = (inp[13]) ? 4'b0000 : node19849;
														assign node19849 = (inp[7]) ? node19851 : 4'b0001;
															assign node19851 = (inp[14]) ? 4'b1001 : node19852;
																assign node19852 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node19857 = (inp[10]) ? node19881 : node19858;
												assign node19858 = (inp[13]) ? node19874 : node19859;
													assign node19859 = (inp[14]) ? node19867 : node19860;
														assign node19860 = (inp[2]) ? node19864 : node19861;
															assign node19861 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19864 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node19867 = (inp[2]) ? node19871 : node19868;
															assign node19868 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node19871 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node19874 = (inp[12]) ? node19876 : 4'b0000;
														assign node19876 = (inp[2]) ? node19878 : 4'b0000;
															assign node19878 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node19881 = (inp[13]) ? 4'b1000 : node19882;
													assign node19882 = (inp[12]) ? node19888 : node19883;
														assign node19883 = (inp[7]) ? 4'b0000 : node19884;
															assign node19884 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node19888 = (inp[7]) ? node19892 : node19889;
															assign node19889 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node19892 = (inp[2]) ? 4'b0000 : 4'b1000;
										assign node19896 = (inp[13]) ? node19946 : node19897;
											assign node19897 = (inp[10]) ? node19931 : node19898;
												assign node19898 = (inp[11]) ? node19918 : node19899;
													assign node19899 = (inp[2]) ? node19909 : node19900;
														assign node19900 = (inp[14]) ? node19904 : node19901;
															assign node19901 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19904 = (inp[12]) ? node19906 : 4'b1000;
																assign node19906 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node19909 = (inp[7]) ? node19915 : node19910;
															assign node19910 = (inp[12]) ? node19912 : 4'b0000;
																assign node19912 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node19915 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node19918 = (inp[7]) ? node19924 : node19919;
														assign node19919 = (inp[2]) ? node19921 : 4'b0000;
															assign node19921 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node19924 = (inp[2]) ? node19928 : node19925;
															assign node19925 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node19928 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node19931 = (inp[11]) ? 4'b0000 : node19932;
													assign node19932 = (inp[7]) ? node19940 : node19933;
														assign node19933 = (inp[14]) ? node19935 : 4'b0000;
															assign node19935 = (inp[12]) ? node19937 : 4'b0001;
																assign node19937 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node19940 = (inp[2]) ? node19942 : 4'b0001;
															assign node19942 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node19946 = (inp[12]) ? node19948 : 4'b0000;
												assign node19948 = (inp[10]) ? 4'b0000 : node19949;
													assign node19949 = (inp[11]) ? 4'b0000 : node19950;
														assign node19950 = (inp[7]) ? node19956 : node19951;
															assign node19951 = (inp[2]) ? 4'b0001 : node19952;
																assign node19952 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node19956 = (inp[14]) ? 4'b0000 : node19957;
																assign node19957 = (inp[2]) ? 4'b0001 : 4'b0000;
					assign node19963 = (inp[6]) ? node19965 : 4'b1000;
						assign node19965 = (inp[5]) ? node20109 : node19966;
							assign node19966 = (inp[3]) ? node19968 : 4'b1000;
								assign node19968 = (inp[2]) ? 4'b1000 : node19969;
									assign node19969 = (inp[4]) ? node20031 : node19970;
										assign node19970 = (inp[7]) ? 4'b1000 : node19971;
											assign node19971 = (inp[13]) ? node19997 : node19972;
												assign node19972 = (inp[10]) ? node19982 : node19973;
													assign node19973 = (inp[1]) ? node19975 : 4'b1000;
														assign node19975 = (inp[12]) ? 4'b1000 : node19976;
															assign node19976 = (inp[11]) ? 4'b0000 : node19977;
																assign node19977 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node19982 = (inp[12]) ? node19994 : node19983;
														assign node19983 = (inp[1]) ? node19989 : node19984;
															assign node19984 = (inp[11]) ? 4'b0001 : node19985;
																assign node19985 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node19989 = (inp[14]) ? node19991 : 4'b0000;
																assign node19991 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node19994 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node19997 = (inp[1]) ? node20013 : node19998;
													assign node19998 = (inp[12]) ? node20008 : node19999;
														assign node19999 = (inp[10]) ? node20003 : node20000;
															assign node20000 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20003 = (inp[14]) ? node20005 : 4'b1001;
																assign node20005 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20008 = (inp[14]) ? node20010 : 4'b0001;
															assign node20010 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node20013 = (inp[10]) ? node20025 : node20014;
														assign node20014 = (inp[12]) ? node20020 : node20015;
															assign node20015 = (inp[11]) ? 4'b1000 : node20016;
																assign node20016 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node20020 = (inp[11]) ? 4'b0000 : node20021;
																assign node20021 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20025 = (inp[14]) ? node20027 : 4'b1000;
															assign node20027 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node20031 = (inp[1]) ? node20071 : node20032;
											assign node20032 = (inp[13]) ? node20054 : node20033;
												assign node20033 = (inp[12]) ? node20047 : node20034;
													assign node20034 = (inp[10]) ? node20042 : node20035;
														assign node20035 = (inp[7]) ? 4'b1000 : node20036;
															assign node20036 = (inp[14]) ? node20038 : 4'b1001;
																assign node20038 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20042 = (inp[14]) ? node20044 : 4'b0001;
															assign node20044 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node20047 = (inp[7]) ? 4'b1000 : node20048;
														assign node20048 = (inp[11]) ? 4'b1001 : node20049;
															assign node20049 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node20054 = (inp[11]) ? node20066 : node20055;
													assign node20055 = (inp[14]) ? node20061 : node20056;
														assign node20056 = (inp[12]) ? 4'b0001 : node20057;
															assign node20057 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node20061 = (inp[12]) ? 4'b0000 : node20062;
															assign node20062 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node20066 = (inp[12]) ? 4'b0001 : node20067;
														assign node20067 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node20071 = (inp[14]) ? node20083 : node20072;
												assign node20072 = (inp[13]) ? node20078 : node20073;
													assign node20073 = (inp[12]) ? node20075 : 4'b0000;
														assign node20075 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node20078 = (inp[10]) ? 4'b1000 : node20079;
														assign node20079 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node20083 = (inp[11]) ? node20097 : node20084;
													assign node20084 = (inp[13]) ? node20092 : node20085;
														assign node20085 = (inp[7]) ? 4'b1000 : node20086;
															assign node20086 = (inp[12]) ? 4'b1001 : node20087;
																assign node20087 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node20092 = (inp[12]) ? 4'b0001 : node20093;
															assign node20093 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node20097 = (inp[13]) ? node20103 : node20098;
														assign node20098 = (inp[10]) ? 4'b0000 : node20099;
															assign node20099 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node20103 = (inp[12]) ? node20105 : 4'b1000;
															assign node20105 = (inp[10]) ? 4'b1000 : 4'b0000;
							assign node20109 = (inp[2]) ? node20573 : node20110;
								assign node20110 = (inp[3]) ? node20344 : node20111;
									assign node20111 = (inp[1]) ? node20221 : node20112;
										assign node20112 = (inp[13]) ? node20176 : node20113;
											assign node20113 = (inp[10]) ? node20137 : node20114;
												assign node20114 = (inp[14]) ? node20120 : node20115;
													assign node20115 = (inp[7]) ? 4'b1001 : node20116;
														assign node20116 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node20120 = (inp[11]) ? node20126 : node20121;
														assign node20121 = (inp[4]) ? node20123 : 4'b1000;
															assign node20123 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node20126 = (inp[12]) ? node20132 : node20127;
															assign node20127 = (inp[4]) ? node20129 : 4'b1001;
																assign node20129 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node20132 = (inp[7]) ? 4'b1001 : node20133;
																assign node20133 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node20137 = (inp[12]) ? node20159 : node20138;
													assign node20138 = (inp[14]) ? node20148 : node20139;
														assign node20139 = (inp[4]) ? node20143 : node20140;
															assign node20140 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node20143 = (inp[7]) ? 4'b0101 : node20144;
																assign node20144 = (inp[11]) ? 4'b1000 : 4'b0001;
														assign node20148 = (inp[4]) ? node20156 : node20149;
															assign node20149 = (inp[7]) ? node20153 : node20150;
																assign node20150 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node20153 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20156 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node20159 = (inp[14]) ? node20165 : node20160;
														assign node20160 = (inp[7]) ? 4'b1001 : node20161;
															assign node20161 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node20165 = (inp[7]) ? node20173 : node20166;
															assign node20166 = (inp[4]) ? node20170 : node20167;
																assign node20167 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node20170 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node20173 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20176 = (inp[4]) ? node20202 : node20177;
												assign node20177 = (inp[7]) ? node20187 : node20178;
													assign node20178 = (inp[10]) ? node20184 : node20179;
														assign node20179 = (inp[14]) ? node20181 : 4'b0101;
															assign node20181 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node20184 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node20187 = (inp[12]) ? node20197 : node20188;
														assign node20188 = (inp[10]) ? node20192 : node20189;
															assign node20189 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20192 = (inp[11]) ? 4'b1001 : node20193;
																assign node20193 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node20197 = (inp[11]) ? 4'b0001 : node20198;
															assign node20198 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node20202 = (inp[11]) ? node20210 : node20203;
													assign node20203 = (inp[10]) ? 4'b0001 : node20204;
														assign node20204 = (inp[7]) ? node20206 : 4'b1001;
															assign node20206 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node20210 = (inp[12]) ? node20214 : node20211;
														assign node20211 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node20214 = (inp[7]) ? node20218 : node20215;
															assign node20215 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node20218 = (inp[10]) ? 4'b0000 : 4'b0101;
										assign node20221 = (inp[11]) ? node20307 : node20222;
											assign node20222 = (inp[14]) ? node20270 : node20223;
												assign node20223 = (inp[4]) ? node20243 : node20224;
													assign node20224 = (inp[7]) ? node20232 : node20225;
														assign node20225 = (inp[13]) ? 4'b1100 : node20226;
															assign node20226 = (inp[10]) ? 4'b0100 : node20227;
																assign node20227 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node20232 = (inp[13]) ? node20238 : node20233;
															assign node20233 = (inp[12]) ? node20235 : 4'b0000;
																assign node20235 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node20238 = (inp[10]) ? 4'b1000 : node20239;
																assign node20239 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20243 = (inp[7]) ? node20259 : node20244;
														assign node20244 = (inp[13]) ? node20252 : node20245;
															assign node20245 = (inp[10]) ? node20249 : node20246;
																assign node20246 = (inp[12]) ? 4'b1100 : 4'b0001;
																assign node20249 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20252 = (inp[10]) ? node20256 : node20253;
																assign node20253 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node20256 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20259 = (inp[13]) ? node20265 : node20260;
															assign node20260 = (inp[12]) ? node20262 : 4'b0100;
																assign node20262 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node20265 = (inp[12]) ? node20267 : 4'b0001;
																assign node20267 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node20270 = (inp[13]) ? node20292 : node20271;
													assign node20271 = (inp[10]) ? node20279 : node20272;
														assign node20272 = (inp[7]) ? 4'b1001 : node20273;
															assign node20273 = (inp[12]) ? 4'b1101 : node20274;
																assign node20274 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node20279 = (inp[12]) ? node20287 : node20280;
															assign node20280 = (inp[4]) ? node20284 : node20281;
																assign node20281 = (inp[7]) ? 4'b0001 : 4'b0101;
																assign node20284 = (inp[7]) ? 4'b0101 : 4'b1001;
															assign node20287 = (inp[4]) ? node20289 : 4'b1001;
																assign node20289 = (inp[7]) ? 4'b1001 : 4'b0001;
													assign node20292 = (inp[10]) ? node20300 : node20293;
														assign node20293 = (inp[7]) ? node20295 : 4'b0101;
															assign node20295 = (inp[4]) ? node20297 : 4'b0001;
																assign node20297 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node20300 = (inp[12]) ? node20302 : 4'b1001;
															assign node20302 = (inp[7]) ? 4'b0001 : node20303;
																assign node20303 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node20307 = (inp[10]) ? node20331 : node20308;
												assign node20308 = (inp[4]) ? node20324 : node20309;
													assign node20309 = (inp[7]) ? node20317 : node20310;
														assign node20310 = (inp[13]) ? node20314 : node20311;
															assign node20311 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node20314 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node20317 = (inp[13]) ? node20321 : node20318;
															assign node20318 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node20321 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20324 = (inp[13]) ? 4'b0000 : node20325;
														assign node20325 = (inp[7]) ? node20327 : 4'b0000;
															assign node20327 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node20331 = (inp[13]) ? node20339 : node20332;
													assign node20332 = (inp[4]) ? node20336 : node20333;
														assign node20333 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20336 = (inp[7]) ? 4'b0100 : 4'b1000;
													assign node20339 = (inp[7]) ? 4'b1000 : node20340;
														assign node20340 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node20344 = (inp[4]) ? node20470 : node20345;
										assign node20345 = (inp[11]) ? node20419 : node20346;
											assign node20346 = (inp[13]) ? node20378 : node20347;
												assign node20347 = (inp[1]) ? node20359 : node20348;
													assign node20348 = (inp[7]) ? node20356 : node20349;
														assign node20349 = (inp[14]) ? 4'b1001 : node20350;
															assign node20350 = (inp[10]) ? 4'b1000 : node20351;
																assign node20351 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node20356 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node20359 = (inp[14]) ? node20369 : node20360;
														assign node20360 = (inp[12]) ? node20362 : 4'b0001;
															assign node20362 = (inp[10]) ? node20366 : node20363;
																assign node20363 = (inp[7]) ? 4'b1001 : 4'b0001;
																assign node20366 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node20369 = (inp[7]) ? node20375 : node20370;
															assign node20370 = (inp[10]) ? node20372 : 4'b0000;
																assign node20372 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node20375 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node20378 = (inp[14]) ? node20398 : node20379;
													assign node20379 = (inp[1]) ? node20391 : node20380;
														assign node20380 = (inp[12]) ? node20386 : node20381;
															assign node20381 = (inp[10]) ? 4'b0000 : node20382;
																assign node20382 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node20386 = (inp[10]) ? node20388 : 4'b0000;
																assign node20388 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node20391 = (inp[12]) ? node20393 : 4'b1000;
															assign node20393 = (inp[10]) ? 4'b0000 : node20394;
																assign node20394 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node20398 = (inp[1]) ? node20410 : node20399;
														assign node20399 = (inp[12]) ? node20405 : node20400;
															assign node20400 = (inp[7]) ? node20402 : 4'b0000;
																assign node20402 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node20405 = (inp[10]) ? node20407 : 4'b0001;
																assign node20407 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node20410 = (inp[10]) ? node20416 : node20411;
															assign node20411 = (inp[12]) ? node20413 : 4'b1000;
																assign node20413 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node20416 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node20419 = (inp[1]) ? node20455 : node20420;
												assign node20420 = (inp[13]) ? node20442 : node20421;
													assign node20421 = (inp[7]) ? node20427 : node20422;
														assign node20422 = (inp[10]) ? 4'b1001 : node20423;
															assign node20423 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node20427 = (inp[14]) ? node20435 : node20428;
															assign node20428 = (inp[12]) ? node20432 : node20429;
																assign node20429 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node20432 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node20435 = (inp[12]) ? node20439 : node20436;
																assign node20436 = (inp[10]) ? 4'b1000 : 4'b0000;
																assign node20439 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node20442 = (inp[14]) ? node20444 : 4'b0000;
														assign node20444 = (inp[12]) ? node20450 : node20445;
															assign node20445 = (inp[7]) ? 4'b1001 : node20446;
																assign node20446 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node20450 = (inp[10]) ? 4'b0000 : node20451;
																assign node20451 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node20455 = (inp[13]) ? node20463 : node20456;
													assign node20456 = (inp[7]) ? 4'b0000 : node20457;
														assign node20457 = (inp[12]) ? 4'b0000 : node20458;
															assign node20458 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node20463 = (inp[12]) ? 4'b1000 : node20464;
														assign node20464 = (inp[7]) ? node20466 : 4'b1000;
															assign node20466 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node20470 = (inp[11]) ? node20554 : node20471;
											assign node20471 = (inp[13]) ? node20523 : node20472;
												assign node20472 = (inp[10]) ? node20500 : node20473;
													assign node20473 = (inp[12]) ? node20487 : node20474;
														assign node20474 = (inp[1]) ? node20480 : node20475;
															assign node20475 = (inp[14]) ? node20477 : 4'b0001;
																assign node20477 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node20480 = (inp[7]) ? node20484 : node20481;
																assign node20481 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node20484 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node20487 = (inp[1]) ? node20493 : node20488;
															assign node20488 = (inp[7]) ? 4'b1000 : node20489;
																assign node20489 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node20493 = (inp[14]) ? node20497 : node20494;
																assign node20494 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node20497 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node20500 = (inp[14]) ? node20514 : node20501;
														assign node20501 = (inp[1]) ? node20507 : node20502;
															assign node20502 = (inp[7]) ? node20504 : 4'b0000;
																assign node20504 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node20507 = (inp[12]) ? node20511 : node20508;
																assign node20508 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node20511 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node20514 = (inp[1]) ? node20520 : node20515;
															assign node20515 = (inp[7]) ? node20517 : 4'b0000;
																assign node20517 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20520 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node20523 = (inp[10]) ? node20545 : node20524;
													assign node20524 = (inp[7]) ? node20536 : node20525;
														assign node20525 = (inp[1]) ? node20531 : node20526;
															assign node20526 = (inp[12]) ? 4'b0000 : node20527;
																assign node20527 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20531 = (inp[12]) ? node20533 : 4'b0001;
																assign node20533 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20536 = (inp[12]) ? 4'b0001 : node20537;
															assign node20537 = (inp[1]) ? node20541 : node20538;
																assign node20538 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node20541 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node20545 = (inp[1]) ? 4'b0000 : node20546;
														assign node20546 = (inp[7]) ? node20548 : 4'b0001;
															assign node20548 = (inp[14]) ? 4'b0000 : node20549;
																assign node20549 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node20554 = (inp[1]) ? 4'b0000 : node20555;
												assign node20555 = (inp[13]) ? node20565 : node20556;
													assign node20556 = (inp[7]) ? 4'b0001 : node20557;
														assign node20557 = (inp[10]) ? node20561 : node20558;
															assign node20558 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20561 = (inp[12]) ? 4'b1000 : 4'b0001;
													assign node20565 = (inp[7]) ? 4'b0000 : node20566;
														assign node20566 = (inp[12]) ? 4'b0000 : node20567;
															assign node20567 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node20573 = (inp[3]) ? node20575 : 4'b1000;
									assign node20575 = (inp[4]) ? node20637 : node20576;
										assign node20576 = (inp[7]) ? 4'b1000 : node20577;
											assign node20577 = (inp[13]) ? node20607 : node20578;
												assign node20578 = (inp[12]) ? node20598 : node20579;
													assign node20579 = (inp[10]) ? node20587 : node20580;
														assign node20580 = (inp[1]) ? node20582 : 4'b1000;
															assign node20582 = (inp[14]) ? node20584 : 4'b0000;
																assign node20584 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node20587 = (inp[1]) ? node20593 : node20588;
															assign node20588 = (inp[14]) ? node20590 : 4'b0001;
																assign node20590 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20593 = (inp[14]) ? node20595 : 4'b0000;
																assign node20595 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node20598 = (inp[10]) ? node20600 : 4'b1000;
														assign node20600 = (inp[1]) ? node20602 : 4'b1000;
															assign node20602 = (inp[14]) ? node20604 : 4'b0000;
																assign node20604 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node20607 = (inp[12]) ? node20623 : node20608;
													assign node20608 = (inp[1]) ? node20616 : node20609;
														assign node20609 = (inp[10]) ? node20611 : 4'b0001;
															assign node20611 = (inp[14]) ? node20613 : 4'b1001;
																assign node20613 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20616 = (inp[14]) ? node20618 : 4'b1000;
															assign node20618 = (inp[11]) ? 4'b1000 : node20619;
																assign node20619 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node20623 = (inp[1]) ? node20629 : node20624;
														assign node20624 = (inp[11]) ? 4'b0001 : node20625;
															assign node20625 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20629 = (inp[10]) ? 4'b1000 : node20630;
															assign node20630 = (inp[11]) ? 4'b0000 : node20631;
																assign node20631 = (inp[14]) ? 4'b0001 : 4'b0000;
										assign node20637 = (inp[13]) ? node20695 : node20638;
											assign node20638 = (inp[1]) ? node20662 : node20639;
												assign node20639 = (inp[10]) ? node20649 : node20640;
													assign node20640 = (inp[7]) ? 4'b1000 : node20641;
														assign node20641 = (inp[12]) ? 4'b1001 : node20642;
															assign node20642 = (inp[11]) ? 4'b0000 : node20643;
																assign node20643 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node20649 = (inp[12]) ? node20659 : node20650;
														assign node20650 = (inp[7]) ? node20654 : node20651;
															assign node20651 = (inp[11]) ? 4'b1000 : 4'b0001;
															assign node20654 = (inp[11]) ? 4'b0001 : node20655;
																assign node20655 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node20659 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node20662 = (inp[11]) ? node20688 : node20663;
													assign node20663 = (inp[7]) ? node20675 : node20664;
														assign node20664 = (inp[10]) ? node20670 : node20665;
															assign node20665 = (inp[12]) ? node20667 : 4'b0001;
																assign node20667 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node20670 = (inp[14]) ? node20672 : 4'b0001;
																assign node20672 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node20675 = (inp[12]) ? node20683 : node20676;
															assign node20676 = (inp[10]) ? node20680 : node20677;
																assign node20677 = (inp[14]) ? 4'b1000 : 4'b0000;
																assign node20680 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node20683 = (inp[10]) ? node20685 : 4'b1000;
																assign node20685 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node20688 = (inp[12]) ? node20690 : 4'b0000;
														assign node20690 = (inp[7]) ? node20692 : 4'b0000;
															assign node20692 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node20695 = (inp[11]) ? node20731 : node20696;
												assign node20696 = (inp[10]) ? node20720 : node20697;
													assign node20697 = (inp[7]) ? node20707 : node20698;
														assign node20698 = (inp[14]) ? node20700 : 4'b0000;
															assign node20700 = (inp[12]) ? node20704 : node20701;
																assign node20701 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node20704 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node20707 = (inp[12]) ? node20713 : node20708;
															assign node20708 = (inp[14]) ? node20710 : 4'b0001;
																assign node20710 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node20713 = (inp[1]) ? node20717 : node20714;
																assign node20714 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node20717 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node20720 = (inp[1]) ? 4'b0000 : node20721;
														assign node20721 = (inp[7]) ? node20727 : node20722;
															assign node20722 = (inp[12]) ? 4'b0000 : node20723;
																assign node20723 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node20727 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node20731 = (inp[1]) ? 4'b0000 : node20732;
													assign node20732 = (inp[7]) ? node20734 : 4'b0000;
														assign node20734 = (inp[10]) ? 4'b0000 : node20735;
															assign node20735 = (inp[12]) ? 4'b0001 : 4'b0000;
			assign node20740 = (inp[15]) ? node24428 : node20741;
				assign node20741 = (inp[6]) ? node21637 : node20742;
					assign node20742 = (inp[0]) ? 4'b0100 : node20743;
						assign node20743 = (inp[5]) ? node21097 : node20744;
							assign node20744 = (inp[2]) ? 4'b0110 : node20745;
								assign node20745 = (inp[3]) ? node20877 : node20746;
									assign node20746 = (inp[4]) ? node20780 : node20747;
										assign node20747 = (inp[7]) ? 4'b0110 : node20748;
											assign node20748 = (inp[13]) ? node20750 : 4'b0110;
												assign node20750 = (inp[10]) ? node20760 : node20751;
													assign node20751 = (inp[12]) ? 4'b0110 : node20752;
														assign node20752 = (inp[1]) ? node20754 : 4'b0110;
															assign node20754 = (inp[11]) ? 4'b0000 : node20755;
																assign node20755 = (inp[14]) ? 4'b0110 : 4'b0000;
													assign node20760 = (inp[12]) ? node20772 : node20761;
														assign node20761 = (inp[1]) ? node20767 : node20762;
															assign node20762 = (inp[14]) ? node20764 : 4'b0001;
																assign node20764 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20767 = (inp[14]) ? node20769 : 4'b0000;
																assign node20769 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node20772 = (inp[1]) ? node20774 : 4'b0110;
															assign node20774 = (inp[11]) ? 4'b0000 : node20775;
																assign node20775 = (inp[14]) ? 4'b0110 : 4'b0000;
										assign node20780 = (inp[7]) ? node20852 : node20781;
											assign node20781 = (inp[1]) ? node20817 : node20782;
												assign node20782 = (inp[13]) ? node20800 : node20783;
													assign node20783 = (inp[14]) ? node20789 : node20784;
														assign node20784 = (inp[12]) ? 4'b0001 : node20785;
															assign node20785 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node20789 = (inp[11]) ? node20795 : node20790;
															assign node20790 = (inp[10]) ? node20792 : 4'b0000;
																assign node20792 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20795 = (inp[10]) ? node20797 : 4'b0001;
																assign node20797 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node20800 = (inp[11]) ? node20812 : node20801;
														assign node20801 = (inp[14]) ? node20807 : node20802;
															assign node20802 = (inp[10]) ? node20804 : 4'b1001;
																assign node20804 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node20807 = (inp[12]) ? 4'b1000 : node20808;
																assign node20808 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node20812 = (inp[12]) ? 4'b1001 : node20813;
															assign node20813 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node20817 = (inp[14]) ? node20829 : node20818;
													assign node20818 = (inp[13]) ? node20824 : node20819;
														assign node20819 = (inp[12]) ? node20821 : 4'b1000;
															assign node20821 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node20824 = (inp[10]) ? 4'b0000 : node20825;
															assign node20825 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node20829 = (inp[11]) ? node20841 : node20830;
														assign node20830 = (inp[13]) ? node20836 : node20831;
															assign node20831 = (inp[10]) ? node20833 : 4'b0001;
																assign node20833 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node20836 = (inp[10]) ? node20838 : 4'b1001;
																assign node20838 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node20841 = (inp[13]) ? node20847 : node20842;
															assign node20842 = (inp[10]) ? 4'b1000 : node20843;
																assign node20843 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node20847 = (inp[12]) ? node20849 : 4'b0000;
																assign node20849 = (inp[10]) ? 4'b0000 : 4'b1000;
											assign node20852 = (inp[13]) ? node20854 : 4'b0110;
												assign node20854 = (inp[10]) ? node20860 : node20855;
													assign node20855 = (inp[12]) ? 4'b0110 : node20856;
														assign node20856 = (inp[1]) ? 4'b0000 : 4'b0110;
													assign node20860 = (inp[12]) ? node20870 : node20861;
														assign node20861 = (inp[1]) ? node20865 : node20862;
															assign node20862 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20865 = (inp[11]) ? 4'b0000 : node20866;
																assign node20866 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node20870 = (inp[1]) ? node20872 : 4'b0110;
															assign node20872 = (inp[11]) ? 4'b0000 : node20873;
																assign node20873 = (inp[14]) ? 4'b0110 : 4'b0000;
									assign node20877 = (inp[4]) ? node20967 : node20878;
										assign node20878 = (inp[1]) ? node20920 : node20879;
											assign node20879 = (inp[13]) ? node20897 : node20880;
												assign node20880 = (inp[10]) ? node20886 : node20881;
													assign node20881 = (inp[14]) ? node20883 : 4'b0001;
														assign node20883 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node20886 = (inp[12]) ? node20892 : node20887;
														assign node20887 = (inp[14]) ? node20889 : 4'b1001;
															assign node20889 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20892 = (inp[11]) ? 4'b0001 : node20893;
															assign node20893 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node20897 = (inp[12]) ? node20915 : node20898;
													assign node20898 = (inp[10]) ? node20904 : node20899;
														assign node20899 = (inp[14]) ? node20901 : 4'b1001;
															assign node20901 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node20904 = (inp[7]) ? node20910 : node20905;
															assign node20905 = (inp[14]) ? node20907 : 4'b0101;
																assign node20907 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node20910 = (inp[14]) ? node20912 : 4'b0001;
																assign node20912 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node20915 = (inp[14]) ? node20917 : 4'b1001;
														assign node20917 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node20920 = (inp[11]) ? node20950 : node20921;
												assign node20921 = (inp[14]) ? node20937 : node20922;
													assign node20922 = (inp[13]) ? node20928 : node20923;
														assign node20923 = (inp[12]) ? node20925 : 4'b1000;
															assign node20925 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node20928 = (inp[7]) ? node20934 : node20929;
															assign node20929 = (inp[10]) ? 4'b0100 : node20930;
																assign node20930 = (inp[12]) ? 4'b1000 : 4'b0100;
															assign node20934 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node20937 = (inp[13]) ? node20943 : node20938;
														assign node20938 = (inp[10]) ? node20940 : 4'b0001;
															assign node20940 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node20943 = (inp[10]) ? node20945 : 4'b1001;
															assign node20945 = (inp[12]) ? 4'b1001 : node20946;
																assign node20946 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node20950 = (inp[13]) ? node20956 : node20951;
													assign node20951 = (inp[10]) ? 4'b1000 : node20952;
														assign node20952 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node20956 = (inp[7]) ? node20962 : node20957;
														assign node20957 = (inp[12]) ? node20959 : 4'b0100;
															assign node20959 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node20962 = (inp[10]) ? 4'b0000 : node20963;
															assign node20963 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node20967 = (inp[7]) ? node21037 : node20968;
											assign node20968 = (inp[1]) ? node21004 : node20969;
												assign node20969 = (inp[11]) ? node20993 : node20970;
													assign node20970 = (inp[14]) ? node20982 : node20971;
														assign node20971 = (inp[13]) ? node20977 : node20972;
															assign node20972 = (inp[10]) ? node20974 : 4'b0101;
																assign node20974 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node20977 = (inp[12]) ? 4'b1101 : node20978;
																assign node20978 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node20982 = (inp[13]) ? node20988 : node20983;
															assign node20983 = (inp[10]) ? node20985 : 4'b0100;
																assign node20985 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node20988 = (inp[10]) ? node20990 : 4'b1100;
																assign node20990 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node20993 = (inp[13]) ? node20999 : node20994;
														assign node20994 = (inp[10]) ? node20996 : 4'b0101;
															assign node20996 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node20999 = (inp[10]) ? node21001 : 4'b1101;
															assign node21001 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node21004 = (inp[11]) ? node21026 : node21005;
													assign node21005 = (inp[14]) ? node21015 : node21006;
														assign node21006 = (inp[10]) ? node21012 : node21007;
															assign node21007 = (inp[13]) ? 4'b1100 : node21008;
																assign node21008 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node21012 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node21015 = (inp[13]) ? node21021 : node21016;
															assign node21016 = (inp[12]) ? 4'b0101 : node21017;
																assign node21017 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node21021 = (inp[12]) ? 4'b1101 : node21022;
																assign node21022 = (inp[10]) ? 4'b0101 : 4'b1101;
													assign node21026 = (inp[13]) ? node21032 : node21027;
														assign node21027 = (inp[12]) ? node21029 : 4'b1100;
															assign node21029 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node21032 = (inp[10]) ? 4'b0100 : node21033;
															assign node21033 = (inp[12]) ? 4'b1100 : 4'b0100;
											assign node21037 = (inp[1]) ? node21067 : node21038;
												assign node21038 = (inp[14]) ? node21050 : node21039;
													assign node21039 = (inp[13]) ? node21045 : node21040;
														assign node21040 = (inp[12]) ? 4'b0001 : node21041;
															assign node21041 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node21045 = (inp[12]) ? 4'b1001 : node21046;
															assign node21046 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node21050 = (inp[11]) ? node21062 : node21051;
														assign node21051 = (inp[13]) ? node21057 : node21052;
															assign node21052 = (inp[12]) ? 4'b0000 : node21053;
																assign node21053 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node21057 = (inp[10]) ? node21059 : 4'b1000;
																assign node21059 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node21062 = (inp[13]) ? node21064 : 4'b0001;
															assign node21064 = (inp[12]) ? 4'b1001 : 4'b0101;
												assign node21067 = (inp[13]) ? node21079 : node21068;
													assign node21068 = (inp[11]) ? node21074 : node21069;
														assign node21069 = (inp[14]) ? 4'b0001 : node21070;
															assign node21070 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21074 = (inp[12]) ? node21076 : 4'b1000;
															assign node21076 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node21079 = (inp[14]) ? node21085 : node21080;
														assign node21080 = (inp[10]) ? 4'b0100 : node21081;
															assign node21081 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node21085 = (inp[11]) ? node21091 : node21086;
															assign node21086 = (inp[12]) ? 4'b1001 : node21087;
																assign node21087 = (inp[10]) ? 4'b0101 : 4'b1001;
															assign node21091 = (inp[10]) ? 4'b0100 : node21092;
																assign node21092 = (inp[12]) ? 4'b1000 : 4'b0100;
							assign node21097 = (inp[3]) ? node21421 : node21098;
								assign node21098 = (inp[2]) ? node21304 : node21099;
									assign node21099 = (inp[4]) ? node21183 : node21100;
										assign node21100 = (inp[1]) ? node21142 : node21101;
											assign node21101 = (inp[13]) ? node21119 : node21102;
												assign node21102 = (inp[14]) ? node21108 : node21103;
													assign node21103 = (inp[10]) ? node21105 : 4'b0101;
														assign node21105 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21108 = (inp[11]) ? node21114 : node21109;
														assign node21109 = (inp[10]) ? node21111 : 4'b0100;
															assign node21111 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node21114 = (inp[12]) ? 4'b0101 : node21115;
															assign node21115 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node21119 = (inp[12]) ? node21137 : node21120;
													assign node21120 = (inp[10]) ? node21126 : node21121;
														assign node21121 = (inp[14]) ? node21123 : 4'b1101;
															assign node21123 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node21126 = (inp[7]) ? node21132 : node21127;
															assign node21127 = (inp[11]) ? 4'b0001 : node21128;
																assign node21128 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21132 = (inp[11]) ? 4'b0101 : node21133;
																assign node21133 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node21137 = (inp[14]) ? node21139 : 4'b1101;
														assign node21139 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node21142 = (inp[14]) ? node21160 : node21143;
												assign node21143 = (inp[13]) ? node21149 : node21144;
													assign node21144 = (inp[12]) ? node21146 : 4'b1100;
														assign node21146 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node21149 = (inp[7]) ? node21155 : node21150;
														assign node21150 = (inp[12]) ? node21152 : 4'b0000;
															assign node21152 = (inp[10]) ? 4'b0000 : 4'b1100;
														assign node21155 = (inp[10]) ? 4'b0100 : node21156;
															assign node21156 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node21160 = (inp[11]) ? node21168 : node21161;
													assign node21161 = (inp[13]) ? 4'b1101 : node21162;
														assign node21162 = (inp[10]) ? node21164 : 4'b0101;
															assign node21164 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21168 = (inp[13]) ? node21174 : node21169;
														assign node21169 = (inp[12]) ? node21171 : 4'b1100;
															assign node21171 = (inp[7]) ? 4'b1100 : 4'b0100;
														assign node21174 = (inp[7]) ? node21180 : node21175;
															assign node21175 = (inp[12]) ? node21177 : 4'b0000;
																assign node21177 = (inp[10]) ? 4'b0000 : 4'b1100;
															assign node21180 = (inp[10]) ? 4'b0100 : 4'b1100;
										assign node21183 = (inp[7]) ? node21243 : node21184;
											assign node21184 = (inp[1]) ? node21216 : node21185;
												assign node21185 = (inp[13]) ? node21199 : node21186;
													assign node21186 = (inp[12]) ? node21194 : node21187;
														assign node21187 = (inp[10]) ? node21189 : 4'b0001;
															assign node21189 = (inp[11]) ? 4'b1001 : node21190;
																assign node21190 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node21194 = (inp[14]) ? node21196 : 4'b0001;
															assign node21196 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21199 = (inp[12]) ? node21211 : node21200;
														assign node21200 = (inp[10]) ? node21206 : node21201;
															assign node21201 = (inp[11]) ? 4'b1001 : node21202;
																assign node21202 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21206 = (inp[11]) ? 4'b0001 : node21207;
																assign node21207 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node21211 = (inp[14]) ? node21213 : 4'b1001;
															assign node21213 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node21216 = (inp[14]) ? node21228 : node21217;
													assign node21217 = (inp[13]) ? node21223 : node21218;
														assign node21218 = (inp[10]) ? 4'b1000 : node21219;
															assign node21219 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21223 = (inp[10]) ? 4'b0000 : node21224;
															assign node21224 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node21228 = (inp[11]) ? node21238 : node21229;
														assign node21229 = (inp[13]) ? node21235 : node21230;
															assign node21230 = (inp[10]) ? node21232 : 4'b0001;
																assign node21232 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node21235 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node21238 = (inp[13]) ? 4'b0000 : node21239;
															assign node21239 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node21243 = (inp[1]) ? node21275 : node21244;
												assign node21244 = (inp[13]) ? node21258 : node21245;
													assign node21245 = (inp[14]) ? node21251 : node21246;
														assign node21246 = (inp[12]) ? 4'b0101 : node21247;
															assign node21247 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node21251 = (inp[11]) ? 4'b0101 : node21252;
															assign node21252 = (inp[10]) ? node21254 : 4'b0100;
																assign node21254 = (inp[12]) ? 4'b0100 : 4'b1100;
													assign node21258 = (inp[12]) ? node21270 : node21259;
														assign node21259 = (inp[10]) ? node21265 : node21260;
															assign node21260 = (inp[14]) ? node21262 : 4'b1101;
																assign node21262 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node21265 = (inp[11]) ? 4'b0001 : node21266;
																assign node21266 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node21270 = (inp[14]) ? node21272 : 4'b1101;
															assign node21272 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node21275 = (inp[13]) ? node21289 : node21276;
													assign node21276 = (inp[10]) ? 4'b1100 : node21277;
														assign node21277 = (inp[12]) ? node21283 : node21278;
															assign node21278 = (inp[14]) ? node21280 : 4'b1100;
																assign node21280 = (inp[11]) ? 4'b1100 : 4'b0101;
															assign node21283 = (inp[14]) ? node21285 : 4'b0100;
																assign node21285 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node21289 = (inp[12]) ? node21295 : node21290;
														assign node21290 = (inp[11]) ? 4'b0000 : node21291;
															assign node21291 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21295 = (inp[10]) ? node21299 : node21296;
															assign node21296 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21299 = (inp[11]) ? 4'b0000 : node21300;
																assign node21300 = (inp[14]) ? 4'b1101 : 4'b0000;
									assign node21304 = (inp[7]) ? node21400 : node21305;
										assign node21305 = (inp[4]) ? node21337 : node21306;
											assign node21306 = (inp[13]) ? node21308 : 4'b0110;
												assign node21308 = (inp[10]) ? node21318 : node21309;
													assign node21309 = (inp[1]) ? node21311 : 4'b0110;
														assign node21311 = (inp[12]) ? 4'b0110 : node21312;
															assign node21312 = (inp[14]) ? node21314 : 4'b0000;
																assign node21314 = (inp[11]) ? 4'b0000 : 4'b0110;
													assign node21318 = (inp[12]) ? node21330 : node21319;
														assign node21319 = (inp[1]) ? node21325 : node21320;
															assign node21320 = (inp[11]) ? 4'b0001 : node21321;
																assign node21321 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21325 = (inp[14]) ? node21327 : 4'b0000;
																assign node21327 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21330 = (inp[1]) ? node21332 : 4'b0110;
															assign node21332 = (inp[11]) ? 4'b0000 : node21333;
																assign node21333 = (inp[14]) ? 4'b0110 : 4'b0000;
											assign node21337 = (inp[1]) ? node21369 : node21338;
												assign node21338 = (inp[13]) ? node21356 : node21339;
													assign node21339 = (inp[10]) ? node21345 : node21340;
														assign node21340 = (inp[14]) ? node21342 : 4'b0001;
															assign node21342 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node21345 = (inp[12]) ? node21351 : node21346;
															assign node21346 = (inp[14]) ? node21348 : 4'b1001;
																assign node21348 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node21351 = (inp[11]) ? 4'b0001 : node21352;
																assign node21352 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node21356 = (inp[14]) ? node21362 : node21357;
														assign node21357 = (inp[10]) ? node21359 : 4'b1001;
															assign node21359 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node21362 = (inp[11]) ? node21364 : 4'b1000;
															assign node21364 = (inp[10]) ? node21366 : 4'b1001;
																assign node21366 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node21369 = (inp[11]) ? node21389 : node21370;
													assign node21370 = (inp[14]) ? node21380 : node21371;
														assign node21371 = (inp[13]) ? node21377 : node21372;
															assign node21372 = (inp[10]) ? 4'b1000 : node21373;
																assign node21373 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node21377 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node21380 = (inp[13]) ? node21384 : node21381;
															assign node21381 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node21384 = (inp[10]) ? node21386 : 4'b1001;
																assign node21386 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node21389 = (inp[13]) ? node21395 : node21390;
														assign node21390 = (inp[10]) ? 4'b1000 : node21391;
															assign node21391 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node21395 = (inp[12]) ? node21397 : 4'b0000;
															assign node21397 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node21400 = (inp[4]) ? node21402 : 4'b0110;
											assign node21402 = (inp[13]) ? node21404 : 4'b0110;
												assign node21404 = (inp[1]) ? node21410 : node21405;
													assign node21405 = (inp[10]) ? node21407 : 4'b0110;
														assign node21407 = (inp[12]) ? 4'b0110 : 4'b0001;
													assign node21410 = (inp[12]) ? node21416 : node21411;
														assign node21411 = (inp[11]) ? 4'b0000 : node21412;
															assign node21412 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21416 = (inp[10]) ? node21418 : 4'b0110;
															assign node21418 = (inp[11]) ? 4'b0000 : 4'b0110;
								assign node21421 = (inp[1]) ? node21531 : node21422;
									assign node21422 = (inp[4]) ? node21464 : node21423;
										assign node21423 = (inp[13]) ? node21441 : node21424;
											assign node21424 = (inp[12]) ? node21436 : node21425;
												assign node21425 = (inp[10]) ? node21431 : node21426;
													assign node21426 = (inp[14]) ? node21428 : 4'b0001;
														assign node21428 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21431 = (inp[14]) ? node21433 : 4'b1001;
														assign node21433 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node21436 = (inp[14]) ? node21438 : 4'b0001;
													assign node21438 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node21441 = (inp[12]) ? node21459 : node21442;
												assign node21442 = (inp[10]) ? node21448 : node21443;
													assign node21443 = (inp[11]) ? 4'b1001 : node21444;
														assign node21444 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node21448 = (inp[7]) ? node21454 : node21449;
														assign node21449 = (inp[11]) ? 4'b0101 : node21450;
															assign node21450 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node21454 = (inp[11]) ? 4'b0001 : node21455;
															assign node21455 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node21459 = (inp[11]) ? 4'b1001 : node21460;
													assign node21460 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node21464 = (inp[7]) ? node21496 : node21465;
											assign node21465 = (inp[13]) ? node21483 : node21466;
												assign node21466 = (inp[14]) ? node21472 : node21467;
													assign node21467 = (inp[10]) ? node21469 : 4'b0101;
														assign node21469 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21472 = (inp[11]) ? node21478 : node21473;
														assign node21473 = (inp[10]) ? node21475 : 4'b0100;
															assign node21475 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node21478 = (inp[12]) ? 4'b0101 : node21479;
															assign node21479 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node21483 = (inp[12]) ? node21491 : node21484;
													assign node21484 = (inp[10]) ? 4'b0101 : node21485;
														assign node21485 = (inp[11]) ? 4'b1101 : node21486;
															assign node21486 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node21491 = (inp[14]) ? node21493 : 4'b1101;
														assign node21493 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node21496 = (inp[13]) ? node21514 : node21497;
												assign node21497 = (inp[10]) ? node21503 : node21498;
													assign node21498 = (inp[14]) ? node21500 : 4'b0001;
														assign node21500 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21503 = (inp[12]) ? node21509 : node21504;
														assign node21504 = (inp[14]) ? node21506 : 4'b1001;
															assign node21506 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node21509 = (inp[11]) ? 4'b0001 : node21510;
															assign node21510 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node21514 = (inp[10]) ? node21520 : node21515;
													assign node21515 = (inp[11]) ? 4'b1001 : node21516;
														assign node21516 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node21520 = (inp[12]) ? node21526 : node21521;
														assign node21521 = (inp[11]) ? 4'b0101 : node21522;
															assign node21522 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node21526 = (inp[11]) ? 4'b1001 : node21527;
															assign node21527 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node21531 = (inp[11]) ? node21601 : node21532;
										assign node21532 = (inp[14]) ? node21566 : node21533;
											assign node21533 = (inp[13]) ? node21551 : node21534;
												assign node21534 = (inp[12]) ? node21540 : node21535;
													assign node21535 = (inp[4]) ? node21537 : 4'b1000;
														assign node21537 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node21540 = (inp[10]) ? node21546 : node21541;
														assign node21541 = (inp[4]) ? node21543 : 4'b0000;
															assign node21543 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21546 = (inp[7]) ? 4'b1000 : node21547;
															assign node21547 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node21551 = (inp[7]) ? node21559 : node21552;
													assign node21552 = (inp[10]) ? 4'b0100 : node21553;
														assign node21553 = (inp[12]) ? node21555 : 4'b0100;
															assign node21555 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node21559 = (inp[4]) ? node21561 : 4'b0000;
														assign node21561 = (inp[12]) ? node21563 : 4'b0100;
															assign node21563 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node21566 = (inp[13]) ? node21584 : node21567;
												assign node21567 = (inp[4]) ? node21573 : node21568;
													assign node21568 = (inp[12]) ? 4'b0001 : node21569;
														assign node21569 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node21573 = (inp[7]) ? node21579 : node21574;
														assign node21574 = (inp[12]) ? 4'b0101 : node21575;
															assign node21575 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node21579 = (inp[12]) ? 4'b0001 : node21580;
															assign node21580 = (inp[10]) ? 4'b1001 : 4'b0001;
												assign node21584 = (inp[10]) ? node21590 : node21585;
													assign node21585 = (inp[4]) ? node21587 : 4'b1001;
														assign node21587 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node21590 = (inp[12]) ? node21596 : node21591;
														assign node21591 = (inp[4]) ? 4'b0101 : node21592;
															assign node21592 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node21596 = (inp[7]) ? 4'b1001 : node21597;
															assign node21597 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node21601 = (inp[13]) ? node21619 : node21602;
											assign node21602 = (inp[10]) ? node21614 : node21603;
												assign node21603 = (inp[12]) ? node21609 : node21604;
													assign node21604 = (inp[7]) ? 4'b1000 : node21605;
														assign node21605 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node21609 = (inp[7]) ? 4'b0000 : node21610;
														assign node21610 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node21614 = (inp[4]) ? node21616 : 4'b1000;
													assign node21616 = (inp[7]) ? 4'b1000 : 4'b1100;
											assign node21619 = (inp[10]) ? node21631 : node21620;
												assign node21620 = (inp[12]) ? node21626 : node21621;
													assign node21621 = (inp[7]) ? node21623 : 4'b0100;
														assign node21623 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node21626 = (inp[4]) ? node21628 : 4'b1000;
														assign node21628 = (inp[7]) ? 4'b1000 : 4'b1100;
												assign node21631 = (inp[7]) ? node21633 : 4'b0100;
													assign node21633 = (inp[4]) ? 4'b0100 : 4'b0000;
					assign node21637 = (inp[5]) ? node22775 : node21638;
						assign node21638 = (inp[0]) ? node22446 : node21639;
							assign node21639 = (inp[11]) ? node22109 : node21640;
								assign node21640 = (inp[3]) ? node21892 : node21641;
									assign node21641 = (inp[4]) ? node21747 : node21642;
										assign node21642 = (inp[13]) ? node21688 : node21643;
											assign node21643 = (inp[12]) ? node21665 : node21644;
												assign node21644 = (inp[10]) ? node21652 : node21645;
													assign node21645 = (inp[1]) ? node21649 : node21646;
														assign node21646 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node21649 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node21652 = (inp[7]) ? node21658 : node21653;
														assign node21653 = (inp[1]) ? 4'b0001 : node21654;
															assign node21654 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node21658 = (inp[14]) ? node21662 : node21659;
															assign node21659 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node21662 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node21665 = (inp[10]) ? node21681 : node21666;
													assign node21666 = (inp[2]) ? node21674 : node21667;
														assign node21667 = (inp[14]) ? node21671 : node21668;
															assign node21668 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node21671 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node21674 = (inp[1]) ? node21678 : node21675;
															assign node21675 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node21678 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node21681 = (inp[1]) ? node21685 : node21682;
														assign node21682 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node21685 = (inp[14]) ? 4'b0101 : 4'b1100;
											assign node21688 = (inp[7]) ? node21720 : node21689;
												assign node21689 = (inp[2]) ? node21701 : node21690;
													assign node21690 = (inp[10]) ? node21696 : node21691;
														assign node21691 = (inp[12]) ? 4'b0001 : node21692;
															assign node21692 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node21696 = (inp[12]) ? 4'b1001 : node21697;
															assign node21697 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node21701 = (inp[14]) ? node21713 : node21702;
														assign node21702 = (inp[1]) ? node21708 : node21703;
															assign node21703 = (inp[10]) ? node21705 : 4'b1101;
																assign node21705 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node21708 = (inp[10]) ? 4'b0000 : node21709;
																assign node21709 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node21713 = (inp[1]) ? 4'b1101 : node21714;
															assign node21714 = (inp[10]) ? node21716 : 4'b1100;
																assign node21716 = (inp[12]) ? 4'b1100 : 4'b0000;
												assign node21720 = (inp[10]) ? node21730 : node21721;
													assign node21721 = (inp[1]) ? node21725 : node21722;
														assign node21722 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node21725 = (inp[14]) ? 4'b1101 : node21726;
															assign node21726 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node21730 = (inp[12]) ? node21740 : node21731;
														assign node21731 = (inp[1]) ? node21735 : node21732;
															assign node21732 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node21735 = (inp[2]) ? node21737 : 4'b0001;
																assign node21737 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node21740 = (inp[1]) ? node21744 : node21741;
															assign node21741 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node21744 = (inp[14]) ? 4'b1101 : 4'b0100;
										assign node21747 = (inp[2]) ? node21783 : node21748;
											assign node21748 = (inp[10]) ? node21766 : node21749;
												assign node21749 = (inp[7]) ? node21761 : node21750;
													assign node21750 = (inp[13]) ? node21756 : node21751;
														assign node21751 = (inp[12]) ? 4'b0001 : node21752;
															assign node21752 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node21756 = (inp[1]) ? node21758 : 4'b0101;
															assign node21758 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21761 = (inp[1]) ? node21763 : 4'b0001;
														assign node21763 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node21766 = (inp[13]) ? node21774 : node21767;
													assign node21767 = (inp[1]) ? node21769 : 4'b1001;
														assign node21769 = (inp[12]) ? 4'b1001 : node21770;
															assign node21770 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node21774 = (inp[12]) ? node21780 : node21775;
														assign node21775 = (inp[1]) ? 4'b0101 : node21776;
															assign node21776 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node21780 = (inp[7]) ? 4'b1001 : 4'b1101;
											assign node21783 = (inp[7]) ? node21835 : node21784;
												assign node21784 = (inp[13]) ? node21808 : node21785;
													assign node21785 = (inp[12]) ? node21801 : node21786;
														assign node21786 = (inp[10]) ? node21794 : node21787;
															assign node21787 = (inp[1]) ? node21791 : node21788;
																assign node21788 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node21791 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node21794 = (inp[1]) ? node21798 : node21795;
																assign node21795 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node21798 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21801 = (inp[1]) ? node21805 : node21802;
															assign node21802 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node21805 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node21808 = (inp[12]) ? node21822 : node21809;
														assign node21809 = (inp[10]) ? node21815 : node21810;
															assign node21810 = (inp[1]) ? 4'b0000 : node21811;
																assign node21811 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21815 = (inp[1]) ? node21819 : node21816;
																assign node21816 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node21819 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node21822 = (inp[10]) ? node21830 : node21823;
															assign node21823 = (inp[1]) ? node21827 : node21824;
																assign node21824 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node21827 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21830 = (inp[14]) ? node21832 : 4'b0000;
																assign node21832 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node21835 = (inp[13]) ? node21861 : node21836;
													assign node21836 = (inp[10]) ? node21846 : node21837;
														assign node21837 = (inp[14]) ? node21843 : node21838;
															assign node21838 = (inp[1]) ? node21840 : 4'b0101;
																assign node21840 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node21843 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node21846 = (inp[12]) ? node21854 : node21847;
															assign node21847 = (inp[1]) ? node21851 : node21848;
																assign node21848 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node21851 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21854 = (inp[1]) ? node21858 : node21855;
																assign node21855 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node21858 = (inp[14]) ? 4'b0101 : 4'b1100;
													assign node21861 = (inp[12]) ? node21877 : node21862;
														assign node21862 = (inp[10]) ? node21870 : node21863;
															assign node21863 = (inp[14]) ? node21867 : node21864;
																assign node21864 = (inp[1]) ? 4'b0000 : 4'b1101;
																assign node21867 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node21870 = (inp[14]) ? node21874 : node21871;
																assign node21871 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node21874 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node21877 = (inp[10]) ? node21885 : node21878;
															assign node21878 = (inp[1]) ? node21882 : node21879;
																assign node21879 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node21882 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node21885 = (inp[14]) ? node21889 : node21886;
																assign node21886 = (inp[1]) ? 4'b0000 : 4'b1101;
																assign node21889 = (inp[1]) ? 4'b1101 : 4'b1100;
									assign node21892 = (inp[2]) ? node22010 : node21893;
										assign node21893 = (inp[4]) ? node21933 : node21894;
											assign node21894 = (inp[10]) ? node21912 : node21895;
												assign node21895 = (inp[13]) ? node21901 : node21896;
													assign node21896 = (inp[1]) ? node21898 : 4'b0101;
														assign node21898 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node21901 = (inp[7]) ? node21907 : node21902;
														assign node21902 = (inp[12]) ? 4'b0001 : node21903;
															assign node21903 = (inp[14]) ? 4'b0001 : 4'b1001;
														assign node21907 = (inp[1]) ? node21909 : 4'b0101;
															assign node21909 = (inp[12]) ? 4'b0101 : 4'b1101;
												assign node21912 = (inp[12]) ? node21928 : node21913;
													assign node21913 = (inp[1]) ? node21919 : node21914;
														assign node21914 = (inp[7]) ? 4'b1101 : node21915;
															assign node21915 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node21919 = (inp[13]) ? node21923 : node21920;
															assign node21920 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node21923 = (inp[14]) ? node21925 : 4'b0001;
																assign node21925 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node21928 = (inp[7]) ? 4'b1101 : node21929;
														assign node21929 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node21933 = (inp[13]) ? node21965 : node21934;
												assign node21934 = (inp[1]) ? node21946 : node21935;
													assign node21935 = (inp[14]) ? node21941 : node21936;
														assign node21936 = (inp[10]) ? 4'b0000 : node21937;
															assign node21937 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node21941 = (inp[10]) ? node21943 : 4'b0001;
															assign node21943 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node21946 = (inp[12]) ? node21954 : node21947;
														assign node21947 = (inp[14]) ? node21949 : 4'b1001;
															assign node21949 = (inp[10]) ? 4'b1000 : node21950;
																assign node21950 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node21954 = (inp[7]) ? node21960 : node21955;
															assign node21955 = (inp[10]) ? 4'b0001 : node21956;
																assign node21956 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21960 = (inp[10]) ? node21962 : 4'b0001;
																assign node21962 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node21965 = (inp[7]) ? node21989 : node21966;
													assign node21966 = (inp[1]) ? node21978 : node21967;
														assign node21967 = (inp[14]) ? node21973 : node21968;
															assign node21968 = (inp[12]) ? 4'b1000 : node21969;
																assign node21969 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node21973 = (inp[12]) ? 4'b0101 : node21974;
																assign node21974 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node21978 = (inp[14]) ? node21984 : node21979;
															assign node21979 = (inp[10]) ? node21981 : 4'b0101;
																assign node21981 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node21984 = (inp[12]) ? node21986 : 4'b0100;
																assign node21986 = (inp[10]) ? 4'b1100 : 4'b0100;
													assign node21989 = (inp[1]) ? node21999 : node21990;
														assign node21990 = (inp[14]) ? node21994 : node21991;
															assign node21991 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node21994 = (inp[10]) ? node21996 : 4'b1001;
																assign node21996 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node21999 = (inp[14]) ? node22005 : node22000;
															assign node22000 = (inp[10]) ? node22002 : 4'b0001;
																assign node22002 = (inp[12]) ? 4'b1001 : 4'b0101;
															assign node22005 = (inp[10]) ? node22007 : 4'b0000;
																assign node22007 = (inp[12]) ? 4'b1000 : 4'b0100;
										assign node22010 = (inp[4]) ? node22072 : node22011;
											assign node22011 = (inp[13]) ? node22037 : node22012;
												assign node22012 = (inp[12]) ? node22028 : node22013;
													assign node22013 = (inp[10]) ? node22021 : node22014;
														assign node22014 = (inp[1]) ? node22018 : node22015;
															assign node22015 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22018 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node22021 = (inp[1]) ? node22025 : node22022;
															assign node22022 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node22025 = (inp[7]) ? 4'b1000 : 4'b0001;
													assign node22028 = (inp[1]) ? node22032 : node22029;
														assign node22029 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node22032 = (inp[14]) ? 4'b0001 : node22033;
															assign node22033 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node22037 = (inp[7]) ? node22049 : node22038;
													assign node22038 = (inp[10]) ? node22044 : node22039;
														assign node22039 = (inp[1]) ? node22041 : 4'b0001;
															assign node22041 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22044 = (inp[12]) ? 4'b1001 : node22045;
															assign node22045 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node22049 = (inp[10]) ? node22059 : node22050;
														assign node22050 = (inp[1]) ? node22054 : node22051;
															assign node22051 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node22054 = (inp[14]) ? 4'b1001 : node22055;
																assign node22055 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22059 = (inp[12]) ? node22065 : node22060;
															assign node22060 = (inp[14]) ? node22062 : 4'b0001;
																assign node22062 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node22065 = (inp[1]) ? node22069 : node22066;
																assign node22066 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node22069 = (inp[14]) ? 4'b1001 : 4'b0000;
											assign node22072 = (inp[7]) ? node22096 : node22073;
												assign node22073 = (inp[13]) ? node22085 : node22074;
													assign node22074 = (inp[10]) ? node22080 : node22075;
														assign node22075 = (inp[12]) ? 4'b0001 : node22076;
															assign node22076 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node22080 = (inp[12]) ? 4'b1001 : node22081;
															assign node22081 = (inp[1]) ? 4'b0101 : 4'b1001;
													assign node22085 = (inp[12]) ? node22093 : node22086;
														assign node22086 = (inp[10]) ? node22090 : node22087;
															assign node22087 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node22090 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node22093 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node22096 = (inp[10]) ? node22102 : node22097;
													assign node22097 = (inp[1]) ? node22099 : 4'b0001;
														assign node22099 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node22102 = (inp[1]) ? node22104 : 4'b1001;
														assign node22104 = (inp[12]) ? 4'b1001 : node22105;
															assign node22105 = (inp[13]) ? 4'b0101 : 4'b0001;
								assign node22109 = (inp[1]) ? node22327 : node22110;
									assign node22110 = (inp[13]) ? node22190 : node22111;
										assign node22111 = (inp[4]) ? node22141 : node22112;
											assign node22112 = (inp[3]) ? node22122 : node22113;
												assign node22113 = (inp[10]) ? node22115 : 4'b0101;
													assign node22115 = (inp[12]) ? 4'b0101 : node22116;
														assign node22116 = (inp[7]) ? 4'b1101 : node22117;
															assign node22117 = (inp[2]) ? 4'b1101 : 4'b0000;
												assign node22122 = (inp[2]) ? node22132 : node22123;
													assign node22123 = (inp[10]) ? node22127 : node22124;
														assign node22124 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node22127 = (inp[12]) ? 4'b1100 : node22128;
															assign node22128 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node22132 = (inp[12]) ? 4'b0001 : node22133;
														assign node22133 = (inp[7]) ? node22137 : node22134;
															assign node22134 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node22137 = (inp[10]) ? 4'b1001 : 4'b0001;
											assign node22141 = (inp[12]) ? node22167 : node22142;
												assign node22142 = (inp[10]) ? node22154 : node22143;
													assign node22143 = (inp[3]) ? node22149 : node22144;
														assign node22144 = (inp[2]) ? node22146 : 4'b1000;
															assign node22146 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node22149 = (inp[2]) ? 4'b1000 : node22150;
															assign node22150 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22154 = (inp[3]) ? node22162 : node22155;
														assign node22155 = (inp[2]) ? node22159 : node22156;
															assign node22156 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node22159 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node22162 = (inp[2]) ? node22164 : 4'b0001;
															assign node22164 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node22167 = (inp[10]) ? node22181 : node22168;
													assign node22168 = (inp[7]) ? node22176 : node22169;
														assign node22169 = (inp[2]) ? node22173 : node22170;
															assign node22170 = (inp[3]) ? 4'b0001 : 4'b0000;
															assign node22173 = (inp[3]) ? 4'b0000 : 4'b0001;
														assign node22176 = (inp[2]) ? node22178 : 4'b0000;
															assign node22178 = (inp[3]) ? 4'b0000 : 4'b0101;
													assign node22181 = (inp[2]) ? node22185 : node22182;
														assign node22182 = (inp[3]) ? 4'b0001 : 4'b1000;
														assign node22185 = (inp[3]) ? 4'b1000 : node22186;
															assign node22186 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node22190 = (inp[3]) ? node22250 : node22191;
											assign node22191 = (inp[2]) ? node22237 : node22192;
												assign node22192 = (inp[4]) ? node22214 : node22193;
													assign node22193 = (inp[7]) ? node22209 : node22194;
														assign node22194 = (inp[14]) ? node22202 : node22195;
															assign node22195 = (inp[10]) ? node22199 : node22196;
																assign node22196 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node22199 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node22202 = (inp[12]) ? node22206 : node22203;
																assign node22203 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node22206 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22209 = (inp[12]) ? 4'b1101 : node22210;
															assign node22210 = (inp[10]) ? 4'b0000 : 4'b1101;
													assign node22214 = (inp[7]) ? node22230 : node22215;
														assign node22215 = (inp[14]) ? node22223 : node22216;
															assign node22216 = (inp[12]) ? node22220 : node22217;
																assign node22217 = (inp[10]) ? 4'b0100 : 4'b1100;
																assign node22220 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node22223 = (inp[12]) ? node22227 : node22224;
																assign node22224 = (inp[10]) ? 4'b0100 : 4'b1100;
																assign node22227 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node22230 = (inp[10]) ? node22234 : node22231;
															assign node22231 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22234 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node22237 = (inp[4]) ? node22239 : 4'b1101;
													assign node22239 = (inp[7]) ? node22245 : node22240;
														assign node22240 = (inp[10]) ? node22242 : 4'b1001;
															assign node22242 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node22245 = (inp[10]) ? node22247 : 4'b1101;
															assign node22247 = (inp[12]) ? 4'b1101 : 4'b0001;
											assign node22250 = (inp[4]) ? node22294 : node22251;
												assign node22251 = (inp[7]) ? node22281 : node22252;
													assign node22252 = (inp[2]) ? node22266 : node22253;
														assign node22253 = (inp[14]) ? node22259 : node22254;
															assign node22254 = (inp[12]) ? 4'b1000 : node22255;
																assign node22255 = (inp[10]) ? 4'b0000 : 4'b1000;
															assign node22259 = (inp[10]) ? node22263 : node22260;
																assign node22260 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node22263 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22266 = (inp[14]) ? node22274 : node22267;
															assign node22267 = (inp[12]) ? node22271 : node22268;
																assign node22268 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node22271 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node22274 = (inp[12]) ? node22278 : node22275;
																assign node22275 = (inp[10]) ? 4'b0000 : 4'b1000;
																assign node22278 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node22281 = (inp[2]) ? node22289 : node22282;
														assign node22282 = (inp[10]) ? node22286 : node22283;
															assign node22283 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node22286 = (inp[12]) ? 4'b1100 : 4'b0000;
														assign node22289 = (inp[10]) ? node22291 : 4'b1001;
															assign node22291 = (inp[12]) ? 4'b1001 : 4'b0000;
												assign node22294 = (inp[2]) ? node22308 : node22295;
													assign node22295 = (inp[7]) ? node22303 : node22296;
														assign node22296 = (inp[12]) ? node22300 : node22297;
															assign node22297 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node22300 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node22303 = (inp[10]) ? 4'b1001 : node22304;
															assign node22304 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node22308 = (inp[7]) ? node22316 : node22309;
														assign node22309 = (inp[10]) ? node22313 : node22310;
															assign node22310 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node22313 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node22316 = (inp[14]) ? node22322 : node22317;
															assign node22317 = (inp[10]) ? 4'b1000 : node22318;
																assign node22318 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22322 = (inp[10]) ? node22324 : 4'b1000;
																assign node22324 = (inp[12]) ? 4'b1000 : 4'b0100;
									assign node22327 = (inp[10]) ? node22405 : node22328;
										assign node22328 = (inp[4]) ? node22364 : node22329;
											assign node22329 = (inp[3]) ? node22349 : node22330;
												assign node22330 = (inp[7]) ? node22342 : node22331;
													assign node22331 = (inp[13]) ? node22335 : node22332;
														assign node22332 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node22335 = (inp[12]) ? node22339 : node22336;
															assign node22336 = (inp[2]) ? 4'b0000 : 4'b1000;
															assign node22339 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node22342 = (inp[12]) ? node22346 : node22343;
														assign node22343 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node22346 = (inp[13]) ? 4'b1100 : 4'b0100;
												assign node22349 = (inp[2]) ? node22355 : node22350;
													assign node22350 = (inp[13]) ? node22352 : 4'b1100;
														assign node22352 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node22355 = (inp[13]) ? node22359 : node22356;
														assign node22356 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22359 = (inp[7]) ? node22361 : 4'b1000;
															assign node22361 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node22364 = (inp[13]) ? node22380 : node22365;
												assign node22365 = (inp[2]) ? node22371 : node22366;
													assign node22366 = (inp[12]) ? 4'b1000 : node22367;
														assign node22367 = (inp[3]) ? 4'b0000 : 4'b1000;
													assign node22371 = (inp[3]) ? 4'b1000 : node22372;
														assign node22372 = (inp[12]) ? node22376 : node22373;
															assign node22373 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node22376 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node22380 = (inp[7]) ? node22392 : node22381;
													assign node22381 = (inp[2]) ? node22387 : node22382;
														assign node22382 = (inp[12]) ? node22384 : 4'b1100;
															assign node22384 = (inp[3]) ? 4'b0100 : 4'b1100;
														assign node22387 = (inp[3]) ? 4'b1100 : node22388;
															assign node22388 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node22392 = (inp[12]) ? node22398 : node22393;
														assign node22393 = (inp[2]) ? node22395 : 4'b1000;
															assign node22395 = (inp[3]) ? 4'b1000 : 4'b0000;
														assign node22398 = (inp[3]) ? node22402 : node22399;
															assign node22399 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node22402 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node22405 = (inp[13]) ? node22433 : node22406;
											assign node22406 = (inp[2]) ? node22420 : node22407;
												assign node22407 = (inp[3]) ? node22415 : node22408;
													assign node22408 = (inp[4]) ? node22412 : node22409;
														assign node22409 = (inp[7]) ? 4'b1100 : 4'b0000;
														assign node22412 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22415 = (inp[4]) ? 4'b1000 : node22416;
														assign node22416 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node22420 = (inp[3]) ? node22426 : node22421;
													assign node22421 = (inp[4]) ? node22423 : 4'b1100;
														assign node22423 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node22426 = (inp[7]) ? node22430 : node22427;
														assign node22427 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node22430 = (inp[4]) ? 4'b0000 : 4'b1000;
											assign node22433 = (inp[4]) ? node22441 : node22434;
												assign node22434 = (inp[7]) ? node22436 : 4'b0000;
													assign node22436 = (inp[3]) ? 4'b0000 : node22437;
														assign node22437 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node22441 = (inp[3]) ? 4'b0100 : node22442;
													assign node22442 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node22446 = (inp[2]) ? 4'b0100 : node22447;
								assign node22447 = (inp[3]) ? node22569 : node22448;
									assign node22448 = (inp[4]) ? node22478 : node22449;
										assign node22449 = (inp[13]) ? node22451 : 4'b0100;
											assign node22451 = (inp[7]) ? 4'b0100 : node22452;
												assign node22452 = (inp[10]) ? node22462 : node22453;
													assign node22453 = (inp[12]) ? 4'b0100 : node22454;
														assign node22454 = (inp[1]) ? node22456 : 4'b0100;
															assign node22456 = (inp[11]) ? 4'b0000 : node22457;
																assign node22457 = (inp[14]) ? 4'b0100 : 4'b0000;
													assign node22462 = (inp[12]) ? node22470 : node22463;
														assign node22463 = (inp[1]) ? 4'b0000 : node22464;
															assign node22464 = (inp[14]) ? node22466 : 4'b0001;
																assign node22466 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node22470 = (inp[1]) ? node22472 : 4'b0100;
															assign node22472 = (inp[11]) ? 4'b0000 : node22473;
																assign node22473 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node22478 = (inp[7]) ? node22540 : node22479;
											assign node22479 = (inp[1]) ? node22511 : node22480;
												assign node22480 = (inp[13]) ? node22498 : node22481;
													assign node22481 = (inp[12]) ? node22493 : node22482;
														assign node22482 = (inp[10]) ? node22488 : node22483;
															assign node22483 = (inp[11]) ? 4'b0001 : node22484;
																assign node22484 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22488 = (inp[14]) ? node22490 : 4'b1001;
																assign node22490 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node22493 = (inp[11]) ? 4'b0001 : node22494;
															assign node22494 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node22498 = (inp[11]) ? node22506 : node22499;
														assign node22499 = (inp[14]) ? 4'b1000 : node22500;
															assign node22500 = (inp[10]) ? node22502 : 4'b1001;
																assign node22502 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node22506 = (inp[10]) ? node22508 : 4'b1001;
															assign node22508 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node22511 = (inp[14]) ? node22523 : node22512;
													assign node22512 = (inp[13]) ? node22518 : node22513;
														assign node22513 = (inp[10]) ? 4'b1000 : node22514;
															assign node22514 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22518 = (inp[10]) ? 4'b0000 : node22519;
															assign node22519 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node22523 = (inp[11]) ? node22533 : node22524;
														assign node22524 = (inp[13]) ? node22530 : node22525;
															assign node22525 = (inp[12]) ? 4'b0001 : node22526;
																assign node22526 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node22530 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node22533 = (inp[13]) ? node22537 : node22534;
															assign node22534 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22537 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node22540 = (inp[13]) ? node22542 : 4'b0100;
												assign node22542 = (inp[12]) ? node22562 : node22543;
													assign node22543 = (inp[10]) ? node22551 : node22544;
														assign node22544 = (inp[1]) ? node22546 : 4'b0100;
															assign node22546 = (inp[14]) ? node22548 : 4'b0000;
																assign node22548 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node22551 = (inp[1]) ? node22557 : node22552;
															assign node22552 = (inp[11]) ? 4'b0001 : node22553;
																assign node22553 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node22557 = (inp[14]) ? node22559 : 4'b0000;
																assign node22559 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node22562 = (inp[1]) ? node22564 : 4'b0100;
														assign node22564 = (inp[10]) ? node22566 : 4'b0100;
															assign node22566 = (inp[11]) ? 4'b0000 : 4'b0100;
									assign node22569 = (inp[7]) ? node22693 : node22570;
										assign node22570 = (inp[4]) ? node22632 : node22571;
											assign node22571 = (inp[1]) ? node22603 : node22572;
												assign node22572 = (inp[14]) ? node22584 : node22573;
													assign node22573 = (inp[13]) ? node22579 : node22574;
														assign node22574 = (inp[10]) ? node22576 : 4'b0001;
															assign node22576 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22579 = (inp[12]) ? 4'b1001 : node22580;
															assign node22580 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node22584 = (inp[11]) ? node22596 : node22585;
														assign node22585 = (inp[13]) ? node22591 : node22586;
															assign node22586 = (inp[10]) ? node22588 : 4'b0000;
																assign node22588 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node22591 = (inp[12]) ? 4'b1000 : node22592;
																assign node22592 = (inp[10]) ? 4'b0100 : 4'b1000;
														assign node22596 = (inp[13]) ? node22600 : node22597;
															assign node22597 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node22600 = (inp[10]) ? 4'b0101 : 4'b1001;
												assign node22603 = (inp[13]) ? node22613 : node22604;
													assign node22604 = (inp[14]) ? node22610 : node22605;
														assign node22605 = (inp[12]) ? node22607 : 4'b1000;
															assign node22607 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22610 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node22613 = (inp[12]) ? node22621 : node22614;
														assign node22614 = (inp[11]) ? 4'b0100 : node22615;
															assign node22615 = (inp[14]) ? node22617 : 4'b0100;
																assign node22617 = (inp[10]) ? 4'b0101 : 4'b1001;
														assign node22621 = (inp[10]) ? node22627 : node22622;
															assign node22622 = (inp[11]) ? 4'b1000 : node22623;
																assign node22623 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node22627 = (inp[14]) ? node22629 : 4'b0100;
																assign node22629 = (inp[11]) ? 4'b0100 : 4'b1001;
											assign node22632 = (inp[1]) ? node22660 : node22633;
												assign node22633 = (inp[11]) ? node22649 : node22634;
													assign node22634 = (inp[14]) ? node22642 : node22635;
														assign node22635 = (inp[13]) ? node22637 : 4'b0101;
															assign node22637 = (inp[12]) ? 4'b1101 : node22638;
																assign node22638 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node22642 = (inp[13]) ? node22644 : 4'b0100;
															assign node22644 = (inp[12]) ? 4'b1100 : node22645;
																assign node22645 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node22649 = (inp[13]) ? node22655 : node22650;
														assign node22650 = (inp[12]) ? 4'b0101 : node22651;
															assign node22651 = (inp[10]) ? 4'b1101 : 4'b0101;
														assign node22655 = (inp[12]) ? 4'b1101 : node22656;
															assign node22656 = (inp[10]) ? 4'b0101 : 4'b1101;
												assign node22660 = (inp[14]) ? node22672 : node22661;
													assign node22661 = (inp[13]) ? node22667 : node22662;
														assign node22662 = (inp[12]) ? node22664 : 4'b1100;
															assign node22664 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node22667 = (inp[10]) ? 4'b0100 : node22668;
															assign node22668 = (inp[12]) ? 4'b1100 : 4'b0100;
													assign node22672 = (inp[11]) ? node22684 : node22673;
														assign node22673 = (inp[13]) ? node22679 : node22674;
															assign node22674 = (inp[12]) ? 4'b0101 : node22675;
																assign node22675 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node22679 = (inp[12]) ? 4'b1101 : node22680;
																assign node22680 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node22684 = (inp[13]) ? node22688 : node22685;
															assign node22685 = (inp[10]) ? 4'b1100 : 4'b0100;
															assign node22688 = (inp[10]) ? 4'b0100 : node22689;
																assign node22689 = (inp[12]) ? 4'b1100 : 4'b0100;
										assign node22693 = (inp[1]) ? node22729 : node22694;
											assign node22694 = (inp[11]) ? node22716 : node22695;
												assign node22695 = (inp[14]) ? node22705 : node22696;
													assign node22696 = (inp[13]) ? node22700 : node22697;
														assign node22697 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node22700 = (inp[12]) ? 4'b1001 : node22701;
															assign node22701 = (inp[10]) ? 4'b0101 : 4'b1001;
													assign node22705 = (inp[13]) ? node22711 : node22706;
														assign node22706 = (inp[12]) ? 4'b0000 : node22707;
															assign node22707 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22711 = (inp[10]) ? node22713 : 4'b1000;
															assign node22713 = (inp[12]) ? 4'b1000 : 4'b0100;
												assign node22716 = (inp[13]) ? node22722 : node22717;
													assign node22717 = (inp[12]) ? 4'b0001 : node22718;
														assign node22718 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node22722 = (inp[10]) ? node22724 : 4'b1001;
														assign node22724 = (inp[12]) ? 4'b1001 : node22725;
															assign node22725 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node22729 = (inp[11]) ? node22757 : node22730;
												assign node22730 = (inp[14]) ? node22744 : node22731;
													assign node22731 = (inp[13]) ? node22737 : node22732;
														assign node22732 = (inp[12]) ? node22734 : 4'b1000;
															assign node22734 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node22737 = (inp[10]) ? node22741 : node22738;
															assign node22738 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node22741 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node22744 = (inp[13]) ? node22750 : node22745;
														assign node22745 = (inp[12]) ? 4'b0001 : node22746;
															assign node22746 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node22750 = (inp[12]) ? 4'b1001 : node22751;
															assign node22751 = (inp[10]) ? node22753 : 4'b1001;
																assign node22753 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node22757 = (inp[13]) ? node22763 : node22758;
													assign node22758 = (inp[10]) ? 4'b1000 : node22759;
														assign node22759 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node22763 = (inp[4]) ? node22769 : node22764;
														assign node22764 = (inp[10]) ? 4'b0000 : node22765;
															assign node22765 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node22769 = (inp[10]) ? 4'b0100 : node22770;
															assign node22770 = (inp[12]) ? 4'b1000 : 4'b0100;
						assign node22775 = (inp[3]) ? node23553 : node22776;
							assign node22776 = (inp[4]) ? node23140 : node22777;
								assign node22777 = (inp[0]) ? node22993 : node22778;
									assign node22778 = (inp[13]) ? node22900 : node22779;
										assign node22779 = (inp[7]) ? node22843 : node22780;
											assign node22780 = (inp[10]) ? node22816 : node22781;
												assign node22781 = (inp[1]) ? node22801 : node22782;
													assign node22782 = (inp[12]) ? node22790 : node22783;
														assign node22783 = (inp[11]) ? node22787 : node22784;
															assign node22784 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node22787 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node22790 = (inp[14]) ? node22796 : node22791;
															assign node22791 = (inp[11]) ? node22793 : 4'b0100;
																assign node22793 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node22796 = (inp[11]) ? node22798 : 4'b0101;
																assign node22798 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node22801 = (inp[11]) ? node22811 : node22802;
														assign node22802 = (inp[2]) ? node22808 : node22803;
															assign node22803 = (inp[12]) ? node22805 : 4'b0000;
																assign node22805 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node22808 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node22811 = (inp[12]) ? node22813 : 4'b0000;
															assign node22813 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node22816 = (inp[2]) ? node22828 : node22817;
													assign node22817 = (inp[1]) ? node22823 : node22818;
														assign node22818 = (inp[12]) ? node22820 : 4'b1000;
															assign node22820 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node22823 = (inp[12]) ? node22825 : 4'b0000;
															assign node22825 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node22828 = (inp[1]) ? node22836 : node22829;
														assign node22829 = (inp[11]) ? 4'b0001 : node22830;
															assign node22830 = (inp[14]) ? node22832 : 4'b0000;
																assign node22832 = (inp[12]) ? 4'b1101 : 4'b0001;
														assign node22836 = (inp[11]) ? 4'b1000 : node22837;
															assign node22837 = (inp[12]) ? node22839 : 4'b1001;
																assign node22839 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node22843 = (inp[11]) ? node22877 : node22844;
												assign node22844 = (inp[2]) ? node22866 : node22845;
													assign node22845 = (inp[10]) ? node22855 : node22846;
														assign node22846 = (inp[1]) ? node22852 : node22847;
															assign node22847 = (inp[12]) ? node22849 : 4'b1100;
																assign node22849 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node22852 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node22855 = (inp[1]) ? node22861 : node22856;
															assign node22856 = (inp[14]) ? node22858 : 4'b0100;
																assign node22858 = (inp[12]) ? 4'b1101 : 4'b0101;
															assign node22861 = (inp[12]) ? node22863 : 4'b0000;
																assign node22863 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node22866 = (inp[10]) ? node22872 : node22867;
														assign node22867 = (inp[1]) ? node22869 : 4'b0101;
															assign node22869 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node22872 = (inp[1]) ? node22874 : 4'b1101;
															assign node22874 = (inp[12]) ? 4'b1101 : 4'b0101;
												assign node22877 = (inp[10]) ? node22891 : node22878;
													assign node22878 = (inp[1]) ? node22886 : node22879;
														assign node22879 = (inp[2]) ? node22883 : node22880;
															assign node22880 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node22883 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node22886 = (inp[12]) ? 4'b1100 : node22887;
															assign node22887 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node22891 = (inp[1]) ? node22897 : node22892;
														assign node22892 = (inp[2]) ? node22894 : 4'b0101;
															assign node22894 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node22897 = (inp[2]) ? 4'b0100 : 4'b0000;
										assign node22900 = (inp[2]) ? node22942 : node22901;
											assign node22901 = (inp[1]) ? node22919 : node22902;
												assign node22902 = (inp[12]) ? node22908 : node22903;
													assign node22903 = (inp[10]) ? node22905 : 4'b1000;
														assign node22905 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node22908 = (inp[11]) ? node22914 : node22909;
														assign node22909 = (inp[7]) ? 4'b0000 : node22910;
															assign node22910 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node22914 = (inp[7]) ? 4'b1000 : node22915;
															assign node22915 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node22919 = (inp[11]) ? node22935 : node22920;
													assign node22920 = (inp[12]) ? node22930 : node22921;
														assign node22921 = (inp[14]) ? node22927 : node22922;
															assign node22922 = (inp[10]) ? 4'b0000 : node22923;
																assign node22923 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node22927 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node22930 = (inp[7]) ? 4'b1000 : node22931;
															assign node22931 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node22935 = (inp[10]) ? node22939 : node22936;
														assign node22936 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node22939 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node22942 = (inp[1]) ? node22970 : node22943;
												assign node22943 = (inp[10]) ? node22963 : node22944;
													assign node22944 = (inp[7]) ? node22954 : node22945;
														assign node22945 = (inp[12]) ? node22951 : node22946;
															assign node22946 = (inp[11]) ? 4'b0001 : node22947;
																assign node22947 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node22951 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node22954 = (inp[12]) ? node22960 : node22955;
															assign node22955 = (inp[11]) ? 4'b0001 : node22956;
																assign node22956 = (inp[14]) ? 4'b0101 : 4'b0000;
															assign node22960 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node22963 = (inp[11]) ? 4'b1001 : node22964;
														assign node22964 = (inp[14]) ? node22966 : 4'b1000;
															assign node22966 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node22970 = (inp[11]) ? node22986 : node22971;
													assign node22971 = (inp[14]) ? node22981 : node22972;
														assign node22972 = (inp[12]) ? node22978 : node22973;
															assign node22973 = (inp[7]) ? 4'b0001 : node22974;
																assign node22974 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node22978 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node22981 = (inp[10]) ? node22983 : 4'b0000;
															assign node22983 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node22986 = (inp[10]) ? node22990 : node22987;
														assign node22987 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node22990 = (inp[7]) ? 4'b0000 : 4'b0100;
									assign node22993 = (inp[2]) ? node23109 : node22994;
										assign node22994 = (inp[13]) ? node23050 : node22995;
											assign node22995 = (inp[1]) ? node23019 : node22996;
												assign node22996 = (inp[10]) ? node23002 : node22997;
													assign node22997 = (inp[14]) ? node22999 : 4'b0101;
														assign node22999 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23002 = (inp[12]) ? node23014 : node23003;
														assign node23003 = (inp[7]) ? node23009 : node23004;
															assign node23004 = (inp[11]) ? 4'b0000 : node23005;
																assign node23005 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node23009 = (inp[14]) ? node23011 : 4'b1101;
																assign node23011 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node23014 = (inp[14]) ? node23016 : 4'b0101;
															assign node23016 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node23019 = (inp[11]) ? node23039 : node23020;
													assign node23020 = (inp[14]) ? node23028 : node23021;
														assign node23021 = (inp[10]) ? node23025 : node23022;
															assign node23022 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node23025 = (inp[12]) ? 4'b1100 : 4'b0001;
														assign node23028 = (inp[7]) ? node23034 : node23029;
															assign node23029 = (inp[12]) ? 4'b0101 : node23030;
																assign node23030 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node23034 = (inp[12]) ? 4'b0101 : node23035;
																assign node23035 = (inp[10]) ? 4'b1101 : 4'b0101;
													assign node23039 = (inp[7]) ? node23045 : node23040;
														assign node23040 = (inp[10]) ? 4'b0000 : node23041;
															assign node23041 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node23045 = (inp[12]) ? node23047 : 4'b1100;
															assign node23047 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node23050 = (inp[7]) ? node23074 : node23051;
												assign node23051 = (inp[11]) ? node23063 : node23052;
													assign node23052 = (inp[10]) ? node23058 : node23053;
														assign node23053 = (inp[12]) ? 4'b0001 : node23054;
															assign node23054 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node23058 = (inp[12]) ? 4'b1001 : node23059;
															assign node23059 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node23063 = (inp[10]) ? node23069 : node23064;
														assign node23064 = (inp[12]) ? node23066 : 4'b1000;
															assign node23066 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node23069 = (inp[1]) ? 4'b0000 : node23070;
															assign node23070 = (inp[12]) ? 4'b1000 : 4'b0000;
												assign node23074 = (inp[10]) ? node23092 : node23075;
													assign node23075 = (inp[1]) ? node23081 : node23076;
														assign node23076 = (inp[11]) ? 4'b1101 : node23077;
															assign node23077 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node23081 = (inp[12]) ? node23087 : node23082;
															assign node23082 = (inp[14]) ? node23084 : 4'b0100;
																assign node23084 = (inp[11]) ? 4'b0100 : 4'b1101;
															assign node23087 = (inp[14]) ? node23089 : 4'b1100;
																assign node23089 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node23092 = (inp[12]) ? node23098 : node23093;
														assign node23093 = (inp[11]) ? 4'b0000 : node23094;
															assign node23094 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node23098 = (inp[14]) ? node23104 : node23099;
															assign node23099 = (inp[1]) ? node23101 : 4'b1101;
																assign node23101 = (inp[11]) ? 4'b0000 : 4'b0100;
															assign node23104 = (inp[11]) ? 4'b1101 : node23105;
																assign node23105 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node23109 = (inp[7]) ? 4'b0100 : node23110;
											assign node23110 = (inp[13]) ? node23112 : 4'b0100;
												assign node23112 = (inp[12]) ? node23132 : node23113;
													assign node23113 = (inp[10]) ? node23121 : node23114;
														assign node23114 = (inp[1]) ? node23116 : 4'b0100;
															assign node23116 = (inp[14]) ? node23118 : 4'b0000;
																assign node23118 = (inp[11]) ? 4'b0000 : 4'b0100;
														assign node23121 = (inp[1]) ? node23127 : node23122;
															assign node23122 = (inp[14]) ? node23124 : 4'b0001;
																assign node23124 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23127 = (inp[11]) ? 4'b0000 : node23128;
																assign node23128 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node23132 = (inp[1]) ? node23134 : 4'b0100;
														assign node23134 = (inp[10]) ? node23136 : 4'b0100;
															assign node23136 = (inp[14]) ? 4'b0100 : 4'b0000;
								assign node23140 = (inp[11]) ? node23410 : node23141;
									assign node23141 = (inp[2]) ? node23257 : node23142;
										assign node23142 = (inp[10]) ? node23202 : node23143;
											assign node23143 = (inp[0]) ? node23177 : node23144;
												assign node23144 = (inp[7]) ? node23156 : node23145;
													assign node23145 = (inp[12]) ? node23149 : node23146;
														assign node23146 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node23149 = (inp[13]) ? 4'b0001 : node23150;
															assign node23150 = (inp[1]) ? node23152 : 4'b0000;
																assign node23152 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node23156 = (inp[1]) ? node23168 : node23157;
														assign node23157 = (inp[13]) ? node23161 : node23158;
															assign node23158 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node23161 = (inp[12]) ? node23165 : node23162;
																assign node23162 = (inp[14]) ? 4'b0100 : 4'b0101;
																assign node23165 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node23168 = (inp[13]) ? 4'b0001 : node23169;
															assign node23169 = (inp[12]) ? node23173 : node23170;
																assign node23170 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node23173 = (inp[14]) ? 4'b1100 : 4'b0000;
												assign node23177 = (inp[1]) ? node23187 : node23178;
													assign node23178 = (inp[7]) ? 4'b0001 : node23179;
														assign node23179 = (inp[13]) ? node23181 : 4'b0001;
															assign node23181 = (inp[12]) ? 4'b0101 : node23182;
																assign node23182 = (inp[14]) ? 4'b0101 : 4'b0000;
													assign node23187 = (inp[12]) ? node23195 : node23188;
														assign node23188 = (inp[7]) ? 4'b1001 : node23189;
															assign node23189 = (inp[13]) ? node23191 : 4'b1001;
																assign node23191 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23195 = (inp[7]) ? 4'b0001 : node23196;
															assign node23196 = (inp[14]) ? node23198 : 4'b0001;
																assign node23198 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node23202 = (inp[1]) ? node23226 : node23203;
												assign node23203 = (inp[13]) ? node23209 : node23204;
													assign node23204 = (inp[0]) ? 4'b1001 : node23205;
														assign node23205 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node23209 = (inp[0]) ? node23217 : node23210;
														assign node23210 = (inp[12]) ? 4'b1001 : node23211;
															assign node23211 = (inp[7]) ? 4'b0001 : node23212;
																assign node23212 = (inp[14]) ? 4'b0101 : 4'b0000;
														assign node23217 = (inp[14]) ? node23221 : node23218;
															assign node23218 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node23221 = (inp[7]) ? 4'b1001 : node23222;
																assign node23222 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node23226 = (inp[13]) ? node23244 : node23227;
													assign node23227 = (inp[7]) ? node23237 : node23228;
														assign node23228 = (inp[0]) ? node23234 : node23229;
															assign node23229 = (inp[14]) ? 4'b0101 : node23230;
																assign node23230 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node23234 = (inp[12]) ? 4'b1001 : 4'b0101;
														assign node23237 = (inp[0]) ? node23241 : node23238;
															assign node23238 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node23241 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node23244 = (inp[12]) ? node23252 : node23245;
														assign node23245 = (inp[0]) ? node23249 : node23246;
															assign node23246 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node23249 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23252 = (inp[14]) ? node23254 : 4'b1001;
															assign node23254 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node23257 = (inp[7]) ? node23355 : node23258;
											assign node23258 = (inp[0]) ? node23302 : node23259;
												assign node23259 = (inp[10]) ? node23279 : node23260;
													assign node23260 = (inp[13]) ? node23272 : node23261;
														assign node23261 = (inp[1]) ? node23267 : node23262;
															assign node23262 = (inp[14]) ? 4'b0101 : node23263;
																assign node23263 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node23267 = (inp[12]) ? node23269 : 4'b0000;
																assign node23269 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node23272 = (inp[1]) ? node23276 : node23273;
															assign node23273 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23276 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node23279 = (inp[13]) ? node23295 : node23280;
														assign node23280 = (inp[14]) ? node23288 : node23281;
															assign node23281 = (inp[1]) ? node23285 : node23282;
																assign node23282 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node23285 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node23288 = (inp[1]) ? node23292 : node23289;
																assign node23289 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node23292 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node23295 = (inp[14]) ? 4'b1001 : node23296;
															assign node23296 = (inp[12]) ? 4'b1000 : node23297;
																assign node23297 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node23302 = (inp[13]) ? node23326 : node23303;
													assign node23303 = (inp[10]) ? node23313 : node23304;
														assign node23304 = (inp[14]) ? node23310 : node23305;
															assign node23305 = (inp[1]) ? node23307 : 4'b0001;
																assign node23307 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23310 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node23313 = (inp[12]) ? node23321 : node23314;
															assign node23314 = (inp[14]) ? node23318 : node23315;
																assign node23315 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node23318 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node23321 = (inp[1]) ? node23323 : 4'b0001;
																assign node23323 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node23326 = (inp[10]) ? node23340 : node23327;
														assign node23327 = (inp[12]) ? node23333 : node23328;
															assign node23328 = (inp[1]) ? 4'b1001 : node23329;
																assign node23329 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23333 = (inp[1]) ? node23337 : node23334;
																assign node23334 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node23337 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node23340 = (inp[12]) ? node23348 : node23341;
															assign node23341 = (inp[14]) ? node23345 : node23342;
																assign node23342 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node23345 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node23348 = (inp[1]) ? node23352 : node23349;
																assign node23349 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node23352 = (inp[14]) ? 4'b1001 : 4'b0000;
											assign node23355 = (inp[0]) ? node23393 : node23356;
												assign node23356 = (inp[13]) ? node23380 : node23357;
													assign node23357 = (inp[10]) ? node23367 : node23358;
														assign node23358 = (inp[1]) ? node23364 : node23359;
															assign node23359 = (inp[14]) ? 4'b0001 : node23360;
																assign node23360 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23364 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node23367 = (inp[14]) ? node23373 : node23368;
															assign node23368 = (inp[1]) ? node23370 : 4'b0100;
																assign node23370 = (inp[12]) ? 4'b0101 : 4'b0000;
															assign node23373 = (inp[1]) ? node23377 : node23374;
																assign node23374 = (inp[12]) ? 4'b1001 : 4'b0101;
																assign node23377 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node23380 = (inp[10]) ? node23386 : node23381;
														assign node23381 = (inp[1]) ? 4'b0000 : node23382;
															assign node23382 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23386 = (inp[12]) ? node23390 : node23387;
															assign node23387 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node23390 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node23393 = (inp[10]) ? node23395 : 4'b0100;
													assign node23395 = (inp[13]) ? node23397 : 4'b0100;
														assign node23397 = (inp[12]) ? node23405 : node23398;
															assign node23398 = (inp[14]) ? node23402 : node23399;
																assign node23399 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node23402 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node23405 = (inp[14]) ? 4'b0100 : node23406;
																assign node23406 = (inp[1]) ? 4'b0000 : 4'b0100;
									assign node23410 = (inp[1]) ? node23498 : node23411;
										assign node23411 = (inp[7]) ? node23461 : node23412;
											assign node23412 = (inp[13]) ? node23438 : node23413;
												assign node23413 = (inp[0]) ? node23425 : node23414;
													assign node23414 = (inp[10]) ? node23420 : node23415;
														assign node23415 = (inp[2]) ? node23417 : 4'b1001;
															assign node23417 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node23420 = (inp[2]) ? 4'b1000 : node23421;
															assign node23421 = (inp[12]) ? 4'b1001 : 4'b0101;
													assign node23425 = (inp[2]) ? node23433 : node23426;
														assign node23426 = (inp[10]) ? node23430 : node23427;
															assign node23427 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23430 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node23433 = (inp[10]) ? node23435 : 4'b0001;
															assign node23435 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node23438 = (inp[10]) ? node23450 : node23439;
													assign node23439 = (inp[0]) ? node23445 : node23440;
														assign node23440 = (inp[12]) ? 4'b1000 : node23441;
															assign node23441 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node23445 = (inp[2]) ? 4'b1001 : node23446;
															assign node23446 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node23450 = (inp[0]) ? node23456 : node23451;
														assign node23451 = (inp[12]) ? 4'b0001 : node23452;
															assign node23452 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node23456 = (inp[2]) ? node23458 : 4'b1001;
															assign node23458 = (inp[12]) ? 4'b1001 : 4'b0001;
											assign node23461 = (inp[0]) ? node23481 : node23462;
												assign node23462 = (inp[13]) ? node23472 : node23463;
													assign node23463 = (inp[2]) ? node23467 : node23464;
														assign node23464 = (inp[10]) ? 4'b0001 : 4'b1100;
														assign node23467 = (inp[10]) ? 4'b0101 : node23468;
															assign node23468 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node23472 = (inp[2]) ? 4'b1000 : node23473;
														assign node23473 = (inp[12]) ? node23477 : node23474;
															assign node23474 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node23477 = (inp[10]) ? 4'b0000 : 4'b0101;
												assign node23481 = (inp[2]) ? node23491 : node23482;
													assign node23482 = (inp[12]) ? node23488 : node23483;
														assign node23483 = (inp[10]) ? node23485 : 4'b1000;
															assign node23485 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node23488 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node23491 = (inp[13]) ? node23493 : 4'b0100;
														assign node23493 = (inp[12]) ? 4'b0100 : node23494;
															assign node23494 = (inp[10]) ? 4'b0001 : 4'b0100;
										assign node23498 = (inp[10]) ? node23538 : node23499;
											assign node23499 = (inp[2]) ? node23511 : node23500;
												assign node23500 = (inp[12]) ? node23502 : 4'b1000;
													assign node23502 = (inp[7]) ? node23506 : node23503;
														assign node23503 = (inp[14]) ? 4'b0000 : 4'b1000;
														assign node23506 = (inp[13]) ? 4'b1000 : node23507;
															assign node23507 = (inp[0]) ? 4'b1000 : 4'b0000;
												assign node23511 = (inp[7]) ? node23525 : node23512;
													assign node23512 = (inp[0]) ? node23518 : node23513;
														assign node23513 = (inp[12]) ? node23515 : 4'b0000;
															assign node23515 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node23518 = (inp[13]) ? node23522 : node23519;
															assign node23519 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23522 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node23525 = (inp[0]) ? node23533 : node23526;
														assign node23526 = (inp[12]) ? node23530 : node23527;
															assign node23527 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node23530 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node23533 = (inp[13]) ? node23535 : 4'b0100;
															assign node23535 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node23538 = (inp[13]) ? 4'b0000 : node23539;
												assign node23539 = (inp[0]) ? node23545 : node23540;
													assign node23540 = (inp[7]) ? node23542 : 4'b0000;
														assign node23542 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node23545 = (inp[2]) ? node23549 : node23546;
														assign node23546 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node23549 = (inp[7]) ? 4'b0100 : 4'b1000;
							assign node23553 = (inp[4]) ? node24033 : node23554;
								assign node23554 = (inp[11]) ? node23858 : node23555;
									assign node23555 = (inp[2]) ? node23705 : node23556;
										assign node23556 = (inp[13]) ? node23640 : node23557;
											assign node23557 = (inp[10]) ? node23607 : node23558;
												assign node23558 = (inp[12]) ? node23586 : node23559;
													assign node23559 = (inp[0]) ? node23573 : node23560;
														assign node23560 = (inp[7]) ? node23566 : node23561;
															assign node23561 = (inp[1]) ? 4'b1000 : node23562;
																assign node23562 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node23566 = (inp[14]) ? node23570 : node23567;
																assign node23567 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node23570 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node23573 = (inp[7]) ? node23581 : node23574;
															assign node23574 = (inp[14]) ? node23578 : node23575;
																assign node23575 = (inp[1]) ? 4'b0000 : 4'b1000;
																assign node23578 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node23581 = (inp[1]) ? node23583 : 4'b1000;
																assign node23583 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node23586 = (inp[7]) ? node23594 : node23587;
														assign node23587 = (inp[0]) ? node23589 : 4'b1000;
															assign node23589 = (inp[1]) ? node23591 : 4'b0001;
																assign node23591 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node23594 = (inp[0]) ? node23602 : node23595;
															assign node23595 = (inp[1]) ? node23599 : node23596;
																assign node23596 = (inp[14]) ? 4'b0001 : 4'b1000;
																assign node23599 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node23602 = (inp[1]) ? 4'b1000 : node23603;
																assign node23603 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node23607 = (inp[1]) ? node23625 : node23608;
													assign node23608 = (inp[0]) ? node23614 : node23609;
														assign node23609 = (inp[12]) ? 4'b1000 : node23610;
															assign node23610 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node23614 = (inp[14]) ? node23620 : node23615;
															assign node23615 = (inp[12]) ? 4'b0000 : node23616;
																assign node23616 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node23620 = (inp[7]) ? 4'b1001 : node23621;
																assign node23621 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23625 = (inp[14]) ? node23631 : node23626;
														assign node23626 = (inp[12]) ? node23628 : 4'b0000;
															assign node23628 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23631 = (inp[0]) ? node23637 : node23632;
															assign node23632 = (inp[12]) ? node23634 : 4'b0001;
																assign node23634 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node23637 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node23640 = (inp[1]) ? node23668 : node23641;
												assign node23641 = (inp[10]) ? node23657 : node23642;
													assign node23642 = (inp[0]) ? node23648 : node23643;
														assign node23643 = (inp[7]) ? node23645 : 4'b1001;
															assign node23645 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23648 = (inp[7]) ? node23654 : node23649;
															assign node23649 = (inp[14]) ? 4'b0000 : node23650;
																assign node23650 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node23654 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23657 = (inp[0]) ? node23663 : node23658;
														assign node23658 = (inp[12]) ? node23660 : 4'b0000;
															assign node23660 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node23663 = (inp[14]) ? node23665 : 4'b0001;
															assign node23665 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node23668 = (inp[0]) ? node23684 : node23669;
													assign node23669 = (inp[10]) ? node23677 : node23670;
														assign node23670 = (inp[7]) ? node23674 : node23671;
															assign node23671 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23674 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node23677 = (inp[14]) ? 4'b0001 : node23678;
															assign node23678 = (inp[7]) ? node23680 : 4'b0001;
																assign node23680 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23684 = (inp[7]) ? node23694 : node23685;
														assign node23685 = (inp[14]) ? node23689 : node23686;
															assign node23686 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node23689 = (inp[10]) ? 4'b1001 : node23690;
																assign node23690 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23694 = (inp[12]) ? node23700 : node23695;
															assign node23695 = (inp[10]) ? node23697 : 4'b0000;
																assign node23697 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node23700 = (inp[10]) ? node23702 : 4'b1000;
																assign node23702 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node23705 = (inp[13]) ? node23783 : node23706;
											assign node23706 = (inp[10]) ? node23738 : node23707;
												assign node23707 = (inp[12]) ? node23723 : node23708;
													assign node23708 = (inp[1]) ? node23716 : node23709;
														assign node23709 = (inp[0]) ? node23713 : node23710;
															assign node23710 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23713 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23716 = (inp[14]) ? 4'b0001 : node23717;
															assign node23717 = (inp[0]) ? 4'b1000 : node23718;
																assign node23718 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node23723 = (inp[1]) ? node23727 : node23724;
														assign node23724 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node23727 = (inp[14]) ? node23733 : node23728;
															assign node23728 = (inp[7]) ? 4'b0000 : node23729;
																assign node23729 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node23733 = (inp[0]) ? 4'b0001 : node23734;
																assign node23734 = (inp[7]) ? 4'b1001 : 4'b0001;
												assign node23738 = (inp[7]) ? node23764 : node23739;
													assign node23739 = (inp[14]) ? node23753 : node23740;
														assign node23740 = (inp[1]) ? node23748 : node23741;
															assign node23741 = (inp[0]) ? node23745 : node23742;
																assign node23742 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node23745 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node23748 = (inp[12]) ? node23750 : 4'b0001;
																assign node23750 = (inp[0]) ? 4'b1000 : 4'b0001;
														assign node23753 = (inp[1]) ? node23761 : node23754;
															assign node23754 = (inp[0]) ? node23758 : node23755;
																assign node23755 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node23758 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node23761 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node23764 = (inp[0]) ? node23770 : node23765;
														assign node23765 = (inp[12]) ? 4'b1001 : node23766;
															assign node23766 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node23770 = (inp[12]) ? node23778 : node23771;
															assign node23771 = (inp[1]) ? node23775 : node23772;
																assign node23772 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node23775 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node23778 = (inp[14]) ? node23780 : 4'b1000;
																assign node23780 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node23783 = (inp[0]) ? node23821 : node23784;
												assign node23784 = (inp[10]) ? node23802 : node23785;
													assign node23785 = (inp[1]) ? node23793 : node23786;
														assign node23786 = (inp[14]) ? node23788 : 4'b0000;
															assign node23788 = (inp[12]) ? node23790 : 4'b0001;
																assign node23790 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node23793 = (inp[7]) ? node23795 : 4'b1000;
															assign node23795 = (inp[12]) ? node23799 : node23796;
																assign node23796 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node23799 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node23802 = (inp[12]) ? node23814 : node23803;
														assign node23803 = (inp[1]) ? node23809 : node23804;
															assign node23804 = (inp[7]) ? 4'b1000 : node23805;
																assign node23805 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node23809 = (inp[14]) ? 4'b1001 : node23810;
																assign node23810 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node23814 = (inp[1]) ? 4'b0001 : node23815;
															assign node23815 = (inp[7]) ? 4'b1000 : node23816;
																assign node23816 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node23821 = (inp[7]) ? node23835 : node23822;
													assign node23822 = (inp[10]) ? node23828 : node23823;
														assign node23823 = (inp[12]) ? 4'b0001 : node23824;
															assign node23824 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node23828 = (inp[12]) ? 4'b1001 : node23829;
															assign node23829 = (inp[1]) ? node23831 : 4'b1001;
																assign node23831 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node23835 = (inp[10]) ? node23845 : node23836;
														assign node23836 = (inp[14]) ? node23842 : node23837;
															assign node23837 = (inp[1]) ? node23839 : 4'b1001;
																assign node23839 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node23842 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node23845 = (inp[12]) ? node23851 : node23846;
															assign node23846 = (inp[14]) ? node23848 : 4'b0001;
																assign node23848 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node23851 = (inp[14]) ? node23855 : node23852;
																assign node23852 = (inp[1]) ? 4'b0000 : 4'b1001;
																assign node23855 = (inp[1]) ? 4'b1001 : 4'b1000;
									assign node23858 = (inp[1]) ? node23972 : node23859;
										assign node23859 = (inp[7]) ? node23911 : node23860;
											assign node23860 = (inp[10]) ? node23886 : node23861;
												assign node23861 = (inp[0]) ? node23873 : node23862;
													assign node23862 = (inp[13]) ? node23868 : node23863;
														assign node23863 = (inp[2]) ? node23865 : 4'b0000;
															assign node23865 = (inp[12]) ? 4'b1001 : 4'b0000;
														assign node23868 = (inp[12]) ? 4'b0000 : node23869;
															assign node23869 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node23873 = (inp[12]) ? node23881 : node23874;
														assign node23874 = (inp[13]) ? node23878 : node23875;
															assign node23875 = (inp[2]) ? 4'b0001 : 4'b1001;
															assign node23878 = (inp[2]) ? 4'b1000 : 4'b0001;
														assign node23881 = (inp[13]) ? node23883 : 4'b0001;
															assign node23883 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node23886 = (inp[0]) ? node23898 : node23887;
													assign node23887 = (inp[2]) ? node23891 : node23888;
														assign node23888 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23891 = (inp[12]) ? node23895 : node23892;
															assign node23892 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node23895 = (inp[13]) ? 4'b1001 : 4'b0000;
													assign node23898 = (inp[2]) ? node23904 : node23899;
														assign node23899 = (inp[13]) ? node23901 : 4'b1000;
															assign node23901 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node23904 = (inp[13]) ? node23908 : node23905;
															assign node23905 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node23908 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node23911 = (inp[10]) ? node23947 : node23912;
												assign node23912 = (inp[2]) ? node23928 : node23913;
													assign node23913 = (inp[13]) ? node23923 : node23914;
														assign node23914 = (inp[14]) ? node23916 : 4'b1001;
															assign node23916 = (inp[0]) ? node23920 : node23917;
																assign node23917 = (inp[12]) ? 4'b1001 : 4'b0001;
																assign node23920 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node23923 = (inp[0]) ? 4'b1000 : node23924;
															assign node23924 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node23928 = (inp[14]) ? node23936 : node23929;
														assign node23929 = (inp[0]) ? node23933 : node23930;
															assign node23930 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node23933 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node23936 = (inp[12]) ? node23942 : node23937;
															assign node23937 = (inp[13]) ? 4'b1001 : node23938;
																assign node23938 = (inp[0]) ? 4'b0001 : 4'b1001;
															assign node23942 = (inp[0]) ? 4'b1001 : node23943;
																assign node23943 = (inp[13]) ? 4'b0001 : 4'b1001;
												assign node23947 = (inp[0]) ? node23959 : node23948;
													assign node23948 = (inp[13]) ? node23954 : node23949;
														assign node23949 = (inp[12]) ? 4'b0000 : node23950;
															assign node23950 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node23954 = (inp[2]) ? node23956 : 4'b1000;
															assign node23956 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node23959 = (inp[12]) ? node23967 : node23960;
														assign node23960 = (inp[2]) ? node23964 : node23961;
															assign node23961 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node23964 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node23967 = (inp[2]) ? node23969 : 4'b0001;
															assign node23969 = (inp[13]) ? 4'b1001 : 4'b0001;
										assign node23972 = (inp[10]) ? node24010 : node23973;
											assign node23973 = (inp[2]) ? node23993 : node23974;
												assign node23974 = (inp[7]) ? node23982 : node23975;
													assign node23975 = (inp[12]) ? node23977 : 4'b0000;
														assign node23977 = (inp[0]) ? node23979 : 4'b0000;
															assign node23979 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node23982 = (inp[12]) ? node23988 : node23983;
														assign node23983 = (inp[0]) ? 4'b0000 : node23984;
															assign node23984 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node23988 = (inp[0]) ? node23990 : 4'b0000;
															assign node23990 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node23993 = (inp[0]) ? node24001 : node23994;
													assign node23994 = (inp[13]) ? 4'b0000 : node23995;
														assign node23995 = (inp[7]) ? node23997 : 4'b1000;
															assign node23997 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node24001 = (inp[13]) ? node24005 : node24002;
														assign node24002 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node24005 = (inp[12]) ? 4'b1000 : node24006;
															assign node24006 = (inp[7]) ? 4'b0000 : 4'b1000;
											assign node24010 = (inp[13]) ? 4'b0000 : node24011;
												assign node24011 = (inp[0]) ? node24027 : node24012;
													assign node24012 = (inp[12]) ? node24020 : node24013;
														assign node24013 = (inp[2]) ? node24017 : node24014;
															assign node24014 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node24017 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node24020 = (inp[2]) ? node24024 : node24021;
															assign node24021 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node24024 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node24027 = (inp[7]) ? node24029 : 4'b0000;
														assign node24029 = (inp[2]) ? 4'b1000 : 4'b0000;
								assign node24033 = (inp[13]) ? node24285 : node24034;
									assign node24034 = (inp[10]) ? node24180 : node24035;
										assign node24035 = (inp[11]) ? node24113 : node24036;
											assign node24036 = (inp[14]) ? node24078 : node24037;
												assign node24037 = (inp[7]) ? node24063 : node24038;
													assign node24038 = (inp[1]) ? node24050 : node24039;
														assign node24039 = (inp[0]) ? node24045 : node24040;
															assign node24040 = (inp[2]) ? node24042 : 4'b0000;
																assign node24042 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node24045 = (inp[12]) ? node24047 : 4'b1000;
																assign node24047 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node24050 = (inp[2]) ? node24058 : node24051;
															assign node24051 = (inp[0]) ? node24055 : node24052;
																assign node24052 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node24055 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node24058 = (inp[0]) ? node24060 : 4'b1000;
																assign node24060 = (inp[12]) ? 4'b1001 : 4'b0000;
													assign node24063 = (inp[0]) ? node24071 : node24064;
														assign node24064 = (inp[12]) ? node24068 : node24065;
															assign node24065 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node24068 = (inp[1]) ? 4'b0000 : 4'b1001;
														assign node24071 = (inp[12]) ? 4'b0001 : node24072;
															assign node24072 = (inp[1]) ? 4'b1001 : node24073;
																assign node24073 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node24078 = (inp[1]) ? node24094 : node24079;
													assign node24079 = (inp[7]) ? node24083 : node24080;
														assign node24080 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node24083 = (inp[0]) ? node24089 : node24084;
															assign node24084 = (inp[12]) ? 4'b1001 : node24085;
																assign node24085 = (inp[2]) ? 4'b1001 : 4'b0001;
															assign node24089 = (inp[12]) ? 4'b0001 : node24090;
																assign node24090 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node24094 = (inp[0]) ? node24108 : node24095;
														assign node24095 = (inp[12]) ? node24103 : node24096;
															assign node24096 = (inp[2]) ? node24100 : node24097;
																assign node24097 = (inp[7]) ? 4'b0001 : 4'b1001;
																assign node24100 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node24103 = (inp[2]) ? node24105 : 4'b0001;
																assign node24105 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24108 = (inp[2]) ? node24110 : 4'b1000;
															assign node24110 = (inp[7]) ? 4'b0001 : 4'b1000;
											assign node24113 = (inp[1]) ? node24155 : node24114;
												assign node24114 = (inp[2]) ? node24136 : node24115;
													assign node24115 = (inp[12]) ? node24129 : node24116;
														assign node24116 = (inp[14]) ? node24124 : node24117;
															assign node24117 = (inp[7]) ? node24121 : node24118;
																assign node24118 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node24121 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node24124 = (inp[0]) ? 4'b0001 : node24125;
																assign node24125 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24129 = (inp[7]) ? node24133 : node24130;
															assign node24130 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node24133 = (inp[0]) ? 4'b1000 : 4'b0000;
													assign node24136 = (inp[12]) ? node24148 : node24137;
														assign node24137 = (inp[14]) ? node24143 : node24138;
															assign node24138 = (inp[0]) ? 4'b1000 : node24139;
																assign node24139 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node24143 = (inp[7]) ? node24145 : 4'b1001;
																assign node24145 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node24148 = (inp[0]) ? node24152 : node24149;
															assign node24149 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node24152 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node24155 = (inp[0]) ? node24169 : node24156;
													assign node24156 = (inp[2]) ? node24162 : node24157;
														assign node24157 = (inp[7]) ? node24159 : 4'b0000;
															assign node24159 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node24162 = (inp[12]) ? node24166 : node24163;
															assign node24163 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node24166 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node24169 = (inp[2]) ? node24175 : node24170;
														assign node24170 = (inp[7]) ? 4'b0000 : node24171;
															assign node24171 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node24175 = (inp[7]) ? node24177 : 4'b0000;
															assign node24177 = (inp[12]) ? 4'b1000 : 4'b0000;
										assign node24180 = (inp[1]) ? node24244 : node24181;
											assign node24181 = (inp[0]) ? node24215 : node24182;
												assign node24182 = (inp[2]) ? node24194 : node24183;
													assign node24183 = (inp[7]) ? node24191 : node24184;
														assign node24184 = (inp[11]) ? 4'b0000 : node24185;
															assign node24185 = (inp[12]) ? node24187 : 4'b0001;
																assign node24187 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node24191 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node24194 = (inp[12]) ? node24202 : node24195;
														assign node24195 = (inp[7]) ? node24197 : 4'b0000;
															assign node24197 = (inp[11]) ? 4'b0000 : node24198;
																assign node24198 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node24202 = (inp[14]) ? node24210 : node24203;
															assign node24203 = (inp[7]) ? node24207 : node24204;
																assign node24204 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node24207 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node24210 = (inp[11]) ? node24212 : 4'b0000;
																assign node24212 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node24215 = (inp[11]) ? node24233 : node24216;
													assign node24216 = (inp[2]) ? node24224 : node24217;
														assign node24217 = (inp[7]) ? node24219 : 4'b0001;
															assign node24219 = (inp[12]) ? 4'b1000 : node24220;
																assign node24220 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24224 = (inp[7]) ? node24228 : node24225;
															assign node24225 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node24228 = (inp[14]) ? node24230 : 4'b0000;
																assign node24230 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node24233 = (inp[2]) ? node24239 : node24234;
														assign node24234 = (inp[12]) ? 4'b0001 : node24235;
															assign node24235 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24239 = (inp[7]) ? 4'b0001 : node24240;
															assign node24240 = (inp[12]) ? 4'b1000 : 4'b0001;
											assign node24244 = (inp[11]) ? 4'b0000 : node24245;
												assign node24245 = (inp[7]) ? node24265 : node24246;
													assign node24246 = (inp[12]) ? node24254 : node24247;
														assign node24247 = (inp[0]) ? node24249 : 4'b0000;
															assign node24249 = (inp[2]) ? 4'b1000 : node24250;
																assign node24250 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node24254 = (inp[0]) ? node24260 : node24255;
															assign node24255 = (inp[2]) ? node24257 : 4'b0001;
																assign node24257 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node24260 = (inp[2]) ? node24262 : 4'b0000;
																assign node24262 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node24265 = (inp[14]) ? node24277 : node24266;
														assign node24266 = (inp[0]) ? node24272 : node24267;
															assign node24267 = (inp[2]) ? node24269 : 4'b0000;
																assign node24269 = (inp[12]) ? 4'b1000 : 4'b0001;
															assign node24272 = (inp[2]) ? node24274 : 4'b0001;
																assign node24274 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node24277 = (inp[0]) ? node24279 : 4'b0001;
															assign node24279 = (inp[12]) ? node24281 : 4'b0000;
																assign node24281 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node24285 = (inp[11]) ? node24391 : node24286;
										assign node24286 = (inp[10]) ? node24344 : node24287;
											assign node24287 = (inp[0]) ? node24317 : node24288;
												assign node24288 = (inp[1]) ? node24304 : node24289;
													assign node24289 = (inp[7]) ? node24299 : node24290;
														assign node24290 = (inp[12]) ? 4'b0001 : node24291;
															assign node24291 = (inp[14]) ? node24295 : node24292;
																assign node24292 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node24295 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node24299 = (inp[2]) ? node24301 : 4'b0000;
															assign node24301 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node24304 = (inp[2]) ? node24310 : node24305;
														assign node24305 = (inp[7]) ? node24307 : 4'b0000;
															assign node24307 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node24310 = (inp[12]) ? node24312 : 4'b0000;
															assign node24312 = (inp[14]) ? 4'b0000 : node24313;
																assign node24313 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node24317 = (inp[1]) ? node24331 : node24318;
													assign node24318 = (inp[7]) ? node24324 : node24319;
														assign node24319 = (inp[14]) ? node24321 : 4'b0000;
															assign node24321 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node24324 = (inp[12]) ? node24326 : 4'b0001;
															assign node24326 = (inp[14]) ? 4'b0000 : node24327;
																assign node24327 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node24331 = (inp[12]) ? node24339 : node24332;
														assign node24332 = (inp[14]) ? 4'b0000 : node24333;
															assign node24333 = (inp[2]) ? 4'b0001 : node24334;
																assign node24334 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24339 = (inp[7]) ? 4'b0001 : node24340;
															assign node24340 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node24344 = (inp[1]) ? 4'b0000 : node24345;
												assign node24345 = (inp[14]) ? node24371 : node24346;
													assign node24346 = (inp[2]) ? node24360 : node24347;
														assign node24347 = (inp[0]) ? node24353 : node24348;
															assign node24348 = (inp[12]) ? 4'b0000 : node24349;
																assign node24349 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node24353 = (inp[12]) ? node24357 : node24354;
																assign node24354 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node24357 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24360 = (inp[0]) ? node24366 : node24361;
															assign node24361 = (inp[7]) ? node24363 : 4'b0000;
																assign node24363 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node24366 = (inp[7]) ? 4'b0000 : node24367;
																assign node24367 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node24371 = (inp[2]) ? node24379 : node24372;
														assign node24372 = (inp[7]) ? 4'b0000 : node24373;
															assign node24373 = (inp[0]) ? node24375 : 4'b0000;
																assign node24375 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node24379 = (inp[12]) ? node24385 : node24380;
															assign node24380 = (inp[0]) ? 4'b0000 : node24381;
																assign node24381 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node24385 = (inp[7]) ? node24387 : 4'b0001;
																assign node24387 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node24391 = (inp[1]) ? 4'b0000 : node24392;
											assign node24392 = (inp[10]) ? 4'b0000 : node24393;
												assign node24393 = (inp[12]) ? node24413 : node24394;
													assign node24394 = (inp[14]) ? node24406 : node24395;
														assign node24395 = (inp[2]) ? node24401 : node24396;
															assign node24396 = (inp[0]) ? node24398 : 4'b0000;
																assign node24398 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node24401 = (inp[7]) ? node24403 : 4'b0000;
																assign node24403 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node24406 = (inp[7]) ? 4'b0000 : node24407;
															assign node24407 = (inp[2]) ? 4'b0000 : node24408;
																assign node24408 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node24413 = (inp[2]) ? node24419 : node24414;
														assign node24414 = (inp[0]) ? 4'b0000 : node24415;
															assign node24415 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node24419 = (inp[7]) ? node24423 : node24420;
															assign node24420 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node24423 = (inp[0]) ? 4'b0001 : 4'b0000;
				assign node24428 = (inp[0]) ? node26654 : node24429;
					assign node24429 = (inp[6]) ? node25077 : node24430;
						assign node24430 = (inp[2]) ? node24948 : node24431;
							assign node24431 = (inp[5]) ? node24553 : node24432;
								assign node24432 = (inp[3]) ? node24434 : 4'b0010;
									assign node24434 = (inp[7]) ? node24520 : node24435;
										assign node24435 = (inp[4]) ? node24465 : node24436;
											assign node24436 = (inp[13]) ? node24438 : 4'b0010;
												assign node24438 = (inp[12]) ? node24456 : node24439;
													assign node24439 = (inp[10]) ? node24447 : node24440;
														assign node24440 = (inp[11]) ? 4'b0000 : node24441;
															assign node24441 = (inp[14]) ? 4'b0010 : node24442;
																assign node24442 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node24447 = (inp[1]) ? node24451 : node24448;
															assign node24448 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24451 = (inp[11]) ? 4'b0000 : node24452;
																assign node24452 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node24456 = (inp[1]) ? node24458 : 4'b0010;
														assign node24458 = (inp[10]) ? node24460 : 4'b0010;
															assign node24460 = (inp[14]) ? node24462 : 4'b0000;
																assign node24462 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node24465 = (inp[1]) ? node24489 : node24466;
												assign node24466 = (inp[13]) ? node24480 : node24467;
													assign node24467 = (inp[10]) ? node24473 : node24468;
														assign node24468 = (inp[11]) ? 4'b0001 : node24469;
															assign node24469 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24473 = (inp[12]) ? 4'b0001 : node24474;
															assign node24474 = (inp[14]) ? node24476 : 4'b1001;
																assign node24476 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node24480 = (inp[12]) ? node24484 : node24481;
														assign node24481 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node24484 = (inp[11]) ? 4'b1001 : node24485;
															assign node24485 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node24489 = (inp[11]) ? node24509 : node24490;
													assign node24490 = (inp[14]) ? node24498 : node24491;
														assign node24491 = (inp[12]) ? node24493 : 4'b1000;
															assign node24493 = (inp[13]) ? 4'b0000 : node24494;
																assign node24494 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node24498 = (inp[13]) ? node24504 : node24499;
															assign node24499 = (inp[10]) ? node24501 : 4'b0001;
																assign node24501 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node24504 = (inp[10]) ? node24506 : 4'b1001;
																assign node24506 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node24509 = (inp[13]) ? node24515 : node24510;
														assign node24510 = (inp[10]) ? 4'b1000 : node24511;
															assign node24511 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node24515 = (inp[12]) ? node24517 : 4'b0000;
															assign node24517 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node24520 = (inp[13]) ? node24522 : 4'b0010;
											assign node24522 = (inp[4]) ? node24524 : 4'b0010;
												assign node24524 = (inp[10]) ? node24534 : node24525;
													assign node24525 = (inp[12]) ? 4'b0010 : node24526;
														assign node24526 = (inp[1]) ? node24528 : 4'b0010;
															assign node24528 = (inp[11]) ? 4'b0000 : node24529;
																assign node24529 = (inp[14]) ? 4'b0010 : 4'b0000;
													assign node24534 = (inp[12]) ? node24546 : node24535;
														assign node24535 = (inp[1]) ? node24541 : node24536;
															assign node24536 = (inp[14]) ? node24538 : 4'b0001;
																assign node24538 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node24541 = (inp[11]) ? 4'b0000 : node24542;
																assign node24542 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node24546 = (inp[1]) ? node24548 : 4'b0010;
															assign node24548 = (inp[14]) ? node24550 : 4'b0000;
																assign node24550 = (inp[11]) ? 4'b0000 : 4'b0010;
								assign node24553 = (inp[1]) ? node24747 : node24554;
									assign node24554 = (inp[13]) ? node24642 : node24555;
										assign node24555 = (inp[3]) ? node24597 : node24556;
											assign node24556 = (inp[4]) ? node24570 : node24557;
												assign node24557 = (inp[10]) ? node24563 : node24558;
													assign node24558 = (inp[14]) ? node24560 : 4'b0001;
														assign node24560 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node24563 = (inp[12]) ? 4'b0001 : node24564;
														assign node24564 = (inp[14]) ? node24566 : 4'b1001;
															assign node24566 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node24570 = (inp[7]) ? node24584 : node24571;
													assign node24571 = (inp[11]) ? node24579 : node24572;
														assign node24572 = (inp[14]) ? 4'b0100 : node24573;
															assign node24573 = (inp[10]) ? node24575 : 4'b0101;
																assign node24575 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node24579 = (inp[10]) ? node24581 : 4'b0101;
															assign node24581 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node24584 = (inp[12]) ? node24592 : node24585;
														assign node24585 = (inp[10]) ? node24587 : 4'b0001;
															assign node24587 = (inp[14]) ? node24589 : 4'b1001;
																assign node24589 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node24592 = (inp[11]) ? 4'b0001 : node24593;
															assign node24593 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node24597 = (inp[10]) ? node24615 : node24598;
												assign node24598 = (inp[4]) ? node24604 : node24599;
													assign node24599 = (inp[11]) ? 4'b0101 : node24600;
														assign node24600 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node24604 = (inp[7]) ? node24610 : node24605;
														assign node24605 = (inp[11]) ? 4'b0001 : node24606;
															assign node24606 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24610 = (inp[11]) ? 4'b0101 : node24611;
															assign node24611 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node24615 = (inp[12]) ? node24629 : node24616;
													assign node24616 = (inp[14]) ? node24622 : node24617;
														assign node24617 = (inp[4]) ? node24619 : 4'b1101;
															assign node24619 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node24622 = (inp[11]) ? node24624 : 4'b1100;
															assign node24624 = (inp[4]) ? node24626 : 4'b1101;
																assign node24626 = (inp[7]) ? 4'b1101 : 4'b1001;
													assign node24629 = (inp[11]) ? node24637 : node24630;
														assign node24630 = (inp[14]) ? node24632 : 4'b0101;
															assign node24632 = (inp[4]) ? node24634 : 4'b0100;
																assign node24634 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node24637 = (inp[4]) ? node24639 : 4'b0101;
															assign node24639 = (inp[7]) ? 4'b0101 : 4'b0001;
										assign node24642 = (inp[14]) ? node24678 : node24643;
											assign node24643 = (inp[12]) ? node24667 : node24644;
												assign node24644 = (inp[10]) ? node24656 : node24645;
													assign node24645 = (inp[3]) ? node24651 : node24646;
														assign node24646 = (inp[7]) ? 4'b1001 : node24647;
															assign node24647 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node24651 = (inp[7]) ? 4'b1101 : node24652;
															assign node24652 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node24656 = (inp[3]) ? node24662 : node24657;
														assign node24657 = (inp[4]) ? 4'b0101 : node24658;
															assign node24658 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node24662 = (inp[7]) ? node24664 : 4'b0001;
															assign node24664 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node24667 = (inp[3]) ? node24673 : node24668;
													assign node24668 = (inp[4]) ? node24670 : 4'b1001;
														assign node24670 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node24673 = (inp[4]) ? node24675 : 4'b1101;
														assign node24675 = (inp[7]) ? 4'b1101 : 4'b1001;
											assign node24678 = (inp[11]) ? node24712 : node24679;
												assign node24679 = (inp[10]) ? node24691 : node24680;
													assign node24680 = (inp[3]) ? node24686 : node24681;
														assign node24681 = (inp[4]) ? node24683 : 4'b1000;
															assign node24683 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node24686 = (inp[7]) ? 4'b1100 : node24687;
															assign node24687 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node24691 = (inp[12]) ? node24703 : node24692;
														assign node24692 = (inp[3]) ? node24698 : node24693;
															assign node24693 = (inp[4]) ? 4'b0100 : node24694;
																assign node24694 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node24698 = (inp[7]) ? node24700 : 4'b0000;
																assign node24700 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node24703 = (inp[3]) ? node24709 : node24704;
															assign node24704 = (inp[4]) ? node24706 : 4'b1000;
																assign node24706 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node24709 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node24712 = (inp[12]) ? node24736 : node24713;
													assign node24713 = (inp[10]) ? node24725 : node24714;
														assign node24714 = (inp[3]) ? node24720 : node24715;
															assign node24715 = (inp[7]) ? 4'b1001 : node24716;
																assign node24716 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node24720 = (inp[4]) ? node24722 : 4'b1101;
																assign node24722 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node24725 = (inp[3]) ? node24731 : node24726;
															assign node24726 = (inp[4]) ? 4'b0101 : node24727;
																assign node24727 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node24731 = (inp[4]) ? 4'b0001 : node24732;
																assign node24732 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node24736 = (inp[3]) ? node24742 : node24737;
														assign node24737 = (inp[7]) ? 4'b1001 : node24738;
															assign node24738 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node24742 = (inp[4]) ? node24744 : 4'b1101;
															assign node24744 = (inp[7]) ? 4'b1101 : 4'b1001;
									assign node24747 = (inp[11]) ? node24877 : node24748;
										assign node24748 = (inp[14]) ? node24806 : node24749;
											assign node24749 = (inp[13]) ? node24779 : node24750;
												assign node24750 = (inp[10]) ? node24768 : node24751;
													assign node24751 = (inp[12]) ? node24759 : node24752;
														assign node24752 = (inp[3]) ? 4'b1100 : node24753;
															assign node24753 = (inp[7]) ? 4'b1000 : node24754;
																assign node24754 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node24759 = (inp[3]) ? node24765 : node24760;
															assign node24760 = (inp[4]) ? node24762 : 4'b0000;
																assign node24762 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node24765 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node24768 = (inp[3]) ? node24774 : node24769;
														assign node24769 = (inp[4]) ? node24771 : 4'b1000;
															assign node24771 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node24774 = (inp[4]) ? node24776 : 4'b1100;
															assign node24776 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node24779 = (inp[10]) ? node24795 : node24780;
													assign node24780 = (inp[12]) ? node24788 : node24781;
														assign node24781 = (inp[3]) ? 4'b0000 : node24782;
															assign node24782 = (inp[4]) ? 4'b0100 : node24783;
																assign node24783 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node24788 = (inp[3]) ? node24790 : 4'b1000;
															assign node24790 = (inp[7]) ? 4'b1100 : node24791;
																assign node24791 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node24795 = (inp[3]) ? node24801 : node24796;
														assign node24796 = (inp[4]) ? 4'b0100 : node24797;
															assign node24797 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node24801 = (inp[4]) ? 4'b0000 : node24802;
															assign node24802 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node24806 = (inp[13]) ? node24842 : node24807;
												assign node24807 = (inp[12]) ? node24831 : node24808;
													assign node24808 = (inp[10]) ? node24820 : node24809;
														assign node24809 = (inp[3]) ? node24815 : node24810;
															assign node24810 = (inp[7]) ? 4'b0001 : node24811;
																assign node24811 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node24815 = (inp[7]) ? 4'b0101 : node24816;
																assign node24816 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node24820 = (inp[3]) ? node24826 : node24821;
															assign node24821 = (inp[7]) ? 4'b1001 : node24822;
																assign node24822 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node24826 = (inp[7]) ? 4'b1101 : node24827;
																assign node24827 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node24831 = (inp[3]) ? node24837 : node24832;
														assign node24832 = (inp[4]) ? node24834 : 4'b0001;
															assign node24834 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node24837 = (inp[7]) ? 4'b0101 : node24838;
															assign node24838 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node24842 = (inp[12]) ? node24866 : node24843;
													assign node24843 = (inp[10]) ? node24855 : node24844;
														assign node24844 = (inp[3]) ? node24850 : node24845;
															assign node24845 = (inp[4]) ? node24847 : 4'b1001;
																assign node24847 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node24850 = (inp[4]) ? node24852 : 4'b1101;
																assign node24852 = (inp[7]) ? 4'b1101 : 4'b1001;
														assign node24855 = (inp[3]) ? node24861 : node24856;
															assign node24856 = (inp[4]) ? 4'b0101 : node24857;
																assign node24857 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node24861 = (inp[4]) ? 4'b0001 : node24862;
																assign node24862 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node24866 = (inp[3]) ? node24872 : node24867;
														assign node24867 = (inp[4]) ? node24869 : 4'b1001;
															assign node24869 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node24872 = (inp[7]) ? 4'b1101 : node24873;
															assign node24873 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node24877 = (inp[13]) ? node24913 : node24878;
											assign node24878 = (inp[3]) ? node24896 : node24879;
												assign node24879 = (inp[10]) ? node24891 : node24880;
													assign node24880 = (inp[12]) ? node24886 : node24881;
														assign node24881 = (inp[7]) ? 4'b1000 : node24882;
															assign node24882 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node24886 = (inp[4]) ? node24888 : 4'b0000;
															assign node24888 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node24891 = (inp[7]) ? 4'b1000 : node24892;
														assign node24892 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node24896 = (inp[7]) ? node24908 : node24897;
													assign node24897 = (inp[4]) ? node24903 : node24898;
														assign node24898 = (inp[10]) ? 4'b1100 : node24899;
															assign node24899 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node24903 = (inp[12]) ? node24905 : 4'b1000;
															assign node24905 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node24908 = (inp[12]) ? node24910 : 4'b1100;
														assign node24910 = (inp[10]) ? 4'b1100 : 4'b0100;
											assign node24913 = (inp[12]) ? node24925 : node24914;
												assign node24914 = (inp[3]) ? node24920 : node24915;
													assign node24915 = (inp[7]) ? node24917 : 4'b0100;
														assign node24917 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node24920 = (inp[7]) ? node24922 : 4'b0000;
														assign node24922 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node24925 = (inp[10]) ? node24937 : node24926;
													assign node24926 = (inp[3]) ? node24932 : node24927;
														assign node24927 = (inp[7]) ? 4'b1000 : node24928;
															assign node24928 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node24932 = (inp[4]) ? node24934 : 4'b1100;
															assign node24934 = (inp[7]) ? 4'b1100 : 4'b1000;
													assign node24937 = (inp[3]) ? node24943 : node24938;
														assign node24938 = (inp[4]) ? 4'b0100 : node24939;
															assign node24939 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node24943 = (inp[7]) ? node24945 : 4'b0000;
															assign node24945 = (inp[4]) ? 4'b0000 : 4'b0100;
							assign node24948 = (inp[3]) ? node24950 : 4'b0010;
								assign node24950 = (inp[5]) ? node24952 : 4'b0010;
									assign node24952 = (inp[4]) ? node24978 : node24953;
										assign node24953 = (inp[7]) ? 4'b0010 : node24954;
											assign node24954 = (inp[13]) ? node24956 : 4'b0010;
												assign node24956 = (inp[10]) ? node24964 : node24957;
													assign node24957 = (inp[1]) ? node24959 : 4'b0010;
														assign node24959 = (inp[11]) ? node24961 : 4'b0010;
															assign node24961 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node24964 = (inp[12]) ? node24970 : node24965;
														assign node24965 = (inp[1]) ? 4'b0000 : node24966;
															assign node24966 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node24970 = (inp[1]) ? node24972 : 4'b0010;
															assign node24972 = (inp[14]) ? node24974 : 4'b0000;
																assign node24974 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node24978 = (inp[7]) ? node25046 : node24979;
											assign node24979 = (inp[1]) ? node25015 : node24980;
												assign node24980 = (inp[11]) ? node25004 : node24981;
													assign node24981 = (inp[14]) ? node24993 : node24982;
														assign node24982 = (inp[13]) ? node24988 : node24983;
															assign node24983 = (inp[10]) ? node24985 : 4'b0001;
																assign node24985 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node24988 = (inp[12]) ? 4'b1001 : node24989;
																assign node24989 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node24993 = (inp[13]) ? node24999 : node24994;
															assign node24994 = (inp[12]) ? 4'b0000 : node24995;
																assign node24995 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node24999 = (inp[12]) ? 4'b1000 : node25000;
																assign node25000 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node25004 = (inp[13]) ? node25010 : node25005;
														assign node25005 = (inp[10]) ? node25007 : 4'b0001;
															assign node25007 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node25010 = (inp[12]) ? 4'b1001 : node25011;
															assign node25011 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node25015 = (inp[11]) ? node25035 : node25016;
													assign node25016 = (inp[14]) ? node25028 : node25017;
														assign node25017 = (inp[13]) ? node25023 : node25018;
															assign node25018 = (inp[12]) ? node25020 : 4'b1000;
																assign node25020 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node25023 = (inp[10]) ? 4'b0000 : node25024;
																assign node25024 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node25028 = (inp[13]) ? node25030 : 4'b0001;
															assign node25030 = (inp[12]) ? 4'b1001 : node25031;
																assign node25031 = (inp[10]) ? 4'b0001 : 4'b1001;
													assign node25035 = (inp[13]) ? node25041 : node25036;
														assign node25036 = (inp[10]) ? 4'b1000 : node25037;
															assign node25037 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node25041 = (inp[10]) ? 4'b0000 : node25042;
															assign node25042 = (inp[12]) ? 4'b1000 : 4'b0000;
											assign node25046 = (inp[13]) ? node25048 : 4'b0010;
												assign node25048 = (inp[10]) ? node25058 : node25049;
													assign node25049 = (inp[12]) ? 4'b0010 : node25050;
														assign node25050 = (inp[1]) ? node25052 : 4'b0010;
															assign node25052 = (inp[11]) ? 4'b0000 : node25053;
																assign node25053 = (inp[14]) ? 4'b0010 : 4'b0000;
													assign node25058 = (inp[12]) ? node25070 : node25059;
														assign node25059 = (inp[1]) ? node25065 : node25060;
															assign node25060 = (inp[14]) ? node25062 : 4'b0001;
																assign node25062 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node25065 = (inp[14]) ? node25067 : 4'b0000;
																assign node25067 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node25070 = (inp[1]) ? node25072 : 4'b0010;
															assign node25072 = (inp[11]) ? 4'b0000 : node25073;
																assign node25073 = (inp[14]) ? 4'b0010 : 4'b0000;
						assign node25077 = (inp[5]) ? node25819 : node25078;
							assign node25078 = (inp[1]) ? node25428 : node25079;
								assign node25079 = (inp[3]) ? node25237 : node25080;
									assign node25080 = (inp[14]) ? node25142 : node25081;
										assign node25081 = (inp[13]) ? node25103 : node25082;
											assign node25082 = (inp[12]) ? node25098 : node25083;
												assign node25083 = (inp[10]) ? node25089 : node25084;
													assign node25084 = (inp[7]) ? 4'b0001 : node25085;
														assign node25085 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node25089 = (inp[4]) ? node25091 : 4'b1001;
														assign node25091 = (inp[7]) ? 4'b1001 : node25092;
															assign node25092 = (inp[11]) ? node25094 : 4'b1101;
																assign node25094 = (inp[2]) ? 4'b1101 : 4'b0000;
												assign node25098 = (inp[7]) ? 4'b0001 : node25099;
													assign node25099 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node25103 = (inp[12]) ? node25127 : node25104;
												assign node25104 = (inp[10]) ? node25112 : node25105;
													assign node25105 = (inp[7]) ? 4'b1001 : node25106;
														assign node25106 = (inp[4]) ? node25108 : 4'b1001;
															assign node25108 = (inp[2]) ? 4'b1101 : 4'b0001;
													assign node25112 = (inp[7]) ? node25120 : node25113;
														assign node25113 = (inp[4]) ? node25115 : 4'b0101;
															assign node25115 = (inp[2]) ? 4'b0101 : node25116;
																assign node25116 = (inp[11]) ? 4'b0000 : 4'b1001;
														assign node25120 = (inp[4]) ? node25122 : 4'b0001;
															assign node25122 = (inp[2]) ? 4'b0101 : node25123;
																assign node25123 = (inp[11]) ? 4'b0000 : 4'b0101;
												assign node25127 = (inp[7]) ? 4'b1001 : node25128;
													assign node25128 = (inp[2]) ? node25138 : node25129;
														assign node25129 = (inp[10]) ? node25135 : node25130;
															assign node25130 = (inp[4]) ? node25132 : 4'b1001;
																assign node25132 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node25135 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node25138 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node25142 = (inp[11]) ? node25184 : node25143;
											assign node25143 = (inp[4]) ? node25157 : node25144;
												assign node25144 = (inp[13]) ? node25150 : node25145;
													assign node25145 = (inp[12]) ? 4'b0000 : node25146;
														assign node25146 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node25150 = (inp[12]) ? 4'b1000 : node25151;
														assign node25151 = (inp[10]) ? node25153 : 4'b1000;
															assign node25153 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node25157 = (inp[7]) ? node25173 : node25158;
													assign node25158 = (inp[13]) ? node25164 : node25159;
														assign node25159 = (inp[10]) ? node25161 : 4'b0100;
															assign node25161 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node25164 = (inp[2]) ? node25168 : node25165;
															assign node25165 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node25168 = (inp[12]) ? 4'b1100 : node25169;
																assign node25169 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node25173 = (inp[13]) ? node25179 : node25174;
														assign node25174 = (inp[12]) ? 4'b0000 : node25175;
															assign node25175 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node25179 = (inp[12]) ? 4'b1000 : node25180;
															assign node25180 = (inp[10]) ? 4'b0100 : 4'b1000;
											assign node25184 = (inp[13]) ? node25202 : node25185;
												assign node25185 = (inp[7]) ? node25197 : node25186;
													assign node25186 = (inp[4]) ? node25192 : node25187;
														assign node25187 = (inp[12]) ? 4'b0001 : node25188;
															assign node25188 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node25192 = (inp[10]) ? node25194 : 4'b0101;
															assign node25194 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node25197 = (inp[10]) ? node25199 : 4'b0001;
														assign node25199 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node25202 = (inp[2]) ? node25222 : node25203;
													assign node25203 = (inp[4]) ? node25209 : node25204;
														assign node25204 = (inp[12]) ? 4'b1001 : node25205;
															assign node25205 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node25209 = (inp[7]) ? node25217 : node25210;
															assign node25210 = (inp[10]) ? node25214 : node25211;
																assign node25211 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node25214 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node25217 = (inp[12]) ? 4'b1001 : node25218;
																assign node25218 = (inp[10]) ? 4'b0000 : 4'b1001;
													assign node25222 = (inp[12]) ? node25232 : node25223;
														assign node25223 = (inp[10]) ? node25227 : node25224;
															assign node25224 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node25227 = (inp[4]) ? 4'b0101 : node25228;
																assign node25228 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node25232 = (inp[4]) ? node25234 : 4'b1001;
															assign node25234 = (inp[7]) ? 4'b1001 : 4'b1101;
									assign node25237 = (inp[10]) ? node25309 : node25238;
										assign node25238 = (inp[2]) ? node25274 : node25239;
											assign node25239 = (inp[11]) ? node25251 : node25240;
												assign node25240 = (inp[4]) ? node25246 : node25241;
													assign node25241 = (inp[13]) ? node25243 : 4'b0001;
														assign node25243 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node25246 = (inp[13]) ? node25248 : 4'b0101;
														assign node25248 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node25251 = (inp[12]) ? node25263 : node25252;
													assign node25252 = (inp[4]) ? node25258 : node25253;
														assign node25253 = (inp[7]) ? 4'b1000 : node25254;
															assign node25254 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node25258 = (inp[7]) ? 4'b1100 : node25259;
															assign node25259 = (inp[13]) ? 4'b0001 : 4'b1100;
													assign node25263 = (inp[4]) ? node25269 : node25264;
														assign node25264 = (inp[13]) ? node25266 : 4'b0000;
															assign node25266 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node25269 = (inp[7]) ? 4'b0100 : node25270;
															assign node25270 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node25274 = (inp[13]) ? node25292 : node25275;
												assign node25275 = (inp[14]) ? node25281 : node25276;
													assign node25276 = (inp[4]) ? node25278 : 4'b0101;
														assign node25278 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node25281 = (inp[11]) ? node25287 : node25282;
														assign node25282 = (inp[7]) ? 4'b0100 : node25283;
															assign node25283 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node25287 = (inp[7]) ? 4'b0101 : node25288;
															assign node25288 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node25292 = (inp[7]) ? node25304 : node25293;
													assign node25293 = (inp[4]) ? node25299 : node25294;
														assign node25294 = (inp[11]) ? 4'b1101 : node25295;
															assign node25295 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node25299 = (inp[11]) ? node25301 : 4'b0001;
															assign node25301 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node25304 = (inp[14]) ? node25306 : 4'b1101;
														assign node25306 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node25309 = (inp[11]) ? node25379 : node25310;
											assign node25310 = (inp[2]) ? node25326 : node25311;
												assign node25311 = (inp[4]) ? node25317 : node25312;
													assign node25312 = (inp[13]) ? node25314 : 4'b1001;
														assign node25314 = (inp[7]) ? 4'b1001 : 4'b1101;
													assign node25317 = (inp[13]) ? node25319 : 4'b1101;
														assign node25319 = (inp[7]) ? 4'b1101 : node25320;
															assign node25320 = (inp[14]) ? node25322 : 4'b1000;
																assign node25322 = (inp[12]) ? 4'b0001 : 4'b1001;
												assign node25326 = (inp[14]) ? node25354 : node25327;
													assign node25327 = (inp[4]) ? node25343 : node25328;
														assign node25328 = (inp[7]) ? node25336 : node25329;
															assign node25329 = (inp[13]) ? node25333 : node25330;
																assign node25330 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node25333 = (inp[12]) ? 4'b1101 : 4'b0001;
															assign node25336 = (inp[13]) ? node25340 : node25337;
																assign node25337 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node25340 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node25343 = (inp[7]) ? node25349 : node25344;
															assign node25344 = (inp[13]) ? 4'b1001 : node25345;
																assign node25345 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node25349 = (inp[13]) ? 4'b0001 : node25350;
																assign node25350 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node25354 = (inp[7]) ? node25364 : node25355;
														assign node25355 = (inp[4]) ? node25359 : node25356;
															assign node25356 = (inp[12]) ? 4'b1100 : 4'b0000;
															assign node25359 = (inp[13]) ? 4'b1001 : node25360;
																assign node25360 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node25364 = (inp[4]) ? node25372 : node25365;
															assign node25365 = (inp[13]) ? node25369 : node25366;
																assign node25366 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node25369 = (inp[12]) ? 4'b1100 : 4'b0100;
															assign node25372 = (inp[13]) ? node25376 : node25373;
																assign node25373 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node25376 = (inp[12]) ? 4'b1100 : 4'b0000;
											assign node25379 = (inp[2]) ? node25403 : node25380;
												assign node25380 = (inp[12]) ? node25392 : node25381;
													assign node25381 = (inp[4]) ? node25387 : node25382;
														assign node25382 = (inp[13]) ? 4'b0100 : node25383;
															assign node25383 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node25387 = (inp[13]) ? 4'b0000 : node25388;
															assign node25388 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node25392 = (inp[4]) ? node25398 : node25393;
														assign node25393 = (inp[13]) ? node25395 : 4'b1000;
															assign node25395 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node25398 = (inp[7]) ? 4'b1100 : node25399;
															assign node25399 = (inp[13]) ? 4'b1001 : 4'b1100;
												assign node25403 = (inp[4]) ? node25413 : node25404;
													assign node25404 = (inp[13]) ? node25408 : node25405;
														assign node25405 = (inp[12]) ? 4'b0101 : 4'b1101;
														assign node25408 = (inp[12]) ? 4'b1101 : node25409;
															assign node25409 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node25413 = (inp[7]) ? node25421 : node25414;
														assign node25414 = (inp[13]) ? node25418 : node25415;
															assign node25415 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node25418 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node25421 = (inp[12]) ? node25425 : node25422;
															assign node25422 = (inp[13]) ? 4'b0000 : 4'b1101;
															assign node25425 = (inp[13]) ? 4'b1101 : 4'b0101;
								assign node25428 = (inp[11]) ? node25708 : node25429;
									assign node25429 = (inp[14]) ? node25581 : node25430;
										assign node25430 = (inp[3]) ? node25482 : node25431;
											assign node25431 = (inp[13]) ? node25449 : node25432;
												assign node25432 = (inp[10]) ? node25444 : node25433;
													assign node25433 = (inp[12]) ? node25439 : node25434;
														assign node25434 = (inp[4]) ? node25436 : 4'b1000;
															assign node25436 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node25439 = (inp[7]) ? 4'b0000 : node25440;
															assign node25440 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node25444 = (inp[7]) ? 4'b1000 : node25445;
														assign node25445 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node25449 = (inp[2]) ? node25471 : node25450;
													assign node25450 = (inp[4]) ? node25458 : node25451;
														assign node25451 = (inp[7]) ? node25453 : 4'b0100;
															assign node25453 = (inp[10]) ? 4'b0000 : node25454;
																assign node25454 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node25458 = (inp[7]) ? node25466 : node25459;
															assign node25459 = (inp[10]) ? node25463 : node25460;
																assign node25460 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node25463 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node25466 = (inp[10]) ? 4'b0001 : node25467;
																assign node25467 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node25471 = (inp[10]) ? node25477 : node25472;
														assign node25472 = (inp[12]) ? 4'b1000 : node25473;
															assign node25473 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25477 = (inp[4]) ? 4'b0100 : node25478;
															assign node25478 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node25482 = (inp[2]) ? node25534 : node25483;
												assign node25483 = (inp[4]) ? node25513 : node25484;
													assign node25484 = (inp[7]) ? node25500 : node25485;
														assign node25485 = (inp[13]) ? node25493 : node25486;
															assign node25486 = (inp[12]) ? node25490 : node25487;
																assign node25487 = (inp[10]) ? 4'b0101 : 4'b1001;
																assign node25490 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node25493 = (inp[10]) ? node25497 : node25494;
																assign node25494 = (inp[12]) ? 4'b0101 : 4'b1101;
																assign node25497 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node25500 = (inp[13]) ? node25508 : node25501;
															assign node25501 = (inp[10]) ? node25505 : node25502;
																assign node25502 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node25505 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node25508 = (inp[10]) ? 4'b1001 : node25509;
																assign node25509 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node25513 = (inp[7]) ? node25525 : node25514;
														assign node25514 = (inp[13]) ? node25522 : node25515;
															assign node25515 = (inp[12]) ? node25519 : node25516;
																assign node25516 = (inp[10]) ? 4'b0001 : 4'b1101;
																assign node25519 = (inp[10]) ? 4'b1101 : 4'b0101;
															assign node25522 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node25525 = (inp[12]) ? node25531 : node25526;
															assign node25526 = (inp[10]) ? node25528 : 4'b1101;
																assign node25528 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node25531 = (inp[10]) ? 4'b1101 : 4'b0101;
												assign node25534 = (inp[4]) ? node25552 : node25535;
													assign node25535 = (inp[13]) ? node25541 : node25536;
														assign node25536 = (inp[12]) ? node25538 : 4'b1100;
															assign node25538 = (inp[10]) ? 4'b1100 : 4'b0100;
														assign node25541 = (inp[7]) ? node25547 : node25542;
															assign node25542 = (inp[12]) ? node25544 : 4'b0000;
																assign node25544 = (inp[10]) ? 4'b0000 : 4'b1100;
															assign node25547 = (inp[12]) ? node25549 : 4'b0100;
																assign node25549 = (inp[10]) ? 4'b0100 : 4'b1100;
													assign node25552 = (inp[7]) ? node25568 : node25553;
														assign node25553 = (inp[13]) ? node25561 : node25554;
															assign node25554 = (inp[12]) ? node25558 : node25555;
																assign node25555 = (inp[10]) ? 4'b0001 : 4'b1000;
																assign node25558 = (inp[10]) ? 4'b1000 : 4'b0000;
															assign node25561 = (inp[12]) ? node25565 : node25562;
																assign node25562 = (inp[10]) ? 4'b0001 : 4'b1001;
																assign node25565 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node25568 = (inp[13]) ? node25574 : node25569;
															assign node25569 = (inp[10]) ? 4'b1100 : node25570;
																assign node25570 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node25574 = (inp[12]) ? node25578 : node25575;
																assign node25575 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node25578 = (inp[10]) ? 4'b0000 : 4'b1100;
										assign node25581 = (inp[13]) ? node25639 : node25582;
											assign node25582 = (inp[12]) ? node25620 : node25583;
												assign node25583 = (inp[10]) ? node25601 : node25584;
													assign node25584 = (inp[2]) ? node25592 : node25585;
														assign node25585 = (inp[3]) ? node25589 : node25586;
															assign node25586 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node25589 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node25592 = (inp[3]) ? node25596 : node25593;
															assign node25593 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node25596 = (inp[4]) ? node25598 : 4'b0101;
																assign node25598 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node25601 = (inp[3]) ? node25613 : node25602;
														assign node25602 = (inp[2]) ? node25608 : node25603;
															assign node25603 = (inp[7]) ? 4'b1001 : node25604;
																assign node25604 = (inp[4]) ? 4'b0001 : 4'b1001;
															assign node25608 = (inp[4]) ? node25610 : 4'b1001;
																assign node25610 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node25613 = (inp[7]) ? node25617 : node25614;
															assign node25614 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node25617 = (inp[2]) ? 4'b1101 : 4'b0001;
												assign node25620 = (inp[4]) ? node25630 : node25621;
													assign node25621 = (inp[2]) ? node25627 : node25622;
														assign node25622 = (inp[10]) ? node25624 : 4'b0001;
															assign node25624 = (inp[3]) ? 4'b1001 : 4'b0001;
														assign node25627 = (inp[3]) ? 4'b0101 : 4'b0001;
													assign node25630 = (inp[7]) ? node25636 : node25631;
														assign node25631 = (inp[3]) ? node25633 : 4'b0101;
															assign node25633 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node25636 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node25639 = (inp[3]) ? node25667 : node25640;
												assign node25640 = (inp[12]) ? node25654 : node25641;
													assign node25641 = (inp[10]) ? node25649 : node25642;
														assign node25642 = (inp[2]) ? node25644 : 4'b1001;
															assign node25644 = (inp[4]) ? node25646 : 4'b1001;
																assign node25646 = (inp[7]) ? 4'b1001 : 4'b1101;
														assign node25649 = (inp[7]) ? node25651 : 4'b0101;
															assign node25651 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node25654 = (inp[2]) ? node25662 : node25655;
														assign node25655 = (inp[10]) ? 4'b1001 : node25656;
															assign node25656 = (inp[7]) ? 4'b1001 : node25657;
																assign node25657 = (inp[4]) ? 4'b0001 : 4'b1001;
														assign node25662 = (inp[4]) ? node25664 : 4'b1001;
															assign node25664 = (inp[7]) ? 4'b1001 : 4'b1101;
												assign node25667 = (inp[4]) ? node25689 : node25668;
													assign node25668 = (inp[2]) ? node25682 : node25669;
														assign node25669 = (inp[7]) ? node25675 : node25670;
															assign node25670 = (inp[10]) ? 4'b1101 : node25671;
																assign node25671 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node25675 = (inp[12]) ? node25679 : node25676;
																assign node25676 = (inp[10]) ? 4'b0101 : 4'b1001;
																assign node25679 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node25682 = (inp[12]) ? 4'b1101 : node25683;
															assign node25683 = (inp[10]) ? node25685 : 4'b1101;
																assign node25685 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node25689 = (inp[7]) ? node25699 : node25690;
														assign node25690 = (inp[2]) ? node25692 : 4'b0000;
															assign node25692 = (inp[10]) ? node25696 : node25693;
																assign node25693 = (inp[12]) ? 4'b0001 : 4'b1001;
																assign node25696 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node25699 = (inp[10]) ? node25705 : node25700;
															assign node25700 = (inp[2]) ? 4'b1101 : node25701;
																assign node25701 = (inp[12]) ? 4'b0101 : 4'b1101;
															assign node25705 = (inp[12]) ? 4'b1101 : 4'b0001;
									assign node25708 = (inp[10]) ? node25778 : node25709;
										assign node25709 = (inp[3]) ? node25741 : node25710;
											assign node25710 = (inp[7]) ? node25732 : node25711;
												assign node25711 = (inp[4]) ? node25719 : node25712;
													assign node25712 = (inp[13]) ? node25716 : node25713;
														assign node25713 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node25716 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node25719 = (inp[2]) ? node25725 : node25720;
														assign node25720 = (inp[13]) ? 4'b1000 : node25721;
															assign node25721 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node25725 = (inp[13]) ? node25729 : node25726;
															assign node25726 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node25729 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node25732 = (inp[13]) ? node25736 : node25733;
													assign node25733 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node25736 = (inp[12]) ? 4'b1000 : node25737;
														assign node25737 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node25741 = (inp[2]) ? node25755 : node25742;
												assign node25742 = (inp[4]) ? node25748 : node25743;
													assign node25743 = (inp[13]) ? node25745 : 4'b1000;
														assign node25745 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node25748 = (inp[7]) ? 4'b1100 : node25749;
														assign node25749 = (inp[13]) ? node25751 : 4'b1100;
															assign node25751 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node25755 = (inp[7]) ? node25769 : node25756;
													assign node25756 = (inp[4]) ? node25764 : node25757;
														assign node25757 = (inp[12]) ? node25761 : node25758;
															assign node25758 = (inp[13]) ? 4'b0000 : 4'b1100;
															assign node25761 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node25764 = (inp[13]) ? 4'b1000 : node25765;
															assign node25765 = (inp[12]) ? 4'b0000 : 4'b1000;
													assign node25769 = (inp[12]) ? node25775 : node25770;
														assign node25770 = (inp[13]) ? node25772 : 4'b1100;
															assign node25772 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node25775 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node25778 = (inp[13]) ? node25800 : node25779;
											assign node25779 = (inp[3]) ? node25787 : node25780;
												assign node25780 = (inp[4]) ? node25782 : 4'b1000;
													assign node25782 = (inp[7]) ? 4'b1000 : node25783;
														assign node25783 = (inp[2]) ? 4'b1100 : 4'b0000;
												assign node25787 = (inp[2]) ? node25795 : node25788;
													assign node25788 = (inp[7]) ? node25792 : node25789;
														assign node25789 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node25792 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node25795 = (inp[4]) ? node25797 : 4'b1100;
														assign node25797 = (inp[7]) ? 4'b1100 : 4'b0000;
											assign node25800 = (inp[4]) ? node25814 : node25801;
												assign node25801 = (inp[2]) ? node25807 : node25802;
													assign node25802 = (inp[3]) ? 4'b0100 : node25803;
														assign node25803 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node25807 = (inp[3]) ? node25811 : node25808;
														assign node25808 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node25811 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node25814 = (inp[3]) ? 4'b0000 : node25815;
													assign node25815 = (inp[2]) ? 4'b0100 : 4'b0000;
							assign node25819 = (inp[3]) ? node26227 : node25820;
								assign node25820 = (inp[11]) ? node26074 : node25821;
									assign node25821 = (inp[2]) ? node25967 : node25822;
										assign node25822 = (inp[13]) ? node25890 : node25823;
											assign node25823 = (inp[7]) ? node25859 : node25824;
												assign node25824 = (inp[10]) ? node25838 : node25825;
													assign node25825 = (inp[1]) ? node25833 : node25826;
														assign node25826 = (inp[14]) ? node25830 : node25827;
															assign node25827 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node25830 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node25833 = (inp[4]) ? node25835 : 4'b1000;
															assign node25835 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node25838 = (inp[12]) ? node25850 : node25839;
														assign node25839 = (inp[1]) ? node25845 : node25840;
															assign node25840 = (inp[4]) ? 4'b1100 : node25841;
																assign node25841 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node25845 = (inp[4]) ? node25847 : 4'b1100;
																assign node25847 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node25850 = (inp[4]) ? 4'b0100 : node25851;
															assign node25851 = (inp[1]) ? node25855 : node25852;
																assign node25852 = (inp[14]) ? 4'b1001 : 4'b0100;
																assign node25855 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node25859 = (inp[4]) ? node25881 : node25860;
													assign node25860 = (inp[1]) ? node25872 : node25861;
														assign node25861 = (inp[14]) ? node25867 : node25862;
															assign node25862 = (inp[10]) ? 4'b0000 : node25863;
																assign node25863 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node25867 = (inp[12]) ? node25869 : 4'b0001;
																assign node25869 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node25872 = (inp[14]) ? node25876 : node25873;
															assign node25873 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node25876 = (inp[12]) ? node25878 : 4'b1000;
																assign node25878 = (inp[10]) ? 4'b0000 : 4'b1000;
													assign node25881 = (inp[1]) ? node25885 : node25882;
														assign node25882 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node25885 = (inp[12]) ? 4'b1000 : node25886;
															assign node25886 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node25890 = (inp[4]) ? node25934 : node25891;
												assign node25891 = (inp[1]) ? node25917 : node25892;
													assign node25892 = (inp[14]) ? node25906 : node25893;
														assign node25893 = (inp[7]) ? node25899 : node25894;
															assign node25894 = (inp[10]) ? node25896 : 4'b1100;
																assign node25896 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node25899 = (inp[12]) ? node25903 : node25900;
																assign node25900 = (inp[10]) ? 4'b1100 : 4'b0100;
																assign node25903 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node25906 = (inp[10]) ? node25910 : node25907;
															assign node25907 = (inp[7]) ? 4'b1001 : 4'b1101;
															assign node25910 = (inp[7]) ? node25914 : node25911;
																assign node25911 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node25914 = (inp[12]) ? 4'b0101 : 4'b1101;
													assign node25917 = (inp[10]) ? node25929 : node25918;
														assign node25918 = (inp[14]) ? node25924 : node25919;
															assign node25919 = (inp[12]) ? 4'b0101 : node25920;
																assign node25920 = (inp[7]) ? 4'b0101 : 4'b0000;
															assign node25924 = (inp[12]) ? 4'b0100 : node25925;
																assign node25925 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node25929 = (inp[12]) ? node25931 : 4'b0000;
															assign node25931 = (inp[7]) ? 4'b1100 : 4'b1000;
												assign node25934 = (inp[1]) ? node25954 : node25935;
													assign node25935 = (inp[12]) ? node25941 : node25936;
														assign node25936 = (inp[14]) ? node25938 : 4'b0001;
															assign node25938 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node25941 = (inp[14]) ? node25947 : node25942;
															assign node25942 = (inp[10]) ? node25944 : 4'b0100;
																assign node25944 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node25947 = (inp[10]) ? node25951 : node25948;
																assign node25948 = (inp[7]) ? 4'b0100 : 4'b1000;
																assign node25951 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node25954 = (inp[14]) ? node25962 : node25955;
														assign node25955 = (inp[10]) ? node25957 : 4'b1000;
															assign node25957 = (inp[7]) ? node25959 : 4'b1001;
																assign node25959 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node25962 = (inp[10]) ? 4'b1001 : node25963;
															assign node25963 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node25967 = (inp[4]) ? node26005 : node25968;
											assign node25968 = (inp[10]) ? node25986 : node25969;
												assign node25969 = (inp[1]) ? node25975 : node25970;
													assign node25970 = (inp[13]) ? node25972 : 4'b0001;
														assign node25972 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node25975 = (inp[12]) ? node25981 : node25976;
														assign node25976 = (inp[7]) ? 4'b1001 : node25977;
															assign node25977 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node25981 = (inp[7]) ? 4'b0001 : node25982;
															assign node25982 = (inp[13]) ? 4'b0101 : 4'b0001;
												assign node25986 = (inp[1]) ? node25992 : node25987;
													assign node25987 = (inp[7]) ? 4'b1001 : node25988;
														assign node25988 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node25992 = (inp[12]) ? node26000 : node25993;
														assign node25993 = (inp[13]) ? node25997 : node25994;
															assign node25994 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node25997 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node26000 = (inp[7]) ? 4'b1001 : node26001;
															assign node26001 = (inp[13]) ? 4'b1101 : 4'b1001;
											assign node26005 = (inp[10]) ? node26043 : node26006;
												assign node26006 = (inp[7]) ? node26028 : node26007;
													assign node26007 = (inp[13]) ? node26017 : node26008;
														assign node26008 = (inp[1]) ? node26014 : node26009;
															assign node26009 = (inp[14]) ? 4'b0001 : node26010;
																assign node26010 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node26014 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node26017 = (inp[14]) ? node26025 : node26018;
															assign node26018 = (inp[12]) ? node26022 : node26019;
																assign node26019 = (inp[1]) ? 4'b0000 : 4'b0100;
																assign node26022 = (inp[1]) ? 4'b0101 : 4'b1000;
															assign node26025 = (inp[1]) ? 4'b0000 : 4'b1001;
													assign node26028 = (inp[13]) ? node26034 : node26029;
														assign node26029 = (inp[12]) ? 4'b0101 : node26030;
															assign node26030 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node26034 = (inp[1]) ? node26040 : node26035;
															assign node26035 = (inp[14]) ? 4'b1001 : node26036;
																assign node26036 = (inp[12]) ? 4'b1000 : 4'b0000;
															assign node26040 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node26043 = (inp[13]) ? node26057 : node26044;
													assign node26044 = (inp[1]) ? node26050 : node26045;
														assign node26045 = (inp[14]) ? node26047 : 4'b0000;
															assign node26047 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node26050 = (inp[12]) ? node26054 : node26051;
															assign node26051 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node26054 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node26057 = (inp[7]) ? node26065 : node26058;
														assign node26058 = (inp[1]) ? node26062 : node26059;
															assign node26059 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node26062 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node26065 = (inp[1]) ? node26069 : node26066;
															assign node26066 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node26069 = (inp[12]) ? node26071 : 4'b0000;
																assign node26071 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node26074 = (inp[1]) ? node26158 : node26075;
										assign node26075 = (inp[4]) ? node26119 : node26076;
											assign node26076 = (inp[2]) ? node26094 : node26077;
												assign node26077 = (inp[13]) ? node26085 : node26078;
													assign node26078 = (inp[10]) ? node26082 : node26079;
														assign node26079 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node26082 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node26085 = (inp[10]) ? node26091 : node26086;
														assign node26086 = (inp[7]) ? 4'b1001 : node26087;
															assign node26087 = (inp[12]) ? 4'b1101 : 4'b0101;
														assign node26091 = (inp[7]) ? 4'b1101 : 4'b1000;
												assign node26094 = (inp[13]) ? node26104 : node26095;
													assign node26095 = (inp[12]) ? node26101 : node26096;
														assign node26096 = (inp[10]) ? node26098 : 4'b1000;
															assign node26098 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node26101 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node26104 = (inp[7]) ? node26112 : node26105;
														assign node26105 = (inp[10]) ? node26109 : node26106;
															assign node26106 = (inp[12]) ? 4'b0100 : 4'b1100;
															assign node26109 = (inp[12]) ? 4'b1100 : 4'b0100;
														assign node26112 = (inp[12]) ? node26116 : node26113;
															assign node26113 = (inp[10]) ? 4'b0100 : 4'b1000;
															assign node26116 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node26119 = (inp[13]) ? node26141 : node26120;
												assign node26120 = (inp[2]) ? node26132 : node26121;
													assign node26121 = (inp[12]) ? node26127 : node26122;
														assign node26122 = (inp[10]) ? node26124 : 4'b1000;
															assign node26124 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node26127 = (inp[7]) ? 4'b1000 : node26128;
															assign node26128 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node26132 = (inp[10]) ? 4'b0001 : node26133;
														assign node26133 = (inp[7]) ? node26137 : node26134;
															assign node26134 = (inp[12]) ? 4'b0001 : 4'b1001;
															assign node26137 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node26141 = (inp[10]) ? node26149 : node26142;
													assign node26142 = (inp[2]) ? node26144 : 4'b0001;
														assign node26144 = (inp[12]) ? 4'b1001 : node26145;
															assign node26145 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node26149 = (inp[7]) ? node26155 : node26150;
														assign node26150 = (inp[12]) ? node26152 : 4'b1000;
															assign node26152 = (inp[2]) ? 4'b1000 : 4'b0000;
														assign node26155 = (inp[2]) ? 4'b1001 : 4'b0001;
										assign node26158 = (inp[13]) ? node26192 : node26159;
											assign node26159 = (inp[2]) ? node26179 : node26160;
												assign node26160 = (inp[10]) ? node26172 : node26161;
													assign node26161 = (inp[7]) ? node26167 : node26162;
														assign node26162 = (inp[12]) ? node26164 : 4'b0100;
															assign node26164 = (inp[4]) ? 4'b0100 : 4'b1000;
														assign node26167 = (inp[12]) ? node26169 : 4'b0000;
															assign node26169 = (inp[4]) ? 4'b0000 : 4'b1000;
													assign node26172 = (inp[7]) ? node26176 : node26173;
														assign node26173 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node26176 = (inp[4]) ? 4'b0100 : 4'b1000;
												assign node26179 = (inp[4]) ? node26185 : node26180;
													assign node26180 = (inp[10]) ? node26182 : 4'b1000;
														assign node26182 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node26185 = (inp[10]) ? 4'b1000 : node26186;
														assign node26186 = (inp[12]) ? node26188 : 4'b0000;
															assign node26188 = (inp[7]) ? 4'b1100 : 4'b1000;
											assign node26192 = (inp[10]) ? node26220 : node26193;
												assign node26193 = (inp[4]) ? node26203 : node26194;
													assign node26194 = (inp[2]) ? node26200 : node26195;
														assign node26195 = (inp[7]) ? node26197 : 4'b0000;
															assign node26197 = (inp[12]) ? 4'b0100 : 4'b1100;
														assign node26200 = (inp[7]) ? 4'b1000 : 4'b1100;
													assign node26203 = (inp[7]) ? node26211 : node26204;
														assign node26204 = (inp[12]) ? node26208 : node26205;
															assign node26205 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node26208 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node26211 = (inp[14]) ? 4'b1000 : node26212;
															assign node26212 = (inp[12]) ? node26216 : node26213;
																assign node26213 = (inp[2]) ? 4'b1000 : 4'b0000;
																assign node26216 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node26220 = (inp[4]) ? 4'b0000 : node26221;
													assign node26221 = (inp[7]) ? node26223 : 4'b0000;
														assign node26223 = (inp[2]) ? 4'b0100 : 4'b0000;
								assign node26227 = (inp[4]) ? node26447 : node26228;
									assign node26228 = (inp[11]) ? node26374 : node26229;
										assign node26229 = (inp[12]) ? node26305 : node26230;
											assign node26230 = (inp[13]) ? node26268 : node26231;
												assign node26231 = (inp[1]) ? node26245 : node26232;
													assign node26232 = (inp[2]) ? node26238 : node26233;
														assign node26233 = (inp[10]) ? node26235 : 4'b1001;
															assign node26235 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node26238 = (inp[10]) ? node26240 : 4'b1000;
															assign node26240 = (inp[7]) ? 4'b1000 : node26241;
																assign node26241 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node26245 = (inp[7]) ? node26257 : node26246;
														assign node26246 = (inp[2]) ? node26252 : node26247;
															assign node26247 = (inp[14]) ? 4'b1000 : node26248;
																assign node26248 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node26252 = (inp[14]) ? 4'b0001 : node26253;
																assign node26253 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node26257 = (inp[2]) ? node26263 : node26258;
															assign node26258 = (inp[10]) ? node26260 : 4'b0001;
																assign node26260 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node26263 = (inp[14]) ? 4'b0001 : node26264;
																assign node26264 = (inp[10]) ? 4'b1000 : 4'b0000;
												assign node26268 = (inp[1]) ? node26290 : node26269;
													assign node26269 = (inp[10]) ? node26283 : node26270;
														assign node26270 = (inp[14]) ? node26278 : node26271;
															assign node26271 = (inp[2]) ? node26275 : node26272;
																assign node26272 = (inp[7]) ? 4'b1000 : 4'b0001;
																assign node26275 = (inp[7]) ? 4'b0001 : 4'b1001;
															assign node26278 = (inp[2]) ? 4'b0000 : node26279;
																assign node26279 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node26283 = (inp[14]) ? 4'b0001 : node26284;
															assign node26284 = (inp[2]) ? 4'b0000 : node26285;
																assign node26285 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node26290 = (inp[10]) ? node26300 : node26291;
														assign node26291 = (inp[2]) ? node26295 : node26292;
															assign node26292 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node26295 = (inp[7]) ? 4'b0001 : node26296;
																assign node26296 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26300 = (inp[7]) ? node26302 : 4'b1000;
															assign node26302 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node26305 = (inp[2]) ? node26349 : node26306;
												assign node26306 = (inp[7]) ? node26328 : node26307;
													assign node26307 = (inp[1]) ? node26317 : node26308;
														assign node26308 = (inp[13]) ? node26310 : 4'b0001;
															assign node26310 = (inp[10]) ? node26314 : node26311;
																assign node26311 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node26314 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node26317 = (inp[10]) ? node26325 : node26318;
															assign node26318 = (inp[13]) ? node26322 : node26319;
																assign node26319 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node26322 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node26325 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node26328 = (inp[1]) ? node26340 : node26329;
														assign node26329 = (inp[14]) ? node26335 : node26330;
															assign node26330 = (inp[13]) ? 4'b0001 : node26331;
																assign node26331 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node26335 = (inp[10]) ? 4'b0001 : node26336;
																assign node26336 = (inp[13]) ? 4'b1000 : 4'b0001;
														assign node26340 = (inp[14]) ? node26346 : node26341;
															assign node26341 = (inp[10]) ? 4'b0001 : node26342;
																assign node26342 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node26346 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node26349 = (inp[13]) ? node26359 : node26350;
													assign node26350 = (inp[10]) ? node26354 : node26351;
														assign node26351 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node26354 = (inp[14]) ? node26356 : 4'b0000;
															assign node26356 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node26359 = (inp[10]) ? node26365 : node26360;
														assign node26360 = (inp[1]) ? 4'b0001 : node26361;
															assign node26361 = (inp[7]) ? 4'b1000 : 4'b0001;
														assign node26365 = (inp[1]) ? node26371 : node26366;
															assign node26366 = (inp[14]) ? 4'b1001 : node26367;
																assign node26367 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node26371 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node26374 = (inp[1]) ? node26420 : node26375;
											assign node26375 = (inp[12]) ? node26399 : node26376;
												assign node26376 = (inp[10]) ? node26386 : node26377;
													assign node26377 = (inp[2]) ? node26383 : node26378;
														assign node26378 = (inp[7]) ? 4'b0000 : node26379;
															assign node26379 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node26383 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node26386 = (inp[2]) ? node26394 : node26387;
														assign node26387 = (inp[14]) ? node26389 : 4'b1001;
															assign node26389 = (inp[7]) ? node26391 : 4'b0000;
																assign node26391 = (inp[13]) ? 4'b0000 : 4'b1001;
														assign node26394 = (inp[7]) ? 4'b0001 : node26395;
															assign node26395 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node26399 = (inp[13]) ? node26409 : node26400;
													assign node26400 = (inp[10]) ? node26402 : 4'b1000;
														assign node26402 = (inp[7]) ? node26406 : node26403;
															assign node26403 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node26406 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node26409 = (inp[7]) ? node26415 : node26410;
														assign node26410 = (inp[2]) ? node26412 : 4'b1001;
															assign node26412 = (inp[10]) ? 4'b0000 : 4'b1000;
														assign node26415 = (inp[2]) ? 4'b0001 : node26416;
															assign node26416 = (inp[10]) ? 4'b1000 : 4'b0000;
											assign node26420 = (inp[10]) ? node26440 : node26421;
												assign node26421 = (inp[13]) ? node26431 : node26422;
													assign node26422 = (inp[2]) ? node26426 : node26423;
														assign node26423 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node26426 = (inp[12]) ? 4'b0000 : node26427;
															assign node26427 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node26431 = (inp[14]) ? 4'b1000 : node26432;
														assign node26432 = (inp[7]) ? node26434 : 4'b1000;
															assign node26434 = (inp[12]) ? 4'b1000 : node26435;
																assign node26435 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node26440 = (inp[13]) ? 4'b0000 : node26441;
													assign node26441 = (inp[2]) ? node26443 : 4'b0000;
														assign node26443 = (inp[7]) ? 4'b1000 : 4'b0000;
									assign node26447 = (inp[13]) ? node26577 : node26448;
										assign node26448 = (inp[1]) ? node26520 : node26449;
											assign node26449 = (inp[12]) ? node26485 : node26450;
												assign node26450 = (inp[2]) ? node26470 : node26451;
													assign node26451 = (inp[7]) ? node26459 : node26452;
														assign node26452 = (inp[10]) ? node26454 : 4'b0001;
															assign node26454 = (inp[11]) ? 4'b0001 : node26455;
																assign node26455 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node26459 = (inp[10]) ? node26465 : node26460;
															assign node26460 = (inp[11]) ? 4'b0000 : node26461;
																assign node26461 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node26465 = (inp[11]) ? 4'b0001 : node26466;
																assign node26466 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node26470 = (inp[7]) ? node26480 : node26471;
														assign node26471 = (inp[11]) ? 4'b1000 : node26472;
															assign node26472 = (inp[10]) ? node26476 : node26473;
																assign node26473 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node26476 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26480 = (inp[11]) ? 4'b0001 : node26481;
															assign node26481 = (inp[14]) ? 4'b0000 : 4'b1000;
												assign node26485 = (inp[10]) ? node26499 : node26486;
													assign node26486 = (inp[11]) ? node26492 : node26487;
														assign node26487 = (inp[7]) ? 4'b1000 : node26488;
															assign node26488 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node26492 = (inp[2]) ? node26496 : node26493;
															assign node26493 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node26496 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node26499 = (inp[7]) ? node26509 : node26500;
														assign node26500 = (inp[2]) ? node26506 : node26501;
															assign node26501 = (inp[11]) ? 4'b1000 : node26502;
																assign node26502 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node26506 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26509 = (inp[2]) ? node26515 : node26510;
															assign node26510 = (inp[11]) ? 4'b0001 : node26511;
																assign node26511 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node26515 = (inp[14]) ? node26517 : 4'b1000;
																assign node26517 = (inp[11]) ? 4'b1000 : 4'b0001;
											assign node26520 = (inp[11]) ? node26552 : node26521;
												assign node26521 = (inp[7]) ? node26533 : node26522;
													assign node26522 = (inp[14]) ? 4'b0000 : node26523;
														assign node26523 = (inp[12]) ? 4'b0001 : node26524;
															assign node26524 = (inp[2]) ? node26528 : node26525;
																assign node26525 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node26528 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node26533 = (inp[2]) ? node26547 : node26534;
														assign node26534 = (inp[12]) ? node26542 : node26535;
															assign node26535 = (inp[10]) ? node26539 : node26536;
																assign node26536 = (inp[14]) ? 4'b0000 : 4'b0001;
																assign node26539 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node26542 = (inp[10]) ? node26544 : 4'b1001;
																assign node26544 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node26547 = (inp[10]) ? 4'b0001 : node26548;
															assign node26548 = (inp[12]) ? 4'b1001 : 4'b0001;
												assign node26552 = (inp[10]) ? 4'b0000 : node26553;
													assign node26553 = (inp[14]) ? node26565 : node26554;
														assign node26554 = (inp[2]) ? node26560 : node26555;
															assign node26555 = (inp[7]) ? 4'b0000 : node26556;
																assign node26556 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node26560 = (inp[7]) ? node26562 : 4'b0000;
																assign node26562 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node26565 = (inp[12]) ? node26571 : node26566;
															assign node26566 = (inp[2]) ? 4'b0000 : node26567;
																assign node26567 = (inp[7]) ? 4'b0000 : 4'b1000;
															assign node26571 = (inp[2]) ? node26573 : 4'b0000;
																assign node26573 = (inp[7]) ? 4'b1000 : 4'b0000;
										assign node26577 = (inp[10]) ? node26633 : node26578;
											assign node26578 = (inp[11]) ? node26620 : node26579;
												assign node26579 = (inp[2]) ? node26601 : node26580;
													assign node26580 = (inp[1]) ? node26590 : node26581;
														assign node26581 = (inp[7]) ? node26587 : node26582;
															assign node26582 = (inp[12]) ? node26584 : 4'b0001;
																assign node26584 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node26587 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node26590 = (inp[7]) ? node26596 : node26591;
															assign node26591 = (inp[14]) ? 4'b0001 : node26592;
																assign node26592 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node26596 = (inp[14]) ? node26598 : 4'b0001;
																assign node26598 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node26601 = (inp[7]) ? node26611 : node26602;
														assign node26602 = (inp[12]) ? 4'b0000 : node26603;
															assign node26603 = (inp[14]) ? node26607 : node26604;
																assign node26604 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node26607 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node26611 = (inp[14]) ? 4'b0001 : node26612;
															assign node26612 = (inp[12]) ? node26616 : node26613;
																assign node26613 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node26616 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node26620 = (inp[1]) ? 4'b0000 : node26621;
													assign node26621 = (inp[7]) ? node26627 : node26622;
														assign node26622 = (inp[12]) ? 4'b0000 : node26623;
															assign node26623 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node26627 = (inp[2]) ? node26629 : 4'b0000;
															assign node26629 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node26633 = (inp[1]) ? 4'b0000 : node26634;
												assign node26634 = (inp[11]) ? 4'b0000 : node26635;
													assign node26635 = (inp[14]) ? node26645 : node26636;
														assign node26636 = (inp[7]) ? 4'b0000 : node26637;
															assign node26637 = (inp[2]) ? node26641 : node26638;
																assign node26638 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node26641 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node26645 = (inp[2]) ? node26647 : 4'b0000;
															assign node26647 = (inp[12]) ? node26649 : 4'b0000;
																assign node26649 = (inp[7]) ? 4'b0001 : 4'b0000;
					assign node26654 = (inp[6]) ? node26656 : 4'b0000;
						assign node26656 = (inp[2]) ? node27184 : node26657;
							assign node26657 = (inp[5]) ? node26759 : node26658;
								assign node26658 = (inp[3]) ? node26660 : 4'b0000;
									assign node26660 = (inp[7]) ? node26740 : node26661;
										assign node26661 = (inp[4]) ? node26679 : node26662;
											assign node26662 = (inp[13]) ? node26664 : 4'b0000;
												assign node26664 = (inp[12]) ? 4'b0000 : node26665;
													assign node26665 = (inp[10]) ? node26667 : 4'b0000;
														assign node26667 = (inp[1]) ? node26673 : node26668;
															assign node26668 = (inp[11]) ? 4'b0001 : node26669;
																assign node26669 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node26673 = (inp[14]) ? node26675 : 4'b0000;
																assign node26675 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node26679 = (inp[1]) ? node26709 : node26680;
												assign node26680 = (inp[13]) ? node26694 : node26681;
													assign node26681 = (inp[14]) ? node26687 : node26682;
														assign node26682 = (inp[10]) ? node26684 : 4'b0001;
															assign node26684 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node26687 = (inp[11]) ? 4'b0001 : node26688;
															assign node26688 = (inp[12]) ? 4'b0000 : node26689;
																assign node26689 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node26694 = (inp[11]) ? node26704 : node26695;
														assign node26695 = (inp[14]) ? node26699 : node26696;
															assign node26696 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node26699 = (inp[10]) ? node26701 : 4'b1000;
																assign node26701 = (inp[12]) ? 4'b1000 : 4'b0000;
														assign node26704 = (inp[12]) ? 4'b1001 : node26705;
															assign node26705 = (inp[10]) ? 4'b0001 : 4'b1001;
												assign node26709 = (inp[14]) ? node26721 : node26710;
													assign node26710 = (inp[13]) ? node26716 : node26711;
														assign node26711 = (inp[12]) ? node26713 : 4'b1000;
															assign node26713 = (inp[10]) ? 4'b1000 : 4'b0000;
														assign node26716 = (inp[10]) ? 4'b0000 : node26717;
															assign node26717 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node26721 = (inp[11]) ? node26731 : node26722;
														assign node26722 = (inp[13]) ? node26728 : node26723;
															assign node26723 = (inp[12]) ? 4'b0001 : node26724;
																assign node26724 = (inp[10]) ? 4'b1001 : 4'b0001;
															assign node26728 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node26731 = (inp[13]) ? node26735 : node26732;
															assign node26732 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node26735 = (inp[12]) ? node26737 : 4'b0000;
																assign node26737 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node26740 = (inp[4]) ? node26742 : 4'b0000;
											assign node26742 = (inp[13]) ? node26744 : 4'b0000;
												assign node26744 = (inp[12]) ? 4'b0000 : node26745;
													assign node26745 = (inp[10]) ? node26747 : 4'b0000;
														assign node26747 = (inp[1]) ? node26753 : node26748;
															assign node26748 = (inp[14]) ? node26750 : 4'b0001;
																assign node26750 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node26753 = (inp[11]) ? 4'b0000 : node26754;
																assign node26754 = (inp[14]) ? 4'b0001 : 4'b0000;
								assign node26759 = (inp[1]) ? node26991 : node26760;
									assign node26760 = (inp[3]) ? node26876 : node26761;
										assign node26761 = (inp[13]) ? node26807 : node26762;
											assign node26762 = (inp[12]) ? node26790 : node26763;
												assign node26763 = (inp[10]) ? node26773 : node26764;
													assign node26764 = (inp[11]) ? node26768 : node26765;
														assign node26765 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26768 = (inp[7]) ? 4'b0001 : node26769;
															assign node26769 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node26773 = (inp[11]) ? node26785 : node26774;
														assign node26774 = (inp[14]) ? node26780 : node26775;
															assign node26775 = (inp[7]) ? 4'b1001 : node26776;
																assign node26776 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node26780 = (inp[4]) ? node26782 : 4'b1000;
																assign node26782 = (inp[7]) ? 4'b1000 : 4'b1100;
														assign node26785 = (inp[7]) ? 4'b1001 : node26786;
															assign node26786 = (inp[4]) ? 4'b0000 : 4'b1001;
												assign node26790 = (inp[7]) ? node26802 : node26791;
													assign node26791 = (inp[4]) ? node26797 : node26792;
														assign node26792 = (inp[14]) ? node26794 : 4'b0001;
															assign node26794 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node26797 = (inp[11]) ? 4'b0101 : node26798;
															assign node26798 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node26802 = (inp[11]) ? 4'b0001 : node26803;
														assign node26803 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node26807 = (inp[12]) ? node26851 : node26808;
												assign node26808 = (inp[10]) ? node26832 : node26809;
													assign node26809 = (inp[14]) ? node26821 : node26810;
														assign node26810 = (inp[11]) ? node26816 : node26811;
															assign node26811 = (inp[4]) ? node26813 : 4'b1001;
																assign node26813 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node26816 = (inp[7]) ? 4'b1001 : node26817;
																assign node26817 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node26821 = (inp[11]) ? node26827 : node26822;
															assign node26822 = (inp[7]) ? 4'b1000 : node26823;
																assign node26823 = (inp[4]) ? 4'b0001 : 4'b1000;
															assign node26827 = (inp[4]) ? node26829 : 4'b1001;
																assign node26829 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node26832 = (inp[4]) ? node26844 : node26833;
														assign node26833 = (inp[7]) ? node26839 : node26834;
															assign node26834 = (inp[14]) ? node26836 : 4'b0101;
																assign node26836 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node26839 = (inp[11]) ? 4'b0001 : node26840;
																assign node26840 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26844 = (inp[11]) ? 4'b0000 : node26845;
															assign node26845 = (inp[7]) ? node26847 : 4'b1001;
																assign node26847 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node26851 = (inp[14]) ? node26861 : node26852;
													assign node26852 = (inp[7]) ? 4'b1001 : node26853;
														assign node26853 = (inp[4]) ? node26855 : 4'b1001;
															assign node26855 = (inp[11]) ? node26857 : 4'b1001;
																assign node26857 = (inp[10]) ? 4'b1000 : 4'b0000;
													assign node26861 = (inp[11]) ? node26869 : node26862;
														assign node26862 = (inp[7]) ? 4'b1000 : node26863;
															assign node26863 = (inp[4]) ? node26865 : 4'b1000;
																assign node26865 = (inp[10]) ? 4'b1001 : 4'b0001;
														assign node26869 = (inp[4]) ? node26871 : 4'b1001;
															assign node26871 = (inp[7]) ? 4'b1001 : node26872;
																assign node26872 = (inp[10]) ? 4'b1000 : 4'b0000;
										assign node26876 = (inp[4]) ? node26926 : node26877;
											assign node26877 = (inp[10]) ? node26901 : node26878;
												assign node26878 = (inp[11]) ? node26890 : node26879;
													assign node26879 = (inp[13]) ? node26881 : 4'b0001;
														assign node26881 = (inp[14]) ? node26887 : node26882;
															assign node26882 = (inp[12]) ? node26884 : 4'b0000;
																assign node26884 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node26887 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node26890 = (inp[13]) ? node26894 : node26891;
														assign node26891 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node26894 = (inp[7]) ? node26898 : node26895;
															assign node26895 = (inp[12]) ? 4'b1001 : 4'b0001;
															assign node26898 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node26901 = (inp[13]) ? node26915 : node26902;
													assign node26902 = (inp[11]) ? node26910 : node26903;
														assign node26903 = (inp[7]) ? 4'b1001 : node26904;
															assign node26904 = (inp[14]) ? node26906 : 4'b0000;
																assign node26906 = (inp[12]) ? 4'b1001 : 4'b0001;
														assign node26910 = (inp[7]) ? node26912 : 4'b0001;
															assign node26912 = (inp[12]) ? 4'b1000 : 4'b0000;
													assign node26915 = (inp[7]) ? node26921 : node26916;
														assign node26916 = (inp[11]) ? 4'b1000 : node26917;
															assign node26917 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node26921 = (inp[11]) ? 4'b1001 : node26922;
															assign node26922 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node26926 = (inp[13]) ? node26960 : node26927;
												assign node26927 = (inp[7]) ? node26945 : node26928;
													assign node26928 = (inp[10]) ? node26940 : node26929;
														assign node26929 = (inp[12]) ? node26935 : node26930;
															assign node26930 = (inp[11]) ? 4'b0000 : node26931;
																assign node26931 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node26935 = (inp[11]) ? 4'b1001 : node26936;
																assign node26936 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node26940 = (inp[11]) ? 4'b0000 : node26941;
															assign node26941 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node26945 = (inp[11]) ? node26955 : node26946;
														assign node26946 = (inp[10]) ? node26950 : node26947;
															assign node26947 = (inp[12]) ? 4'b0000 : 4'b1000;
															assign node26950 = (inp[12]) ? node26952 : 4'b0001;
																assign node26952 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node26955 = (inp[12]) ? node26957 : 4'b1000;
															assign node26957 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node26960 = (inp[10]) ? node26976 : node26961;
													assign node26961 = (inp[14]) ? node26971 : node26962;
														assign node26962 = (inp[7]) ? node26966 : node26963;
															assign node26963 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node26966 = (inp[11]) ? node26968 : 4'b0001;
																assign node26968 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node26971 = (inp[12]) ? node26973 : 4'b0000;
															assign node26973 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node26976 = (inp[11]) ? 4'b0000 : node26977;
														assign node26977 = (inp[14]) ? node26983 : node26978;
															assign node26978 = (inp[12]) ? node26980 : 4'b0000;
																assign node26980 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node26983 = (inp[7]) ? node26987 : node26984;
																assign node26984 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node26987 = (inp[12]) ? 4'b0000 : 4'b0001;
									assign node26991 = (inp[11]) ? node27121 : node26992;
										assign node26992 = (inp[3]) ? node27058 : node26993;
											assign node26993 = (inp[14]) ? node27031 : node26994;
												assign node26994 = (inp[7]) ? node27018 : node26995;
													assign node26995 = (inp[4]) ? node27005 : node26996;
														assign node26996 = (inp[12]) ? node26998 : 4'b0100;
															assign node26998 = (inp[10]) ? node27002 : node26999;
																assign node26999 = (inp[13]) ? 4'b1000 : 4'b0000;
																assign node27002 = (inp[13]) ? 4'b0100 : 4'b1000;
														assign node27005 = (inp[13]) ? node27013 : node27006;
															assign node27006 = (inp[10]) ? node27010 : node27007;
																assign node27007 = (inp[12]) ? 4'b0100 : 4'b1100;
																assign node27010 = (inp[12]) ? 4'b1100 : 4'b0001;
															assign node27013 = (inp[10]) ? 4'b1001 : node27014;
																assign node27014 = (inp[12]) ? 4'b0001 : 4'b1001;
													assign node27018 = (inp[13]) ? node27024 : node27019;
														assign node27019 = (inp[10]) ? 4'b1000 : node27020;
															assign node27020 = (inp[12]) ? 4'b0000 : 4'b1000;
														assign node27024 = (inp[12]) ? 4'b1000 : node27025;
															assign node27025 = (inp[4]) ? node27027 : 4'b0000;
																assign node27027 = (inp[10]) ? 4'b0001 : 4'b0100;
												assign node27031 = (inp[13]) ? node27049 : node27032;
													assign node27032 = (inp[10]) ? node27038 : node27033;
														assign node27033 = (inp[4]) ? node27035 : 4'b0001;
															assign node27035 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node27038 = (inp[12]) ? node27044 : node27039;
															assign node27039 = (inp[4]) ? node27041 : 4'b1001;
																assign node27041 = (inp[7]) ? 4'b1001 : 4'b0001;
															assign node27044 = (inp[7]) ? 4'b0001 : node27045;
																assign node27045 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node27049 = (inp[10]) ? node27051 : 4'b1001;
														assign node27051 = (inp[12]) ? 4'b1001 : node27052;
															assign node27052 = (inp[7]) ? 4'b0001 : node27053;
																assign node27053 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node27058 = (inp[13]) ? node27108 : node27059;
												assign node27059 = (inp[4]) ? node27079 : node27060;
													assign node27060 = (inp[12]) ? node27070 : node27061;
														assign node27061 = (inp[7]) ? node27067 : node27062;
															assign node27062 = (inp[10]) ? node27064 : 4'b1001;
																assign node27064 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node27067 = (inp[10]) ? 4'b0001 : 4'b1001;
														assign node27070 = (inp[7]) ? node27076 : node27071;
															assign node27071 = (inp[10]) ? node27073 : 4'b0001;
																assign node27073 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node27076 = (inp[10]) ? 4'b1001 : 4'b0001;
													assign node27079 = (inp[12]) ? node27093 : node27080;
														assign node27080 = (inp[10]) ? node27086 : node27081;
															assign node27081 = (inp[7]) ? node27083 : 4'b0001;
																assign node27083 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node27086 = (inp[14]) ? node27090 : node27087;
																assign node27087 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node27090 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node27093 = (inp[14]) ? node27101 : node27094;
															assign node27094 = (inp[7]) ? node27098 : node27095;
																assign node27095 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node27098 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node27101 = (inp[7]) ? node27105 : node27102;
																assign node27102 = (inp[10]) ? 4'b1000 : 4'b0001;
																assign node27105 = (inp[10]) ? 4'b0000 : 4'b1000;
												assign node27108 = (inp[4]) ? 4'b0000 : node27109;
													assign node27109 = (inp[10]) ? node27113 : node27110;
														assign node27110 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node27113 = (inp[12]) ? node27115 : 4'b0000;
															assign node27115 = (inp[14]) ? 4'b1000 : node27116;
																assign node27116 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node27121 = (inp[13]) ? node27159 : node27122;
											assign node27122 = (inp[4]) ? node27142 : node27123;
												assign node27123 = (inp[10]) ? node27137 : node27124;
													assign node27124 = (inp[7]) ? node27132 : node27125;
														assign node27125 = (inp[12]) ? node27129 : node27126;
															assign node27126 = (inp[3]) ? 4'b0000 : 4'b1000;
															assign node27129 = (inp[3]) ? 4'b1000 : 4'b0000;
														assign node27132 = (inp[12]) ? node27134 : 4'b1000;
															assign node27134 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node27137 = (inp[3]) ? node27139 : 4'b1000;
														assign node27139 = (inp[7]) ? 4'b0000 : 4'b1000;
												assign node27142 = (inp[10]) ? node27154 : node27143;
													assign node27143 = (inp[12]) ? node27149 : node27144;
														assign node27144 = (inp[7]) ? 4'b1000 : node27145;
															assign node27145 = (inp[3]) ? 4'b0000 : 4'b1100;
														assign node27149 = (inp[7]) ? 4'b0000 : node27150;
															assign node27150 = (inp[3]) ? 4'b1000 : 4'b0100;
													assign node27154 = (inp[3]) ? 4'b0000 : node27155;
														assign node27155 = (inp[7]) ? 4'b1000 : 4'b0000;
											assign node27159 = (inp[10]) ? node27177 : node27160;
												assign node27160 = (inp[3]) ? node27170 : node27161;
													assign node27161 = (inp[12]) ? 4'b1000 : node27162;
														assign node27162 = (inp[7]) ? node27166 : node27163;
															assign node27163 = (inp[4]) ? 4'b1000 : 4'b0100;
															assign node27166 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node27170 = (inp[7]) ? node27172 : 4'b0000;
														assign node27172 = (inp[4]) ? 4'b0000 : node27173;
															assign node27173 = (inp[12]) ? 4'b0000 : 4'b1000;
												assign node27177 = (inp[3]) ? 4'b0000 : node27178;
													assign node27178 = (inp[4]) ? 4'b0000 : node27179;
														assign node27179 = (inp[7]) ? 4'b0000 : 4'b0100;
							assign node27184 = (inp[5]) ? node27186 : 4'b0000;
								assign node27186 = (inp[3]) ? node27188 : 4'b0000;
									assign node27188 = (inp[7]) ? node27268 : node27189;
										assign node27189 = (inp[4]) ? node27207 : node27190;
											assign node27190 = (inp[10]) ? node27192 : 4'b0000;
												assign node27192 = (inp[13]) ? node27194 : 4'b0000;
													assign node27194 = (inp[12]) ? 4'b0000 : node27195;
														assign node27195 = (inp[1]) ? node27201 : node27196;
															assign node27196 = (inp[14]) ? node27198 : 4'b0001;
																assign node27198 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node27201 = (inp[11]) ? 4'b0000 : node27202;
																assign node27202 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node27207 = (inp[1]) ? node27245 : node27208;
												assign node27208 = (inp[10]) ? node27224 : node27209;
													assign node27209 = (inp[13]) ? node27215 : node27210;
														assign node27210 = (inp[14]) ? node27212 : 4'b0001;
															assign node27212 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node27215 = (inp[11]) ? node27221 : node27216;
															assign node27216 = (inp[12]) ? 4'b0001 : node27217;
																assign node27217 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node27221 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node27224 = (inp[13]) ? node27236 : node27225;
														assign node27225 = (inp[12]) ? node27231 : node27226;
															assign node27226 = (inp[11]) ? 4'b0000 : node27227;
																assign node27227 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node27231 = (inp[11]) ? 4'b0001 : node27232;
																assign node27232 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node27236 = (inp[11]) ? 4'b0000 : node27237;
															assign node27237 = (inp[12]) ? node27241 : node27238;
																assign node27238 = (inp[14]) ? 4'b0001 : 4'b0000;
																assign node27241 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node27245 = (inp[11]) ? node27261 : node27246;
													assign node27246 = (inp[13]) ? node27256 : node27247;
														assign node27247 = (inp[14]) ? 4'b0001 : node27248;
															assign node27248 = (inp[10]) ? node27252 : node27249;
																assign node27249 = (inp[12]) ? 4'b0000 : 4'b1000;
																assign node27252 = (inp[12]) ? 4'b1000 : 4'b0001;
														assign node27256 = (inp[10]) ? 4'b0000 : node27257;
															assign node27257 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node27261 = (inp[10]) ? 4'b0000 : node27262;
														assign node27262 = (inp[12]) ? 4'b0000 : node27263;
															assign node27263 = (inp[13]) ? 4'b0000 : 4'b1000;
										assign node27268 = (inp[10]) ? node27270 : 4'b0000;
											assign node27270 = (inp[13]) ? node27272 : 4'b0000;
												assign node27272 = (inp[1]) ? 4'b0000 : node27273;
													assign node27273 = (inp[4]) ? node27275 : 4'b0000;
														assign node27275 = (inp[14]) ? 4'b0000 : node27276;
															assign node27276 = (inp[11]) ? 4'b0000 : node27277;
																assign node27277 = (inp[12]) ? 4'b0000 : 4'b0001;

endmodule