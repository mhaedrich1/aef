module dtc_split75_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node685;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node720;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node860;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node873;
	wire [3-1:0] node875;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node944;
	wire [3-1:0] node946;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node981;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1015;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1101;
	wire [3-1:0] node1104;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1111;
	wire [3-1:0] node1114;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1121;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1143;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1155;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1210;
	wire [3-1:0] node1212;
	wire [3-1:0] node1213;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1230;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1248;
	wire [3-1:0] node1251;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1282;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1294;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1321;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1329;
	wire [3-1:0] node1331;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1356;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1367;
	wire [3-1:0] node1370;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1384;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1389;
	wire [3-1:0] node1392;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1400;
	wire [3-1:0] node1403;
	wire [3-1:0] node1404;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1417;
	wire [3-1:0] node1423;
	wire [3-1:0] node1425;
	wire [3-1:0] node1426;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1436;
	wire [3-1:0] node1439;
	wire [3-1:0] node1441;
	wire [3-1:0] node1445;
	wire [3-1:0] node1446;
	wire [3-1:0] node1448;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1461;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1472;
	wire [3-1:0] node1474;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1480;
	wire [3-1:0] node1481;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1501;
	wire [3-1:0] node1504;
	wire [3-1:0] node1505;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1514;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1519;
	wire [3-1:0] node1520;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1535;
	wire [3-1:0] node1536;
	wire [3-1:0] node1539;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1547;
	wire [3-1:0] node1548;
	wire [3-1:0] node1551;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1584;
	wire [3-1:0] node1587;
	wire [3-1:0] node1588;
	wire [3-1:0] node1590;
	wire [3-1:0] node1593;
	wire [3-1:0] node1596;
	wire [3-1:0] node1597;
	wire [3-1:0] node1598;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1604;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1614;
	wire [3-1:0] node1615;
	wire [3-1:0] node1619;
	wire [3-1:0] node1620;
	wire [3-1:0] node1621;
	wire [3-1:0] node1622;
	wire [3-1:0] node1626;
	wire [3-1:0] node1627;
	wire [3-1:0] node1632;
	wire [3-1:0] node1633;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1647;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1654;
	wire [3-1:0] node1657;
	wire [3-1:0] node1659;
	wire [3-1:0] node1662;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1677;
	wire [3-1:0] node1678;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1690;
	wire [3-1:0] node1693;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1704;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1709;
	wire [3-1:0] node1711;
	wire [3-1:0] node1712;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1720;
	wire [3-1:0] node1723;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1728;
	wire [3-1:0] node1729;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1742;
	wire [3-1:0] node1743;
	wire [3-1:0] node1745;
	wire [3-1:0] node1747;
	wire [3-1:0] node1750;
	wire [3-1:0] node1751;
	wire [3-1:0] node1754;
	wire [3-1:0] node1757;
	wire [3-1:0] node1758;
	wire [3-1:0] node1759;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1767;
	wire [3-1:0] node1770;
	wire [3-1:0] node1771;
	wire [3-1:0] node1772;
	wire [3-1:0] node1774;
	wire [3-1:0] node1777;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1790;
	wire [3-1:0] node1791;
	wire [3-1:0] node1792;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1799;
	wire [3-1:0] node1800;
	wire [3-1:0] node1801;
	wire [3-1:0] node1803;
	wire [3-1:0] node1805;
	wire [3-1:0] node1808;
	wire [3-1:0] node1809;
	wire [3-1:0] node1810;
	wire [3-1:0] node1814;
	wire [3-1:0] node1816;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1825;
	wire [3-1:0] node1828;
	wire [3-1:0] node1831;
	wire [3-1:0] node1833;
	wire [3-1:0] node1836;
	wire [3-1:0] node1838;
	wire [3-1:0] node1840;
	wire [3-1:0] node1841;
	wire [3-1:0] node1845;
	wire [3-1:0] node1846;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1852;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1857;
	wire [3-1:0] node1860;
	wire [3-1:0] node1863;
	wire [3-1:0] node1866;
	wire [3-1:0] node1867;
	wire [3-1:0] node1868;
	wire [3-1:0] node1872;
	wire [3-1:0] node1873;
	wire [3-1:0] node1874;
	wire [3-1:0] node1878;
	wire [3-1:0] node1881;
	wire [3-1:0] node1882;
	wire [3-1:0] node1883;
	wire [3-1:0] node1884;
	wire [3-1:0] node1886;
	wire [3-1:0] node1889;
	wire [3-1:0] node1891;
	wire [3-1:0] node1894;
	wire [3-1:0] node1896;
	wire [3-1:0] node1897;
	wire [3-1:0] node1901;
	wire [3-1:0] node1902;
	wire [3-1:0] node1903;
	wire [3-1:0] node1904;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1912;
	wire [3-1:0] node1915;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1924;
	wire [3-1:0] node1925;
	wire [3-1:0] node1926;
	wire [3-1:0] node1927;
	wire [3-1:0] node1928;
	wire [3-1:0] node1929;
	wire [3-1:0] node1930;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1935;
	wire [3-1:0] node1936;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1943;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1951;
	wire [3-1:0] node1953;
	wire [3-1:0] node1956;
	wire [3-1:0] node1957;
	wire [3-1:0] node1958;
	wire [3-1:0] node1959;
	wire [3-1:0] node1963;
	wire [3-1:0] node1964;
	wire [3-1:0] node1968;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1973;
	wire [3-1:0] node1974;
	wire [3-1:0] node1978;
	wire [3-1:0] node1980;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1985;
	wire [3-1:0] node1986;
	wire [3-1:0] node1987;
	wire [3-1:0] node1990;
	wire [3-1:0] node1993;
	wire [3-1:0] node1994;
	wire [3-1:0] node1999;
	wire [3-1:0] node2001;
	wire [3-1:0] node2002;
	wire [3-1:0] node2003;
	wire [3-1:0] node2006;
	wire [3-1:0] node2009;
	wire [3-1:0] node2012;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2015;
	wire [3-1:0] node2016;
	wire [3-1:0] node2017;
	wire [3-1:0] node2020;
	wire [3-1:0] node2022;
	wire [3-1:0] node2025;
	wire [3-1:0] node2027;
	wire [3-1:0] node2030;
	wire [3-1:0] node2031;
	wire [3-1:0] node2033;
	wire [3-1:0] node2035;
	wire [3-1:0] node2038;
	wire [3-1:0] node2039;
	wire [3-1:0] node2042;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2047;
	wire [3-1:0] node2048;
	wire [3-1:0] node2052;
	wire [3-1:0] node2053;
	wire [3-1:0] node2055;
	wire [3-1:0] node2059;
	wire [3-1:0] node2060;
	wire [3-1:0] node2061;
	wire [3-1:0] node2064;
	wire [3-1:0] node2066;
	wire [3-1:0] node2069;
	wire [3-1:0] node2070;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2076;
	wire [3-1:0] node2077;
	wire [3-1:0] node2079;
	wire [3-1:0] node2081;
	wire [3-1:0] node2084;
	wire [3-1:0] node2087;
	wire [3-1:0] node2088;
	wire [3-1:0] node2089;
	wire [3-1:0] node2091;
	wire [3-1:0] node2094;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2102;
	wire [3-1:0] node2106;
	wire [3-1:0] node2107;
	wire [3-1:0] node2109;
	wire [3-1:0] node2110;
	wire [3-1:0] node2111;
	wire [3-1:0] node2117;
	wire [3-1:0] node2118;
	wire [3-1:0] node2119;
	wire [3-1:0] node2120;
	wire [3-1:0] node2121;
	wire [3-1:0] node2123;
	wire [3-1:0] node2124;
	wire [3-1:0] node2129;
	wire [3-1:0] node2130;
	wire [3-1:0] node2132;
	wire [3-1:0] node2134;
	wire [3-1:0] node2136;
	wire [3-1:0] node2139;
	wire [3-1:0] node2140;
	wire [3-1:0] node2142;
	wire [3-1:0] node2145;
	wire [3-1:0] node2146;
	wire [3-1:0] node2149;
	wire [3-1:0] node2152;
	wire [3-1:0] node2153;
	wire [3-1:0] node2155;
	wire [3-1:0] node2156;
	wire [3-1:0] node2158;
	wire [3-1:0] node2160;
	wire [3-1:0] node2163;
	wire [3-1:0] node2167;
	wire [3-1:0] node2168;
	wire [3-1:0] node2169;
	wire [3-1:0] node2171;
	wire [3-1:0] node2172;
	wire [3-1:0] node2174;
	wire [3-1:0] node2177;
	wire [3-1:0] node2179;
	wire [3-1:0] node2182;
	wire [3-1:0] node2183;
	wire [3-1:0] node2184;
	wire [3-1:0] node2186;
	wire [3-1:0] node2189;
	wire [3-1:0] node2191;
	wire [3-1:0] node2192;
	wire [3-1:0] node2196;
	wire [3-1:0] node2197;
	wire [3-1:0] node2199;
	wire [3-1:0] node2202;
	wire [3-1:0] node2203;
	wire [3-1:0] node2204;
	wire [3-1:0] node2207;
	wire [3-1:0] node2211;
	wire [3-1:0] node2212;
	wire [3-1:0] node2213;
	wire [3-1:0] node2214;
	wire [3-1:0] node2215;
	wire [3-1:0] node2218;
	wire [3-1:0] node2221;
	wire [3-1:0] node2223;
	wire [3-1:0] node2226;
	wire [3-1:0] node2227;
	wire [3-1:0] node2228;
	wire [3-1:0] node2229;
	wire [3-1:0] node2233;
	wire [3-1:0] node2236;
	wire [3-1:0] node2237;
	wire [3-1:0] node2240;
	wire [3-1:0] node2242;
	wire [3-1:0] node2245;
	wire [3-1:0] node2246;
	wire [3-1:0] node2247;
	wire [3-1:0] node2248;
	wire [3-1:0] node2250;
	wire [3-1:0] node2253;
	wire [3-1:0] node2256;
	wire [3-1:0] node2259;
	wire [3-1:0] node2260;
	wire [3-1:0] node2261;
	wire [3-1:0] node2265;
	wire [3-1:0] node2266;
	wire [3-1:0] node2268;
	wire [3-1:0] node2272;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2275;
	wire [3-1:0] node2276;
	wire [3-1:0] node2277;
	wire [3-1:0] node2278;
	wire [3-1:0] node2283;
	wire [3-1:0] node2285;
	wire [3-1:0] node2286;
	wire [3-1:0] node2288;
	wire [3-1:0] node2289;
	wire [3-1:0] node2294;
	wire [3-1:0] node2295;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2302;
	wire [3-1:0] node2303;
	wire [3-1:0] node2305;
	wire [3-1:0] node2308;
	wire [3-1:0] node2309;
	wire [3-1:0] node2310;
	wire [3-1:0] node2315;
	wire [3-1:0] node2317;
	wire [3-1:0] node2319;
	wire [3-1:0] node2320;
	wire [3-1:0] node2321;
	wire [3-1:0] node2323;
	wire [3-1:0] node2324;
	wire [3-1:0] node2330;
	wire [3-1:0] node2331;
	wire [3-1:0] node2332;
	wire [3-1:0] node2334;
	wire [3-1:0] node2336;
	wire [3-1:0] node2337;
	wire [3-1:0] node2341;
	wire [3-1:0] node2342;
	wire [3-1:0] node2343;
	wire [3-1:0] node2344;
	wire [3-1:0] node2345;
	wire [3-1:0] node2349;
	wire [3-1:0] node2352;
	wire [3-1:0] node2353;
	wire [3-1:0] node2354;
	wire [3-1:0] node2358;
	wire [3-1:0] node2359;
	wire [3-1:0] node2362;
	wire [3-1:0] node2364;
	wire [3-1:0] node2367;
	wire [3-1:0] node2369;
	wire [3-1:0] node2370;
	wire [3-1:0] node2372;
	wire [3-1:0] node2374;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2380;
	wire [3-1:0] node2381;
	wire [3-1:0] node2382;
	wire [3-1:0] node2385;
	wire [3-1:0] node2388;
	wire [3-1:0] node2389;
	wire [3-1:0] node2390;
	wire [3-1:0] node2392;
	wire [3-1:0] node2396;
	wire [3-1:0] node2397;
	wire [3-1:0] node2398;
	wire [3-1:0] node2402;
	wire [3-1:0] node2403;
	wire [3-1:0] node2406;
	wire [3-1:0] node2409;
	wire [3-1:0] node2410;
	wire [3-1:0] node2411;
	wire [3-1:0] node2412;
	wire [3-1:0] node2413;
	wire [3-1:0] node2417;
	wire [3-1:0] node2418;
	wire [3-1:0] node2422;
	wire [3-1:0] node2423;
	wire [3-1:0] node2424;
	wire [3-1:0] node2427;
	wire [3-1:0] node2431;
	wire [3-1:0] node2432;
	wire [3-1:0] node2433;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2441;
	wire [3-1:0] node2442;
	wire [3-1:0] node2443;
	wire [3-1:0] node2446;
	wire [3-1:0] node2450;
	wire [3-1:0] node2451;
	wire [3-1:0] node2452;
	wire [3-1:0] node2453;
	wire [3-1:0] node2457;
	wire [3-1:0] node2458;
	wire [3-1:0] node2460;
	wire [3-1:0] node2461;
	wire [3-1:0] node2464;
	wire [3-1:0] node2467;
	wire [3-1:0] node2468;
	wire [3-1:0] node2472;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2475;
	wire [3-1:0] node2477;
	wire [3-1:0] node2480;
	wire [3-1:0] node2481;
	wire [3-1:0] node2485;
	wire [3-1:0] node2487;
	wire [3-1:0] node2488;
	wire [3-1:0] node2492;
	wire [3-1:0] node2493;
	wire [3-1:0] node2494;
	wire [3-1:0] node2495;
	wire [3-1:0] node2498;
	wire [3-1:0] node2502;
	wire [3-1:0] node2504;
	wire [3-1:0] node2505;

	assign outp = (inp[0]) ? node1068 : node1;
		assign node1 = (inp[6]) ? node81 : node2;
			assign node2 = (inp[3]) ? node14 : node3;
				assign node3 = (inp[4]) ? node5 : 3'b011;
					assign node5 = (inp[7]) ? node7 : 3'b011;
						assign node7 = (inp[8]) ? node9 : 3'b111;
							assign node9 = (inp[1]) ? node11 : 3'b111;
								assign node11 = (inp[2]) ? 3'b011 : 3'b111;
				assign node14 = (inp[7]) ? node16 : 3'b111;
					assign node16 = (inp[9]) ? 3'b111 : node17;
						assign node17 = (inp[1]) ? node25 : node18;
							assign node18 = (inp[2]) ? node20 : 3'b111;
								assign node20 = (inp[8]) ? node22 : 3'b111;
									assign node22 = (inp[4]) ? 3'b111 : 3'b011;
							assign node25 = (inp[4]) ? node67 : node26;
								assign node26 = (inp[5]) ? node52 : node27;
									assign node27 = (inp[11]) ? node41 : node28;
										assign node28 = (inp[10]) ? node36 : node29;
											assign node29 = (inp[8]) ? node33 : node30;
												assign node30 = (inp[2]) ? 3'b001 : 3'b101;
												assign node33 = (inp[2]) ? 3'b101 : 3'b001;
											assign node36 = (inp[8]) ? node38 : 3'b001;
												assign node38 = (inp[2]) ? 3'b001 : 3'b101;
										assign node41 = (inp[2]) ? node47 : node42;
											assign node42 = (inp[10]) ? 3'b001 : node43;
												assign node43 = (inp[8]) ? 3'b001 : 3'b101;
											assign node47 = (inp[10]) ? 3'b101 : node48;
												assign node48 = (inp[8]) ? 3'b101 : 3'b001;
									assign node52 = (inp[8]) ? node60 : node53;
										assign node53 = (inp[2]) ? node57 : node54;
											assign node54 = (inp[10]) ? 3'b111 : 3'b011;
											assign node57 = (inp[10]) ? 3'b001 : 3'b101;
										assign node60 = (inp[10]) ? node64 : node61;
											assign node61 = (inp[2]) ? 3'b001 : 3'b101;
											assign node64 = (inp[2]) ? 3'b101 : 3'b001;
								assign node67 = (inp[2]) ? node73 : node68;
									assign node68 = (inp[8]) ? node70 : 3'b111;
										assign node70 = (inp[5]) ? 3'b111 : 3'b011;
									assign node73 = (inp[5]) ? node77 : node74;
										assign node74 = (inp[8]) ? 3'b101 : 3'b011;
										assign node77 = (inp[8]) ? 3'b011 : 3'b111;
			assign node81 = (inp[7]) ? node571 : node82;
				assign node82 = (inp[3]) ? node336 : node83;
					assign node83 = (inp[4]) ? node223 : node84;
						assign node84 = (inp[1]) ? node160 : node85;
							assign node85 = (inp[9]) ? node115 : node86;
								assign node86 = (inp[5]) ? node100 : node87;
									assign node87 = (inp[8]) ? 3'b101 : node88;
										assign node88 = (inp[11]) ? node94 : node89;
											assign node89 = (inp[2]) ? 3'b001 : node90;
												assign node90 = (inp[10]) ? 3'b001 : 3'b101;
											assign node94 = (inp[2]) ? 3'b101 : node95;
												assign node95 = (inp[10]) ? 3'b101 : 3'b001;
									assign node100 = (inp[8]) ? node106 : node101;
										assign node101 = (inp[2]) ? node103 : 3'b101;
											assign node103 = (inp[10]) ? 3'b001 : 3'b101;
										assign node106 = (inp[11]) ? 3'b001 : node107;
											assign node107 = (inp[2]) ? node111 : node108;
												assign node108 = (inp[10]) ? 3'b001 : 3'b101;
												assign node111 = (inp[10]) ? 3'b101 : 3'b001;
								assign node115 = (inp[10]) ? node139 : node116;
									assign node116 = (inp[11]) ? node130 : node117;
										assign node117 = (inp[5]) ? node123 : node118;
											assign node118 = (inp[8]) ? 3'b001 : node119;
												assign node119 = (inp[2]) ? 3'b001 : 3'b101;
											assign node123 = (inp[8]) ? node127 : node124;
												assign node124 = (inp[2]) ? 3'b101 : 3'b001;
												assign node127 = (inp[2]) ? 3'b001 : 3'b101;
										assign node130 = (inp[2]) ? node134 : node131;
											assign node131 = (inp[5]) ? 3'b001 : 3'b101;
											assign node134 = (inp[8]) ? node136 : 3'b101;
												assign node136 = (inp[5]) ? 3'b101 : 3'b001;
									assign node139 = (inp[8]) ? node147 : node140;
										assign node140 = (inp[5]) ? 3'b001 : node141;
											assign node141 = (inp[2]) ? node143 : 3'b001;
												assign node143 = (inp[11]) ? 3'b001 : 3'b101;
										assign node147 = (inp[11]) ? node155 : node148;
											assign node148 = (inp[2]) ? node152 : node149;
												assign node149 = (inp[5]) ? 3'b001 : 3'b101;
												assign node152 = (inp[5]) ? 3'b101 : 3'b001;
											assign node155 = (inp[5]) ? 3'b001 : node156;
												assign node156 = (inp[2]) ? 3'b101 : 3'b001;
							assign node160 = (inp[8]) ? node190 : node161;
								assign node161 = (inp[11]) ? node177 : node162;
									assign node162 = (inp[9]) ? 3'b101 : node163;
										assign node163 = (inp[2]) ? node169 : node164;
											assign node164 = (inp[10]) ? node166 : 3'b101;
												assign node166 = (inp[5]) ? 3'b101 : 3'b001;
											assign node169 = (inp[10]) ? node173 : node170;
												assign node170 = (inp[5]) ? 3'b101 : 3'b001;
												assign node173 = (inp[5]) ? 3'b001 : 3'b101;
									assign node177 = (inp[10]) ? node183 : node178;
										assign node178 = (inp[2]) ? node180 : 3'b001;
											assign node180 = (inp[5]) ? 3'b101 : 3'b001;
										assign node183 = (inp[2]) ? node185 : 3'b101;
											assign node185 = (inp[9]) ? 3'b001 : node186;
												assign node186 = (inp[5]) ? 3'b001 : 3'b101;
								assign node190 = (inp[2]) ? node210 : node191;
									assign node191 = (inp[10]) ? node205 : node192;
										assign node192 = (inp[9]) ? node200 : node193;
											assign node193 = (inp[5]) ? node197 : node194;
												assign node194 = (inp[11]) ? 3'b101 : 3'b001;
												assign node197 = (inp[11]) ? 3'b001 : 3'b101;
											assign node200 = (inp[11]) ? 3'b101 : node201;
												assign node201 = (inp[5]) ? 3'b101 : 3'b001;
										assign node205 = (inp[11]) ? 3'b001 : node206;
											assign node206 = (inp[5]) ? 3'b001 : 3'b101;
									assign node210 = (inp[10]) ? node218 : node211;
										assign node211 = (inp[5]) ? 3'b010 : node212;
											assign node212 = (inp[11]) ? node214 : 3'b110;
												assign node214 = (inp[9]) ? 3'b010 : 3'b110;
										assign node218 = (inp[11]) ? 3'b110 : node219;
											assign node219 = (inp[5]) ? 3'b110 : 3'b010;
						assign node223 = (inp[9]) ? node285 : node224;
							assign node224 = (inp[1]) ? node254 : node225;
								assign node225 = (inp[2]) ? node241 : node226;
									assign node226 = (inp[8]) ? node236 : node227;
										assign node227 = (inp[11]) ? node229 : 3'b101;
											assign node229 = (inp[10]) ? node233 : node230;
												assign node230 = (inp[5]) ? 3'b011 : 3'b001;
												assign node233 = (inp[5]) ? 3'b111 : 3'b101;
										assign node236 = (inp[10]) ? 3'b001 : node237;
											assign node237 = (inp[5]) ? 3'b101 : 3'b001;
									assign node241 = (inp[8]) ? node247 : node242;
										assign node242 = (inp[5]) ? node244 : 3'b001;
											assign node244 = (inp[10]) ? 3'b011 : 3'b001;
										assign node247 = (inp[10]) ? 3'b101 : node248;
											assign node248 = (inp[5]) ? 3'b001 : node249;
												assign node249 = (inp[11]) ? 3'b011 : 3'b111;
								assign node254 = (inp[10]) ? node268 : node255;
									assign node255 = (inp[5]) ? node261 : node256;
										assign node256 = (inp[8]) ? 3'b011 : node257;
											assign node257 = (inp[2]) ? 3'b011 : 3'b111;
										assign node261 = (inp[8]) ? node265 : node262;
											assign node262 = (inp[2]) ? 3'b011 : 3'b111;
											assign node265 = (inp[2]) ? 3'b101 : 3'b111;
									assign node268 = (inp[8]) ? node278 : node269;
										assign node269 = (inp[2]) ? node271 : 3'b001;
											assign node271 = (inp[5]) ? node275 : node272;
												assign node272 = (inp[11]) ? 3'b101 : 3'b001;
												assign node275 = (inp[11]) ? 3'b001 : 3'b101;
										assign node278 = (inp[11]) ? node280 : 3'b011;
											assign node280 = (inp[5]) ? node282 : 3'b011;
												assign node282 = (inp[2]) ? 3'b111 : 3'b001;
							assign node285 = (inp[1]) ? node295 : node286;
								assign node286 = (inp[2]) ? node288 : 3'b111;
									assign node288 = (inp[10]) ? node290 : 3'b011;
										assign node290 = (inp[5]) ? 3'b111 : node291;
											assign node291 = (inp[8]) ? 3'b011 : 3'b111;
								assign node295 = (inp[2]) ? node313 : node296;
									assign node296 = (inp[10]) ? node306 : node297;
										assign node297 = (inp[8]) ? node301 : node298;
											assign node298 = (inp[5]) ? 3'b101 : 3'b001;
											assign node301 = (inp[5]) ? node303 : 3'b111;
												assign node303 = (inp[11]) ? 3'b001 : 3'b011;
										assign node306 = (inp[11]) ? node308 : 3'b111;
											assign node308 = (inp[5]) ? node310 : 3'b011;
												assign node310 = (inp[8]) ? 3'b011 : 3'b111;
									assign node313 = (inp[10]) ? node325 : node314;
										assign node314 = (inp[8]) ? node318 : node315;
											assign node315 = (inp[5]) ? 3'b101 : 3'b001;
											assign node318 = (inp[11]) ? node322 : node319;
												assign node319 = (inp[5]) ? 3'b111 : 3'b101;
												assign node322 = (inp[5]) ? 3'b001 : 3'b111;
										assign node325 = (inp[8]) ? node331 : node326;
											assign node326 = (inp[11]) ? node328 : 3'b101;
												assign node328 = (inp[5]) ? 3'b011 : 3'b101;
											assign node331 = (inp[11]) ? node333 : 3'b001;
												assign node333 = (inp[5]) ? 3'b101 : 3'b001;
					assign node336 = (inp[1]) ? node416 : node337;
						assign node337 = (inp[5]) ? node377 : node338;
							assign node338 = (inp[8]) ? node358 : node339;
								assign node339 = (inp[2]) ? node341 : 3'b111;
									assign node341 = (inp[11]) ? node351 : node342;
										assign node342 = (inp[10]) ? node346 : node343;
											assign node343 = (inp[4]) ? 3'b011 : 3'b101;
											assign node346 = (inp[4]) ? 3'b111 : node347;
												assign node347 = (inp[9]) ? 3'b111 : 3'b011;
										assign node351 = (inp[9]) ? 3'b111 : node352;
											assign node352 = (inp[10]) ? 3'b111 : node353;
												assign node353 = (inp[4]) ? 3'b111 : 3'b011;
								assign node358 = (inp[4]) ? node370 : node359;
									assign node359 = (inp[11]) ? node367 : node360;
										assign node360 = (inp[2]) ? 3'b111 : node361;
											assign node361 = (inp[9]) ? 3'b111 : node362;
												assign node362 = (inp[10]) ? 3'b011 : 3'b111;
										assign node367 = (inp[10]) ? 3'b011 : 3'b101;
									assign node370 = (inp[11]) ? node372 : 3'b101;
										assign node372 = (inp[10]) ? 3'b101 : node373;
											assign node373 = (inp[2]) ? 3'b001 : 3'b101;
							assign node377 = (inp[9]) ? node407 : node378;
								assign node378 = (inp[4]) ? node400 : node379;
									assign node379 = (inp[2]) ? node389 : node380;
										assign node380 = (inp[10]) ? node386 : node381;
											assign node381 = (inp[11]) ? 3'b111 : node382;
												assign node382 = (inp[8]) ? 3'b011 : 3'b111;
											assign node386 = (inp[11]) ? 3'b011 : 3'b111;
										assign node389 = (inp[10]) ? node395 : node390;
											assign node390 = (inp[8]) ? node392 : 3'b011;
												assign node392 = (inp[11]) ? 3'b011 : 3'b101;
											assign node395 = (inp[8]) ? node397 : 3'b111;
												assign node397 = (inp[11]) ? 3'b111 : 3'b011;
									assign node400 = (inp[10]) ? 3'b111 : node401;
										assign node401 = (inp[11]) ? 3'b111 : node402;
											assign node402 = (inp[8]) ? 3'b011 : 3'b111;
								assign node407 = (inp[8]) ? node409 : 3'b111;
									assign node409 = (inp[11]) ? 3'b111 : node410;
										assign node410 = (inp[10]) ? 3'b111 : node411;
											assign node411 = (inp[2]) ? 3'b011 : 3'b111;
						assign node416 = (inp[9]) ? node492 : node417;
							assign node417 = (inp[5]) ? node457 : node418;
								assign node418 = (inp[8]) ? node436 : node419;
									assign node419 = (inp[4]) ? node429 : node420;
										assign node420 = (inp[11]) ? node424 : node421;
											assign node421 = (inp[2]) ? 3'b110 : 3'b101;
											assign node424 = (inp[2]) ? 3'b001 : node425;
												assign node425 = (inp[10]) ? 3'b110 : 3'b001;
										assign node429 = (inp[2]) ? node433 : node430;
											assign node430 = (inp[10]) ? 3'b001 : 3'b101;
											assign node433 = (inp[10]) ? 3'b101 : 3'b001;
									assign node436 = (inp[2]) ? node446 : node437;
										assign node437 = (inp[4]) ? node441 : node438;
											assign node438 = (inp[10]) ? 3'b010 : 3'b110;
											assign node441 = (inp[11]) ? 3'b001 : node442;
												assign node442 = (inp[10]) ? 3'b101 : 3'b001;
										assign node446 = (inp[4]) ? node452 : node447;
											assign node447 = (inp[10]) ? node449 : 3'b010;
												assign node449 = (inp[11]) ? 3'b001 : 3'b110;
											assign node452 = (inp[11]) ? 3'b110 : node453;
												assign node453 = (inp[10]) ? 3'b010 : 3'b110;
								assign node457 = (inp[2]) ? node473 : node458;
									assign node458 = (inp[4]) ? node468 : node459;
										assign node459 = (inp[10]) ? node463 : node460;
											assign node460 = (inp[8]) ? 3'b001 : 3'b101;
											assign node463 = (inp[8]) ? node465 : 3'b010;
												assign node465 = (inp[11]) ? 3'b110 : 3'b101;
										assign node468 = (inp[8]) ? 3'b001 : node469;
											assign node469 = (inp[10]) ? 3'b111 : 3'b011;
									assign node473 = (inp[10]) ? node487 : node474;
										assign node474 = (inp[11]) ? node480 : node475;
											assign node475 = (inp[8]) ? 3'b001 : node476;
												assign node476 = (inp[4]) ? 3'b101 : 3'b001;
											assign node480 = (inp[8]) ? node484 : node481;
												assign node481 = (inp[4]) ? 3'b101 : 3'b001;
												assign node484 = (inp[4]) ? 3'b001 : 3'b101;
										assign node487 = (inp[4]) ? 3'b101 : node488;
											assign node488 = (inp[8]) ? 3'b001 : 3'b101;
							assign node492 = (inp[4]) ? node532 : node493;
								assign node493 = (inp[8]) ? node511 : node494;
									assign node494 = (inp[2]) ? node500 : node495;
										assign node495 = (inp[5]) ? 3'b111 : node496;
											assign node496 = (inp[10]) ? 3'b111 : 3'b101;
										assign node500 = (inp[5]) ? node508 : node501;
											assign node501 = (inp[11]) ? node505 : node502;
												assign node502 = (inp[10]) ? 3'b001 : 3'b011;
												assign node505 = (inp[10]) ? 3'b011 : 3'b001;
											assign node508 = (inp[10]) ? 3'b111 : 3'b101;
									assign node511 = (inp[10]) ? node525 : node512;
										assign node512 = (inp[2]) ? node520 : node513;
											assign node513 = (inp[5]) ? node517 : node514;
												assign node514 = (inp[11]) ? 3'b001 : 3'b011;
												assign node517 = (inp[11]) ? 3'b111 : 3'b101;
											assign node520 = (inp[5]) ? node522 : 3'b101;
												assign node522 = (inp[11]) ? 3'b001 : 3'b011;
										assign node525 = (inp[11]) ? 3'b011 : node526;
											assign node526 = (inp[5]) ? 3'b001 : node527;
												assign node527 = (inp[2]) ? 3'b111 : 3'b001;
								assign node532 = (inp[10]) ? node554 : node533;
									assign node533 = (inp[8]) ? node539 : node534;
										assign node534 = (inp[2]) ? 3'b011 : node535;
											assign node535 = (inp[5]) ? 3'b011 : 3'b111;
										assign node539 = (inp[11]) ? node547 : node540;
											assign node540 = (inp[2]) ? node544 : node541;
												assign node541 = (inp[5]) ? 3'b111 : 3'b011;
												assign node544 = (inp[5]) ? 3'b011 : 3'b111;
											assign node547 = (inp[5]) ? node551 : node548;
												assign node548 = (inp[2]) ? 3'b111 : 3'b011;
												assign node551 = (inp[2]) ? 3'b011 : 3'b111;
									assign node554 = (inp[2]) ? node562 : node555;
										assign node555 = (inp[8]) ? node559 : node556;
											assign node556 = (inp[5]) ? 3'b101 : 3'b001;
											assign node559 = (inp[11]) ? 3'b001 : 3'b011;
										assign node562 = (inp[11]) ? node568 : node563;
											assign node563 = (inp[5]) ? node565 : 3'b011;
												assign node565 = (inp[8]) ? 3'b111 : 3'b011;
											assign node568 = (inp[5]) ? 3'b011 : 3'b111;
				assign node571 = (inp[3]) ? node797 : node572;
					assign node572 = (inp[9]) ? node666 : node573;
						assign node573 = (inp[4]) ? node603 : node574;
							assign node574 = (inp[1]) ? 3'b000 : node575;
								assign node575 = (inp[11]) ? node585 : node576;
									assign node576 = (inp[8]) ? node582 : node577;
										assign node577 = (inp[5]) ? node579 : 3'b100;
											assign node579 = (inp[2]) ? 3'b100 : 3'b000;
										assign node582 = (inp[5]) ? 3'b100 : 3'b000;
									assign node585 = (inp[2]) ? node593 : node586;
										assign node586 = (inp[5]) ? node590 : node587;
											assign node587 = (inp[8]) ? 3'b000 : 3'b100;
											assign node590 = (inp[10]) ? 3'b100 : 3'b000;
										assign node593 = (inp[8]) ? node595 : 3'b000;
											assign node595 = (inp[10]) ? node599 : node596;
												assign node596 = (inp[5]) ? 3'b100 : 3'b000;
												assign node599 = (inp[5]) ? 3'b000 : 3'b100;
							assign node603 = (inp[1]) ? node645 : node604;
								assign node604 = (inp[2]) ? node624 : node605;
									assign node605 = (inp[10]) ? node615 : node606;
										assign node606 = (inp[8]) ? node610 : node607;
											assign node607 = (inp[5]) ? 3'b011 : 3'b111;
											assign node610 = (inp[11]) ? 3'b111 : node611;
												assign node611 = (inp[5]) ? 3'b110 : 3'b010;
										assign node615 = (inp[11]) ? 3'b011 : node616;
											assign node616 = (inp[8]) ? node620 : node617;
												assign node617 = (inp[5]) ? 3'b101 : 3'b001;
												assign node620 = (inp[5]) ? 3'b001 : 3'b111;
									assign node624 = (inp[10]) ? node632 : node625;
										assign node625 = (inp[8]) ? node629 : node626;
											assign node626 = (inp[5]) ? 3'b110 : 3'b010;
											assign node629 = (inp[5]) ? 3'b010 : 3'b100;
										assign node632 = (inp[11]) ? node638 : node633;
											assign node633 = (inp[5]) ? 3'b110 : node634;
												assign node634 = (inp[8]) ? 3'b010 : 3'b110;
											assign node638 = (inp[8]) ? node642 : node639;
												assign node639 = (inp[5]) ? 3'b001 : 3'b111;
												assign node642 = (inp[5]) ? 3'b111 : 3'b110;
								assign node645 = (inp[10]) ? node655 : node646;
									assign node646 = (inp[2]) ? 3'b000 : node647;
										assign node647 = (inp[11]) ? 3'b000 : node648;
											assign node648 = (inp[5]) ? node650 : 3'b100;
												assign node650 = (inp[8]) ? 3'b100 : 3'b000;
									assign node655 = (inp[5]) ? node657 : 3'b100;
										assign node657 = (inp[2]) ? node663 : node658;
											assign node658 = (inp[8]) ? node660 : 3'b010;
												assign node660 = (inp[11]) ? 3'b010 : 3'b100;
											assign node663 = (inp[8]) ? 3'b100 : 3'b000;
						assign node666 = (inp[1]) ? node738 : node667;
							assign node667 = (inp[4]) ? node709 : node668;
								assign node668 = (inp[10]) ? node690 : node669;
									assign node669 = (inp[2]) ? node679 : node670;
										assign node670 = (inp[5]) ? node676 : node671;
											assign node671 = (inp[8]) ? 3'b000 : node672;
												assign node672 = (inp[11]) ? 3'b101 : 3'b100;
											assign node676 = (inp[8]) ? 3'b101 : 3'b011;
										assign node679 = (inp[8]) ? node685 : node680;
											assign node680 = (inp[11]) ? 3'b100 : node681;
												assign node681 = (inp[5]) ? 3'b100 : 3'b000;
											assign node685 = (inp[5]) ? node687 : 3'b010;
												assign node687 = (inp[11]) ? 3'b100 : 3'b000;
									assign node690 = (inp[5]) ? node700 : node691;
										assign node691 = (inp[2]) ? node695 : node692;
											assign node692 = (inp[8]) ? 3'b001 : 3'b101;
											assign node695 = (inp[8]) ? 3'b110 : node696;
												assign node696 = (inp[11]) ? 3'b001 : 3'b100;
										assign node700 = (inp[2]) ? node704 : node701;
											assign node701 = (inp[8]) ? 3'b101 : 3'b011;
											assign node704 = (inp[11]) ? node706 : 3'b001;
												assign node706 = (inp[8]) ? 3'b001 : 3'b101;
								assign node709 = (inp[5]) ? node725 : node710;
									assign node710 = (inp[2]) ? node718 : node711;
										assign node711 = (inp[8]) ? node713 : 3'b101;
											assign node713 = (inp[10]) ? 3'b101 : node714;
												assign node714 = (inp[11]) ? 3'b101 : 3'b001;
										assign node718 = (inp[8]) ? node720 : 3'b001;
											assign node720 = (inp[10]) ? node722 : 3'b101;
												assign node722 = (inp[11]) ? 3'b101 : 3'b001;
									assign node725 = (inp[10]) ? node733 : node726;
										assign node726 = (inp[8]) ? node730 : node727;
											assign node727 = (inp[2]) ? 3'b111 : 3'b001;
											assign node730 = (inp[2]) ? 3'b001 : 3'b101;
										assign node733 = (inp[11]) ? 3'b011 : node734;
											assign node734 = (inp[8]) ? 3'b101 : 3'b011;
							assign node738 = (inp[8]) ? node768 : node739;
								assign node739 = (inp[5]) ? node757 : node740;
									assign node740 = (inp[4]) ? node750 : node741;
										assign node741 = (inp[2]) ? node743 : 3'b110;
											assign node743 = (inp[11]) ? node747 : node744;
												assign node744 = (inp[10]) ? 3'b100 : 3'b000;
												assign node747 = (inp[10]) ? 3'b010 : 3'b100;
										assign node750 = (inp[2]) ? node754 : node751;
											assign node751 = (inp[10]) ? 3'b001 : 3'b110;
											assign node754 = (inp[10]) ? 3'b110 : 3'b010;
									assign node757 = (inp[2]) ? node763 : node758;
										assign node758 = (inp[4]) ? node760 : 3'b001;
											assign node760 = (inp[10]) ? 3'b101 : 3'b110;
										assign node763 = (inp[4]) ? node765 : 3'b110;
											assign node765 = (inp[10]) ? 3'b001 : 3'b011;
								assign node768 = (inp[2]) ? node780 : node769;
									assign node769 = (inp[5]) ? node775 : node770;
										assign node770 = (inp[4]) ? node772 : 3'b010;
											assign node772 = (inp[10]) ? 3'b110 : 3'b010;
										assign node775 = (inp[10]) ? node777 : 3'b110;
											assign node777 = (inp[4]) ? 3'b001 : 3'b110;
									assign node780 = (inp[4]) ? node790 : node781;
										assign node781 = (inp[10]) ? node785 : node782;
											assign node782 = (inp[5]) ? 3'b100 : 3'b010;
											assign node785 = (inp[11]) ? node787 : 3'b100;
												assign node787 = (inp[5]) ? 3'b010 : 3'b100;
										assign node790 = (inp[5]) ? node794 : node791;
											assign node791 = (inp[10]) ? 3'b010 : 3'b100;
											assign node794 = (inp[10]) ? 3'b110 : 3'b010;
					assign node797 = (inp[1]) ? node925 : node798;
						assign node798 = (inp[9]) ? node878 : node799;
							assign node799 = (inp[4]) ? node845 : node800;
								assign node800 = (inp[2]) ? node820 : node801;
									assign node801 = (inp[10]) ? node809 : node802;
										assign node802 = (inp[5]) ? node804 : 3'b001;
											assign node804 = (inp[11]) ? 3'b101 : node805;
												assign node805 = (inp[8]) ? 3'b001 : 3'b101;
										assign node809 = (inp[8]) ? node815 : node810;
											assign node810 = (inp[5]) ? 3'b011 : node811;
												assign node811 = (inp[11]) ? 3'b011 : 3'b101;
											assign node815 = (inp[5]) ? node817 : 3'b101;
												assign node817 = (inp[11]) ? 3'b011 : 3'b101;
									assign node820 = (inp[5]) ? node834 : node821;
										assign node821 = (inp[8]) ? node829 : node822;
											assign node822 = (inp[10]) ? node826 : node823;
												assign node823 = (inp[11]) ? 3'b010 : 3'b110;
												assign node826 = (inp[11]) ? 3'b110 : 3'b010;
											assign node829 = (inp[10]) ? 3'b001 : node830;
												assign node830 = (inp[11]) ? 3'b110 : 3'b010;
										assign node834 = (inp[11]) ? node842 : node835;
											assign node835 = (inp[8]) ? node839 : node836;
												assign node836 = (inp[10]) ? 3'b110 : 3'b001;
												assign node839 = (inp[10]) ? 3'b001 : 3'b110;
											assign node842 = (inp[8]) ? 3'b101 : 3'b001;
								assign node845 = (inp[11]) ? node865 : node846;
									assign node846 = (inp[8]) ? node858 : node847;
										assign node847 = (inp[5]) ? node853 : node848;
											assign node848 = (inp[2]) ? node850 : 3'b011;
												assign node850 = (inp[10]) ? 3'b101 : 3'b001;
											assign node853 = (inp[2]) ? node855 : 3'b101;
												assign node855 = (inp[10]) ? 3'b011 : 3'b111;
										assign node858 = (inp[2]) ? node860 : 3'b011;
											assign node860 = (inp[5]) ? node862 : 3'b001;
												assign node862 = (inp[10]) ? 3'b101 : 3'b001;
									assign node865 = (inp[8]) ? node871 : node866;
										assign node866 = (inp[10]) ? node868 : 3'b111;
											assign node868 = (inp[5]) ? 3'b101 : 3'b111;
										assign node871 = (inp[5]) ? node873 : 3'b011;
											assign node873 = (inp[2]) ? node875 : 3'b111;
												assign node875 = (inp[10]) ? 3'b011 : 3'b111;
							assign node878 = (inp[4]) ? node914 : node879;
								assign node879 = (inp[10]) ? node907 : node880;
									assign node880 = (inp[11]) ? node894 : node881;
										assign node881 = (inp[2]) ? node887 : node882;
											assign node882 = (inp[8]) ? node884 : 3'b011;
												assign node884 = (inp[5]) ? 3'b011 : 3'b101;
											assign node887 = (inp[8]) ? node891 : node888;
												assign node888 = (inp[5]) ? 3'b011 : 3'b101;
												assign node891 = (inp[5]) ? 3'b101 : 3'b001;
										assign node894 = (inp[2]) ? node902 : node895;
											assign node895 = (inp[5]) ? node899 : node896;
												assign node896 = (inp[8]) ? 3'b011 : 3'b111;
												assign node899 = (inp[8]) ? 3'b111 : 3'b101;
											assign node902 = (inp[5]) ? 3'b011 : node903;
												assign node903 = (inp[8]) ? 3'b101 : 3'b011;
									assign node907 = (inp[11]) ? 3'b111 : node908;
										assign node908 = (inp[5]) ? node910 : 3'b011;
											assign node910 = (inp[2]) ? 3'b011 : 3'b111;
								assign node914 = (inp[2]) ? node916 : 3'b111;
									assign node916 = (inp[10]) ? 3'b111 : node917;
										assign node917 = (inp[11]) ? node921 : node918;
											assign node918 = (inp[5]) ? 3'b011 : 3'b111;
											assign node921 = (inp[5]) ? 3'b111 : 3'b011;
						assign node925 = (inp[9]) ? node1005 : node926;
							assign node926 = (inp[4]) ? node972 : node927;
								assign node927 = (inp[5]) ? node949 : node928;
									assign node928 = (inp[8]) ? node938 : node929;
										assign node929 = (inp[10]) ? node935 : node930;
											assign node930 = (inp[11]) ? 3'b110 : node931;
												assign node931 = (inp[2]) ? 3'b100 : 3'b010;
											assign node935 = (inp[2]) ? 3'b010 : 3'b001;
										assign node938 = (inp[10]) ? node944 : node939;
											assign node939 = (inp[11]) ? 3'b000 : node940;
												assign node940 = (inp[2]) ? 3'b000 : 3'b100;
											assign node944 = (inp[11]) ? node946 : 3'b000;
												assign node946 = (inp[2]) ? 3'b010 : 3'b110;
									assign node949 = (inp[2]) ? node959 : node950;
										assign node950 = (inp[10]) ? node956 : node951;
											assign node951 = (inp[8]) ? node953 : 3'b110;
												assign node953 = (inp[11]) ? 3'b110 : 3'b010;
											assign node956 = (inp[8]) ? 3'b110 : 3'b001;
										assign node959 = (inp[11]) ? node965 : node960;
											assign node960 = (inp[8]) ? 3'b010 : node961;
												assign node961 = (inp[10]) ? 3'b110 : 3'b010;
											assign node965 = (inp[10]) ? node969 : node966;
												assign node966 = (inp[8]) ? 3'b110 : 3'b010;
												assign node969 = (inp[8]) ? 3'b010 : 3'b110;
								assign node972 = (inp[2]) ? node990 : node973;
									assign node973 = (inp[8]) ? node981 : node974;
										assign node974 = (inp[10]) ? node976 : 3'b001;
											assign node976 = (inp[11]) ? 3'b101 : node977;
												assign node977 = (inp[5]) ? 3'b101 : 3'b001;
										assign node981 = (inp[5]) ? node983 : 3'b110;
											assign node983 = (inp[11]) ? node987 : node984;
												assign node984 = (inp[10]) ? 3'b001 : 3'b110;
												assign node987 = (inp[10]) ? 3'b101 : 3'b001;
									assign node990 = (inp[10]) ? node998 : node991;
										assign node991 = (inp[8]) ? node993 : 3'b110;
											assign node993 = (inp[11]) ? node995 : 3'b010;
												assign node995 = (inp[5]) ? 3'b110 : 3'b010;
										assign node998 = (inp[11]) ? 3'b001 : node999;
											assign node999 = (inp[5]) ? node1001 : 3'b110;
												assign node1001 = (inp[8]) ? 3'b110 : 3'b001;
							assign node1005 = (inp[4]) ? node1041 : node1006;
								assign node1006 = (inp[10]) ? node1022 : node1007;
									assign node1007 = (inp[2]) ? node1015 : node1008;
										assign node1008 = (inp[11]) ? 3'b101 : node1009;
											assign node1009 = (inp[5]) ? 3'b110 : node1010;
												assign node1010 = (inp[8]) ? 3'b110 : 3'b001;
										assign node1015 = (inp[11]) ? node1017 : 3'b010;
											assign node1017 = (inp[8]) ? 3'b110 : node1018;
												assign node1018 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1022 = (inp[2]) ? node1028 : node1023;
										assign node1023 = (inp[8]) ? 3'b101 : node1024;
											assign node1024 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1028 = (inp[11]) ? node1036 : node1029;
											assign node1029 = (inp[5]) ? node1033 : node1030;
												assign node1030 = (inp[8]) ? 3'b110 : 3'b001;
												assign node1033 = (inp[8]) ? 3'b001 : 3'b000;
											assign node1036 = (inp[8]) ? 3'b001 : node1037;
												assign node1037 = (inp[5]) ? 3'b100 : 3'b101;
								assign node1041 = (inp[2]) ? node1057 : node1042;
									assign node1042 = (inp[10]) ? node1054 : node1043;
										assign node1043 = (inp[8]) ? node1049 : node1044;
											assign node1044 = (inp[5]) ? 3'b011 : node1045;
												assign node1045 = (inp[11]) ? 3'b011 : 3'b101;
											assign node1049 = (inp[11]) ? node1051 : 3'b101;
												assign node1051 = (inp[5]) ? 3'b011 : 3'b101;
										assign node1054 = (inp[5]) ? 3'b111 : 3'b011;
									assign node1057 = (inp[10]) ? node1065 : node1058;
										assign node1058 = (inp[8]) ? node1060 : 3'b101;
											assign node1060 = (inp[5]) ? node1062 : 3'b001;
												assign node1062 = (inp[11]) ? 3'b101 : 3'b001;
										assign node1065 = (inp[5]) ? 3'b011 : 3'b101;
		assign node1068 = (inp[6]) ? node1924 : node1069;
			assign node1069 = (inp[3]) ? node1477 : node1070;
				assign node1070 = (inp[4]) ? node1286 : node1071;
					assign node1071 = (inp[9]) ? node1205 : node1072;
						assign node1072 = (inp[7]) ? node1146 : node1073;
							assign node1073 = (inp[8]) ? node1107 : node1074;
								assign node1074 = (inp[10]) ? node1084 : node1075;
									assign node1075 = (inp[1]) ? node1079 : node1076;
										assign node1076 = (inp[2]) ? 3'b100 : 3'b110;
										assign node1079 = (inp[11]) ? 3'b100 : node1080;
											assign node1080 = (inp[5]) ? 3'b100 : 3'b000;
									assign node1084 = (inp[11]) ? node1098 : node1085;
										assign node1085 = (inp[5]) ? node1091 : node1086;
											assign node1086 = (inp[1]) ? 3'b100 : node1087;
												assign node1087 = (inp[2]) ? 3'b100 : 3'b010;
											assign node1091 = (inp[1]) ? node1095 : node1092;
												assign node1092 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1095 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1098 = (inp[1]) ? node1104 : node1099;
											assign node1099 = (inp[2]) ? node1101 : 3'b110;
												assign node1101 = (inp[5]) ? 3'b110 : 3'b010;
											assign node1104 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1107 = (inp[2]) ? node1119 : node1108;
									assign node1108 = (inp[1]) ? node1114 : node1109;
										assign node1109 = (inp[5]) ? node1111 : 3'b010;
											assign node1111 = (inp[11]) ? 3'b110 : 3'b010;
										assign node1114 = (inp[11]) ? node1116 : 3'b000;
											assign node1116 = (inp[10]) ? 3'b010 : 3'b100;
									assign node1119 = (inp[10]) ? node1133 : node1120;
										assign node1120 = (inp[1]) ? node1126 : node1121;
											assign node1121 = (inp[5]) ? node1123 : 3'b100;
												assign node1123 = (inp[11]) ? 3'b010 : 3'b100;
											assign node1126 = (inp[11]) ? node1130 : node1127;
												assign node1127 = (inp[5]) ? 3'b110 : 3'b010;
												assign node1130 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1133 = (inp[1]) ? node1139 : node1134;
											assign node1134 = (inp[11]) ? node1136 : 3'b100;
												assign node1136 = (inp[5]) ? 3'b010 : 3'b100;
											assign node1139 = (inp[5]) ? node1143 : node1140;
												assign node1140 = (inp[11]) ? 3'b000 : 3'b100;
												assign node1143 = (inp[11]) ? 3'b100 : 3'b000;
							assign node1146 = (inp[1]) ? node1178 : node1147;
								assign node1147 = (inp[2]) ? node1163 : node1148;
									assign node1148 = (inp[8]) ? node1158 : node1149;
										assign node1149 = (inp[5]) ? node1155 : node1150;
											assign node1150 = (inp[10]) ? 3'b100 : node1151;
												assign node1151 = (inp[11]) ? 3'b000 : 3'b100;
											assign node1155 = (inp[10]) ? 3'b110 : 3'b100;
										assign node1158 = (inp[10]) ? 3'b000 : node1159;
											assign node1159 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1163 = (inp[8]) ? node1171 : node1164;
										assign node1164 = (inp[10]) ? node1168 : node1165;
											assign node1165 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1168 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1171 = (inp[10]) ? 3'b100 : node1172;
											assign node1172 = (inp[11]) ? node1174 : 3'b110;
												assign node1174 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1178 = (inp[10]) ? node1188 : node1179;
									assign node1179 = (inp[2]) ? node1185 : node1180;
										assign node1180 = (inp[5]) ? 3'b110 : node1181;
											assign node1181 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1185 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1188 = (inp[8]) ? node1198 : node1189;
										assign node1189 = (inp[2]) ? node1191 : 3'b000;
											assign node1191 = (inp[5]) ? node1195 : node1192;
												assign node1192 = (inp[11]) ? 3'b100 : 3'b000;
												assign node1195 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1198 = (inp[5]) ? node1200 : 3'b010;
											assign node1200 = (inp[2]) ? 3'b110 : node1201;
												assign node1201 = (inp[11]) ? 3'b000 : 3'b010;
						assign node1205 = (inp[1]) ? node1217 : node1206;
							assign node1206 = (inp[7]) ? node1208 : 3'b110;
								assign node1208 = (inp[2]) ? node1210 : 3'b110;
									assign node1210 = (inp[10]) ? node1212 : 3'b010;
										assign node1212 = (inp[5]) ? 3'b110 : node1213;
											assign node1213 = (inp[8]) ? 3'b010 : 3'b110;
							assign node1217 = (inp[7]) ? node1255 : node1218;
								assign node1218 = (inp[5]) ? node1244 : node1219;
									assign node1219 = (inp[10]) ? node1233 : node1220;
										assign node1220 = (inp[2]) ? node1226 : node1221;
											assign node1221 = (inp[8]) ? 3'b010 : node1222;
												assign node1222 = (inp[11]) ? 3'b110 : 3'b010;
											assign node1226 = (inp[8]) ? node1230 : node1227;
												assign node1227 = (inp[11]) ? 3'b010 : 3'b100;
												assign node1230 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1233 = (inp[2]) ? node1239 : node1234;
											assign node1234 = (inp[8]) ? node1236 : 3'b110;
												assign node1236 = (inp[11]) ? 3'b110 : 3'b010;
											assign node1239 = (inp[11]) ? 3'b010 : node1240;
												assign node1240 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1244 = (inp[10]) ? 3'b110 : node1245;
										assign node1245 = (inp[2]) ? node1251 : node1246;
											assign node1246 = (inp[8]) ? node1248 : 3'b110;
												assign node1248 = (inp[11]) ? 3'b110 : 3'b010;
											assign node1251 = (inp[11]) ? 3'b010 : 3'b100;
								assign node1255 = (inp[8]) ? node1271 : node1256;
									assign node1256 = (inp[5]) ? node1266 : node1257;
										assign node1257 = (inp[2]) ? node1263 : node1258;
											assign node1258 = (inp[10]) ? 3'b000 : node1259;
												assign node1259 = (inp[11]) ? 3'b000 : 3'b010;
											assign node1263 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1266 = (inp[10]) ? node1268 : 3'b100;
											assign node1268 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1271 = (inp[10]) ? node1277 : node1272;
										assign node1272 = (inp[11]) ? 3'b110 : node1273;
											assign node1273 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1277 = (inp[2]) ? 3'b000 : node1278;
											assign node1278 = (inp[5]) ? node1282 : node1279;
												assign node1279 = (inp[11]) ? 3'b100 : 3'b110;
												assign node1282 = (inp[11]) ? 3'b010 : 3'b000;
					assign node1286 = (inp[1]) ? node1410 : node1287;
						assign node1287 = (inp[7]) ? node1359 : node1288;
							assign node1288 = (inp[8]) ? node1324 : node1289;
								assign node1289 = (inp[9]) ? node1309 : node1290;
									assign node1290 = (inp[10]) ? node1298 : node1291;
										assign node1291 = (inp[11]) ? 3'b110 : node1292;
											assign node1292 = (inp[5]) ? node1294 : 3'b110;
												assign node1294 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1298 = (inp[2]) ? node1304 : node1299;
											assign node1299 = (inp[5]) ? 3'b110 : node1300;
												assign node1300 = (inp[11]) ? 3'b110 : 3'b001;
											assign node1304 = (inp[11]) ? 3'b001 : node1305;
												assign node1305 = (inp[5]) ? 3'b001 : 3'b110;
									assign node1309 = (inp[10]) ? node1319 : node1310;
										assign node1310 = (inp[2]) ? node1316 : node1311;
											assign node1311 = (inp[11]) ? 3'b001 : node1312;
												assign node1312 = (inp[5]) ? 3'b001 : 3'b110;
											assign node1316 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1319 = (inp[2]) ? node1321 : 3'b110;
											assign node1321 = (inp[11]) ? 3'b001 : 3'b110;
								assign node1324 = (inp[11]) ? node1334 : node1325;
									assign node1325 = (inp[10]) ? node1329 : node1326;
										assign node1326 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1329 = (inp[2]) ? node1331 : 3'b001;
											assign node1331 = (inp[9]) ? 3'b001 : 3'b110;
									assign node1334 = (inp[9]) ? node1344 : node1335;
										assign node1335 = (inp[2]) ? node1337 : 3'b110;
											assign node1337 = (inp[5]) ? node1341 : node1338;
												assign node1338 = (inp[10]) ? 3'b110 : 3'b001;
												assign node1341 = (inp[10]) ? 3'b001 : 3'b110;
										assign node1344 = (inp[2]) ? node1352 : node1345;
											assign node1345 = (inp[5]) ? node1349 : node1346;
												assign node1346 = (inp[10]) ? 3'b001 : 3'b110;
												assign node1349 = (inp[10]) ? 3'b110 : 3'b001;
											assign node1352 = (inp[5]) ? node1356 : node1353;
												assign node1353 = (inp[10]) ? 3'b110 : 3'b001;
												assign node1356 = (inp[10]) ? 3'b001 : 3'b110;
							assign node1359 = (inp[5]) ? node1379 : node1360;
								assign node1360 = (inp[2]) ? node1370 : node1361;
									assign node1361 = (inp[8]) ? node1365 : node1362;
										assign node1362 = (inp[10]) ? 3'b101 : 3'b001;
										assign node1365 = (inp[10]) ? node1367 : 3'b101;
											assign node1367 = (inp[11]) ? 3'b101 : 3'b001;
									assign node1370 = (inp[8]) ? node1374 : node1371;
										assign node1371 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1374 = (inp[10]) ? node1376 : 3'b001;
											assign node1376 = (inp[9]) ? 3'b101 : 3'b001;
								assign node1379 = (inp[8]) ? node1387 : node1380;
									assign node1380 = (inp[2]) ? node1384 : node1381;
										assign node1381 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1384 = (inp[10]) ? 3'b101 : 3'b001;
									assign node1387 = (inp[9]) ? node1395 : node1388;
										assign node1388 = (inp[2]) ? node1392 : node1389;
											assign node1389 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1392 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1395 = (inp[11]) ? node1403 : node1396;
											assign node1396 = (inp[10]) ? node1400 : node1397;
												assign node1397 = (inp[2]) ? 3'b101 : 3'b001;
												assign node1400 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1403 = (inp[2]) ? node1407 : node1404;
												assign node1404 = (inp[10]) ? 3'b101 : 3'b001;
												assign node1407 = (inp[10]) ? 3'b001 : 3'b101;
						assign node1410 = (inp[9]) ? node1430 : node1411;
							assign node1411 = (inp[7]) ? node1423 : node1412;
								assign node1412 = (inp[2]) ? 3'b001 : node1413;
									assign node1413 = (inp[8]) ? 3'b001 : node1414;
										assign node1414 = (inp[10]) ? node1416 : 3'b001;
											assign node1416 = (inp[5]) ? 3'b110 : node1417;
												assign node1417 = (inp[11]) ? 3'b110 : 3'b001;
								assign node1423 = (inp[5]) ? node1425 : 3'b000;
									assign node1425 = (inp[8]) ? 3'b000 : node1426;
										assign node1426 = (inp[2]) ? 3'b000 : 3'b001;
							assign node1430 = (inp[7]) ? node1464 : node1431;
								assign node1431 = (inp[11]) ? node1445 : node1432;
									assign node1432 = (inp[2]) ? 3'b001 : node1433;
										assign node1433 = (inp[8]) ? node1439 : node1434;
											assign node1434 = (inp[5]) ? node1436 : 3'b001;
												assign node1436 = (inp[10]) ? 3'b110 : 3'b001;
											assign node1439 = (inp[10]) ? node1441 : 3'b110;
												assign node1441 = (inp[5]) ? 3'b001 : 3'b110;
									assign node1445 = (inp[8]) ? node1451 : node1446;
										assign node1446 = (inp[10]) ? node1448 : 3'b110;
											assign node1448 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1451 = (inp[2]) ? node1457 : node1452;
											assign node1452 = (inp[10]) ? 3'b001 : node1453;
												assign node1453 = (inp[5]) ? 3'b001 : 3'b110;
											assign node1457 = (inp[5]) ? node1461 : node1458;
												assign node1458 = (inp[10]) ? 3'b110 : 3'b001;
												assign node1461 = (inp[10]) ? 3'b001 : 3'b110;
								assign node1464 = (inp[8]) ? node1472 : node1465;
									assign node1465 = (inp[2]) ? node1469 : node1466;
										assign node1466 = (inp[5]) ? 3'b001 : 3'b110;
										assign node1469 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1472 = (inp[2]) ? node1474 : 3'b110;
										assign node1474 = (inp[5]) ? 3'b010 : 3'b100;
				assign node1477 = (inp[7]) ? node1671 : node1478;
					assign node1478 = (inp[1]) ? node1530 : node1479;
						assign node1479 = (inp[9]) ? node1517 : node1480;
							assign node1480 = (inp[4]) ? node1498 : node1481;
								assign node1481 = (inp[2]) ? node1483 : 3'b111;
									assign node1483 = (inp[10]) ? 3'b111 : node1484;
										assign node1484 = (inp[5]) ? node1492 : node1485;
											assign node1485 = (inp[8]) ? node1489 : node1486;
												assign node1486 = (inp[11]) ? 3'b111 : 3'b011;
												assign node1489 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1492 = (inp[11]) ? 3'b111 : node1493;
												assign node1493 = (inp[8]) ? 3'b011 : 3'b111;
								assign node1498 = (inp[2]) ? node1504 : node1499;
									assign node1499 = (inp[8]) ? node1501 : 3'b111;
										assign node1501 = (inp[11]) ? 3'b111 : 3'b011;
									assign node1504 = (inp[8]) ? node1512 : node1505;
										assign node1505 = (inp[11]) ? node1509 : node1506;
											assign node1506 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1509 = (inp[5]) ? 3'b111 : 3'b011;
										assign node1512 = (inp[5]) ? node1514 : 3'b101;
											assign node1514 = (inp[11]) ? 3'b011 : 3'b101;
							assign node1517 = (inp[4]) ? 3'b111 : node1518;
								assign node1518 = (inp[10]) ? 3'b111 : node1519;
									assign node1519 = (inp[5]) ? 3'b111 : node1520;
										assign node1520 = (inp[2]) ? node1522 : 3'b111;
											assign node1522 = (inp[8]) ? 3'b011 : node1523;
												assign node1523 = (inp[11]) ? 3'b111 : 3'b011;
						assign node1530 = (inp[9]) ? node1596 : node1531;
							assign node1531 = (inp[4]) ? node1567 : node1532;
								assign node1532 = (inp[8]) ? node1554 : node1533;
									assign node1533 = (inp[5]) ? node1547 : node1534;
										assign node1534 = (inp[11]) ? node1542 : node1535;
											assign node1535 = (inp[10]) ? node1539 : node1536;
												assign node1536 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1539 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1542 = (inp[2]) ? 3'b010 : node1543;
												assign node1543 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1547 = (inp[2]) ? node1551 : node1548;
											assign node1548 = (inp[10]) ? 3'b111 : 3'b011;
											assign node1551 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1554 = (inp[5]) ? node1560 : node1555;
										assign node1555 = (inp[10]) ? 3'b000 : node1556;
											assign node1556 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1560 = (inp[10]) ? node1564 : node1561;
											assign node1561 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1564 = (inp[11]) ? 3'b110 : 3'b010;
								assign node1567 = (inp[2]) ? node1579 : node1568;
									assign node1568 = (inp[10]) ? node1574 : node1569;
										assign node1569 = (inp[11]) ? 3'b101 : node1570;
											assign node1570 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1574 = (inp[5]) ? 3'b011 : node1575;
											assign node1575 = (inp[8]) ? 3'b001 : 3'b101;
									assign node1579 = (inp[5]) ? node1587 : node1580;
										assign node1580 = (inp[10]) ? node1584 : node1581;
											assign node1581 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1584 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1587 = (inp[10]) ? node1593 : node1588;
											assign node1588 = (inp[8]) ? node1590 : 3'b001;
												assign node1590 = (inp[11]) ? 3'b011 : 3'b110;
											assign node1593 = (inp[8]) ? 3'b101 : 3'b111;
							assign node1596 = (inp[2]) ? node1632 : node1597;
								assign node1597 = (inp[4]) ? node1619 : node1598;
									assign node1598 = (inp[10]) ? node1614 : node1599;
										assign node1599 = (inp[11]) ? node1607 : node1600;
											assign node1600 = (inp[5]) ? node1604 : node1601;
												assign node1601 = (inp[8]) ? 3'b011 : 3'b111;
												assign node1604 = (inp[8]) ? 3'b111 : 3'b011;
											assign node1607 = (inp[5]) ? node1611 : node1608;
												assign node1608 = (inp[8]) ? 3'b011 : 3'b111;
												assign node1611 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1614 = (inp[8]) ? 3'b011 : node1615;
											assign node1615 = (inp[5]) ? 3'b111 : 3'b011;
									assign node1619 = (inp[10]) ? 3'b111 : node1620;
										assign node1620 = (inp[8]) ? node1626 : node1621;
											assign node1621 = (inp[5]) ? 3'b111 : node1622;
												assign node1622 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1626 = (inp[5]) ? 3'b011 : node1627;
												assign node1627 = (inp[11]) ? 3'b011 : 3'b111;
								assign node1632 = (inp[4]) ? node1650 : node1633;
									assign node1633 = (inp[5]) ? node1643 : node1634;
										assign node1634 = (inp[10]) ? node1638 : node1635;
											assign node1635 = (inp[8]) ? 3'b111 : 3'b001;
											assign node1638 = (inp[11]) ? 3'b101 : node1639;
												assign node1639 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1643 = (inp[10]) ? node1647 : node1644;
											assign node1644 = (inp[8]) ? 3'b001 : 3'b101;
											assign node1647 = (inp[8]) ? 3'b101 : 3'b011;
									assign node1650 = (inp[10]) ? node1662 : node1651;
										assign node1651 = (inp[5]) ? node1657 : node1652;
											assign node1652 = (inp[11]) ? node1654 : 3'b101;
												assign node1654 = (inp[8]) ? 3'b101 : 3'b011;
											assign node1657 = (inp[8]) ? node1659 : 3'b011;
												assign node1659 = (inp[11]) ? 3'b011 : 3'b101;
										assign node1662 = (inp[8]) ? node1664 : 3'b111;
											assign node1664 = (inp[11]) ? node1668 : node1665;
												assign node1665 = (inp[5]) ? 3'b011 : 3'b111;
												assign node1668 = (inp[5]) ? 3'b111 : 3'b011;
					assign node1671 = (inp[9]) ? node1797 : node1672;
						assign node1672 = (inp[4]) ? node1740 : node1673;
							assign node1673 = (inp[5]) ? node1707 : node1674;
								assign node1674 = (inp[1]) ? node1688 : node1675;
									assign node1675 = (inp[2]) ? node1683 : node1676;
										assign node1676 = (inp[10]) ? 3'b000 : node1677;
											assign node1677 = (inp[8]) ? 3'b110 : node1678;
												assign node1678 = (inp[11]) ? 3'b000 : 3'b110;
										assign node1683 = (inp[10]) ? 3'b110 : node1684;
											assign node1684 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1688 = (inp[8]) ? node1698 : node1689;
										assign node1689 = (inp[11]) ? node1693 : node1690;
											assign node1690 = (inp[2]) ? 3'b100 : 3'b010;
											assign node1693 = (inp[10]) ? node1695 : 3'b010;
												assign node1695 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1698 = (inp[11]) ? node1700 : 3'b000;
											assign node1700 = (inp[10]) ? node1704 : node1701;
												assign node1701 = (inp[2]) ? 3'b000 : 3'b100;
												assign node1704 = (inp[2]) ? 3'b100 : 3'b010;
								assign node1707 = (inp[1]) ? node1723 : node1708;
									assign node1708 = (inp[2]) ? node1716 : node1709;
										assign node1709 = (inp[8]) ? node1711 : 3'b001;
											assign node1711 = (inp[10]) ? 3'b000 : node1712;
												assign node1712 = (inp[11]) ? 3'b000 : 3'b110;
										assign node1716 = (inp[8]) ? node1720 : node1717;
											assign node1717 = (inp[10]) ? 3'b000 : 3'b110;
											assign node1720 = (inp[10]) ? 3'b110 : 3'b010;
									assign node1723 = (inp[10]) ? node1733 : node1724;
										assign node1724 = (inp[2]) ? node1728 : node1725;
											assign node1725 = (inp[11]) ? 3'b010 : 3'b100;
											assign node1728 = (inp[11]) ? 3'b100 : node1729;
												assign node1729 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1733 = (inp[11]) ? 3'b010 : node1734;
											assign node1734 = (inp[8]) ? 3'b100 : node1735;
												assign node1735 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1740 = (inp[1]) ? node1770 : node1741;
								assign node1741 = (inp[8]) ? node1757 : node1742;
									assign node1742 = (inp[2]) ? node1750 : node1743;
										assign node1743 = (inp[11]) ? node1745 : 3'b101;
											assign node1745 = (inp[5]) ? node1747 : 3'b001;
												assign node1747 = (inp[10]) ? 3'b111 : 3'b011;
										assign node1750 = (inp[10]) ? node1754 : node1751;
											assign node1751 = (inp[11]) ? 3'b101 : 3'b001;
											assign node1754 = (inp[5]) ? 3'b011 : 3'b001;
									assign node1757 = (inp[2]) ? node1763 : node1758;
										assign node1758 = (inp[10]) ? 3'b001 : node1759;
											assign node1759 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1763 = (inp[5]) ? node1767 : node1764;
											assign node1764 = (inp[10]) ? 3'b100 : 3'b110;
											assign node1767 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1770 = (inp[10]) ? node1780 : node1771;
									assign node1771 = (inp[2]) ? node1777 : node1772;
										assign node1772 = (inp[8]) ? node1774 : 3'b110;
											assign node1774 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1777 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1780 = (inp[8]) ? node1790 : node1781;
										assign node1781 = (inp[2]) ? node1785 : node1782;
											assign node1782 = (inp[11]) ? 3'b001 : 3'b011;
											assign node1785 = (inp[5]) ? 3'b001 : node1786;
												assign node1786 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1790 = (inp[2]) ? 3'b010 : node1791;
											assign node1791 = (inp[5]) ? 3'b011 : node1792;
												assign node1792 = (inp[11]) ? 3'b011 : 3'b010;
						assign node1797 = (inp[1]) ? node1845 : node1798;
							assign node1798 = (inp[4]) ? node1836 : node1799;
								assign node1799 = (inp[2]) ? node1819 : node1800;
									assign node1800 = (inp[10]) ? node1808 : node1801;
										assign node1801 = (inp[8]) ? node1803 : 3'b011;
											assign node1803 = (inp[5]) ? node1805 : 3'b101;
												assign node1805 = (inp[11]) ? 3'b011 : 3'b101;
										assign node1808 = (inp[8]) ? node1814 : node1809;
											assign node1809 = (inp[11]) ? 3'b111 : node1810;
												assign node1810 = (inp[5]) ? 3'b111 : 3'b011;
											assign node1814 = (inp[5]) ? node1816 : 3'b011;
												assign node1816 = (inp[11]) ? 3'b111 : 3'b011;
									assign node1819 = (inp[10]) ? node1823 : node1820;
										assign node1820 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1823 = (inp[5]) ? node1831 : node1824;
											assign node1824 = (inp[11]) ? node1828 : node1825;
												assign node1825 = (inp[8]) ? 3'b001 : 3'b101;
												assign node1828 = (inp[8]) ? 3'b101 : 3'b011;
											assign node1831 = (inp[8]) ? node1833 : 3'b011;
												assign node1833 = (inp[11]) ? 3'b011 : 3'b101;
								assign node1836 = (inp[2]) ? node1838 : 3'b111;
									assign node1838 = (inp[10]) ? node1840 : 3'b011;
										assign node1840 = (inp[5]) ? 3'b111 : node1841;
											assign node1841 = (inp[8]) ? 3'b011 : 3'b111;
							assign node1845 = (inp[10]) ? node1881 : node1846;
								assign node1846 = (inp[2]) ? node1866 : node1847;
									assign node1847 = (inp[8]) ? node1855 : node1848;
										assign node1848 = (inp[5]) ? node1852 : node1849;
											assign node1849 = (inp[11]) ? 3'b001 : 3'b010;
											assign node1852 = (inp[4]) ? 3'b101 : 3'b001;
										assign node1855 = (inp[5]) ? node1863 : node1856;
											assign node1856 = (inp[4]) ? node1860 : node1857;
												assign node1857 = (inp[11]) ? 3'b110 : 3'b010;
												assign node1860 = (inp[11]) ? 3'b110 : 3'b111;
											assign node1863 = (inp[11]) ? 3'b001 : 3'b110;
									assign node1866 = (inp[4]) ? node1872 : node1867;
										assign node1867 = (inp[11]) ? 3'b110 : node1868;
											assign node1868 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1872 = (inp[5]) ? node1878 : node1873;
											assign node1873 = (inp[11]) ? 3'b110 : node1874;
												assign node1874 = (inp[8]) ? 3'b101 : 3'b110;
											assign node1878 = (inp[8]) ? 3'b001 : 3'b101;
								assign node1881 = (inp[4]) ? node1901 : node1882;
									assign node1882 = (inp[2]) ? node1894 : node1883;
										assign node1883 = (inp[11]) ? node1889 : node1884;
											assign node1884 = (inp[8]) ? node1886 : 3'b001;
												assign node1886 = (inp[5]) ? 3'b001 : 3'b100;
											assign node1889 = (inp[8]) ? node1891 : 3'b101;
												assign node1891 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1894 = (inp[5]) ? node1896 : 3'b110;
											assign node1896 = (inp[11]) ? 3'b001 : node1897;
												assign node1897 = (inp[8]) ? 3'b110 : 3'b001;
									assign node1901 = (inp[2]) ? node1915 : node1902;
										assign node1902 = (inp[8]) ? node1908 : node1903;
											assign node1903 = (inp[5]) ? 3'b111 : node1904;
												assign node1904 = (inp[11]) ? 3'b011 : 3'b001;
											assign node1908 = (inp[5]) ? node1912 : node1909;
												assign node1909 = (inp[11]) ? 3'b101 : 3'b111;
												assign node1912 = (inp[11]) ? 3'b011 : 3'b001;
										assign node1915 = (inp[5]) ? node1919 : node1916;
											assign node1916 = (inp[8]) ? 3'b001 : 3'b101;
											assign node1919 = (inp[8]) ? 3'b101 : node1920;
												assign node1920 = (inp[11]) ? 3'b011 : 3'b101;
			assign node1924 = (inp[1]) ? node2272 : node1925;
				assign node1925 = (inp[7]) ? node2117 : node1926;
					assign node1926 = (inp[9]) ? node2012 : node1927;
						assign node1927 = (inp[2]) ? node1983 : node1928;
							assign node1928 = (inp[4]) ? node1956 : node1929;
								assign node1929 = (inp[3]) ? node1951 : node1930;
									assign node1930 = (inp[5]) ? node1940 : node1931;
										assign node1931 = (inp[10]) ? node1935 : node1932;
											assign node1932 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1935 = (inp[11]) ? 3'b010 : node1936;
												assign node1936 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1940 = (inp[11]) ? node1946 : node1941;
											assign node1941 = (inp[8]) ? node1943 : 3'b010;
												assign node1943 = (inp[10]) ? 3'b010 : 3'b110;
											assign node1946 = (inp[8]) ? 3'b010 : node1947;
												assign node1947 = (inp[10]) ? 3'b110 : 3'b010;
									assign node1951 = (inp[8]) ? node1953 : 3'b010;
										assign node1953 = (inp[5]) ? 3'b010 : 3'b100;
								assign node1956 = (inp[3]) ? node1968 : node1957;
									assign node1957 = (inp[10]) ? node1963 : node1958;
										assign node1958 = (inp[5]) ? 3'b100 : node1959;
											assign node1959 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1963 = (inp[5]) ? 3'b101 : node1964;
											assign node1964 = (inp[8]) ? 3'b110 : 3'b101;
									assign node1968 = (inp[5]) ? node1978 : node1969;
										assign node1969 = (inp[8]) ? node1973 : node1970;
											assign node1970 = (inp[10]) ? 3'b010 : 3'b110;
											assign node1973 = (inp[11]) ? 3'b010 : node1974;
												assign node1974 = (inp[10]) ? 3'b110 : 3'b010;
										assign node1978 = (inp[8]) ? node1980 : 3'b101;
											assign node1980 = (inp[10]) ? 3'b010 : 3'b110;
							assign node1983 = (inp[4]) ? node1999 : node1984;
								assign node1984 = (inp[3]) ? 3'b100 : node1985;
									assign node1985 = (inp[5]) ? node1993 : node1986;
										assign node1986 = (inp[8]) ? node1990 : node1987;
											assign node1987 = (inp[10]) ? 3'b100 : 3'b000;
											assign node1990 = (inp[10]) ? 3'b000 : 3'b110;
										assign node1993 = (inp[10]) ? 3'b010 : node1994;
											assign node1994 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1999 = (inp[3]) ? node2001 : 3'b110;
									assign node2001 = (inp[8]) ? node2009 : node2002;
										assign node2002 = (inp[5]) ? node2006 : node2003;
											assign node2003 = (inp[10]) ? 3'b110 : 3'b010;
											assign node2006 = (inp[10]) ? 3'b010 : 3'b110;
										assign node2009 = (inp[5]) ? 3'b010 : 3'b100;
						assign node2012 = (inp[3]) ? node2074 : node2013;
							assign node2013 = (inp[8]) ? node2045 : node2014;
								assign node2014 = (inp[5]) ? node2030 : node2015;
									assign node2015 = (inp[2]) ? node2025 : node2016;
										assign node2016 = (inp[4]) ? node2020 : node2017;
											assign node2017 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2020 = (inp[11]) ? node2022 : 3'b000;
												assign node2022 = (inp[10]) ? 3'b001 : 3'b000;
										assign node2025 = (inp[10]) ? node2027 : 3'b000;
											assign node2027 = (inp[4]) ? 3'b110 : 3'b100;
									assign node2030 = (inp[10]) ? node2038 : node2031;
										assign node2031 = (inp[11]) ? node2033 : 3'b100;
											assign node2033 = (inp[4]) ? node2035 : 3'b100;
												assign node2035 = (inp[2]) ? 3'b110 : 3'b100;
										assign node2038 = (inp[2]) ? node2042 : node2039;
											assign node2039 = (inp[4]) ? 3'b101 : 3'b110;
											assign node2042 = (inp[4]) ? 3'b110 : 3'b010;
								assign node2045 = (inp[5]) ? node2059 : node2046;
									assign node2046 = (inp[2]) ? node2052 : node2047;
										assign node2047 = (inp[4]) ? 3'b110 : node2048;
											assign node2048 = (inp[10]) ? 3'b110 : 3'b010;
										assign node2052 = (inp[4]) ? 3'b010 : node2053;
											assign node2053 = (inp[10]) ? node2055 : 3'b110;
												assign node2055 = (inp[11]) ? 3'b100 : 3'b000;
									assign node2059 = (inp[2]) ? node2069 : node2060;
										assign node2060 = (inp[4]) ? node2064 : node2061;
											assign node2061 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2064 = (inp[10]) ? node2066 : 3'b000;
												assign node2066 = (inp[11]) ? 3'b001 : 3'b000;
										assign node2069 = (inp[4]) ? 3'b110 : node2070;
											assign node2070 = (inp[10]) ? 3'b100 : 3'b000;
							assign node2074 = (inp[4]) ? node2106 : node2075;
								assign node2075 = (inp[2]) ? node2087 : node2076;
									assign node2076 = (inp[5]) ? node2084 : node2077;
										assign node2077 = (inp[8]) ? node2079 : 3'b101;
											assign node2079 = (inp[11]) ? node2081 : 3'b000;
												assign node2081 = (inp[10]) ? 3'b001 : 3'b000;
										assign node2084 = (inp[8]) ? 3'b101 : 3'b011;
									assign node2087 = (inp[10]) ? node2097 : node2088;
										assign node2088 = (inp[8]) ? node2094 : node2089;
											assign node2089 = (inp[5]) ? node2091 : 3'b100;
												assign node2091 = (inp[11]) ? 3'b000 : 3'b100;
											assign node2094 = (inp[5]) ? 3'b000 : 3'b010;
										assign node2097 = (inp[8]) ? 3'b100 : node2098;
											assign node2098 = (inp[5]) ? node2102 : node2099;
												assign node2099 = (inp[11]) ? 3'b001 : 3'b100;
												assign node2102 = (inp[11]) ? 3'b101 : 3'b001;
								assign node2106 = (inp[2]) ? 3'b101 : node2107;
									assign node2107 = (inp[10]) ? node2109 : 3'b101;
										assign node2109 = (inp[5]) ? 3'b111 : node2110;
											assign node2110 = (inp[8]) ? 3'b101 : node2111;
												assign node2111 = (inp[11]) ? 3'b111 : 3'b101;
					assign node2117 = (inp[3]) ? node2167 : node2118;
						assign node2118 = (inp[2]) ? node2152 : node2119;
							assign node2119 = (inp[9]) ? node2129 : node2120;
								assign node2120 = (inp[4]) ? 3'b000 : node2121;
									assign node2121 = (inp[10]) ? node2123 : 3'b000;
										assign node2123 = (inp[11]) ? 3'b100 : node2124;
											assign node2124 = (inp[5]) ? 3'b100 : 3'b000;
								assign node2129 = (inp[4]) ? node2139 : node2130;
									assign node2130 = (inp[10]) ? node2132 : 3'b000;
										assign node2132 = (inp[8]) ? node2134 : 3'b100;
											assign node2134 = (inp[11]) ? node2136 : 3'b000;
												assign node2136 = (inp[5]) ? 3'b100 : 3'b000;
									assign node2139 = (inp[10]) ? node2145 : node2140;
										assign node2140 = (inp[8]) ? node2142 : 3'b100;
											assign node2142 = (inp[5]) ? 3'b100 : 3'b000;
										assign node2145 = (inp[8]) ? node2149 : node2146;
											assign node2146 = (inp[5]) ? 3'b110 : 3'b010;
											assign node2149 = (inp[5]) ? 3'b010 : 3'b100;
							assign node2152 = (inp[8]) ? 3'b000 : node2153;
								assign node2153 = (inp[9]) ? node2155 : 3'b000;
									assign node2155 = (inp[5]) ? node2163 : node2156;
										assign node2156 = (inp[4]) ? node2158 : 3'b000;
											assign node2158 = (inp[10]) ? node2160 : 3'b000;
												assign node2160 = (inp[11]) ? 3'b100 : 3'b000;
										assign node2163 = (inp[10]) ? 3'b000 : 3'b010;
						assign node2167 = (inp[9]) ? node2211 : node2168;
							assign node2168 = (inp[4]) ? node2182 : node2169;
								assign node2169 = (inp[10]) ? node2171 : 3'b000;
									assign node2171 = (inp[2]) ? node2177 : node2172;
										assign node2172 = (inp[5]) ? node2174 : 3'b100;
											assign node2174 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2177 = (inp[5]) ? node2179 : 3'b000;
											assign node2179 = (inp[8]) ? 3'b000 : 3'b100;
								assign node2182 = (inp[8]) ? node2196 : node2183;
									assign node2183 = (inp[2]) ? node2189 : node2184;
										assign node2184 = (inp[11]) ? node2186 : 3'b010;
											assign node2186 = (inp[5]) ? 3'b110 : 3'b010;
										assign node2189 = (inp[10]) ? node2191 : 3'b100;
											assign node2191 = (inp[11]) ? 3'b010 : node2192;
												assign node2192 = (inp[5]) ? 3'b010 : 3'b100;
									assign node2196 = (inp[5]) ? node2202 : node2197;
										assign node2197 = (inp[2]) ? node2199 : 3'b100;
											assign node2199 = (inp[10]) ? 3'b100 : 3'b000;
										assign node2202 = (inp[2]) ? 3'b100 : node2203;
											assign node2203 = (inp[11]) ? node2207 : node2204;
												assign node2204 = (inp[10]) ? 3'b010 : 3'b100;
												assign node2207 = (inp[10]) ? 3'b110 : 3'b010;
							assign node2211 = (inp[2]) ? node2245 : node2212;
								assign node2212 = (inp[8]) ? node2226 : node2213;
									assign node2213 = (inp[10]) ? node2221 : node2214;
										assign node2214 = (inp[5]) ? node2218 : node2215;
											assign node2215 = (inp[4]) ? 3'b001 : 3'b011;
											assign node2218 = (inp[4]) ? 3'b001 : 3'b101;
										assign node2221 = (inp[11]) ? node2223 : 3'b101;
											assign node2223 = (inp[4]) ? 3'b101 : 3'b001;
									assign node2226 = (inp[4]) ? node2236 : node2227;
										assign node2227 = (inp[10]) ? node2233 : node2228;
											assign node2228 = (inp[5]) ? 3'b010 : node2229;
												assign node2229 = (inp[11]) ? 3'b010 : 3'b100;
											assign node2233 = (inp[11]) ? 3'b110 : 3'b010;
										assign node2236 = (inp[10]) ? node2240 : node2237;
											assign node2237 = (inp[11]) ? 3'b001 : 3'b110;
											assign node2240 = (inp[5]) ? node2242 : 3'b001;
												assign node2242 = (inp[11]) ? 3'b101 : 3'b001;
								assign node2245 = (inp[10]) ? node2259 : node2246;
									assign node2246 = (inp[4]) ? node2256 : node2247;
										assign node2247 = (inp[5]) ? node2253 : node2248;
											assign node2248 = (inp[8]) ? node2250 : 3'b100;
												assign node2250 = (inp[11]) ? 3'b100 : 3'b000;
											assign node2253 = (inp[8]) ? 3'b100 : 3'b000;
										assign node2256 = (inp[11]) ? 3'b110 : 3'b010;
									assign node2259 = (inp[4]) ? node2265 : node2260;
										assign node2260 = (inp[8]) ? 3'b010 : node2261;
											assign node2261 = (inp[5]) ? 3'b110 : 3'b010;
										assign node2265 = (inp[5]) ? 3'b001 : node2266;
											assign node2266 = (inp[8]) ? node2268 : 3'b110;
												assign node2268 = (inp[11]) ? 3'b110 : 3'b010;
				assign node2272 = (inp[3]) ? node2330 : node2273;
					assign node2273 = (inp[2]) ? node2315 : node2274;
						assign node2274 = (inp[9]) ? node2294 : node2275;
							assign node2275 = (inp[4]) ? node2283 : node2276;
								assign node2276 = (inp[8]) ? 3'b000 : node2277;
									assign node2277 = (inp[7]) ? 3'b000 : node2278;
										assign node2278 = (inp[5]) ? 3'b100 : 3'b000;
								assign node2283 = (inp[10]) ? node2285 : 3'b000;
									assign node2285 = (inp[7]) ? 3'b000 : node2286;
										assign node2286 = (inp[5]) ? node2288 : 3'b000;
											assign node2288 = (inp[11]) ? 3'b010 : node2289;
												assign node2289 = (inp[8]) ? 3'b000 : 3'b010;
							assign node2294 = (inp[4]) ? node2302 : node2295;
								assign node2295 = (inp[8]) ? 3'b000 : node2296;
									assign node2296 = (inp[7]) ? 3'b000 : node2297;
										assign node2297 = (inp[5]) ? 3'b100 : 3'b000;
								assign node2302 = (inp[5]) ? node2308 : node2303;
									assign node2303 = (inp[8]) ? node2305 : 3'b000;
										assign node2305 = (inp[7]) ? 3'b000 : 3'b100;
									assign node2308 = (inp[8]) ? 3'b000 : node2309;
										assign node2309 = (inp[7]) ? 3'b100 : node2310;
											assign node2310 = (inp[10]) ? 3'b010 : 3'b000;
						assign node2315 = (inp[9]) ? node2317 : 3'b000;
							assign node2317 = (inp[4]) ? node2319 : 3'b000;
								assign node2319 = (inp[7]) ? 3'b000 : node2320;
									assign node2320 = (inp[8]) ? 3'b000 : node2321;
										assign node2321 = (inp[10]) ? node2323 : 3'b000;
											assign node2323 = (inp[5]) ? 3'b100 : node2324;
												assign node2324 = (inp[11]) ? 3'b100 : 3'b000;
					assign node2330 = (inp[9]) ? node2378 : node2331;
						assign node2331 = (inp[4]) ? node2341 : node2332;
							assign node2332 = (inp[5]) ? node2334 : 3'b000;
								assign node2334 = (inp[7]) ? node2336 : 3'b000;
									assign node2336 = (inp[8]) ? 3'b000 : node2337;
										assign node2337 = (inp[2]) ? 3'b000 : 3'b010;
							assign node2341 = (inp[7]) ? node2367 : node2342;
								assign node2342 = (inp[5]) ? node2352 : node2343;
									assign node2343 = (inp[11]) ? node2349 : node2344;
										assign node2344 = (inp[2]) ? 3'b000 : node2345;
											assign node2345 = (inp[8]) ? 3'b000 : 3'b100;
										assign node2349 = (inp[8]) ? 3'b100 : 3'b010;
									assign node2352 = (inp[8]) ? node2358 : node2353;
										assign node2353 = (inp[10]) ? 3'b010 : node2354;
											assign node2354 = (inp[2]) ? 3'b100 : 3'b010;
										assign node2358 = (inp[11]) ? node2362 : node2359;
											assign node2359 = (inp[2]) ? 3'b000 : 3'b100;
											assign node2362 = (inp[2]) ? node2364 : 3'b010;
												assign node2364 = (inp[10]) ? 3'b100 : 3'b000;
								assign node2367 = (inp[10]) ? node2369 : 3'b000;
									assign node2369 = (inp[2]) ? 3'b000 : node2370;
										assign node2370 = (inp[8]) ? node2372 : 3'b100;
											assign node2372 = (inp[5]) ? node2374 : 3'b000;
												assign node2374 = (inp[11]) ? 3'b100 : 3'b000;
						assign node2378 = (inp[7]) ? node2450 : node2379;
							assign node2379 = (inp[2]) ? node2409 : node2380;
								assign node2380 = (inp[4]) ? node2388 : node2381;
									assign node2381 = (inp[5]) ? node2385 : node2382;
										assign node2382 = (inp[8]) ? 3'b010 : 3'b110;
										assign node2385 = (inp[8]) ? 3'b110 : 3'b001;
									assign node2388 = (inp[5]) ? node2396 : node2389;
										assign node2389 = (inp[11]) ? 3'b001 : node2390;
											assign node2390 = (inp[10]) ? node2392 : 3'b001;
												assign node2392 = (inp[8]) ? 3'b101 : 3'b001;
										assign node2396 = (inp[11]) ? node2402 : node2397;
											assign node2397 = (inp[10]) ? 3'b001 : node2398;
												assign node2398 = (inp[8]) ? 3'b101 : 3'b001;
											assign node2402 = (inp[10]) ? node2406 : node2403;
												assign node2403 = (inp[8]) ? 3'b101 : 3'b001;
												assign node2406 = (inp[8]) ? 3'b001 : 3'b101;
								assign node2409 = (inp[10]) ? node2431 : node2410;
									assign node2410 = (inp[8]) ? node2422 : node2411;
										assign node2411 = (inp[5]) ? node2417 : node2412;
											assign node2412 = (inp[4]) ? 3'b010 : node2413;
												assign node2413 = (inp[11]) ? 3'b100 : 3'b000;
											assign node2417 = (inp[4]) ? 3'b110 : node2418;
												assign node2418 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2422 = (inp[11]) ? 3'b100 : node2423;
											assign node2423 = (inp[4]) ? node2427 : node2424;
												assign node2424 = (inp[5]) ? 3'b000 : 3'b010;
												assign node2427 = (inp[5]) ? 3'b010 : 3'b100;
									assign node2431 = (inp[5]) ? node2441 : node2432;
										assign node2432 = (inp[4]) ? node2436 : node2433;
											assign node2433 = (inp[11]) ? 3'b010 : 3'b100;
											assign node2436 = (inp[11]) ? 3'b110 : node2437;
												assign node2437 = (inp[8]) ? 3'b010 : 3'b110;
										assign node2441 = (inp[4]) ? 3'b001 : node2442;
											assign node2442 = (inp[8]) ? node2446 : node2443;
												assign node2443 = (inp[11]) ? 3'b110 : 3'b010;
												assign node2446 = (inp[11]) ? 3'b010 : 3'b100;
							assign node2450 = (inp[4]) ? node2472 : node2451;
								assign node2451 = (inp[10]) ? node2457 : node2452;
									assign node2452 = (inp[8]) ? 3'b000 : node2453;
										assign node2453 = (inp[2]) ? 3'b000 : 3'b010;
									assign node2457 = (inp[8]) ? node2467 : node2458;
										assign node2458 = (inp[11]) ? node2460 : 3'b100;
											assign node2460 = (inp[2]) ? node2464 : node2461;
												assign node2461 = (inp[5]) ? 3'b010 : 3'b100;
												assign node2464 = (inp[5]) ? 3'b100 : 3'b000;
										assign node2467 = (inp[2]) ? 3'b000 : node2468;
											assign node2468 = (inp[5]) ? 3'b100 : 3'b000;
								assign node2472 = (inp[10]) ? node2492 : node2473;
									assign node2473 = (inp[2]) ? node2485 : node2474;
										assign node2474 = (inp[5]) ? node2480 : node2475;
											assign node2475 = (inp[11]) ? node2477 : 3'b100;
												assign node2477 = (inp[8]) ? 3'b100 : 3'b010;
											assign node2480 = (inp[11]) ? 3'b010 : node2481;
												assign node2481 = (inp[8]) ? 3'b100 : 3'b010;
										assign node2485 = (inp[11]) ? node2487 : 3'b000;
											assign node2487 = (inp[5]) ? 3'b100 : node2488;
												assign node2488 = (inp[8]) ? 3'b000 : 3'b100;
									assign node2492 = (inp[2]) ? node2502 : node2493;
										assign node2493 = (inp[5]) ? 3'b110 : node2494;
											assign node2494 = (inp[11]) ? node2498 : node2495;
												assign node2495 = (inp[8]) ? 3'b100 : 3'b010;
												assign node2498 = (inp[8]) ? 3'b010 : 3'b110;
										assign node2502 = (inp[8]) ? node2504 : 3'b010;
											assign node2504 = (inp[11]) ? 3'b010 : node2505;
												assign node2505 = (inp[5]) ? 3'b100 : 3'b000;

endmodule