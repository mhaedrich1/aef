module dtc_split25_bm74 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node114;

	assign outp = (inp[0]) ? node56 : node1;
		assign node1 = (inp[6]) ? node25 : node2;
			assign node2 = (inp[3]) ? node18 : node3;
				assign node3 = (inp[9]) ? node11 : node4;
					assign node4 = (inp[1]) ? node8 : node5;
						assign node5 = (inp[7]) ? 3'b111 : 3'b111;
						assign node8 = (inp[7]) ? 3'b001 : 3'b111;
					assign node11 = (inp[2]) ? node15 : node12;
						assign node12 = (inp[4]) ? 3'b111 : 3'b111;
						assign node15 = (inp[1]) ? 3'b111 : 3'b111;
				assign node18 = (inp[9]) ? 3'b111 : node19;
					assign node19 = (inp[1]) ? node21 : 3'b111;
						assign node21 = (inp[7]) ? 3'b111 : 3'b111;
			assign node25 = (inp[3]) ? node41 : node26;
				assign node26 = (inp[1]) ? node34 : node27;
					assign node27 = (inp[7]) ? node31 : node28;
						assign node28 = (inp[4]) ? 3'b111 : 3'b001;
						assign node31 = (inp[4]) ? 3'b001 : 3'b110;
					assign node34 = (inp[9]) ? node38 : node35;
						assign node35 = (inp[7]) ? 3'b000 : 3'b010;
						assign node38 = (inp[10]) ? 3'b000 : 3'b010;
				assign node41 = (inp[1]) ? node49 : node42;
					assign node42 = (inp[9]) ? node46 : node43;
						assign node43 = (inp[5]) ? 3'b111 : 3'b001;
						assign node46 = (inp[4]) ? 3'b111 : 3'b111;
					assign node49 = (inp[8]) ? node53 : node50;
						assign node50 = (inp[2]) ? 3'b101 : 3'b111;
						assign node53 = (inp[9]) ? 3'b101 : 3'b001;
		assign node56 = (inp[6]) ? node88 : node57;
			assign node57 = (inp[3]) ? node73 : node58;
				assign node58 = (inp[1]) ? node66 : node59;
					assign node59 = (inp[7]) ? node63 : node60;
						assign node60 = (inp[9]) ? 3'b101 : 3'b101;
						assign node63 = (inp[9]) ? 3'b100 : 3'b100;
					assign node66 = (inp[9]) ? node70 : node67;
						assign node67 = (inp[7]) ? 3'b000 : 3'b000;
						assign node70 = (inp[4]) ? 3'b000 : 3'b100;
				assign node73 = (inp[9]) ? node81 : node74;
					assign node74 = (inp[7]) ? node78 : node75;
						assign node75 = (inp[1]) ? 3'b001 : 3'b011;
						assign node78 = (inp[1]) ? 3'b010 : 3'b001;
					assign node81 = (inp[1]) ? node85 : node82;
						assign node82 = (inp[5]) ? 3'b111 : 3'b111;
						assign node85 = (inp[8]) ? 3'b001 : 3'b101;
			assign node88 = (inp[3]) ? node102 : node89;
				assign node89 = (inp[1]) ? node97 : node90;
					assign node90 = (inp[9]) ? node94 : node91;
						assign node91 = (inp[7]) ? 3'b000 : 3'b000;
						assign node94 = (inp[4]) ? 3'b100 : 3'b000;
					assign node97 = (inp[2]) ? 3'b000 : node98;
						assign node98 = (inp[5]) ? 3'b000 : 3'b000;
				assign node102 = (inp[7]) ? node110 : node103;
					assign node103 = (inp[9]) ? node107 : node104;
						assign node104 = (inp[1]) ? 3'b000 : 3'b110;
						assign node107 = (inp[1]) ? 3'b010 : 3'b101;
					assign node110 = (inp[1]) ? node114 : node111;
						assign node111 = (inp[10]) ? 3'b100 : 3'b000;
						assign node114 = (inp[9]) ? 3'b000 : 3'b000;

endmodule